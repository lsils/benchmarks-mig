module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 ;
  assign n61 = x23 & x24 ;
  assign n62 = x25 & n61 ;
  assign n63 = x27 & x28 ;
  assign n64 = x29 & n63 ;
  assign n65 = n62 & n64 ;
  assign n66 = x0 & x1 ;
  assign n67 = x6 & x7 ;
  assign n68 = x4 & x5 ;
  assign n69 = x2 & x3 ;
  assign n70 = ( ~n67 & n68 ) | ( ~n67 & n69 ) | ( n68 & n69 ) ;
  assign n71 = ( ~x8 & n67 ) | ( ~x8 & n70 ) | ( n67 & n70 ) ;
  assign n72 = ( x8 & ~n66 ) | ( x8 & n71 ) | ( ~n66 & n71 ) ;
  assign n73 = n66 & n72 ;
  assign n74 = x9 & x11 ;
  assign n75 = ( x11 & n73 ) | ( x11 & n74 ) | ( n73 & n74 ) ;
  assign n76 = x14 & x15 ;
  assign n77 = x19 & x20 ;
  assign n78 = x17 & n77 ;
  assign n79 = n76 & n78 ;
  assign n80 = ( ~n65 & n75 ) | ( ~n65 & n79 ) | ( n75 & n79 ) ;
  assign n81 = n65 & n80 ;
  assign n82 = x26 | n62 ;
  assign n83 = x21 | x22 ;
  assign n84 = x12 | x13 ;
  assign n85 = x11 | n84 ;
  assign n86 = x9 | x10 ;
  assign n87 = x1 | x2 ;
  assign n88 = x5 | x6 ;
  assign n89 = x7 | x8 ;
  assign n90 = ( ~n87 & n88 ) | ( ~n87 & n89 ) | ( n88 & n89 ) ;
  assign n91 = x3 | x4 ;
  assign n92 = ( ~n87 & n90 ) | ( ~n87 & n91 ) | ( n90 & n91 ) ;
  assign n93 = n87 | n92 ;
  assign n94 = ( x10 & n86 ) | ( x10 & n93 ) | ( n86 & n93 ) ;
  assign n95 = ( n84 & n85 ) | ( n84 & n94 ) | ( n85 & n94 ) ;
  assign n96 = n79 & n95 ;
  assign n97 = ( x16 & n78 ) | ( x16 & n96 ) | ( n78 & n96 ) ;
  assign n98 = ( x18 & n77 ) | ( x18 & n97 ) | ( n77 & n97 ) ;
  assign n99 = n83 | n98 ;
  assign n100 = ( x26 & n82 ) | ( x26 & n99 ) | ( n82 & n99 ) ;
  assign n101 = n81 & ~n100 ;
  assign n102 = x57 & x58 ;
  assign n103 = x59 & n102 ;
  assign n104 = x48 | x56 ;
  assign n105 = x43 | x46 ;
  assign n106 = n104 | n105 ;
  assign n107 = x40 | x42 ;
  assign n108 = x33 | x34 ;
  assign n109 = x35 | x36 ;
  assign n110 = x37 | x38 ;
  assign n111 = ( ~n107 & n109 ) | ( ~n107 & n110 ) | ( n109 & n110 ) ;
  assign n112 = ( ~n107 & n108 ) | ( ~n107 & n111 ) | ( n108 & n111 ) ;
  assign n113 = n107 | n112 ;
  assign n114 = x31 | x32 ;
  assign n115 = ~x0 & x30 ;
  assign n116 = x51 | x52 ;
  assign n117 = ( x30 & ~n115 ) | ( x30 & n116 ) | ( ~n115 & n116 ) ;
  assign n118 = n114 | n117 ;
  assign n119 = ( ~n106 & n113 ) | ( ~n106 & n118 ) | ( n113 & n118 ) ;
  assign n120 = n106 | n119 ;
  assign n121 = ( x0 & n103 ) | ( x0 & n115 ) | ( n103 & n115 ) ;
  assign n122 = ( n103 & n120 ) | ( n103 & n121 ) | ( n120 & n121 ) ;
  assign n123 = n81 & n122 ;
  assign n124 = x53 & x54 ;
  assign n125 = x55 & n124 ;
  assign n126 = x49 & x50 ;
  assign n127 = x44 & x45 ;
  assign n128 = n126 & n127 ;
  assign n129 = x31 & x32 ;
  assign n130 = ( n115 & ~n125 ) | ( n115 & n129 ) | ( ~n125 & n129 ) ;
  assign n131 = ( ~n125 & n128 ) | ( ~n125 & n130 ) | ( n128 & n130 ) ;
  assign n132 = n125 & n131 ;
  assign n133 = x48 & n126 ;
  assign n134 = x39 | n107 ;
  assign n135 = ( x41 & x42 ) | ( x41 & n134 ) | ( x42 & n134 ) ;
  assign n136 = x43 & n127 ;
  assign n137 = ( n127 & n135 ) | ( n127 & n136 ) | ( n135 & n136 ) ;
  assign n138 = x46 & x47 ;
  assign n139 = ( x47 & n137 ) | ( x47 & n138 ) | ( n137 & n138 ) ;
  assign n140 = ( n126 & n133 ) | ( n126 & n139 ) | ( n133 & n139 ) ;
  assign n141 = n116 | n140 ;
  assign n142 = x56 | n125 ;
  assign n143 = ( x56 & n141 ) | ( x56 & n142 ) | ( n141 & n142 ) ;
  assign n144 = x33 & x34 ;
  assign n145 = x35 & x36 ;
  assign n146 = x37 & x38 ;
  assign n147 = x41 & x47 ;
  assign n148 = ( ~n144 & n146 ) | ( ~n144 & n147 ) | ( n146 & n147 ) ;
  assign n149 = ( ~n144 & n145 ) | ( ~n144 & n148 ) | ( n145 & n148 ) ;
  assign n150 = n144 & n149 ;
  assign n151 = n132 & ~n150 ;
  assign n152 = ( n132 & n143 ) | ( n132 & ~n151 ) | ( n143 & ~n151 ) ;
  assign n153 = n123 & n152 ;
  assign n154 = ( n64 & n100 ) | ( n64 & n153 ) | ( n100 & n153 ) ;
  assign n155 = n103 & n120 ;
  assign n156 = n143 & n155 ;
  assign n157 = n101 & n156 ;
  assign y0 = ~n101 ;
  assign y1 = ~n154 ;
  assign y2 = n157 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
