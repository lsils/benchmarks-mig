module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 ;
  assign n33 = x1 & x2 ;
  assign n34 = ( x0 & ~x2 ) | ( x0 & n33 ) | ( ~x2 & n33 ) ;
  assign n35 = ( ~x1 & n33 ) | ( ~x1 & n34 ) | ( n33 & n34 ) ;
  assign n36 = x0 & ~n35 ;
  assign n37 = ( x23 & x24 ) | ( x23 & ~x26 ) | ( x24 & ~x26 ) ;
  assign n38 = ( x25 & ~x26 ) | ( x25 & n37 ) | ( ~x26 & n37 ) ;
  assign n39 = x24 & x25 ;
  assign n40 = x23 & ~x26 ;
  assign n41 = n39 & n40 ;
  assign n42 = x29 | x30 ;
  assign n43 = ~x27 & x28 ;
  assign n44 = ~n42 & n43 ;
  assign n45 = n41 & n44 ;
  assign n46 = x27 & x28 ;
  assign n47 = x29 & x30 ;
  assign n48 = n46 & n47 ;
  assign n49 = x23 | x26 ;
  assign n50 = n39 & ~n49 ;
  assign n51 = n48 & n50 ;
  assign n52 = n45 | n51 ;
  assign n53 = x27 | x28 ;
  assign n54 = n42 | n53 ;
  assign n55 = n41 & ~n54 ;
  assign n56 = x24 | x25 ;
  assign n57 = n40 & ~n56 ;
  assign n58 = x29 & ~x30 ;
  assign n59 = n46 & n58 ;
  assign n60 = n57 & n59 ;
  assign n61 = n55 | n60 ;
  assign n62 = n52 | n61 ;
  assign n63 = ~x23 & x26 ;
  assign n64 = ~n56 & n63 ;
  assign n65 = x24 & ~x25 ;
  assign n66 = n40 & n65 ;
  assign n67 = n41 & n48 ;
  assign n68 = n66 | n67 ;
  assign n69 = ( n48 & n64 ) | ( n48 & n68 ) | ( n64 & n68 ) ;
  assign n70 = ~x24 & x25 ;
  assign n71 = x23 & x26 ;
  assign n72 = n70 & n71 ;
  assign n73 = n43 & n47 ;
  assign n74 = n72 & n73 ;
  assign n75 = ~n49 & n65 ;
  assign n76 = n48 & n75 ;
  assign n77 = n74 | n76 ;
  assign n78 = n49 | n56 ;
  assign n79 = n48 & ~n78 ;
  assign n80 = n39 & n71 ;
  assign n81 = n73 & n80 ;
  assign n82 = n79 | n81 ;
  assign n83 = ~n49 & n70 ;
  assign n84 = n40 & n70 ;
  assign n85 = n48 & n84 ;
  assign n86 = ( n40 & ~n56 ) | ( n40 & n85 ) | ( ~n56 & n85 ) ;
  assign n87 = ( n48 & n83 ) | ( n48 & n86 ) | ( n83 & n86 ) ;
  assign n88 = n82 | n87 ;
  assign n89 = ( ~n69 & n77 ) | ( ~n69 & n88 ) | ( n77 & n88 ) ;
  assign n90 = n69 | n89 ;
  assign n91 = n59 & n75 ;
  assign n92 = n59 & n66 ;
  assign n93 = n91 | n92 ;
  assign n94 = ( ~n62 & n90 ) | ( ~n62 & n93 ) | ( n90 & n93 ) ;
  assign n95 = n62 | n94 ;
  assign n96 = ~x29 & x30 ;
  assign n97 = n46 & n96 ;
  assign n98 = n63 & n70 ;
  assign n99 = ( n80 & n97 ) | ( n80 & n98 ) | ( n97 & n98 ) ;
  assign n100 = n47 & ~n53 ;
  assign n101 = n84 & n100 ;
  assign n102 = n39 & n63 ;
  assign n103 = n97 & n102 ;
  assign n104 = n83 & n100 ;
  assign n105 = n103 | n104 ;
  assign n106 = ( ~n99 & n101 ) | ( ~n99 & n105 ) | ( n101 & n105 ) ;
  assign n107 = n99 | n106 ;
  assign n108 = x27 & ~x28 ;
  assign n109 = n96 & n108 ;
  assign n110 = ( n50 & n84 ) | ( n50 & n109 ) | ( n84 & n109 ) ;
  assign n111 = n57 & n100 ;
  assign n112 = n50 & ~n54 ;
  assign n113 = n111 | n112 ;
  assign n114 = n110 | n113 ;
  assign n115 = ~n54 & n84 ;
  assign n116 = n43 & n96 ;
  assign n117 = n72 & n116 ;
  assign n118 = n115 | n117 ;
  assign n119 = n47 & n108 ;
  assign n120 = n98 & n119 ;
  assign n121 = ( n98 & n116 ) | ( n98 & n120 ) | ( n116 & n120 ) ;
  assign n122 = n58 & n108 ;
  assign n123 = n64 & n122 ;
  assign n124 = ~n54 & n80 ;
  assign n125 = ( ~n121 & n123 ) | ( ~n121 & n124 ) | ( n123 & n124 ) ;
  assign n126 = n121 | n125 ;
  assign n127 = ( ~n114 & n118 ) | ( ~n114 & n126 ) | ( n118 & n126 ) ;
  assign n128 = n114 | n127 ;
  assign n129 = ~n56 & n71 ;
  assign n130 = ( n44 & n48 ) | ( n44 & n129 ) | ( n48 & n129 ) ;
  assign n131 = n66 & n109 ;
  assign n132 = n41 & n116 ;
  assign n133 = n131 | n132 ;
  assign n134 = n130 | n133 ;
  assign n135 = n59 & n84 ;
  assign n136 = ~n53 & n58 ;
  assign n137 = ~n78 & n136 ;
  assign n138 = ( n41 & n84 ) | ( n41 & n122 ) | ( n84 & n122 ) ;
  assign n139 = n137 | n138 ;
  assign n140 = n135 | n139 ;
  assign n141 = n134 | n140 ;
  assign n142 = n84 & n119 ;
  assign n143 = ( n119 & n129 ) | ( n119 & n142 ) | ( n129 & n142 ) ;
  assign n144 = n44 & ~n78 ;
  assign n145 = ~n42 & n108 ;
  assign n146 = n80 & n145 ;
  assign n147 = n144 | n146 ;
  assign n148 = n83 & n109 ;
  assign n149 = ~n53 & n96 ;
  assign n150 = n41 & n149 ;
  assign n151 = n148 | n150 ;
  assign n152 = n65 & n71 ;
  assign n153 = n116 & n152 ;
  assign n154 = n151 | n153 ;
  assign n155 = n147 | n154 ;
  assign n156 = n143 | n155 ;
  assign n157 = ( ~n128 & n141 ) | ( ~n128 & n156 ) | ( n141 & n156 ) ;
  assign n158 = n128 | n157 ;
  assign n159 = ( n59 & n64 ) | ( n59 & n149 ) | ( n64 & n149 ) ;
  assign n160 = ~n42 & n46 ;
  assign n161 = ( n75 & n149 ) | ( n75 & n160 ) | ( n149 & n160 ) ;
  assign n162 = n159 | n161 ;
  assign n163 = n83 & n160 ;
  assign n164 = n41 & n109 ;
  assign n165 = n163 | n164 ;
  assign n166 = n63 & n65 ;
  assign n167 = n48 & n166 ;
  assign n168 = ~n78 & n100 ;
  assign n169 = n167 | n168 ;
  assign n170 = n102 & n160 ;
  assign n171 = n57 & n136 ;
  assign n172 = n170 | n171 ;
  assign n173 = n50 & n149 ;
  assign n174 = n64 & n119 ;
  assign n175 = n173 | n174 ;
  assign n176 = n119 & n166 ;
  assign n177 = n50 & n145 ;
  assign n178 = n176 | n177 ;
  assign n179 = ( ~n172 & n175 ) | ( ~n172 & n178 ) | ( n175 & n178 ) ;
  assign n180 = ( ~n169 & n172 ) | ( ~n169 & n179 ) | ( n172 & n179 ) ;
  assign n181 = n169 | n180 ;
  assign n182 = ( ~n162 & n165 ) | ( ~n162 & n181 ) | ( n165 & n181 ) ;
  assign n183 = n162 | n182 ;
  assign n184 = ( n107 & n158 ) | ( n107 & ~n183 ) | ( n158 & ~n183 ) ;
  assign n185 = n50 & n116 ;
  assign n186 = n102 & n119 ;
  assign n187 = n185 | n186 ;
  assign n188 = n109 & n129 ;
  assign n189 = n102 & n145 ;
  assign n190 = n188 | n189 ;
  assign n191 = n187 | n190 ;
  assign n192 = n66 & n160 ;
  assign n193 = n50 & n122 ;
  assign n194 = n192 | n193 ;
  assign n195 = n119 & n152 ;
  assign n196 = n50 & n59 ;
  assign n197 = ~n54 & n64 ;
  assign n198 = n196 | n197 ;
  assign n199 = n195 | n198 ;
  assign n200 = ( ~n191 & n194 ) | ( ~n191 & n199 ) | ( n194 & n199 ) ;
  assign n201 = n191 | n200 ;
  assign n202 = n41 & n145 ;
  assign n203 = n83 & n149 ;
  assign n204 = n202 | n203 ;
  assign n205 = n64 & n109 ;
  assign n206 = n72 & n136 ;
  assign n207 = ~n78 & n145 ;
  assign n208 = n206 | n207 ;
  assign n209 = ( ~n204 & n205 ) | ( ~n204 & n208 ) | ( n205 & n208 ) ;
  assign n210 = n204 | n209 ;
  assign n211 = n122 & n129 ;
  assign n212 = n66 & n149 ;
  assign n213 = n211 | n212 ;
  assign n214 = ( n41 & n59 ) | ( n41 & n83 ) | ( n59 & n83 ) ;
  assign n215 = n116 & n166 ;
  assign n216 = n43 & n58 ;
  assign n217 = n129 & n216 ;
  assign n218 = n54 | n78 ;
  assign n219 = ~n217 & n218 ;
  assign n220 = ~n215 & n219 ;
  assign n221 = ( n213 & ~n214 ) | ( n213 & n220 ) | ( ~n214 & n220 ) ;
  assign n222 = ( n210 & ~n213 ) | ( n210 & n221 ) | ( ~n213 & n221 ) ;
  assign n223 = ~n210 & n222 ;
  assign n224 = n41 & n119 ;
  assign n225 = n84 & n149 ;
  assign n226 = n224 | n225 ;
  assign n227 = n116 & n129 ;
  assign n228 = n50 & n119 ;
  assign n229 = n227 | n228 ;
  assign n230 = n44 & n64 ;
  assign n231 = n66 & n100 ;
  assign n232 = n230 | n231 ;
  assign n233 = n72 & n119 ;
  assign n234 = n64 & n136 ;
  assign n235 = n233 | n234 ;
  assign n236 = n232 | n235 ;
  assign n237 = ( n226 & ~n229 ) | ( n226 & n236 ) | ( ~n229 & n236 ) ;
  assign n238 = n75 & n100 ;
  assign n239 = n64 & n116 ;
  assign n240 = n97 & n152 ;
  assign n241 = n72 & n97 ;
  assign n242 = n80 & n160 ;
  assign n243 = n241 | n242 ;
  assign n244 = n240 | n243 ;
  assign n245 = ( ~n238 & n239 ) | ( ~n238 & n244 ) | ( n239 & n244 ) ;
  assign n246 = n238 | n245 ;
  assign n247 = ( n229 & ~n237 ) | ( n229 & n246 ) | ( ~n237 & n246 ) ;
  assign n248 = n237 | n247 ;
  assign n249 = ( n201 & n223 ) | ( n201 & ~n248 ) | ( n223 & ~n248 ) ;
  assign n250 = ~n201 & n249 ;
  assign n251 = ( ~n183 & n184 ) | ( ~n183 & n250 ) | ( n184 & n250 ) ;
  assign n252 = ~n184 & n251 ;
  assign n253 = ( n44 & n152 ) | ( n44 & n166 ) | ( n152 & n166 ) ;
  assign n254 = n72 & n160 ;
  assign n255 = n64 & n145 ;
  assign n256 = n254 | n255 ;
  assign n257 = n253 | n256 ;
  assign n258 = n102 & n116 ;
  assign n259 = n50 & n100 ;
  assign n260 = n258 | n259 ;
  assign n261 = ~n54 & n72 ;
  assign n262 = n109 & n152 ;
  assign n263 = n261 | n262 ;
  assign n264 = n260 | n263 ;
  assign n265 = n80 & n116 ;
  assign n266 = n73 & n102 ;
  assign n267 = n84 & n145 ;
  assign n268 = n266 | n267 ;
  assign n269 = n265 | n268 ;
  assign n270 = ( n257 & ~n264 ) | ( n257 & n269 ) | ( ~n264 & n269 ) ;
  assign n271 = ( n50 & n66 ) | ( n50 & n216 ) | ( n66 & n216 ) ;
  assign n272 = n50 & n160 ;
  assign n273 = n66 & n119 ;
  assign n274 = n272 | n273 ;
  assign n275 = ( n64 & n83 ) | ( n64 & n216 ) | ( n83 & n216 ) ;
  assign n276 = ( n271 & ~n274 ) | ( n271 & n275 ) | ( ~n274 & n275 ) ;
  assign n277 = n57 & n149 ;
  assign n278 = ( n84 & n160 ) | ( n84 & n216 ) | ( n160 & n216 ) ;
  assign n279 = n277 | n278 ;
  assign n280 = ( n274 & ~n276 ) | ( n274 & n279 ) | ( ~n276 & n279 ) ;
  assign n281 = n276 | n280 ;
  assign n282 = ( n264 & ~n270 ) | ( n264 & n281 ) | ( ~n270 & n281 ) ;
  assign n283 = n270 | n282 ;
  assign n284 = ( n95 & n252 ) | ( n95 & n283 ) | ( n252 & n283 ) ;
  assign n285 = n41 & n216 ;
  assign n286 = n136 & n152 ;
  assign n287 = n285 | n286 ;
  assign n288 = ( n98 & n136 ) | ( n98 & n166 ) | ( n136 & n166 ) ;
  assign n289 = n287 | n288 ;
  assign n290 = n83 & n119 ;
  assign n291 = n129 & n136 ;
  assign n292 = n290 | n291 ;
  assign n293 = n44 & n75 ;
  assign n294 = n122 & n166 ;
  assign n295 = n73 & n98 ;
  assign n296 = n294 | n295 ;
  assign n297 = n293 | n296 ;
  assign n298 = ~n54 & n102 ;
  assign n299 = n122 & n152 ;
  assign n300 = n44 & n57 ;
  assign n301 = n109 & n166 ;
  assign n302 = n129 & n149 ;
  assign n303 = n301 | n302 ;
  assign n304 = n300 | n303 ;
  assign n305 = n299 | n304 ;
  assign n306 = ( ~n297 & n298 ) | ( ~n297 & n305 ) | ( n298 & n305 ) ;
  assign n307 = n297 | n306 ;
  assign n308 = ( ~n289 & n292 ) | ( ~n289 & n307 ) | ( n292 & n307 ) ;
  assign n309 = n289 | n308 ;
  assign n310 = ( n252 & n284 ) | ( n252 & ~n309 ) | ( n284 & ~n309 ) ;
  assign n311 = ~n284 & n310 ;
  assign n312 = ~n54 & n83 ;
  assign n313 = n111 | n240 ;
  assign n314 = n312 | n313 ;
  assign n315 = ( n80 & n100 ) | ( n80 & n166 ) | ( n100 & n166 ) ;
  assign n316 = n100 & n102 ;
  assign n317 = n75 & n119 ;
  assign n318 = n316 | n317 ;
  assign n319 = n315 | n318 ;
  assign n320 = n100 & n152 ;
  assign n321 = n290 | n320 ;
  assign n322 = n143 | n321 ;
  assign n323 = ( n119 & n152 ) | ( n119 & n228 ) | ( n152 & n228 ) ;
  assign n324 = ( ~n319 & n322 ) | ( ~n319 & n323 ) | ( n322 & n323 ) ;
  assign n325 = n319 | n324 ;
  assign n326 = ( n54 & ~n57 ) | ( n54 & n78 ) | ( ~n57 & n78 ) ;
  assign n327 = ( ~n78 & n119 ) | ( ~n78 & n273 ) | ( n119 & n273 ) ;
  assign n328 = n98 & n100 ;
  assign n329 = n64 & n100 ;
  assign n330 = n176 | n329 ;
  assign n331 = n72 & n100 ;
  assign n332 = n224 | n331 ;
  assign n333 = n330 | n332 ;
  assign n334 = n174 | n333 ;
  assign n335 = ( ~n327 & n328 ) | ( ~n327 & n334 ) | ( n328 & n334 ) ;
  assign n336 = n327 | n335 ;
  assign n337 = n100 & n129 ;
  assign n338 = n57 & n119 ;
  assign n339 = n337 | n338 ;
  assign n340 = ( ~n54 & n66 ) | ( ~n54 & n75 ) | ( n66 & n75 ) ;
  assign n341 = ( ~n336 & n339 ) | ( ~n336 & n340 ) | ( n339 & n340 ) ;
  assign n342 = n336 | n341 ;
  assign n343 = ( n325 & n326 ) | ( n325 & ~n342 ) | ( n326 & ~n342 ) ;
  assign n344 = ~n325 & n343 ;
  assign n345 = ~n314 & n344 ;
  assign n346 = ( n50 & n73 ) | ( n50 & n84 ) | ( n73 & n84 ) ;
  assign n347 = ( n73 & n75 ) | ( n73 & n166 ) | ( n75 & n166 ) ;
  assign n348 = n57 & n73 ;
  assign n349 = n120 | n348 ;
  assign n350 = ( ~n346 & n347 ) | ( ~n346 & n349 ) | ( n347 & n349 ) ;
  assign n351 = n346 | n350 ;
  assign n352 = n73 & n129 ;
  assign n353 = n80 & n119 ;
  assign n354 = n352 | n353 ;
  assign n355 = ( n66 & n73 ) | ( n66 & ~n78 ) | ( n73 & ~n78 ) ;
  assign n356 = n64 & n73 ;
  assign n357 = ( n73 & n83 ) | ( n73 & n356 ) | ( n83 & n356 ) ;
  assign n358 = ( ~n354 & n355 ) | ( ~n354 & n357 ) | ( n355 & n357 ) ;
  assign n359 = n354 | n358 ;
  assign n360 = n41 & n73 ;
  assign n361 = n73 & n152 ;
  assign n362 = n186 | n361 ;
  assign n363 = ( n233 & ~n360 ) | ( n233 & n362 ) | ( ~n360 & n362 ) ;
  assign n364 = n360 | n363 ;
  assign n365 = ( ~n351 & n359 ) | ( ~n351 & n364 ) | ( n359 & n364 ) ;
  assign n366 = n351 | n365 ;
  assign n367 = n41 & n100 ;
  assign n368 = n241 | n367 ;
  assign n369 = ( n50 & ~n78 ) | ( n50 & n100 ) | ( ~n78 & n100 ) ;
  assign n370 = ( n66 & n75 ) | ( n66 & n100 ) | ( n75 & n100 ) ;
  assign n371 = n369 | n370 ;
  assign n372 = n107 | n371 ;
  assign n373 = n368 | n372 ;
  assign n374 = ( n345 & n366 ) | ( n345 & n373 ) | ( n366 & n373 ) ;
  assign n375 = n345 & ~n374 ;
  assign n376 = ( n57 & n75 ) | ( n57 & n109 ) | ( n75 & n109 ) ;
  assign n377 = ( n41 & n59 ) | ( n41 & n84 ) | ( n59 & n84 ) ;
  assign n378 = ( n50 & n59 ) | ( n50 & n377 ) | ( n59 & n377 ) ;
  assign n379 = ( n57 & n59 ) | ( n57 & n66 ) | ( n59 & n66 ) ;
  assign n380 = ( n59 & n75 ) | ( n59 & n379 ) | ( n75 & n379 ) ;
  assign n381 = n378 | n380 ;
  assign n382 = ( n59 & n64 ) | ( n59 & n83 ) | ( n64 & n83 ) ;
  assign n383 = ( n50 & n57 ) | ( n50 & n149 ) | ( n57 & n149 ) ;
  assign n384 = ( n98 & n129 ) | ( n98 & n149 ) | ( n129 & n149 ) ;
  assign n385 = n383 | n384 ;
  assign n386 = ( n64 & n102 ) | ( n64 & n149 ) | ( n102 & n149 ) ;
  assign n387 = ( ~n78 & n149 ) | ( ~n78 & n166 ) | ( n149 & n166 ) ;
  assign n388 = ( n41 & n75 ) | ( n41 & n149 ) | ( n75 & n149 ) ;
  assign n389 = ( n80 & n149 ) | ( n80 & n152 ) | ( n149 & n152 ) ;
  assign n390 = n388 | n389 ;
  assign n391 = ( n225 & ~n387 ) | ( n225 & n390 ) | ( ~n387 & n390 ) ;
  assign n392 = n387 | n391 ;
  assign n393 = ( n66 & n83 ) | ( n66 & n149 ) | ( n83 & n149 ) ;
  assign n394 = n72 & n149 ;
  assign n395 = n59 & n80 ;
  assign n396 = n394 | n395 ;
  assign n397 = ( ~n392 & n393 ) | ( ~n392 & n396 ) | ( n393 & n396 ) ;
  assign n398 = n392 | n397 ;
  assign n399 = ( ~n385 & n386 ) | ( ~n385 & n398 ) | ( n386 & n398 ) ;
  assign n400 = n385 | n399 ;
  assign n401 = ( n59 & n129 ) | ( n59 & n152 ) | ( n129 & n152 ) ;
  assign n402 = ( n59 & n98 ) | ( n59 & n102 ) | ( n98 & n102 ) ;
  assign n403 = ( n59 & n72 ) | ( n59 & n166 ) | ( n72 & n166 ) ;
  assign n404 = n402 | n403 ;
  assign n405 = ( ~n400 & n401 ) | ( ~n400 & n404 ) | ( n401 & n404 ) ;
  assign n406 = n400 | n405 ;
  assign n407 = ( ~n381 & n382 ) | ( ~n381 & n406 ) | ( n382 & n406 ) ;
  assign n408 = n381 | n407 ;
  assign n409 = ( n41 & n129 ) | ( n41 & n145 ) | ( n129 & n145 ) ;
  assign n410 = ~x25 & n63 ;
  assign n411 = ( n50 & n145 ) | ( n50 & n410 ) | ( n145 & n410 ) ;
  assign n412 = n409 | n411 ;
  assign n413 = n267 | n412 ;
  assign n414 = n408 | n413 ;
  assign n415 = n376 | n414 ;
  assign n416 = ( n64 & n83 ) | ( n64 & n136 ) | ( n83 & n136 ) ;
  assign n417 = ( n50 & n72 ) | ( n50 & n136 ) | ( n72 & n136 ) ;
  assign n418 = n416 | n417 ;
  assign n419 = ( n98 & n136 ) | ( n98 & n152 ) | ( n136 & n152 ) ;
  assign n420 = ( n41 & n84 ) | ( n41 & n136 ) | ( n84 & n136 ) ;
  assign n421 = ( n80 & n136 ) | ( n80 & n420 ) | ( n136 & n420 ) ;
  assign n422 = ( n66 & n129 ) | ( n66 & n136 ) | ( n129 & n136 ) ;
  assign n423 = n137 | n242 ;
  assign n424 = ( ~n172 & n422 ) | ( ~n172 & n423 ) | ( n422 & n423 ) ;
  assign n425 = ( n172 & ~n421 ) | ( n172 & n424 ) | ( ~n421 & n424 ) ;
  assign n426 = n421 | n425 ;
  assign n427 = ( ~n418 & n419 ) | ( ~n418 & n426 ) | ( n419 & n426 ) ;
  assign n428 = n418 | n427 ;
  assign n429 = n189 | n300 ;
  assign n430 = ( n66 & n75 ) | ( n66 & n122 ) | ( n75 & n122 ) ;
  assign n431 = n429 | n430 ;
  assign n432 = n147 | n431 ;
  assign n433 = n57 & n122 ;
  assign n434 = n293 | n433 ;
  assign n435 = n102 & n136 ;
  assign n436 = ( ~n78 & n83 ) | ( ~n78 & n122 ) | ( n83 & n122 ) ;
  assign n437 = n435 | n436 ;
  assign n438 = ( ~n432 & n434 ) | ( ~n432 & n437 ) | ( n434 & n437 ) ;
  assign n439 = n432 | n438 ;
  assign n440 = n44 & n66 ;
  assign n441 = ( n44 & n50 ) | ( n44 & n83 ) | ( n50 & n83 ) ;
  assign n442 = n440 | n441 ;
  assign n443 = ( ~n428 & n439 ) | ( ~n428 & n442 ) | ( n439 & n442 ) ;
  assign n444 = n72 & n145 ;
  assign n445 = n75 & n136 ;
  assign n446 = n444 | n445 ;
  assign n447 = n44 & n84 ;
  assign n448 = n136 & n166 ;
  assign n449 = n447 | n448 ;
  assign n450 = ( n98 & n145 ) | ( n98 & n152 ) | ( n145 & n152 ) ;
  assign n451 = ( ~n446 & n449 ) | ( ~n446 & n450 ) | ( n449 & n450 ) ;
  assign n452 = n446 | n451 ;
  assign n453 = ( n428 & ~n443 ) | ( n428 & n452 ) | ( ~n443 & n452 ) ;
  assign n454 = n443 | n453 ;
  assign n455 = ~n78 & n109 ;
  assign n456 = n254 | n455 ;
  assign n457 = ( ~n376 & n454 ) | ( ~n376 & n456 ) | ( n454 & n456 ) ;
  assign n458 = ( n375 & n415 ) | ( n375 & n457 ) | ( n415 & n457 ) ;
  assign n459 = n375 & ~n458 ;
  assign n460 = ( n38 & n311 ) | ( n38 & n459 ) | ( n311 & n459 ) ;
  assign n461 = ( ~n38 & n311 ) | ( ~n38 & n459 ) | ( n311 & n459 ) ;
  assign n462 = ( n38 & ~n460 ) | ( n38 & n461 ) | ( ~n460 & n461 ) ;
  assign n463 = ( n50 & ~n54 ) | ( n50 & n84 ) | ( ~n54 & n84 ) ;
  assign n464 = n296 | n463 ;
  assign n465 = n72 & n122 ;
  assign n466 = ( n50 & n122 ) | ( n50 & n152 ) | ( n122 & n152 ) ;
  assign n467 = ( n266 & ~n465 ) | ( n266 & n466 ) | ( ~n465 & n466 ) ;
  assign n468 = n465 | n467 ;
  assign n469 = ( ~n56 & n71 ) | ( ~n56 & n123 ) | ( n71 & n123 ) ;
  assign n470 = ( n98 & n122 ) | ( n98 & n469 ) | ( n122 & n469 ) ;
  assign n471 = ( ~n464 & n468 ) | ( ~n464 & n470 ) | ( n468 & n470 ) ;
  assign n472 = n464 | n471 ;
  assign n473 = n95 | n472 ;
  assign n474 = n101 | n317 ;
  assign n475 = n402 | n474 ;
  assign n476 = n262 | n382 ;
  assign n477 = ( n232 & ~n475 ) | ( n232 & n476 ) | ( ~n475 & n476 ) ;
  assign n478 = n475 | n477 ;
  assign n479 = n57 & n116 ;
  assign n480 = n137 | n331 ;
  assign n481 = n479 | n480 ;
  assign n482 = n48 & n102 ;
  assign n483 = n50 & n109 ;
  assign n484 = n482 | n483 ;
  assign n485 = ~n78 & n216 ;
  assign n486 = ( n328 & ~n484 ) | ( n328 & n485 ) | ( ~n484 & n485 ) ;
  assign n487 = n484 | n486 ;
  assign n488 = n44 & n98 ;
  assign n489 = n102 & n109 ;
  assign n490 = n313 | n489 ;
  assign n491 = n488 | n490 ;
  assign n492 = n80 & n109 ;
  assign n493 = n83 & n136 ;
  assign n494 = n492 | n493 ;
  assign n495 = ( n196 & ~n491 ) | ( n196 & n494 ) | ( ~n491 & n494 ) ;
  assign n496 = n491 | n495 ;
  assign n497 = ( ~n481 & n487 ) | ( ~n481 & n496 ) | ( n487 & n496 ) ;
  assign n498 = n481 | n497 ;
  assign n499 = n177 | n205 ;
  assign n500 = n75 & n216 ;
  assign n501 = n339 | n500 ;
  assign n502 = ( n243 & ~n499 ) | ( n243 & n501 ) | ( ~n499 & n501 ) ;
  assign n503 = n499 | n502 ;
  assign n504 = ( n48 & n98 ) | ( n48 & n166 ) | ( n98 & n166 ) ;
  assign n505 = n57 & n216 ;
  assign n506 = n504 | n505 ;
  assign n507 = ~n54 & n166 ;
  assign n508 = ( n445 & ~n506 ) | ( n445 & n507 ) | ( ~n506 & n507 ) ;
  assign n509 = n506 | n508 ;
  assign n510 = n503 | n509 ;
  assign n511 = ( n478 & n498 ) | ( n478 & ~n510 ) | ( n498 & ~n510 ) ;
  assign n512 = n48 & n152 ;
  assign n513 = n202 | n512 ;
  assign n514 = n98 & n109 ;
  assign n515 = n513 | n514 ;
  assign n516 = n301 | n395 ;
  assign n517 = n59 & n166 ;
  assign n518 = n320 | n517 ;
  assign n519 = n66 & n136 ;
  assign n520 = ( n41 & n75 ) | ( n41 & n100 ) | ( n75 & n100 ) ;
  assign n521 = n519 | n520 ;
  assign n522 = ( ~n516 & n518 ) | ( ~n516 & n521 ) | ( n518 & n521 ) ;
  assign n523 = n48 & n80 ;
  assign n524 = n104 | n523 ;
  assign n525 = n255 | n524 ;
  assign n526 = ( n516 & ~n522 ) | ( n516 & n525 ) | ( ~n522 & n525 ) ;
  assign n527 = n522 | n526 ;
  assign n528 = n59 & n72 ;
  assign n529 = n75 & n116 ;
  assign n530 = n528 | n529 ;
  assign n531 = ( ~n515 & n527 ) | ( ~n515 & n530 ) | ( n527 & n530 ) ;
  assign n532 = n515 | n531 ;
  assign n533 = n172 | n253 ;
  assign n534 = n59 & n152 ;
  assign n535 = n316 | n534 ;
  assign n536 = ~n78 & n119 ;
  assign n537 = n84 & n109 ;
  assign n538 = n536 | n537 ;
  assign n539 = n535 | n538 ;
  assign n540 = ~n54 & n129 ;
  assign n541 = n103 | n540 ;
  assign n542 = ( n70 & n71 ) | ( n70 & n148 ) | ( n71 & n148 ) ;
  assign n543 = ( n66 & n109 ) | ( n66 & n542 ) | ( n109 & n542 ) ;
  assign n544 = n48 & n72 ;
  assign n545 = n100 & n166 ;
  assign n546 = n544 | n545 ;
  assign n547 = ( ~n541 & n543 ) | ( ~n541 & n546 ) | ( n543 & n546 ) ;
  assign n548 = n541 | n547 ;
  assign n549 = n59 & n129 ;
  assign n550 = n102 & n122 ;
  assign n551 = n549 | n550 ;
  assign n552 = n130 | n551 ;
  assign n553 = ( ~n539 & n548 ) | ( ~n539 & n552 ) | ( n548 & n552 ) ;
  assign n554 = n539 | n553 ;
  assign n555 = ( n50 & n64 ) | ( n50 & n100 ) | ( n64 & n100 ) ;
  assign n556 = n41 | n145 ;
  assign n557 = ( n109 & n129 ) | ( n109 & n556 ) | ( n129 & n556 ) ;
  assign n558 = ( n377 & ~n555 ) | ( n377 & n557 ) | ( ~n555 & n557 ) ;
  assign n559 = n555 | n558 ;
  assign n560 = ( ~n533 & n554 ) | ( ~n533 & n559 ) | ( n554 & n559 ) ;
  assign n561 = n533 | n560 ;
  assign n562 = ~n78 & n116 ;
  assign n563 = n168 | n197 ;
  assign n564 = n562 | n563 ;
  assign n565 = n80 & n100 ;
  assign n566 = ~n78 & n149 ;
  assign n567 = n80 & n122 ;
  assign n568 = n99 | n567 ;
  assign n569 = n566 | n568 ;
  assign n570 = ( ~n564 & n565 ) | ( ~n564 & n569 ) | ( n565 & n569 ) ;
  assign n571 = n564 | n570 ;
  assign n572 = ( ~n532 & n561 ) | ( ~n532 & n571 ) | ( n561 & n571 ) ;
  assign n573 = n532 | n572 ;
  assign n574 = ( n510 & ~n511 ) | ( n510 & n573 ) | ( ~n511 & n573 ) ;
  assign n575 = n511 | n574 ;
  assign n576 = n44 & n102 ;
  assign n577 = n444 | n576 ;
  assign n578 = ( ~n254 & n267 ) | ( ~n254 & n577 ) | ( n267 & n577 ) ;
  assign n579 = n254 | n578 ;
  assign n580 = ( ~n54 & n98 ) | ( ~n54 & n152 ) | ( n98 & n152 ) ;
  assign n581 = n83 & n116 ;
  assign n582 = ~n78 & n160 ;
  assign n583 = n581 | n582 ;
  assign n584 = ( ~n579 & n580 ) | ( ~n579 & n583 ) | ( n580 & n583 ) ;
  assign n585 = n579 | n584 ;
  assign n586 = n84 & n116 ;
  assign n587 = n44 & n72 ;
  assign n588 = n138 | n587 ;
  assign n589 = n586 | n588 ;
  assign n590 = n66 & n116 ;
  assign n591 = n57 & n160 ;
  assign n592 = n84 & n136 ;
  assign n593 = ( ~n590 & n591 ) | ( ~n590 & n592 ) | ( n591 & n592 ) ;
  assign n594 = n590 | n593 ;
  assign n595 = n145 & n166 ;
  assign n596 = ( n41 & n50 ) | ( n41 & n136 ) | ( n50 & n136 ) ;
  assign n597 = n595 | n596 ;
  assign n598 = n594 | n597 ;
  assign n599 = n44 & n80 ;
  assign n600 = n450 | n599 ;
  assign n601 = n598 | n600 ;
  assign n602 = ( ~n585 & n589 ) | ( ~n585 & n601 ) | ( n589 & n601 ) ;
  assign n603 = n585 | n602 ;
  assign n604 = ( ~n473 & n575 ) | ( ~n473 & n603 ) | ( n575 & n603 ) ;
  assign n605 = n473 | n604 ;
  assign n606 = ( ~x31 & n58 ) | ( ~x31 & n96 ) | ( n58 & n96 ) ;
  assign n607 = x31 & n47 ;
  assign n608 = n435 | n567 ;
  assign n609 = n149 & n152 ;
  assign n610 = n565 | n609 ;
  assign n611 = n608 | n610 ;
  assign n612 = n286 | n447 ;
  assign n613 = n59 & ~n78 ;
  assign n614 = n225 | n613 ;
  assign n615 = ( n142 & n255 ) | ( n142 & ~n614 ) | ( n255 & ~n614 ) ;
  assign n616 = n614 | n615 ;
  assign n617 = ( ~n378 & n546 ) | ( ~n378 & n616 ) | ( n546 & n616 ) ;
  assign n618 = ( n376 & n378 ) | ( n376 & ~n617 ) | ( n378 & ~n617 ) ;
  assign n619 = n617 | n618 ;
  assign n620 = ( ~n611 & n612 ) | ( ~n611 & n619 ) | ( n612 & n619 ) ;
  assign n621 = n611 | n620 ;
  assign n622 = ( n98 & n145 ) | ( n98 & n160 ) | ( n145 & n160 ) ;
  assign n623 = ( n448 & ~n621 ) | ( n448 & n622 ) | ( ~n621 & n622 ) ;
  assign n624 = n621 | n623 ;
  assign n625 = n258 | n294 ;
  assign n626 = n208 | n590 ;
  assign n627 = n625 | n626 ;
  assign n628 = ( n50 & n116 ) | ( n50 & n152 ) | ( n116 & n152 ) ;
  assign n629 = n159 | n628 ;
  assign n630 = ( n57 & ~n78 ) | ( n57 & n216 ) | ( ~n78 & n216 ) ;
  assign n631 = n197 | n630 ;
  assign n632 = n582 | n631 ;
  assign n633 = n92 | n331 ;
  assign n634 = n170 | n633 ;
  assign n635 = ( ~n629 & n632 ) | ( ~n629 & n634 ) | ( n632 & n634 ) ;
  assign n636 = n629 | n635 ;
  assign n637 = ( n98 & n102 ) | ( n98 & n149 ) | ( n102 & n149 ) ;
  assign n638 = n44 & n83 ;
  assign n639 = n132 | n638 ;
  assign n640 = n637 | n639 ;
  assign n641 = n98 & n122 ;
  assign n642 = n129 & n145 ;
  assign n643 = n581 | n642 ;
  assign n644 = ( ~n504 & n641 ) | ( ~n504 & n643 ) | ( n641 & n643 ) ;
  assign n645 = ( n55 & n504 ) | ( n55 & ~n644 ) | ( n504 & ~n644 ) ;
  assign n646 = n644 | n645 ;
  assign n647 = ( n75 & n145 ) | ( n75 & n160 ) | ( n145 & n160 ) ;
  assign n648 = ( n41 & n100 ) | ( n41 & n129 ) | ( n100 & n129 ) ;
  assign n649 = n647 | n648 ;
  assign n650 = ( ~n640 & n646 ) | ( ~n640 & n649 ) | ( n646 & n649 ) ;
  assign n651 = n640 | n650 ;
  assign n652 = ( n627 & ~n636 ) | ( n627 & n651 ) | ( ~n636 & n651 ) ;
  assign n653 = n80 & n149 ;
  assign n654 = n455 | n653 ;
  assign n655 = n59 & n83 ;
  assign n656 = n482 | n655 ;
  assign n657 = n48 & n129 ;
  assign n658 = n137 | n657 ;
  assign n659 = ( ~n654 & n656 ) | ( ~n654 & n658 ) | ( n656 & n658 ) ;
  assign n660 = n654 | n659 ;
  assign n661 = n48 & n64 ;
  assign n662 = n75 & n97 ;
  assign n663 = n224 | n662 ;
  assign n664 = n661 | n663 ;
  assign n665 = ( n80 & n116 ) | ( n80 & n166 ) | ( n116 & n166 ) ;
  assign n666 = n160 & n166 ;
  assign n667 = n218 & ~n666 ;
  assign n668 = ( n664 & ~n665 ) | ( n664 & n667 ) | ( ~n665 & n667 ) ;
  assign n669 = ~n664 & n668 ;
  assign n670 = ( ~n292 & n660 ) | ( ~n292 & n669 ) | ( n660 & n669 ) ;
  assign n671 = ~n660 & n670 ;
  assign n672 = ( ~n636 & n652 ) | ( ~n636 & n671 ) | ( n652 & n671 ) ;
  assign n673 = ~n652 & n672 ;
  assign n674 = n91 | n599 ;
  assign n675 = n98 & n116 ;
  assign n676 = n173 | n675 ;
  assign n677 = ( n117 & ~n674 ) | ( n117 & n676 ) | ( ~n674 & n676 ) ;
  assign n678 = n674 | n677 ;
  assign n679 = ( n48 & n80 ) | ( n48 & n152 ) | ( n80 & n152 ) ;
  assign n680 = x25 & n71 ;
  assign n681 = n216 & ~n680 ;
  assign n682 = ( n216 & n679 ) | ( n216 & ~n681 ) | ( n679 & ~n681 ) ;
  assign n683 = n678 | n682 ;
  assign n684 = n227 | n394 ;
  assign n685 = n102 & n216 ;
  assign n686 = n242 | n685 ;
  assign n687 = n684 | n686 ;
  assign n688 = ( n57 & n119 ) | ( n57 & n160 ) | ( n119 & n160 ) ;
  assign n689 = ~n78 & n122 ;
  assign n690 = n254 | n689 ;
  assign n691 = n57 & n97 ;
  assign n692 = n320 | n691 ;
  assign n693 = n690 | n692 ;
  assign n694 = n688 | n693 ;
  assign n695 = ( ~n682 & n687 ) | ( ~n682 & n694 ) | ( n687 & n694 ) ;
  assign n696 = n119 & n129 ;
  assign n697 = n145 & n152 ;
  assign n698 = n696 | n697 ;
  assign n699 = n318 | n698 ;
  assign n700 = ( ~n54 & n57 ) | ( ~n54 & n59 ) | ( n57 & n59 ) ;
  assign n701 = n239 | n700 ;
  assign n702 = n174 | n595 ;
  assign n703 = n293 | n536 ;
  assign n704 = ( ~n701 & n702 ) | ( ~n701 & n703 ) | ( n702 & n703 ) ;
  assign n705 = n701 | n704 ;
  assign n706 = ( n80 & n98 ) | ( n80 & n136 ) | ( n98 & n136 ) ;
  assign n707 = ( n176 & n500 ) | ( n176 & ~n706 ) | ( n500 & ~n706 ) ;
  assign n708 = n706 | n707 ;
  assign n709 = ( ~n699 & n705 ) | ( ~n699 & n708 ) | ( n705 & n708 ) ;
  assign n710 = n699 | n709 ;
  assign n711 = ( n683 & n695 ) | ( n683 & ~n710 ) | ( n695 & ~n710 ) ;
  assign n712 = n124 | n587 ;
  assign n713 = n152 & n160 ;
  assign n714 = ( n150 & ~n712 ) | ( n150 & n713 ) | ( ~n712 & n713 ) ;
  assign n715 = n712 | n714 ;
  assign n716 = n112 | n440 ;
  assign n717 = n44 | n48 ;
  assign n718 = ( n50 & n716 ) | ( n50 & n717 ) | ( n716 & n717 ) ;
  assign n719 = n57 & n145 ;
  assign n720 = n195 | n719 ;
  assign n721 = n540 | n550 ;
  assign n722 = n720 | n721 ;
  assign n723 = n228 | n329 ;
  assign n724 = ( n302 & n576 ) | ( n302 & ~n723 ) | ( n576 & ~n723 ) ;
  assign n725 = n723 | n724 ;
  assign n726 = n67 | n328 ;
  assign n727 = n586 | n726 ;
  assign n728 = ( ~n722 & n725 ) | ( ~n722 & n727 ) | ( n725 & n727 ) ;
  assign n729 = n722 | n728 ;
  assign n730 = ( n72 & n122 ) | ( n72 & n152 ) | ( n122 & n152 ) ;
  assign n731 = n259 | n730 ;
  assign n732 = ~n78 & n97 ;
  assign n733 = n529 | n732 ;
  assign n734 = n149 & n166 ;
  assign n735 = ( n273 & ~n733 ) | ( n273 & n734 ) | ( ~n733 & n734 ) ;
  assign n736 = n733 | n735 ;
  assign n737 = ( ~n718 & n731 ) | ( ~n718 & n736 ) | ( n731 & n736 ) ;
  assign n738 = n729 | n737 ;
  assign n739 = ( ~n715 & n718 ) | ( ~n715 & n738 ) | ( n718 & n738 ) ;
  assign n740 = n715 | n739 ;
  assign n741 = ( n710 & ~n711 ) | ( n710 & n740 ) | ( ~n711 & n740 ) ;
  assign n742 = n711 | n741 ;
  assign n743 = ( n624 & n673 ) | ( n624 & ~n742 ) | ( n673 & ~n742 ) ;
  assign n744 = ~n624 & n743 ;
  assign n745 = n112 | n545 ;
  assign n746 = n75 & n122 ;
  assign n747 = ( n75 & n216 ) | ( n75 & n746 ) | ( n216 & n746 ) ;
  assign n748 = n745 | n747 ;
  assign n749 = n173 | n523 ;
  assign n750 = n91 | n174 ;
  assign n751 = n749 | n750 ;
  assign n752 = n748 | n751 ;
  assign n753 = n73 & n84 ;
  assign n754 = n48 | n64 ;
  assign n755 = ( n44 & n152 ) | ( n44 & n754 ) | ( n152 & n754 ) ;
  assign n756 = n753 | n755 ;
  assign n757 = ( n48 & n129 ) | ( n48 & n136 ) | ( n129 & n136 ) ;
  assign n758 = n197 | n757 ;
  assign n759 = n83 & n97 ;
  assign n760 = n59 & n64 ;
  assign n761 = n759 | n760 ;
  assign n762 = n50 & n216 ;
  assign n763 = n186 | n762 ;
  assign n764 = n98 & n136 ;
  assign n765 = ( n254 & ~n763 ) | ( n254 & n764 ) | ( ~n763 & n764 ) ;
  assign n766 = n763 | n765 ;
  assign n767 = ( ~n758 & n761 ) | ( ~n758 & n766 ) | ( n761 & n766 ) ;
  assign n768 = ( ~n756 & n758 ) | ( ~n756 & n767 ) | ( n758 & n767 ) ;
  assign n769 = n534 | n662 ;
  assign n770 = ( n124 & ~n766 ) | ( n124 & n769 ) | ( ~n766 & n769 ) ;
  assign n771 = n756 | n770 ;
  assign n772 = n768 | n771 ;
  assign n773 = n519 | n732 ;
  assign n774 = n294 | n773 ;
  assign n775 = n50 & n136 ;
  assign n776 = n638 | n775 ;
  assign n777 = n98 & n145 ;
  assign n778 = n195 | n266 ;
  assign n779 = ( ~n776 & n777 ) | ( ~n776 & n778 ) | ( n777 & n778 ) ;
  assign n780 = n776 | n779 ;
  assign n781 = n196 | n586 ;
  assign n782 = ( n41 & n80 ) | ( n41 & n136 ) | ( n80 & n136 ) ;
  assign n783 = n66 & n145 ;
  assign n784 = ( ~n781 & n782 ) | ( ~n781 & n783 ) | ( n782 & n783 ) ;
  assign n785 = n781 | n784 ;
  assign n786 = n73 & n83 ;
  assign n787 = ( n202 & ~n485 ) | ( n202 & n786 ) | ( ~n485 & n786 ) ;
  assign n788 = n485 | n787 ;
  assign n789 = n207 | n685 ;
  assign n790 = n723 | n789 ;
  assign n791 = n479 | n641 ;
  assign n792 = ( n80 & n100 ) | ( n80 & n395 ) | ( n100 & n395 ) ;
  assign n793 = ( ~n790 & n791 ) | ( ~n790 & n792 ) | ( n791 & n792 ) ;
  assign n794 = n790 | n793 ;
  assign n795 = n44 & n129 ;
  assign n796 = n80 & n216 ;
  assign n797 = n402 | n796 ;
  assign n798 = n795 | n797 ;
  assign n799 = ( ~n788 & n794 ) | ( ~n788 & n798 ) | ( n794 & n798 ) ;
  assign n800 = n788 | n799 ;
  assign n801 = ( ~n780 & n785 ) | ( ~n780 & n800 ) | ( n785 & n800 ) ;
  assign n802 = n780 | n801 ;
  assign n803 = ( ~n751 & n774 ) | ( ~n751 & n802 ) | ( n774 & n802 ) ;
  assign n804 = ( ~n752 & n772 ) | ( ~n752 & n803 ) | ( n772 & n803 ) ;
  assign n805 = n752 | n804 ;
  assign n806 = n102 & n149 ;
  assign n807 = n117 | n806 ;
  assign n808 = n360 | n807 ;
  assign n809 = n203 | n227 ;
  assign n810 = n44 & n50 ;
  assign n811 = n168 | n810 ;
  assign n812 = n317 | n811 ;
  assign n813 = n809 | n812 ;
  assign n814 = n188 | n231 ;
  assign n815 = n76 | n153 ;
  assign n816 = ( ~n135 & n144 ) | ( ~n135 & n211 ) | ( n144 & n211 ) ;
  assign n817 = n135 | n816 ;
  assign n818 = ( ~n814 & n815 ) | ( ~n814 & n817 ) | ( n815 & n817 ) ;
  assign n819 = n814 | n818 ;
  assign n820 = ( ~n808 & n813 ) | ( ~n808 & n819 ) | ( n813 & n819 ) ;
  assign n821 = n808 | n820 ;
  assign n822 = ( n75 & n109 ) | ( n75 & n680 ) | ( n109 & n680 ) ;
  assign n823 = ( n48 & n84 ) | ( n48 & n115 ) | ( n84 & n115 ) ;
  assign n824 = n50 & n97 ;
  assign n825 = ( n331 & ~n823 ) | ( n331 & n824 ) | ( ~n823 & n824 ) ;
  assign n826 = n823 | n825 ;
  assign n827 = n361 | n455 ;
  assign n828 = n150 | n827 ;
  assign n829 = ( n102 & n136 ) | ( n102 & n166 ) | ( n136 & n166 ) ;
  assign n830 = n286 | n595 ;
  assign n831 = n265 | n830 ;
  assign n832 = ( n262 & ~n829 ) | ( n262 & n831 ) | ( ~n829 & n831 ) ;
  assign n833 = ( ~n828 & n829 ) | ( ~n828 & n832 ) | ( n829 & n832 ) ;
  assign n834 = ( ~n826 & n828 ) | ( ~n826 & n833 ) | ( n828 & n833 ) ;
  assign n835 = n826 | n834 ;
  assign n836 = n55 | n592 ;
  assign n837 = n142 | n689 ;
  assign n838 = n75 & n160 ;
  assign n839 = n152 & n216 ;
  assign n840 = n277 | n839 ;
  assign n841 = n838 | n840 ;
  assign n842 = ( ~n836 & n837 ) | ( ~n836 & n841 ) | ( n837 & n841 ) ;
  assign n843 = ( ~n835 & n836 ) | ( ~n835 & n842 ) | ( n836 & n842 ) ;
  assign n844 = n835 | n843 ;
  assign n845 = ( ~n821 & n822 ) | ( ~n821 & n844 ) | ( n822 & n844 ) ;
  assign n846 = n821 | n845 ;
  assign n847 = n177 | n505 ;
  assign n848 = n189 | n536 ;
  assign n849 = n847 | n848 ;
  assign n850 = n661 | n713 ;
  assign n851 = n83 & n145 ;
  assign n852 = n241 | n851 ;
  assign n853 = ( n238 & n272 ) | ( n238 & ~n852 ) | ( n272 & ~n852 ) ;
  assign n854 = n852 | n853 ;
  assign n855 = n348 | n642 ;
  assign n856 = n41 & n160 ;
  assign n857 = n356 | n856 ;
  assign n858 = ( ~n854 & n855 ) | ( ~n854 & n857 ) | ( n855 & n857 ) ;
  assign n859 = n854 | n858 ;
  assign n860 = ( ~n849 & n850 ) | ( ~n849 & n859 ) | ( n850 & n859 ) ;
  assign n861 = n849 | n860 ;
  assign n862 = n576 | n609 ;
  assign n863 = n299 | n862 ;
  assign n864 = n240 | n549 ;
  assign n865 = n48 & n83 ;
  assign n866 = n101 | n206 ;
  assign n867 = n133 | n866 ;
  assign n868 = ( ~n864 & n865 ) | ( ~n864 & n867 ) | ( n865 & n867 ) ;
  assign n869 = n864 | n868 ;
  assign n870 = ( ~n861 & n863 ) | ( ~n861 & n869 ) | ( n863 & n869 ) ;
  assign n871 = n861 | n870 ;
  assign n872 = ( ~n805 & n846 ) | ( ~n805 & n871 ) | ( n846 & n871 ) ;
  assign n873 = n84 & n216 ;
  assign n874 = n103 | n873 ;
  assign n875 = n488 | n874 ;
  assign n876 = n66 & n122 ;
  assign n877 = n164 | n367 ;
  assign n878 = n73 & n166 ;
  assign n879 = ( n590 & ~n877 ) | ( n590 & n878 ) | ( ~n877 & n878 ) ;
  assign n880 = n877 | n879 ;
  assign n881 = ( ~n875 & n876 ) | ( ~n875 & n880 ) | ( n876 & n880 ) ;
  assign n882 = n875 | n881 ;
  assign n883 = n384 | n434 ;
  assign n884 = n273 | n537 ;
  assign n885 = n48 & n98 ;
  assign n886 = n166 & n216 ;
  assign n887 = n885 | n886 ;
  assign n888 = n97 & n129 ;
  assign n889 = n599 | n888 ;
  assign n890 = n98 & n160 ;
  assign n891 = n298 | n890 ;
  assign n892 = ( ~n887 & n889 ) | ( ~n887 & n891 ) | ( n889 & n891 ) ;
  assign n893 = ( ~n884 & n887 ) | ( ~n884 & n892 ) | ( n887 & n892 ) ;
  assign n894 = n884 | n893 ;
  assign n895 = n48 & n57 ;
  assign n896 = n285 | n416 ;
  assign n897 = n895 | n896 ;
  assign n898 = ( ~n883 & n894 ) | ( ~n883 & n897 ) | ( n894 & n897 ) ;
  assign n899 = n883 | n898 ;
  assign n900 = ( ~n871 & n882 ) | ( ~n871 & n899 ) | ( n882 & n899 ) ;
  assign n901 = ( ~n805 & n872 ) | ( ~n805 & n900 ) | ( n872 & n900 ) ;
  assign n902 = n805 | n901 ;
  assign n903 = n104 | n696 ;
  assign n904 = ( n48 & n75 ) | ( n48 & n102 ) | ( n75 & n102 ) ;
  assign n905 = n316 | n440 ;
  assign n906 = ( n662 & ~n904 ) | ( n662 & n905 ) | ( ~n904 & n905 ) ;
  assign n907 = ( n505 & n904 ) | ( n505 & ~n906 ) | ( n904 & ~n906 ) ;
  assign n908 = n906 | n907 ;
  assign n909 = ( n791 & ~n903 ) | ( n791 & n908 ) | ( ~n903 & n908 ) ;
  assign n910 = n903 | n909 ;
  assign n911 = n562 | n786 ;
  assign n912 = ~n54 & n57 ;
  assign n913 = n734 | n912 ;
  assign n914 = n690 | n913 ;
  assign n915 = n911 | n914 ;
  assign n916 = n331 | n356 ;
  assign n917 = n64 & n149 ;
  assign n918 = n164 | n917 ;
  assign n919 = ( n48 & n72 ) | ( n48 & n84 ) | ( n72 & n84 ) ;
  assign n920 = n258 | n697 ;
  assign n921 = n98 & n216 ;
  assign n922 = n48 & n66 ;
  assign n923 = n921 | n922 ;
  assign n924 = ( ~n544 & n920 ) | ( ~n544 & n923 ) | ( n920 & n923 ) ;
  assign n925 = n919 | n924 ;
  assign n926 = ( ~n915 & n918 ) | ( ~n915 & n925 ) | ( n918 & n925 ) ;
  assign n927 = n916 | n926 ;
  assign n928 = n75 & n149 ;
  assign n929 = ( n119 & n136 ) | ( n119 & n152 ) | ( n136 & n152 ) ;
  assign n930 = n928 | n929 ;
  assign n931 = n176 | n492 ;
  assign n932 = n489 | n851 ;
  assign n933 = n41 & n136 ;
  assign n934 = ( n239 & ~n932 ) | ( n239 & n933 ) | ( ~n932 & n933 ) ;
  assign n935 = n932 | n934 ;
  assign n936 = ( ~n930 & n931 ) | ( ~n930 & n935 ) | ( n931 & n935 ) ;
  assign n937 = ( ~n927 & n930 ) | ( ~n927 & n936 ) | ( n930 & n936 ) ;
  assign n938 = n927 | n937 ;
  assign n939 = ( ~n910 & n915 ) | ( ~n910 & n938 ) | ( n915 & n938 ) ;
  assign n940 = n910 | n939 ;
  assign n941 = n97 & n166 ;
  assign n942 = n137 | n941 ;
  assign n943 = n55 | n211 ;
  assign n944 = n942 | n943 ;
  assign n945 = ( n44 & n57 ) | ( n44 & n80 ) | ( n57 & n80 ) ;
  assign n946 = n196 | n402 ;
  assign n947 = n41 & n122 ;
  assign n948 = ( n764 & ~n946 ) | ( n764 & n947 ) | ( ~n946 & n947 ) ;
  assign n949 = n946 | n948 ;
  assign n950 = ( ~n944 & n945 ) | ( ~n944 & n949 ) | ( n945 & n949 ) ;
  assign n951 = n944 | n950 ;
  assign n952 = n64 & n160 ;
  assign n953 = n81 | n952 ;
  assign n954 = ( n609 & n890 ) | ( n609 & ~n953 ) | ( n890 & ~n953 ) ;
  assign n955 = n953 | n954 ;
  assign n956 = n80 & n136 ;
  assign n957 = n865 | n956 ;
  assign n958 = n639 | n957 ;
  assign n959 = n240 | n328 ;
  assign n960 = ~n54 & n152 ;
  assign n961 = n205 | n960 ;
  assign n962 = n959 | n961 ;
  assign n963 = n285 | n653 ;
  assign n964 = ( n773 & ~n962 ) | ( n773 & n963 ) | ( ~n962 & n963 ) ;
  assign n965 = n962 | n964 ;
  assign n966 = ( ~n955 & n958 ) | ( ~n955 & n965 ) | ( n958 & n965 ) ;
  assign n967 = ( n951 & n955 ) | ( n951 & ~n966 ) | ( n955 & ~n966 ) ;
  assign n968 = n123 | n185 ;
  assign n969 = n261 | n968 ;
  assign n970 = ( n642 & n876 ) | ( n642 & ~n969 ) | ( n876 & ~n969 ) ;
  assign n971 = n969 | n970 ;
  assign n972 = n174 | n488 ;
  assign n973 = n101 | n972 ;
  assign n974 = n809 | n973 ;
  assign n975 = n346 | n465 ;
  assign n976 = n895 | n975 ;
  assign n977 = n41 & n59 ;
  assign n978 = n188 | n523 ;
  assign n979 = ( n302 & ~n977 ) | ( n302 & n978 ) | ( ~n977 & n978 ) ;
  assign n980 = n977 | n979 ;
  assign n981 = n234 | n839 ;
  assign n982 = ( n376 & ~n980 ) | ( n376 & n981 ) | ( ~n980 & n981 ) ;
  assign n983 = n980 | n982 ;
  assign n984 = n207 | n565 ;
  assign n985 = n66 & n73 ;
  assign n986 = ( n212 & ~n984 ) | ( n212 & n985 ) | ( ~n984 & n985 ) ;
  assign n987 = n984 | n986 ;
  assign n988 = ( ~n976 & n983 ) | ( ~n976 & n987 ) | ( n983 & n987 ) ;
  assign n989 = n976 | n988 ;
  assign n990 = ~n54 & n66 ;
  assign n991 = n613 | n990 ;
  assign n992 = n83 & n122 ;
  assign n993 = n455 | n992 ;
  assign n994 = n991 | n993 ;
  assign n995 = n75 & n145 ;
  assign n996 = n111 | n995 ;
  assign n997 = ( n692 & ~n994 ) | ( n692 & n996 ) | ( ~n994 & n996 ) ;
  assign n998 = n994 | n997 ;
  assign n999 = ( ~n974 & n989 ) | ( ~n974 & n998 ) | ( n989 & n998 ) ;
  assign n1000 = ( ~n971 & n974 ) | ( ~n971 & n999 ) | ( n974 & n999 ) ;
  assign n1001 = n41 & n97 ;
  assign n1002 = n500 | n1001 ;
  assign n1003 = n536 | n1002 ;
  assign n1004 = n971 | n1003 ;
  assign n1005 = n79 | n202 ;
  assign n1006 = n777 | n810 ;
  assign n1007 = n1005 | n1006 ;
  assign n1008 = ( n64 & n97 ) | ( n64 & n129 ) | ( n97 & n129 ) ;
  assign n1009 = n360 | n760 ;
  assign n1010 = ( ~n1007 & n1008 ) | ( ~n1007 & n1009 ) | ( n1008 & n1009 ) ;
  assign n1011 = n1007 | n1010 ;
  assign n1012 = n540 | n762 ;
  assign n1013 = ( n50 & n160 ) | ( n50 & n483 ) | ( n160 & n483 ) ;
  assign n1014 = n1012 | n1013 ;
  assign n1015 = ( ~n1003 & n1011 ) | ( ~n1003 & n1014 ) | ( n1011 & n1014 ) ;
  assign n1016 = ( ~n1000 & n1004 ) | ( ~n1000 & n1015 ) | ( n1004 & n1015 ) ;
  assign n1017 = n1000 | n1016 ;
  assign n1018 = ( n966 & ~n967 ) | ( n966 & n1017 ) | ( ~n967 & n1017 ) ;
  assign n1019 = n967 | n1018 ;
  assign n1020 = n60 | n231 ;
  assign n1021 = ( n84 & n115 ) | ( n84 & n160 ) | ( n115 & n160 ) ;
  assign n1022 = n1020 | n1021 ;
  assign n1023 = n242 | n528 ;
  assign n1024 = n238 | n265 ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = ( n59 & n75 ) | ( n59 & n160 ) | ( n75 & n160 ) ;
  assign n1027 = n73 & n75 ;
  assign n1028 = ( n493 & ~n1026 ) | ( n493 & n1027 ) | ( ~n1026 & n1027 ) ;
  assign n1029 = n1026 | n1028 ;
  assign n1030 = ( n1022 & ~n1025 ) | ( n1022 & n1029 ) | ( ~n1025 & n1029 ) ;
  assign n1031 = n129 & n160 ;
  assign n1032 = n189 | n1031 ;
  assign n1033 = n224 | n1032 ;
  assign n1034 = ( n298 & n795 ) | ( n298 & ~n1033 ) | ( n795 & ~n1033 ) ;
  assign n1035 = n1033 | n1034 ;
  assign n1036 = ( n1025 & ~n1030 ) | ( n1025 & n1035 ) | ( ~n1030 & n1035 ) ;
  assign n1037 = n1030 | n1036 ;
  assign n1038 = ( ~n940 & n1019 ) | ( ~n940 & n1037 ) | ( n1019 & n1037 ) ;
  assign n1039 = n940 | n1038 ;
  assign n1040 = ( ~x26 & n902 ) | ( ~x26 & n1039 ) | ( n902 & n1039 ) ;
  assign n1041 = ( n57 & n216 ) | ( n57 & n912 ) | ( n216 & n912 ) ;
  assign n1042 = ( n500 & n696 ) | ( n500 & ~n1041 ) | ( n696 & ~n1041 ) ;
  assign n1043 = n1041 | n1042 ;
  assign n1044 = n44 & n152 ;
  assign n1045 = n338 | n1044 ;
  assign n1046 = ( n196 & n234 ) | ( n196 & ~n1045 ) | ( n234 & ~n1045 ) ;
  assign n1047 = n1045 | n1046 ;
  assign n1048 = n57 & n109 ;
  assign n1049 = n218 & ~n1048 ;
  assign n1050 = n146 | n865 ;
  assign n1051 = n1049 & ~n1050 ;
  assign n1052 = ( n1043 & ~n1047 ) | ( n1043 & n1051 ) | ( ~n1047 & n1051 ) ;
  assign n1053 = ~n1043 & n1052 ;
  assign n1054 = n775 | n922 ;
  assign n1055 = n298 | n1054 ;
  assign n1056 = ( n85 & n86 ) | ( n85 & n145 ) | ( n86 & n145 ) ;
  assign n1057 = ( ~n78 & n149 ) | ( ~n78 & n216 ) | ( n149 & n216 ) ;
  assign n1058 = n1056 | n1057 ;
  assign n1059 = n97 & n98 ;
  assign n1060 = n290 | n1059 ;
  assign n1061 = n115 | n217 ;
  assign n1062 = n77 | n138 ;
  assign n1063 = ( n665 & ~n1061 ) | ( n665 & n1062 ) | ( ~n1061 & n1062 ) ;
  assign n1064 = n1061 | n1063 ;
  assign n1065 = ( ~n1058 & n1060 ) | ( ~n1058 & n1064 ) | ( n1060 & n1064 ) ;
  assign n1066 = n1058 | n1065 ;
  assign n1067 = n202 | n592 ;
  assign n1068 = n98 & n149 ;
  assign n1069 = ( n856 & ~n1067 ) | ( n856 & n1068 ) | ( ~n1067 & n1068 ) ;
  assign n1070 = n1067 | n1069 ;
  assign n1071 = ( ~n1055 & n1066 ) | ( ~n1055 & n1070 ) | ( n1066 & n1070 ) ;
  assign n1072 = n111 | n1031 ;
  assign n1073 = ( n301 & n488 ) | ( n301 & ~n1072 ) | ( n488 & ~n1072 ) ;
  assign n1074 = n1072 | n1073 ;
  assign n1075 = ( n1055 & ~n1071 ) | ( n1055 & n1074 ) | ( ~n1071 & n1074 ) ;
  assign n1076 = n1071 | n1075 ;
  assign n1077 = n92 | n300 ;
  assign n1078 = n277 | n295 ;
  assign n1079 = n241 | n697 ;
  assign n1080 = n1078 | n1079 ;
  assign n1081 = n1077 | n1080 ;
  assign n1082 = n75 & n109 ;
  assign n1083 = n193 | n1082 ;
  assign n1084 = n79 | n273 ;
  assign n1085 = ( n72 & ~n78 ) | ( n72 & n136 ) | ( ~n78 & n136 ) ;
  assign n1086 = ( n75 & n100 ) | ( n75 & n149 ) | ( n100 & n149 ) ;
  assign n1087 = n455 | n1086 ;
  assign n1088 = ( ~n1084 & n1085 ) | ( ~n1084 & n1087 ) | ( n1085 & n1087 ) ;
  assign n1089 = n1084 | n1088 ;
  assign n1090 = ( ~n1081 & n1083 ) | ( ~n1081 & n1089 ) | ( n1083 & n1089 ) ;
  assign n1091 = n1081 | n1090 ;
  assign n1092 = ( n64 & n102 ) | ( n64 & n160 ) | ( n102 & n160 ) ;
  assign n1093 = n197 | n1092 ;
  assign n1094 = n476 | n1093 ;
  assign n1095 = n396 | n1006 ;
  assign n1096 = n44 & n166 ;
  assign n1097 = n312 | n1096 ;
  assign n1098 = n242 | n895 ;
  assign n1099 = ( n50 & n75 ) | ( n50 & n145 ) | ( n75 & n145 ) ;
  assign n1100 = n806 | n1099 ;
  assign n1101 = ( ~n1097 & n1098 ) | ( ~n1097 & n1100 ) | ( n1098 & n1100 ) ;
  assign n1102 = n1097 | n1101 ;
  assign n1103 = n393 | n782 ;
  assign n1104 = ( ~n1095 & n1102 ) | ( ~n1095 & n1103 ) | ( n1102 & n1103 ) ;
  assign n1105 = n1095 | n1104 ;
  assign n1106 = ( n817 & ~n1094 ) | ( n817 & n1105 ) | ( ~n1094 & n1105 ) ;
  assign n1107 = n1094 | n1106 ;
  assign n1108 = ( n1076 & ~n1091 ) | ( n1076 & n1107 ) | ( ~n1091 & n1107 ) ;
  assign n1109 = n1053 & ~n1108 ;
  assign n1110 = n80 & n97 ;
  assign n1111 = ( n123 & ~n837 ) | ( n123 & n1110 ) | ( ~n837 & n1110 ) ;
  assign n1112 = n837 | n1111 ;
  assign n1113 = ( n73 & n102 ) | ( n73 & n129 ) | ( n102 & n129 ) ;
  assign n1114 = ( n702 & ~n1112 ) | ( n702 & n1113 ) | ( ~n1112 & n1113 ) ;
  assign n1115 = n1112 | n1114 ;
  assign n1116 = ~n54 & n98 ;
  assign n1117 = n567 | n1116 ;
  assign n1118 = n117 | n317 ;
  assign n1119 = ( n721 & ~n1117 ) | ( n721 & n1118 ) | ( ~n1117 & n1118 ) ;
  assign n1120 = n1117 | n1119 ;
  assign n1121 = n224 | n732 ;
  assign n1122 = ( n64 & n98 ) | ( n64 & n216 ) | ( n98 & n216 ) ;
  assign n1123 = n323 | n1122 ;
  assign n1124 = ( n514 & ~n1121 ) | ( n514 & n1123 ) | ( ~n1121 & n1123 ) ;
  assign n1125 = n1121 | n1124 ;
  assign n1126 = n1120 | n1125 ;
  assign n1127 = n1115 | n1126 ;
  assign n1128 = n231 | n582 ;
  assign n1129 = n447 | n479 ;
  assign n1130 = n1128 | n1129 ;
  assign n1131 = n838 | n878 ;
  assign n1132 = n562 | n591 ;
  assign n1133 = n101 | n675 ;
  assign n1134 = n105 | n1133 ;
  assign n1135 = n1132 | n1134 ;
  assign n1136 = n168 | n662 ;
  assign n1137 = n653 | n931 ;
  assign n1138 = ( ~n1135 & n1136 ) | ( ~n1135 & n1137 ) | ( n1136 & n1137 ) ;
  assign n1139 = n1135 | n1138 ;
  assign n1140 = ( ~n1130 & n1131 ) | ( ~n1130 & n1139 ) | ( n1131 & n1139 ) ;
  assign n1141 = n1130 | n1140 ;
  assign n1142 = ( n258 & n839 ) | ( n258 & ~n977 ) | ( n839 & ~n977 ) ;
  assign n1143 = n977 | n1142 ;
  assign n1144 = n81 | n691 ;
  assign n1145 = n267 | n435 ;
  assign n1146 = n1144 | n1145 ;
  assign n1147 = ( ~n261 & n361 ) | ( ~n261 & n886 ) | ( n361 & n886 ) ;
  assign n1148 = n261 | n1147 ;
  assign n1149 = ( n72 & n102 ) | ( n72 & n109 ) | ( n102 & n109 ) ;
  assign n1150 = n153 | n1149 ;
  assign n1151 = ( ~n1143 & n1148 ) | ( ~n1143 & n1150 ) | ( n1148 & n1150 ) ;
  assign n1152 = ( ~n1143 & n1146 ) | ( ~n1143 & n1151 ) | ( n1146 & n1151 ) ;
  assign n1153 = n1143 | n1152 ;
  assign n1154 = ( ~n1127 & n1141 ) | ( ~n1127 & n1153 ) | ( n1141 & n1153 ) ;
  assign n1155 = n1127 | n1154 ;
  assign n1156 = ( n1091 & n1109 ) | ( n1091 & n1155 ) | ( n1109 & n1155 ) ;
  assign n1157 = n1109 & ~n1156 ;
  assign n1158 = ( n109 & n129 ) | ( n109 & n166 ) | ( n129 & n166 ) ;
  assign n1159 = ( n80 & n98 ) | ( n80 & n109 ) | ( n98 & n109 ) ;
  assign n1160 = n205 | n1159 ;
  assign n1161 = ( n479 & ~n1158 ) | ( n479 & n1160 ) | ( ~n1158 & n1160 ) ;
  assign n1162 = n1158 | n1161 ;
  assign n1163 = n164 | n562 ;
  assign n1164 = ( n102 & n109 ) | ( n102 & n152 ) | ( n109 & n152 ) ;
  assign n1165 = ( n110 & n543 ) | ( n110 & ~n1164 ) | ( n543 & ~n1164 ) ;
  assign n1166 = n1164 | n1165 ;
  assign n1167 = ( ~n1162 & n1163 ) | ( ~n1162 & n1166 ) | ( n1163 & n1166 ) ;
  assign n1168 = n1162 | n1167 ;
  assign n1169 = n72 & n216 ;
  assign n1170 = n177 | n1169 ;
  assign n1171 = n64 & n216 ;
  assign n1172 = n582 | n1171 ;
  assign n1173 = n255 | n581 ;
  assign n1174 = n529 | n576 ;
  assign n1175 = ( ~n1172 & n1173 ) | ( ~n1172 & n1174 ) | ( n1173 & n1174 ) ;
  assign n1176 = ( ~n271 & n1172 ) | ( ~n271 & n1175 ) | ( n1172 & n1175 ) ;
  assign n1177 = n271 | n1176 ;
  assign n1178 = n482 | n599 ;
  assign n1179 = ( n75 & ~n78 ) | ( n75 & n97 ) | ( ~n78 & n97 ) ;
  assign n1180 = ( n291 & ~n1096 ) | ( n291 & n1179 ) | ( ~n1096 & n1179 ) ;
  assign n1181 = n1096 | n1180 ;
  assign n1182 = ( n287 & ~n1178 ) | ( n287 & n1181 ) | ( ~n1178 & n1181 ) ;
  assign n1183 = n1178 | n1182 ;
  assign n1184 = ( n1170 & ~n1177 ) | ( n1170 & n1183 ) | ( ~n1177 & n1183 ) ;
  assign n1185 = n493 | n839 ;
  assign n1186 = n288 | n1185 ;
  assign n1187 = ( n1177 & ~n1184 ) | ( n1177 & n1186 ) | ( ~n1184 & n1186 ) ;
  assign n1188 = n1184 | n1187 ;
  assign n1189 = ( n72 & n84 ) | ( n72 & n116 ) | ( n84 & n116 ) ;
  assign n1190 = ( n64 & n102 ) | ( n64 & n116 ) | ( n102 & n116 ) ;
  assign n1191 = n691 | n1190 ;
  assign n1192 = ( n628 & ~n1189 ) | ( n628 & n1191 ) | ( ~n1189 & n1191 ) ;
  assign n1193 = n1189 | n1192 ;
  assign n1194 = ( n665 & n675 ) | ( n665 & ~n1193 ) | ( n675 & ~n1193 ) ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = ( n84 & n129 ) | ( n84 & n216 ) | ( n129 & n216 ) ;
  assign n1197 = n130 | n1196 ;
  assign n1198 = n1195 | n1197 ;
  assign n1199 = n921 | n1044 ;
  assign n1200 = n598 | n1199 ;
  assign n1201 = ( n41 & n132 ) | ( n41 & n145 ) | ( n132 & n145 ) ;
  assign n1202 = ( n44 & n64 ) | ( n44 & n98 ) | ( n64 & n98 ) ;
  assign n1203 = ( n234 & ~n1201 ) | ( n234 & n1202 ) | ( ~n1201 & n1202 ) ;
  assign n1204 = n1201 | n1203 ;
  assign n1205 = ( n83 & n102 ) | ( n83 & n216 ) | ( n102 & n216 ) ;
  assign n1206 = ( n44 & n48 ) | ( n44 & n72 ) | ( n48 & n72 ) ;
  assign n1207 = n1205 | n1206 ;
  assign n1208 = n227 | n886 ;
  assign n1209 = n1207 | n1208 ;
  assign n1210 = ( ~n1200 & n1204 ) | ( ~n1200 & n1209 ) | ( n1204 & n1209 ) ;
  assign n1211 = n1200 | n1210 ;
  assign n1212 = ( n66 & n75 ) | ( n66 & n136 ) | ( n75 & n136 ) ;
  assign n1213 = n504 | n679 ;
  assign n1214 = ( n642 & ~n1212 ) | ( n642 & n1213 ) | ( ~n1212 & n1213 ) ;
  assign n1215 = n1212 | n1214 ;
  assign n1216 = ( ~n1195 & n1211 ) | ( ~n1195 & n1215 ) | ( n1211 & n1215 ) ;
  assign n1217 = ( ~n1188 & n1198 ) | ( ~n1188 & n1216 ) | ( n1198 & n1216 ) ;
  assign n1218 = n1188 | n1217 ;
  assign n1219 = n1168 | n1218 ;
  assign n1220 = n507 | n796 ;
  assign n1221 = n423 | n1220 ;
  assign n1222 = ( ~n54 & n72 ) | ( ~n54 & n129 ) | ( n72 & n129 ) ;
  assign n1223 = n613 | n1222 ;
  assign n1224 = ( n580 & n1221 ) | ( n580 & ~n1223 ) | ( n1221 & ~n1223 ) ;
  assign n1225 = n84 & n97 ;
  assign n1226 = n824 | n1008 ;
  assign n1227 = n1225 | n1226 ;
  assign n1228 = ( n1223 & ~n1224 ) | ( n1223 & n1227 ) | ( ~n1224 & n1227 ) ;
  assign n1229 = n1224 | n1228 ;
  assign n1230 = n218 & ~n380 ;
  assign n1231 = ( ~n54 & n57 ) | ( ~n54 & n102 ) | ( n57 & n102 ) ;
  assign n1232 = n1230 & ~n1231 ;
  assign n1233 = ~n1002 & n1232 ;
  assign n1234 = n172 | n450 ;
  assign n1235 = n567 | n759 ;
  assign n1236 = n630 | n1235 ;
  assign n1237 = n66 & n97 ;
  assign n1238 = ( n197 & ~n444 ) | ( n197 & n550 ) | ( ~n444 & n550 ) ;
  assign n1239 = ( n444 & ~n1237 ) | ( n444 & n1238 ) | ( ~n1237 & n1238 ) ;
  assign n1240 = n1237 | n1239 ;
  assign n1241 = ( ~n1234 & n1236 ) | ( ~n1234 & n1240 ) | ( n1236 & n1240 ) ;
  assign n1242 = n1234 | n1241 ;
  assign n1243 = ( n376 & n1233 ) | ( n376 & n1242 ) | ( n1233 & n1242 ) ;
  assign n1244 = n1233 & ~n1243 ;
  assign n1245 = ( n1219 & ~n1229 ) | ( n1219 & n1244 ) | ( ~n1229 & n1244 ) ;
  assign n1246 = ~n1219 & n1245 ;
  assign n1247 = ( x29 & x31 ) | ( x29 & ~n96 ) | ( x31 & ~n96 ) ;
  assign n1248 = ( x31 & n58 ) | ( x31 & n96 ) | ( n58 & n96 ) ;
  assign n1249 = ( ~x31 & n47 ) | ( ~x31 & n1248 ) | ( n47 & n1248 ) ;
  assign n1250 = ( ~x29 & n1247 ) | ( ~x29 & n1249 ) | ( n1247 & n1249 ) ;
  assign n1251 = ~n1246 & n1250 ;
  assign n1252 = n208 | n376 ;
  assign n1253 = n312 | n719 ;
  assign n1254 = ( n66 & n83 ) | ( n66 & n160 ) | ( n83 & n160 ) ;
  assign n1255 = n340 | n1254 ;
  assign n1256 = ( n41 & n75 ) | ( n41 & n160 ) | ( n75 & n160 ) ;
  assign n1257 = n124 | n1256 ;
  assign n1258 = n290 | n941 ;
  assign n1259 = ( n285 & ~n956 ) | ( n285 & n1258 ) | ( ~n956 & n1258 ) ;
  assign n1260 = n956 | n1259 ;
  assign n1261 = ( ~n1255 & n1257 ) | ( ~n1255 & n1260 ) | ( n1257 & n1260 ) ;
  assign n1262 = n1255 | n1261 ;
  assign n1263 = ( ~n1252 & n1253 ) | ( ~n1252 & n1262 ) | ( n1253 & n1262 ) ;
  assign n1264 = n1252 | n1263 ;
  assign n1265 = n439 | n575 ;
  assign n1266 = ( n281 & ~n1264 ) | ( n281 & n1265 ) | ( ~n1264 & n1265 ) ;
  assign n1267 = n1264 | n1266 ;
  assign n1268 = n607 & n1267 ;
  assign n1269 = n1251 | n1268 ;
  assign n1270 = n45 | n138 ;
  assign n1271 = n412 | n454 ;
  assign n1272 = ( n472 & n1270 ) | ( n472 & ~n1271 ) | ( n1270 & ~n1271 ) ;
  assign n1273 = n51 | n90 ;
  assign n1274 = n55 | n1273 ;
  assign n1275 = x28 & n96 ;
  assign n1276 = ( n41 & n75 ) | ( n41 & n1275 ) | ( n75 & n1275 ) ;
  assign n1277 = n227 | n1048 ;
  assign n1278 = n732 | n1277 ;
  assign n1279 = n1276 | n1278 ;
  assign n1280 = n941 | n1082 ;
  assign n1281 = ( n66 & n83 ) | ( n66 & n1275 ) | ( n83 & n1275 ) ;
  assign n1282 = n1280 | n1281 ;
  assign n1283 = ( n1227 & ~n1279 ) | ( n1227 & n1282 ) | ( ~n1279 & n1282 ) ;
  assign n1284 = ( ~n1195 & n1279 ) | ( ~n1195 & n1283 ) | ( n1279 & n1283 ) ;
  assign n1285 = ( n1168 & n1195 ) | ( n1168 & ~n1284 ) | ( n1195 & ~n1284 ) ;
  assign n1286 = n1284 | n1285 ;
  assign n1287 = ( n375 & n1274 ) | ( n375 & ~n1286 ) | ( n1274 & ~n1286 ) ;
  assign n1288 = ~n1274 & n1287 ;
  assign n1289 = ( ~n1271 & n1272 ) | ( ~n1271 & n1288 ) | ( n1272 & n1288 ) ;
  assign n1290 = ~n1272 & n1289 ;
  assign n1291 = n606 & n1290 ;
  assign n1292 = ( n606 & n1269 ) | ( n606 & ~n1291 ) | ( n1269 & ~n1291 ) ;
  assign n1293 = n576 | n786 ;
  assign n1294 = ( n540 & n952 ) | ( n540 & ~n1293 ) | ( n952 & ~n1293 ) ;
  assign n1295 = n1293 | n1294 ;
  assign n1296 = ( n348 & n353 ) | ( n348 & ~n990 ) | ( n353 & ~n990 ) ;
  assign n1297 = n990 | n1296 ;
  assign n1298 = ( n66 & n83 ) | ( n66 & n116 ) | ( n83 & n116 ) ;
  assign n1299 = ( n73 & n84 ) | ( n73 & n116 ) | ( n84 & n116 ) ;
  assign n1300 = n505 | n1299 ;
  assign n1301 = ( n887 & ~n1298 ) | ( n887 & n1300 ) | ( ~n1298 & n1300 ) ;
  assign n1302 = n1298 | n1301 ;
  assign n1303 = ( ~n1295 & n1297 ) | ( ~n1295 & n1302 ) | ( n1297 & n1302 ) ;
  assign n1304 = n1295 | n1303 ;
  assign n1305 = n252 & ~n1304 ;
  assign n1306 = n1031 | n1169 ;
  assign n1307 = n440 | n1306 ;
  assign n1308 = n587 | n839 ;
  assign n1309 = n517 | n1308 ;
  assign n1310 = ( n421 & ~n1307 ) | ( n421 & n1309 ) | ( ~n1307 & n1309 ) ;
  assign n1311 = n1307 | n1310 ;
  assign n1312 = n697 | n1116 ;
  assign n1313 = n73 & ~n78 ;
  assign n1314 = n567 | n1313 ;
  assign n1315 = n544 | n775 ;
  assign n1316 = ( ~n1312 & n1314 ) | ( ~n1312 & n1315 ) | ( n1314 & n1315 ) ;
  assign n1317 = n1312 | n1316 ;
  assign n1318 = ( n482 & ~n679 ) | ( n482 & n941 ) | ( ~n679 & n941 ) ;
  assign n1319 = n679 | n1318 ;
  assign n1320 = n595 | n985 ;
  assign n1321 = ( n376 & ~n1319 ) | ( n376 & n1320 ) | ( ~n1319 & n1320 ) ;
  assign n1322 = n1319 | n1321 ;
  assign n1323 = n435 | n666 ;
  assign n1324 = ( n75 & n98 ) | ( n75 & n216 ) | ( n98 & n216 ) ;
  assign n1325 = ( n66 & n75 ) | ( n66 & n145 ) | ( n75 & n145 ) ;
  assign n1326 = n960 | n1325 ;
  assign n1327 = ( ~n78 & n122 ) | ( ~n78 & n216 ) | ( n122 & n216 ) ;
  assign n1328 = ( ~n1324 & n1326 ) | ( ~n1324 & n1327 ) | ( n1326 & n1327 ) ;
  assign n1329 = n1324 | n1328 ;
  assign n1330 = ( ~n54 & n73 ) | ( ~n54 & n75 ) | ( n73 & n75 ) ;
  assign n1331 = ( n551 & n638 ) | ( n551 & ~n1330 ) | ( n638 & ~n1330 ) ;
  assign n1332 = n1330 | n1331 ;
  assign n1333 = ( ~n1323 & n1329 ) | ( ~n1323 & n1332 ) | ( n1329 & n1332 ) ;
  assign n1334 = ( ~n1322 & n1323 ) | ( ~n1322 & n1333 ) | ( n1323 & n1333 ) ;
  assign n1335 = ( ~n1317 & n1322 ) | ( ~n1317 & n1334 ) | ( n1322 & n1334 ) ;
  assign n1336 = n1317 | n1335 ;
  assign n1337 = ( n1305 & n1311 ) | ( n1305 & n1336 ) | ( n1311 & n1336 ) ;
  assign n1338 = n1305 & ~n1337 ;
  assign n1339 = n206 | n512 ;
  assign n1340 = n586 | n1339 ;
  assign n1341 = n50 & n73 ;
  assign n1342 = ( n567 & ~n1068 ) | ( n567 & n1341 ) | ( ~n1068 & n1341 ) ;
  assign n1343 = n1068 | n1342 ;
  assign n1344 = ( n368 & ~n1340 ) | ( n368 & n1343 ) | ( ~n1340 & n1343 ) ;
  assign n1345 = ( n1173 & ~n1340 ) | ( n1173 & n1344 ) | ( ~n1340 & n1344 ) ;
  assign n1346 = ~n54 & n75 ;
  assign n1347 = n177 | n1346 ;
  assign n1348 = n228 | n440 ;
  assign n1349 = ( n1110 & ~n1347 ) | ( n1110 & n1348 ) | ( ~n1347 & n1348 ) ;
  assign n1350 = n1347 | n1349 ;
  assign n1351 = n142 | n839 ;
  assign n1352 = ( n75 & n136 ) | ( n75 & n149 ) | ( n136 & n149 ) ;
  assign n1353 = n261 | n1352 ;
  assign n1354 = ( n217 & n230 ) | ( n217 & ~n1353 ) | ( n230 & ~n1353 ) ;
  assign n1355 = n1353 | n1354 ;
  assign n1356 = ( n149 & n166 ) | ( n149 & n216 ) | ( n166 & n216 ) ;
  assign n1357 = ( n916 & ~n1355 ) | ( n916 & n1356 ) | ( ~n1355 & n1356 ) ;
  assign n1358 = n1355 | n1357 ;
  assign n1359 = ( ~n1350 & n1351 ) | ( ~n1350 & n1358 ) | ( n1351 & n1358 ) ;
  assign n1360 = n1350 | n1359 ;
  assign n1361 = ( n1340 & ~n1345 ) | ( n1340 & n1360 ) | ( ~n1345 & n1360 ) ;
  assign n1362 = n1345 | n1361 ;
  assign n1363 = n124 | n851 ;
  assign n1364 = n590 | n1363 ;
  assign n1365 = n59 & n98 ;
  assign n1366 = n72 & n109 ;
  assign n1367 = ( ~n1363 & n1365 ) | ( ~n1363 & n1366 ) | ( n1365 & n1366 ) ;
  assign n1368 = ( n662 & ~n1364 ) | ( n662 & n1367 ) | ( ~n1364 & n1367 ) ;
  assign n1369 = n1364 | n1368 ;
  assign n1370 = n329 | n959 ;
  assign n1371 = n952 | n960 ;
  assign n1372 = ( n195 & n545 ) | ( n195 & ~n1371 ) | ( n545 & ~n1371 ) ;
  assign n1373 = n1371 | n1372 ;
  assign n1374 = ( n838 & ~n1370 ) | ( n838 & n1373 ) | ( ~n1370 & n1373 ) ;
  assign n1375 = n1370 | n1374 ;
  assign n1376 = n84 & n160 ;
  assign n1377 = n167 | n1376 ;
  assign n1378 = n449 | n1377 ;
  assign n1379 = n203 | n1378 ;
  assign n1380 = n361 | n466 ;
  assign n1381 = ( n75 & n98 ) | ( n75 & n109 ) | ( n98 & n109 ) ;
  assign n1382 = ( ~n1379 & n1380 ) | ( ~n1379 & n1381 ) | ( n1380 & n1381 ) ;
  assign n1383 = n1379 | n1382 ;
  assign n1384 = ( n1369 & ~n1375 ) | ( n1369 & n1383 ) | ( ~n1375 & n1383 ) ;
  assign n1385 = ( n599 & n874 ) | ( n599 & ~n890 ) | ( n874 & ~n890 ) ;
  assign n1386 = n890 | n1385 ;
  assign n1387 = n1048 | n1096 ;
  assign n1388 = n74 | n582 ;
  assign n1389 = n259 | n1388 ;
  assign n1390 = n1387 | n1389 ;
  assign n1391 = ( n170 & n262 ) | ( n170 & ~n777 ) | ( n262 & ~n777 ) ;
  assign n1392 = n777 | n1391 ;
  assign n1393 = ( ~n1386 & n1390 ) | ( ~n1386 & n1392 ) | ( n1390 & n1392 ) ;
  assign n1394 = n1386 | n1393 ;
  assign n1395 = ( n1375 & ~n1384 ) | ( n1375 & n1394 ) | ( ~n1384 & n1394 ) ;
  assign n1396 = n1384 | n1395 ;
  assign n1397 = n485 | n696 ;
  assign n1398 = ( n352 & n613 ) | ( n352 & ~n1397 ) | ( n613 & ~n1397 ) ;
  assign n1399 = n1397 | n1398 ;
  assign n1400 = n258 | n775 ;
  assign n1401 = n435 | n878 ;
  assign n1402 = ( ~n1399 & n1400 ) | ( ~n1399 & n1401 ) | ( n1400 & n1401 ) ;
  assign n1403 = n1399 | n1402 ;
  assign n1404 = n422 | n732 ;
  assign n1405 = n592 | n691 ;
  assign n1406 = ( n1023 & ~n1404 ) | ( n1023 & n1405 ) | ( ~n1404 & n1405 ) ;
  assign n1407 = n1404 | n1406 ;
  assign n1408 = n360 | n523 ;
  assign n1409 = ( ~n54 & n145 ) | ( ~n54 & n166 ) | ( n145 & n166 ) ;
  assign n1410 = ( n239 & ~n995 ) | ( n239 & n1409 ) | ( ~n995 & n1409 ) ;
  assign n1411 = n995 | n1410 ;
  assign n1412 = ( n133 & ~n1408 ) | ( n133 & n1411 ) | ( ~n1408 & n1411 ) ;
  assign n1413 = n1408 | n1412 ;
  assign n1414 = ( ~n1403 & n1407 ) | ( ~n1403 & n1413 ) | ( n1407 & n1413 ) ;
  assign n1415 = n1403 | n1414 ;
  assign n1416 = n1396 | n1415 ;
  assign n1417 = ( n48 & n72 ) | ( n48 & n129 ) | ( n72 & n129 ) ;
  assign n1418 = n295 | n482 ;
  assign n1419 = ( n266 & ~n1417 ) | ( n266 & n1418 ) | ( ~n1417 & n1418 ) ;
  assign n1420 = n1417 | n1419 ;
  assign n1421 = ( n66 & n97 ) | ( n66 & n216 ) | ( n97 & n216 ) ;
  assign n1422 = n429 | n1421 ;
  assign n1423 = n433 | n796 ;
  assign n1424 = ( n294 & ~n1205 ) | ( n294 & n1423 ) | ( ~n1205 & n1423 ) ;
  assign n1425 = n1205 | n1424 ;
  assign n1426 = n550 | n655 ;
  assign n1427 = n941 | n1426 ;
  assign n1428 = ( ~n1422 & n1425 ) | ( ~n1422 & n1427 ) | ( n1425 & n1427 ) ;
  assign n1429 = n1422 | n1428 ;
  assign n1430 = n115 | n587 ;
  assign n1431 = ( n197 & ~n378 ) | ( n197 & n1430 ) | ( ~n378 & n1430 ) ;
  assign n1432 = n378 | n1431 ;
  assign n1433 = ( ~n1420 & n1429 ) | ( ~n1420 & n1432 ) | ( n1429 & n1432 ) ;
  assign n1434 = n1420 | n1433 ;
  assign n1435 = ( n98 & n119 ) | ( n98 & n166 ) | ( n119 & n166 ) ;
  assign n1436 = n185 | n885 ;
  assign n1437 = n1435 | n1436 ;
  assign n1438 = n224 | n337 ;
  assign n1439 = ( n265 & n320 ) | ( n265 & ~n1438 ) | ( n320 & ~n1438 ) ;
  assign n1440 = n1438 | n1439 ;
  assign n1441 = n713 | n746 ;
  assign n1442 = n534 | n1441 ;
  assign n1443 = ( ~n1437 & n1440 ) | ( ~n1437 & n1442 ) | ( n1440 & n1442 ) ;
  assign n1444 = n1437 | n1443 ;
  assign n1445 = ( n66 & n149 ) | ( n66 & n160 ) | ( n149 & n160 ) ;
  assign n1446 = n148 | n1445 ;
  assign n1447 = n489 | n1031 ;
  assign n1448 = ( ~n609 & n1059 ) | ( ~n609 & n1447 ) | ( n1059 & n1447 ) ;
  assign n1449 = n609 | n1448 ;
  assign n1450 = n84 & n122 ;
  assign n1451 = ( n174 & n303 ) | ( n174 & ~n1450 ) | ( n303 & ~n1450 ) ;
  assign n1452 = n1450 | n1451 ;
  assign n1453 = ( ~n1446 & n1449 ) | ( ~n1446 & n1452 ) | ( n1449 & n1452 ) ;
  assign n1454 = n1446 | n1453 ;
  assign n1455 = ( ~n1434 & n1444 ) | ( ~n1434 & n1454 ) | ( n1444 & n1454 ) ;
  assign n1456 = ( ~n1415 & n1434 ) | ( ~n1415 & n1455 ) | ( n1434 & n1455 ) ;
  assign n1457 = ( ~n1362 & n1416 ) | ( ~n1362 & n1456 ) | ( n1416 & n1456 ) ;
  assign n1458 = n1362 | n1457 ;
  assign n1459 = n382 | n855 ;
  assign n1460 = n581 | n592 ;
  assign n1461 = n1387 | n1460 ;
  assign n1462 = n301 | n353 ;
  assign n1463 = n895 | n1462 ;
  assign n1464 = ( ~n1459 & n1461 ) | ( ~n1459 & n1463 ) | ( n1461 & n1463 ) ;
  assign n1465 = ( ~n54 & n84 ) | ( ~n54 & n98 ) | ( n84 & n98 ) ;
  assign n1466 = n732 | n1465 ;
  assign n1467 = ( n1459 & n1464 ) | ( n1459 & ~n1466 ) | ( n1464 & ~n1466 ) ;
  assign n1468 = n102 | n149 ;
  assign n1469 = ( n48 & n166 ) | ( n48 & n1468 ) | ( n166 & n1468 ) ;
  assign n1470 = n538 | n782 ;
  assign n1471 = n1469 | n1470 ;
  assign n1472 = n142 | n759 ;
  assign n1473 = n294 | n302 ;
  assign n1474 = ( ~n1471 & n1472 ) | ( ~n1471 & n1473 ) | ( n1472 & n1473 ) ;
  assign n1475 = n1471 | n1474 ;
  assign n1476 = n111 | n492 ;
  assign n1477 = n66 & n216 ;
  assign n1478 = ( n433 & n441 ) | ( n433 & ~n1477 ) | ( n441 & ~n1477 ) ;
  assign n1479 = n1477 | n1478 ;
  assign n1480 = ( ~n111 & n272 ) | ( ~n111 & n1479 ) | ( n272 & n1479 ) ;
  assign n1481 = n233 | n1450 ;
  assign n1482 = n1480 | n1481 ;
  assign n1483 = n254 | n576 ;
  assign n1484 = n757 | n1483 ;
  assign n1485 = ( ~n1476 & n1482 ) | ( ~n1476 & n1484 ) | ( n1482 & n1484 ) ;
  assign n1486 = n1476 | n1485 ;
  assign n1487 = n599 | n783 ;
  assign n1488 = n360 | n1044 ;
  assign n1489 = n329 | n921 ;
  assign n1490 = n1488 | n1489 ;
  assign n1491 = n1487 | n1490 ;
  assign n1492 = n447 | n1313 ;
  assign n1493 = n227 | n947 ;
  assign n1494 = n91 | n215 ;
  assign n1495 = n1493 | n1494 ;
  assign n1496 = n226 | n1347 ;
  assign n1497 = n61 | n367 ;
  assign n1498 = n806 | n1497 ;
  assign n1499 = ( ~n1495 & n1496 ) | ( ~n1495 & n1498 ) | ( n1496 & n1498 ) ;
  assign n1500 = n1495 | n1499 ;
  assign n1501 = ( ~n1491 & n1492 ) | ( ~n1491 & n1500 ) | ( n1492 & n1500 ) ;
  assign n1502 = n1491 | n1501 ;
  assign n1503 = ( ~n1475 & n1486 ) | ( ~n1475 & n1502 ) | ( n1486 & n1502 ) ;
  assign n1504 = n1475 | n1503 ;
  assign n1505 = ( n1466 & ~n1467 ) | ( n1466 & n1504 ) | ( ~n1467 & n1504 ) ;
  assign n1506 = n1467 | n1505 ;
  assign n1507 = n352 | n928 ;
  assign n1508 = ( n146 & n312 ) | ( n146 & ~n1507 ) | ( n312 & ~n1507 ) ;
  assign n1509 = n1507 | n1508 ;
  assign n1510 = ( n75 & n136 ) | ( n75 & n145 ) | ( n136 & n145 ) ;
  assign n1511 = n76 | n641 ;
  assign n1512 = ( ~n54 & n152 ) | ( ~n54 & n160 ) | ( n152 & n160 ) ;
  assign n1513 = ( ~n1510 & n1511 ) | ( ~n1510 & n1512 ) | ( n1511 & n1512 ) ;
  assign n1514 = n1510 | n1513 ;
  assign n1515 = n81 | n1082 ;
  assign n1516 = n170 | n1225 ;
  assign n1517 = n885 | n1516 ;
  assign n1518 = ( n450 & n535 ) | ( n450 & ~n1517 ) | ( n535 & ~n1517 ) ;
  assign n1519 = n1517 | n1518 ;
  assign n1520 = ( ~n1514 & n1515 ) | ( ~n1514 & n1519 ) | ( n1515 & n1519 ) ;
  assign n1521 = n1514 | n1520 ;
  assign n1522 = n356 | n922 ;
  assign n1523 = n337 | n762 ;
  assign n1524 = ( n260 & ~n1522 ) | ( n260 & n1523 ) | ( ~n1522 & n1523 ) ;
  assign n1525 = n1522 | n1524 ;
  assign n1526 = n83 & n216 ;
  assign n1527 = ( n586 & ~n1024 ) | ( n586 & n1526 ) | ( ~n1024 & n1526 ) ;
  assign n1528 = n1024 | n1527 ;
  assign n1529 = ( ~n1521 & n1525 ) | ( ~n1521 & n1528 ) | ( n1525 & n1528 ) ;
  assign n1530 = ( n97 & n98 ) | ( n97 & n152 ) | ( n98 & n152 ) ;
  assign n1531 = n189 | n1530 ;
  assign n1532 = n267 | n567 ;
  assign n1533 = n135 | n562 ;
  assign n1534 = n444 | n796 ;
  assign n1535 = ( ~n263 & n1533 ) | ( ~n263 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1536 = n263 | n1535 ;
  assign n1537 = ( n878 & ~n1532 ) | ( n878 & n1536 ) | ( ~n1532 & n1536 ) ;
  assign n1538 = n1532 | n1537 ;
  assign n1539 = ( ~n1521 & n1531 ) | ( ~n1521 & n1538 ) | ( n1531 & n1538 ) ;
  assign n1540 = n1521 | n1539 ;
  assign n1541 = ( ~n1509 & n1529 ) | ( ~n1509 & n1540 ) | ( n1529 & n1540 ) ;
  assign n1542 = n1509 | n1541 ;
  assign n1543 = n512 | n876 ;
  assign n1544 = n217 | n719 ;
  assign n1545 = ( n175 & ~n1543 ) | ( n175 & n1544 ) | ( ~n1543 & n1544 ) ;
  assign n1546 = n1543 | n1545 ;
  assign n1547 = n544 | n590 ;
  assign n1548 = n851 | n1341 ;
  assign n1549 = n550 | n952 ;
  assign n1550 = n168 | n1549 ;
  assign n1551 = ( n685 & ~n1548 ) | ( n685 & n1550 ) | ( ~n1548 & n1550 ) ;
  assign n1552 = n1548 | n1551 ;
  assign n1553 = ( ~n1546 & n1547 ) | ( ~n1546 & n1552 ) | ( n1547 & n1552 ) ;
  assign n1554 = n1546 | n1553 ;
  assign n1555 = ( ~n1506 & n1542 ) | ( ~n1506 & n1554 ) | ( n1542 & n1554 ) ;
  assign n1556 = n59 & n102 ;
  assign n1557 = ( n1005 & n1376 ) | ( n1005 & ~n1556 ) | ( n1376 & ~n1556 ) ;
  assign n1558 = n1556 | n1557 ;
  assign n1559 = n595 | n838 ;
  assign n1560 = n164 | n1559 ;
  assign n1561 = ( n50 & n102 ) | ( n50 & n119 ) | ( n102 & n119 ) ;
  assign n1562 = ( ~n912 & n941 ) | ( ~n912 & n1561 ) | ( n941 & n1561 ) ;
  assign n1563 = n912 | n1562 ;
  assign n1564 = n286 | n565 ;
  assign n1565 = n396 | n1564 ;
  assign n1566 = ( ~n1560 & n1563 ) | ( ~n1560 & n1565 ) | ( n1563 & n1565 ) ;
  assign n1567 = ( ~n1558 & n1560 ) | ( ~n1558 & n1566 ) | ( n1560 & n1566 ) ;
  assign n1568 = n1558 | n1567 ;
  assign n1569 = ( n64 & n122 ) | ( n64 & n255 ) | ( n122 & n255 ) ;
  assign n1570 = n1085 | n1569 ;
  assign n1571 = ( ~n483 & n505 ) | ( ~n483 & n1570 ) | ( n505 & n1570 ) ;
  assign n1572 = ( n197 & n483 ) | ( n197 & ~n1571 ) | ( n483 & ~n1571 ) ;
  assign n1573 = n1571 | n1572 ;
  assign n1574 = ( ~n1554 & n1568 ) | ( ~n1554 & n1573 ) | ( n1568 & n1573 ) ;
  assign n1575 = ( ~n1506 & n1555 ) | ( ~n1506 & n1574 ) | ( n1555 & n1574 ) ;
  assign n1576 = n1506 | n1575 ;
  assign n1577 = n369 | n691 ;
  assign n1578 = n131 | n1577 ;
  assign n1579 = n1053 & ~n1578 ;
  assign n1580 = ( n368 & n550 ) | ( n368 & ~n1027 ) | ( n550 & ~n1027 ) ;
  assign n1581 = n1027 | n1580 ;
  assign n1582 = n193 | n362 ;
  assign n1583 = n293 | n360 ;
  assign n1584 = n153 | n1583 ;
  assign n1585 = ( n685 & ~n1582 ) | ( n685 & n1584 ) | ( ~n1582 & n1584 ) ;
  assign n1586 = n1582 | n1585 ;
  assign n1587 = ( ~n1578 & n1581 ) | ( ~n1578 & n1586 ) | ( n1581 & n1586 ) ;
  assign n1588 = n465 | n514 ;
  assign n1589 = n163 | n534 ;
  assign n1590 = n225 | n992 ;
  assign n1591 = ( ~n1588 & n1589 ) | ( ~n1588 & n1590 ) | ( n1589 & n1590 ) ;
  assign n1592 = n1588 | n1591 ;
  assign n1593 = n231 | n1341 ;
  assign n1594 = n592 | n746 ;
  assign n1595 = ( ~n54 & n83 ) | ( ~n54 & n102 ) | ( n83 & n102 ) ;
  assign n1596 = n189 | n1595 ;
  assign n1597 = ( ~n1593 & n1594 ) | ( ~n1593 & n1596 ) | ( n1594 & n1596 ) ;
  assign n1598 = n1593 | n1597 ;
  assign n1599 = ( n48 & n80 ) | ( n48 & n129 ) | ( n80 & n129 ) ;
  assign n1600 = ( n50 & n97 ) | ( n50 & n160 ) | ( n97 & n160 ) ;
  assign n1601 = ( ~n402 & n1472 ) | ( ~n402 & n1600 ) | ( n1472 & n1600 ) ;
  assign n1602 = ( n402 & ~n1599 ) | ( n402 & n1601 ) | ( ~n1599 & n1601 ) ;
  assign n1603 = n1599 | n1602 ;
  assign n1604 = ( ~n1592 & n1598 ) | ( ~n1592 & n1603 ) | ( n1598 & n1603 ) ;
  assign n1605 = n1592 | n1604 ;
  assign n1606 = ( n1579 & n1587 ) | ( n1579 & n1605 ) | ( n1587 & n1605 ) ;
  assign n1607 = n1579 & ~n1606 ;
  assign n1608 = n233 | n895 ;
  assign n1609 = ( n512 & n666 ) | ( n512 & ~n1608 ) | ( n666 & ~n1608 ) ;
  assign n1610 = n1608 | n1609 ;
  assign n1611 = n285 | n493 ;
  assign n1612 = n51 | n295 ;
  assign n1613 = n590 | n1612 ;
  assign n1614 = n185 | n537 ;
  assign n1615 = ( n302 & n713 ) | ( n302 & ~n1614 ) | ( n713 & ~n1614 ) ;
  assign n1616 = n1614 | n1615 ;
  assign n1617 = ( ~n1610 & n1613 ) | ( ~n1610 & n1616 ) | ( n1613 & n1616 ) ;
  assign n1618 = ( ~n1610 & n1611 ) | ( ~n1610 & n1617 ) | ( n1611 & n1617 ) ;
  assign n1619 = n1610 | n1618 ;
  assign n1620 = n440 | n947 ;
  assign n1621 = n55 | n545 ;
  assign n1622 = ( n995 & ~n1620 ) | ( n995 & n1621 ) | ( ~n1620 & n1621 ) ;
  assign n1623 = n1620 | n1622 ;
  assign n1624 = ( n57 & n116 ) | ( n57 & n160 ) | ( n116 & n160 ) ;
  assign n1625 = n810 | n856 ;
  assign n1626 = ( n66 & n122 ) | ( n66 & n149 ) | ( n122 & n149 ) ;
  assign n1627 = ( ~n1624 & n1625 ) | ( ~n1624 & n1626 ) | ( n1625 & n1626 ) ;
  assign n1628 = n1624 | n1627 ;
  assign n1629 = ( n1619 & ~n1623 ) | ( n1619 & n1628 ) | ( ~n1623 & n1628 ) ;
  assign n1630 = n301 | n675 ;
  assign n1631 = n104 | n795 ;
  assign n1632 = n92 | n167 ;
  assign n1633 = ( n81 & n587 ) | ( n81 & ~n1632 ) | ( n587 & ~n1632 ) ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = ( n1630 & ~n1631 ) | ( n1630 & n1634 ) | ( ~n1631 & n1634 ) ;
  assign n1636 = n655 | n1169 ;
  assign n1637 = ( n59 & ~n78 ) | ( n59 & n149 ) | ( ~n78 & n149 ) ;
  assign n1638 = ( n961 & ~n1636 ) | ( n961 & n1637 ) | ( ~n1636 & n1637 ) ;
  assign n1639 = n1636 | n1638 ;
  assign n1640 = ( n1631 & ~n1635 ) | ( n1631 & n1639 ) | ( ~n1635 & n1639 ) ;
  assign n1641 = n1635 | n1640 ;
  assign n1642 = ( n1623 & ~n1629 ) | ( n1623 & n1641 ) | ( ~n1629 & n1641 ) ;
  assign n1643 = n1629 | n1642 ;
  assign n1644 = n242 | n1001 ;
  assign n1645 = n549 | n1644 ;
  assign n1646 = n79 | n170 ;
  assign n1647 = n931 | n1646 ;
  assign n1648 = n1645 | n1647 ;
  assign n1649 = n60 | n318 ;
  assign n1650 = n390 | n1450 ;
  assign n1651 = n1649 | n1650 ;
  assign n1652 = n581 | n985 ;
  assign n1653 = n444 | n941 ;
  assign n1654 = ( n1012 & ~n1652 ) | ( n1012 & n1653 ) | ( ~n1652 & n1653 ) ;
  assign n1655 = n1652 | n1654 ;
  assign n1656 = ( n1056 & ~n1648 ) | ( n1056 & n1655 ) | ( ~n1648 & n1655 ) ;
  assign n1657 = ( n1648 & ~n1651 ) | ( n1648 & n1656 ) | ( ~n1651 & n1656 ) ;
  assign n1658 = n228 | n258 ;
  assign n1659 = n684 | n1658 ;
  assign n1660 = ( n66 & n166 ) | ( n66 & n216 ) | ( n166 & n216 ) ;
  assign n1661 = n596 | n1660 ;
  assign n1662 = n320 | n641 ;
  assign n1663 = ( n1487 & ~n1661 ) | ( n1487 & n1662 ) | ( ~n1661 & n1662 ) ;
  assign n1664 = n1661 | n1663 ;
  assign n1665 = ( ~n1056 & n1659 ) | ( ~n1056 & n1664 ) | ( n1659 & n1664 ) ;
  assign n1666 = n1651 | n1665 ;
  assign n1667 = n1657 | n1666 ;
  assign n1668 = ( n1607 & n1643 ) | ( n1607 & n1667 ) | ( n1643 & n1667 ) ;
  assign n1669 = n1607 & ~n1668 ;
  assign n1670 = n226 | n1436 ;
  assign n1671 = n137 | n1044 ;
  assign n1672 = n795 | n1397 ;
  assign n1673 = ( n549 & ~n1671 ) | ( n549 & n1672 ) | ( ~n1671 & n1672 ) ;
  assign n1674 = n1671 | n1673 ;
  assign n1675 = n113 | n151 ;
  assign n1676 = ( ~n1670 & n1674 ) | ( ~n1670 & n1675 ) | ( n1674 & n1675 ) ;
  assign n1677 = n1670 | n1676 ;
  assign n1678 = n231 | n433 ;
  assign n1679 = n267 | n921 ;
  assign n1680 = n338 | n956 ;
  assign n1681 = ( ~n1678 & n1679 ) | ( ~n1678 & n1680 ) | ( n1679 & n1680 ) ;
  assign n1682 = n1678 | n1681 ;
  assign n1683 = n1056 | n1624 ;
  assign n1684 = ( n913 & n963 ) | ( n913 & ~n1683 ) | ( n963 & ~n1683 ) ;
  assign n1685 = n1683 | n1684 ;
  assign n1686 = ( ~n1677 & n1682 ) | ( ~n1677 & n1685 ) | ( n1682 & n1685 ) ;
  assign n1687 = n1677 | n1686 ;
  assign n1688 = n625 | n837 ;
  assign n1689 = n171 | n465 ;
  assign n1690 = n316 | n666 ;
  assign n1691 = n1689 | n1690 ;
  assign n1692 = n64 & n97 ;
  assign n1693 = n76 | n1692 ;
  assign n1694 = n394 | n483 ;
  assign n1695 = n60 | n353 ;
  assign n1696 = ( ~n1693 & n1694 ) | ( ~n1693 & n1695 ) | ( n1694 & n1695 ) ;
  assign n1697 = n1693 | n1696 ;
  assign n1698 = ( ~n1688 & n1691 ) | ( ~n1688 & n1697 ) | ( n1691 & n1697 ) ;
  assign n1699 = n528 | n609 ;
  assign n1700 = n356 | n1699 ;
  assign n1701 = ( n59 & n102 ) | ( n59 & n149 ) | ( n102 & n149 ) ;
  assign n1702 = n565 | n1701 ;
  assign n1703 = ( n1600 & ~n1700 ) | ( n1600 & n1702 ) | ( ~n1700 & n1702 ) ;
  assign n1704 = ( n1312 & n1700 ) | ( n1312 & ~n1703 ) | ( n1700 & ~n1703 ) ;
  assign n1705 = n1703 | n1704 ;
  assign n1706 = ( n1688 & ~n1698 ) | ( n1688 & n1705 ) | ( ~n1698 & n1705 ) ;
  assign n1707 = n1698 | n1706 ;
  assign n1708 = n168 | n440 ;
  assign n1709 = n300 | n1708 ;
  assign n1710 = n153 | n212 ;
  assign n1711 = n529 | n764 ;
  assign n1712 = n286 | n1711 ;
  assign n1713 = ( ~n1709 & n1710 ) | ( ~n1709 & n1712 ) | ( n1710 & n1712 ) ;
  assign n1714 = n1709 | n1713 ;
  assign n1715 = n455 | n917 ;
  assign n1716 = n537 | n1341 ;
  assign n1717 = n1715 | n1716 ;
  assign n1718 = n146 | n217 ;
  assign n1719 = n523 | n1225 ;
  assign n1720 = n786 | n1477 ;
  assign n1721 = n1426 | n1720 ;
  assign n1722 = n81 | n493 ;
  assign n1723 = ( ~n1719 & n1721 ) | ( ~n1719 & n1722 ) | ( n1721 & n1722 ) ;
  assign n1724 = n1719 | n1723 ;
  assign n1725 = ( ~n1717 & n1718 ) | ( ~n1717 & n1724 ) | ( n1718 & n1724 ) ;
  assign n1726 = n1717 | n1725 ;
  assign n1727 = ( ~n54 & n66 ) | ( ~n54 & n119 ) | ( n66 & n119 ) ;
  assign n1728 = n947 | n1727 ;
  assign n1729 = n867 | n1728 ;
  assign n1730 = n1726 | n1729 ;
  assign n1731 = n79 | n760 ;
  assign n1732 = n135 | n265 ;
  assign n1733 = ( ~n435 & n836 ) | ( ~n435 & n1732 ) | ( n836 & n1732 ) ;
  assign n1734 = ( n435 & ~n1731 ) | ( n435 & n1733 ) | ( ~n1731 & n1733 ) ;
  assign n1735 = n1731 | n1734 ;
  assign n1736 = n67 | n230 ;
  assign n1737 = n233 | n865 ;
  assign n1738 = n1736 | n1737 ;
  assign n1739 = n173 | n1027 ;
  assign n1740 = ( n384 & n757 ) | ( n384 & ~n1739 ) | ( n757 & ~n1739 ) ;
  assign n1741 = n1739 | n1740 ;
  assign n1742 = n218 & ~n685 ;
  assign n1743 = ( n1738 & ~n1741 ) | ( n1738 & n1742 ) | ( ~n1741 & n1742 ) ;
  assign n1744 = ~n1738 & n1743 ;
  assign n1745 = ( n1729 & ~n1735 ) | ( n1729 & n1744 ) | ( ~n1735 & n1744 ) ;
  assign n1746 = ( n1714 & ~n1730 ) | ( n1714 & n1745 ) | ( ~n1730 & n1745 ) ;
  assign n1747 = ~n1714 & n1746 ;
  assign n1748 = ( n1396 & ~n1707 ) | ( n1396 & n1747 ) | ( ~n1707 & n1747 ) ;
  assign n1749 = ( ~n1396 & n1687 ) | ( ~n1396 & n1748 ) | ( n1687 & n1748 ) ;
  assign n1750 = ~n1687 & n1749 ;
  assign n1751 = n255 | n266 ;
  assign n1752 = n224 | n1751 ;
  assign n1753 = ( n50 & n97 ) | ( n50 & n145 ) | ( n97 & n145 ) ;
  assign n1754 = ( n59 & n72 ) | ( n59 & n109 ) | ( n72 & n109 ) ;
  assign n1755 = n1006 | n1754 ;
  assign n1756 = ( ~n1752 & n1753 ) | ( ~n1752 & n1755 ) | ( n1753 & n1755 ) ;
  assign n1757 = n1752 | n1756 ;
  assign n1758 = n117 | n922 ;
  assign n1759 = n1144 | n1758 ;
  assign n1760 = ( n80 & n83 ) | ( n80 & n136 ) | ( n83 & n136 ) ;
  assign n1761 = ( n83 & n119 ) | ( n83 & n166 ) | ( n119 & n166 ) ;
  assign n1762 = n230 | n1761 ;
  assign n1763 = n132 | n259 ;
  assign n1764 = ( ~n1760 & n1762 ) | ( ~n1760 & n1763 ) | ( n1762 & n1763 ) ;
  assign n1765 = n1760 | n1764 ;
  assign n1766 = ( n111 & n174 ) | ( n111 & ~n538 ) | ( n174 & ~n538 ) ;
  assign n1767 = n538 | n1766 ;
  assign n1768 = ( ~n1759 & n1765 ) | ( ~n1759 & n1767 ) | ( n1765 & n1767 ) ;
  assign n1769 = n1759 | n1768 ;
  assign n1770 = n285 | n562 ;
  assign n1771 = ( n142 & n566 ) | ( n142 & ~n1770 ) | ( n566 & ~n1770 ) ;
  assign n1772 = n1770 | n1771 ;
  assign n1773 = n544 | n1363 ;
  assign n1774 = n1313 | n1510 ;
  assign n1775 = n540 | n1774 ;
  assign n1776 = ( ~n1772 & n1773 ) | ( ~n1772 & n1775 ) | ( n1773 & n1775 ) ;
  assign n1777 = n1772 | n1776 ;
  assign n1778 = n1769 | n1777 ;
  assign n1779 = n189 | n395 ;
  assign n1780 = n1171 | n1779 ;
  assign n1781 = n60 | n272 ;
  assign n1782 = n576 | n775 ;
  assign n1783 = n98 & ~n717 ;
  assign n1784 = ( n98 & n1782 ) | ( n98 & ~n1783 ) | ( n1782 & ~n1783 ) ;
  assign n1785 = ( n203 & ~n1781 ) | ( n203 & n1784 ) | ( ~n1781 & n1784 ) ;
  assign n1786 = n1781 | n1785 ;
  assign n1787 = ( ~n1777 & n1780 ) | ( ~n1777 & n1786 ) | ( n1780 & n1786 ) ;
  assign n1788 = ( ~n1757 & n1778 ) | ( ~n1757 & n1787 ) | ( n1778 & n1787 ) ;
  assign n1789 = n1757 | n1788 ;
  assign n1790 = n91 | n137 ;
  assign n1791 = n857 | n1790 ;
  assign n1792 = n1365 | n1526 ;
  assign n1793 = n195 | n507 ;
  assign n1794 = ( ~n368 & n449 ) | ( ~n368 & n1024 ) | ( n449 & n1024 ) ;
  assign n1795 = ( n368 & ~n1793 ) | ( n368 & n1794 ) | ( ~n1793 & n1794 ) ;
  assign n1796 = n1793 | n1795 ;
  assign n1797 = ( ~n1791 & n1792 ) | ( ~n1791 & n1796 ) | ( n1792 & n1796 ) ;
  assign n1798 = n225 | n719 ;
  assign n1799 = n211 | n1595 ;
  assign n1800 = n338 | n689 ;
  assign n1801 = ( ~n1798 & n1799 ) | ( ~n1798 & n1800 ) | ( n1799 & n1800 ) ;
  assign n1802 = n1798 | n1801 ;
  assign n1803 = ( n1791 & n1797 ) | ( n1791 & ~n1802 ) | ( n1797 & ~n1802 ) ;
  assign n1804 = n483 | n655 ;
  assign n1805 = ( n661 & n1563 ) | ( n661 & ~n1804 ) | ( n1563 & ~n1804 ) ;
  assign n1806 = n1804 | n1805 ;
  assign n1807 = n789 | n1523 ;
  assign n1808 = n196 | n466 ;
  assign n1809 = ( ~n193 & n517 ) | ( ~n193 & n1808 ) | ( n517 & n1808 ) ;
  assign n1810 = n1559 | n1809 ;
  assign n1811 = ( n83 & n109 ) | ( n83 & n166 ) | ( n109 & n166 ) ;
  assign n1812 = ( n590 & ~n1810 ) | ( n590 & n1811 ) | ( ~n1810 & n1811 ) ;
  assign n1813 = n1810 | n1812 ;
  assign n1814 = n273 | n642 ;
  assign n1815 = ( n163 & n215 ) | ( n163 & ~n1814 ) | ( n215 & ~n1814 ) ;
  assign n1816 = n1814 | n1815 ;
  assign n1817 = ( ~n1807 & n1813 ) | ( ~n1807 & n1816 ) | ( n1813 & n1816 ) ;
  assign n1818 = n1807 | n1817 ;
  assign n1819 = ( ~n589 & n1806 ) | ( ~n589 & n1818 ) | ( n1806 & n1818 ) ;
  assign n1820 = n589 | n1819 ;
  assign n1821 = ( n1802 & ~n1803 ) | ( n1802 & n1820 ) | ( ~n1803 & n1820 ) ;
  assign n1822 = n1803 | n1821 ;
  assign n1823 = ( n75 & n119 ) | ( n75 & n129 ) | ( n119 & n129 ) ;
  assign n1824 = n131 | n1823 ;
  assign n1825 = ( n83 & n102 ) | ( n83 & n122 ) | ( n102 & n122 ) ;
  assign n1826 = n1660 | n1825 ;
  assign n1827 = n242 | n1826 ;
  assign n1828 = ( n202 & n1116 ) | ( n202 & ~n1827 ) | ( n1116 & ~n1827 ) ;
  assign n1829 = n1827 | n1828 ;
  assign n1830 = n120 | n352 ;
  assign n1831 = n591 | n1830 ;
  assign n1832 = ( n1002 & n1197 ) | ( n1002 & ~n1831 ) | ( n1197 & ~n1831 ) ;
  assign n1833 = n1831 | n1832 ;
  assign n1834 = ( n1824 & n1829 ) | ( n1824 & ~n1833 ) | ( n1829 & ~n1833 ) ;
  assign n1835 = n197 | n340 ;
  assign n1836 = ( n112 & ~n291 ) | ( n112 & n1835 ) | ( ~n291 & n1835 ) ;
  assign n1837 = n291 | n1836 ;
  assign n1838 = n212 | n759 ;
  assign n1839 = n188 | n353 ;
  assign n1840 = ( n1009 & ~n1737 ) | ( n1009 & n1839 ) | ( ~n1737 & n1839 ) ;
  assign n1841 = ( n1737 & ~n1838 ) | ( n1737 & n1840 ) | ( ~n1838 & n1840 ) ;
  assign n1842 = n1838 | n1841 ;
  assign n1843 = ( n1564 & n1593 ) | ( n1564 & ~n1842 ) | ( n1593 & ~n1842 ) ;
  assign n1844 = n1842 | n1843 ;
  assign n1845 = ( n103 & n329 ) | ( n103 & ~n1423 ) | ( n329 & ~n1423 ) ;
  assign n1846 = n1423 | n1845 ;
  assign n1847 = ( ~n1837 & n1844 ) | ( ~n1837 & n1846 ) | ( n1844 & n1846 ) ;
  assign n1848 = n1837 | n1847 ;
  assign n1849 = ( n1833 & ~n1834 ) | ( n1833 & n1848 ) | ( ~n1834 & n1848 ) ;
  assign n1850 = n1834 | n1849 ;
  assign n1851 = ( ~n1789 & n1822 ) | ( ~n1789 & n1850 ) | ( n1822 & n1850 ) ;
  assign n1852 = n1789 | n1851 ;
  assign n1853 = ( n41 & n136 ) | ( n41 & n149 ) | ( n136 & n149 ) ;
  assign n1854 = n595 | n1853 ;
  assign n1855 = ( n500 & n1110 ) | ( n500 & ~n1854 ) | ( n1110 & ~n1854 ) ;
  assign n1856 = n1854 | n1855 ;
  assign n1857 = n92 | n215 ;
  assign n1858 = ( n173 & n753 ) | ( n173 & ~n1857 ) | ( n753 & ~n1857 ) ;
  assign n1859 = n1857 | n1858 ;
  assign n1860 = n298 | n876 ;
  assign n1861 = n301 | n338 ;
  assign n1862 = ( ~n1859 & n1860 ) | ( ~n1859 & n1861 ) | ( n1860 & n1861 ) ;
  assign n1863 = n1859 | n1862 ;
  assign n1864 = n186 | n395 ;
  assign n1865 = n367 | n1096 ;
  assign n1866 = ( n647 & ~n1864 ) | ( n647 & n1865 ) | ( ~n1864 & n1865 ) ;
  assign n1867 = n1864 | n1866 ;
  assign n1868 = ( ~n1856 & n1863 ) | ( ~n1856 & n1867 ) | ( n1863 & n1867 ) ;
  assign n1869 = n317 | n1225 ;
  assign n1870 = ( ~n54 & n57 ) | ( ~n54 & n129 ) | ( n57 & n129 ) ;
  assign n1871 = n1306 | n1870 ;
  assign n1872 = ( n1711 & n1790 ) | ( n1711 & ~n1871 ) | ( n1790 & ~n1871 ) ;
  assign n1873 = n1871 | n1872 ;
  assign n1874 = ( n507 & ~n1869 ) | ( n507 & n1873 ) | ( ~n1869 & n1873 ) ;
  assign n1875 = n1869 | n1874 ;
  assign n1876 = ( n1856 & ~n1868 ) | ( n1856 & n1875 ) | ( ~n1868 & n1875 ) ;
  assign n1877 = n1868 | n1876 ;
  assign n1878 = n402 | n1515 ;
  assign n1879 = n1692 | n1736 ;
  assign n1880 = ( n44 & n72 ) | ( n44 & n97 ) | ( n72 & n97 ) ;
  assign n1881 = n197 | n1880 ;
  assign n1882 = ( ~n1878 & n1879 ) | ( ~n1878 & n1881 ) | ( n1879 & n1881 ) ;
  assign n1883 = n1878 | n1882 ;
  assign n1884 = n206 | n488 ;
  assign n1885 = ( n153 & n259 ) | ( n153 & ~n1884 ) | ( n259 & ~n1884 ) ;
  assign n1886 = n1884 | n1885 ;
  assign n1887 = n320 | n1376 ;
  assign n1888 = ( n1511 & ~n1886 ) | ( n1511 & n1887 ) | ( ~n1886 & n1887 ) ;
  assign n1889 = n1886 | n1888 ;
  assign n1890 = n466 | n1547 ;
  assign n1891 = n192 | n662 ;
  assign n1892 = n483 | n952 ;
  assign n1893 = n786 | n917 ;
  assign n1894 = ( ~n1718 & n1892 ) | ( ~n1718 & n1893 ) | ( n1892 & n1893 ) ;
  assign n1895 = ( n1718 & ~n1891 ) | ( n1718 & n1894 ) | ( ~n1891 & n1894 ) ;
  assign n1896 = n1891 | n1895 ;
  assign n1897 = n45 | n352 ;
  assign n1898 = n523 | n1897 ;
  assign n1899 = ( ~n1890 & n1896 ) | ( ~n1890 & n1898 ) | ( n1896 & n1898 ) ;
  assign n1900 = n1890 | n1899 ;
  assign n1901 = ( ~n1883 & n1889 ) | ( ~n1883 & n1900 ) | ( n1889 & n1900 ) ;
  assign n1902 = n170 | n353 ;
  assign n1903 = ( n84 & n98 ) | ( n84 & n109 ) | ( n98 & n109 ) ;
  assign n1904 = ( n886 & ~n1902 ) | ( n886 & n1903 ) | ( ~n1902 & n1903 ) ;
  assign n1905 = n1902 | n1904 ;
  assign n1906 = ( n393 & n608 ) | ( n393 & ~n1905 ) | ( n608 & ~n1905 ) ;
  assign n1907 = n1905 | n1906 ;
  assign n1908 = n104 | n1277 ;
  assign n1909 = n1078 | n1313 ;
  assign n1910 = ( n1907 & n1908 ) | ( n1907 & ~n1909 ) | ( n1908 & ~n1909 ) ;
  assign n1911 = n315 | n691 ;
  assign n1912 = n240 | n536 ;
  assign n1913 = n1589 | n1912 ;
  assign n1914 = n74 | n796 ;
  assign n1915 = n824 | n865 ;
  assign n1916 = n499 | n513 ;
  assign n1917 = ( ~n1914 & n1915 ) | ( ~n1914 & n1916 ) | ( n1915 & n1916 ) ;
  assign n1918 = n1914 | n1917 ;
  assign n1919 = ( ~n1911 & n1913 ) | ( ~n1911 & n1918 ) | ( n1913 & n1918 ) ;
  assign n1920 = n1911 | n1919 ;
  assign n1921 = ( n1909 & ~n1910 ) | ( n1909 & n1920 ) | ( ~n1910 & n1920 ) ;
  assign n1922 = n1910 | n1921 ;
  assign n1923 = ( n1486 & ~n1883 ) | ( n1486 & n1922 ) | ( ~n1883 & n1922 ) ;
  assign n1924 = n1883 | n1923 ;
  assign n1925 = ( ~n1877 & n1901 ) | ( ~n1877 & n1924 ) | ( n1901 & n1924 ) ;
  assign n1926 = n1877 | n1925 ;
  assign n1927 = n263 | n1435 ;
  assign n1928 = n873 | n1116 ;
  assign n1929 = n1110 | n1450 ;
  assign n1930 = ( n750 & ~n1914 ) | ( n750 & n1929 ) | ( ~n1914 & n1929 ) ;
  assign n1931 = ( n1914 & ~n1928 ) | ( n1914 & n1930 ) | ( ~n1928 & n1930 ) ;
  assign n1932 = n1928 | n1931 ;
  assign n1933 = n285 | n435 ;
  assign n1934 = ( n259 & n810 ) | ( n259 & ~n1933 ) | ( n810 & ~n1933 ) ;
  assign n1935 = n1933 | n1934 ;
  assign n1936 = ( ~n1927 & n1932 ) | ( ~n1927 & n1935 ) | ( n1932 & n1935 ) ;
  assign n1937 = n1927 | n1936 ;
  assign n1938 = n512 | n775 ;
  assign n1939 = n111 | n587 ;
  assign n1940 = n211 | n613 ;
  assign n1941 = n1569 | n1940 ;
  assign n1942 = ( ~n1938 & n1939 ) | ( ~n1938 & n1941 ) | ( n1939 & n1941 ) ;
  assign n1943 = n1938 | n1942 ;
  assign n1944 = ( n866 & n1366 ) | ( n866 & ~n1711 ) | ( n1366 & ~n1711 ) ;
  assign n1945 = n1711 | n1944 ;
  assign n1946 = n960 | n1365 ;
  assign n1947 = ( ~n78 & n97 ) | ( ~n78 & n116 ) | ( n97 & n116 ) ;
  assign n1948 = n565 | n1947 ;
  assign n1949 = ( n173 & n227 ) | ( n173 & ~n1948 ) | ( n227 & ~n1948 ) ;
  assign n1950 = n1948 | n1949 ;
  assign n1951 = ( n75 & n149 ) | ( n75 & n1082 ) | ( n149 & n1082 ) ;
  assign n1952 = ( ~n1946 & n1950 ) | ( ~n1946 & n1951 ) | ( n1950 & n1951 ) ;
  assign n1953 = ( ~n1945 & n1946 ) | ( ~n1945 & n1952 ) | ( n1946 & n1952 ) ;
  assign n1954 = ( ~n1943 & n1945 ) | ( ~n1943 & n1953 ) | ( n1945 & n1953 ) ;
  assign n1955 = n1943 | n1954 ;
  assign n1956 = ( n671 & n1937 ) | ( n671 & ~n1955 ) | ( n1937 & ~n1955 ) ;
  assign n1957 = ~n1937 & n1956 ;
  assign n1958 = ( n50 & n83 ) | ( n50 & n109 ) | ( n83 & n109 ) ;
  assign n1959 = ( n759 & n886 ) | ( n759 & ~n1958 ) | ( n886 & ~n1958 ) ;
  assign n1960 = n1958 | n1959 ;
  assign n1961 = n267 | n507 ;
  assign n1962 = ( n177 & n230 ) | ( n177 & ~n1961 ) | ( n230 & ~n1961 ) ;
  assign n1963 = n1961 | n1962 ;
  assign n1964 = n164 | n566 ;
  assign n1965 = ( n857 & ~n978 ) | ( n857 & n1964 ) | ( ~n978 & n1964 ) ;
  assign n1966 = n978 | n1965 ;
  assign n1967 = n51 | n168 ;
  assign n1968 = ( ~n1079 & n1122 ) | ( ~n1079 & n1967 ) | ( n1122 & n1967 ) ;
  assign n1969 = n1079 | n1968 ;
  assign n1970 = ( n1113 & ~n1966 ) | ( n1113 & n1969 ) | ( ~n1966 & n1969 ) ;
  assign n1971 = n1966 | n1970 ;
  assign n1972 = ( n1960 & ~n1963 ) | ( n1960 & n1971 ) | ( ~n1963 & n1971 ) ;
  assign n1973 = n1645 | n1972 ;
  assign n1974 = ( n75 & n100 ) | ( n75 & n166 ) | ( n100 & n166 ) ;
  assign n1975 = n1320 | n1974 ;
  assign n1976 = n514 | n734 ;
  assign n1977 = n103 | n1169 ;
  assign n1978 = n277 | n1977 ;
  assign n1979 = n205 | n933 ;
  assign n1980 = n567 | n1979 ;
  assign n1981 = n76 | n395 ;
  assign n1982 = ( n272 & n947 ) | ( n272 & ~n1981 ) | ( n947 & ~n1981 ) ;
  assign n1983 = n1981 | n1982 ;
  assign n1984 = ( ~n1978 & n1980 ) | ( ~n1978 & n1983 ) | ( n1980 & n1983 ) ;
  assign n1985 = n1978 | n1984 ;
  assign n1986 = ( ~n1975 & n1976 ) | ( ~n1975 & n1985 ) | ( n1976 & n1985 ) ;
  assign n1987 = n1975 | n1986 ;
  assign n1988 = ( n1963 & ~n1973 ) | ( n1963 & n1987 ) | ( ~n1973 & n1987 ) ;
  assign n1989 = n1973 | n1988 ;
  assign n1990 = n646 | n729 ;
  assign n1991 = ( n66 & n119 ) | ( n66 & n145 ) | ( n119 & n145 ) ;
  assign n1992 = ( n941 & n1710 ) | ( n941 & ~n1991 ) | ( n1710 & ~n1991 ) ;
  assign n1993 = n1991 | n1992 ;
  assign n1994 = ( n294 & n485 ) | ( n294 & ~n1773 ) | ( n485 & ~n1773 ) ;
  assign n1995 = n1773 | n1994 ;
  assign n1996 = ( ~n1990 & n1993 ) | ( ~n1990 & n1995 ) | ( n1993 & n1995 ) ;
  assign n1997 = n1990 | n1996 ;
  assign n1998 = n312 | n488 ;
  assign n1999 = n1205 | n1998 ;
  assign n2000 = n197 | n753 ;
  assign n2001 = ( n59 & n84 ) | ( n59 & n136 ) | ( n84 & n136 ) ;
  assign n2002 = ( n80 & n119 ) | ( n80 & n129 ) | ( n119 & n129 ) ;
  assign n2003 = ( n225 & n824 ) | ( n225 & ~n2002 ) | ( n824 & ~n2002 ) ;
  assign n2004 = n2002 | n2003 ;
  assign n2005 = ( ~n2000 & n2001 ) | ( ~n2000 & n2004 ) | ( n2001 & n2004 ) ;
  assign n2006 = n2000 | n2005 ;
  assign n2007 = ( n448 & ~n500 ) | ( n448 & n582 ) | ( ~n500 & n582 ) ;
  assign n2008 = n500 | n2007 ;
  assign n2009 = ( ~n1999 & n2006 ) | ( ~n1999 & n2008 ) | ( n2006 & n2008 ) ;
  assign n2010 = n1999 | n2009 ;
  assign n2011 = n952 | n1313 ;
  assign n2012 = n361 | n895 ;
  assign n2013 = ( n172 & ~n2011 ) | ( n172 & n2012 ) | ( ~n2011 & n2012 ) ;
  assign n2014 = ( n837 & n2011 ) | ( n837 & ~n2013 ) | ( n2011 & ~n2013 ) ;
  assign n2015 = n2013 | n2014 ;
  assign n2016 = ( n98 & n152 ) | ( n98 & n160 ) | ( n152 & n160 ) ;
  assign n2017 = ( n517 & n1531 ) | ( n517 & ~n2016 ) | ( n1531 & ~n2016 ) ;
  assign n2018 = n2016 | n2017 ;
  assign n2019 = ( ~n2010 & n2015 ) | ( ~n2010 & n2018 ) | ( n2015 & n2018 ) ;
  assign n2020 = ( ~n1997 & n2010 ) | ( ~n1997 & n2019 ) | ( n2010 & n2019 ) ;
  assign n2021 = n1997 | n2020 ;
  assign n2022 = ( n1957 & n1989 ) | ( n1957 & n2021 ) | ( n1989 & n2021 ) ;
  assign n2023 = n1957 & ~n2022 ;
  assign n2024 = n419 | n1009 ;
  assign n2025 = n1146 | n1774 ;
  assign n2026 = ( n527 & ~n2024 ) | ( n527 & n2025 ) | ( ~n2024 & n2025 ) ;
  assign n2027 = n1612 | n1835 ;
  assign n2028 = n1692 | n2027 ;
  assign n2029 = n215 | n550 ;
  assign n2030 = ( n196 & n234 ) | ( n196 & ~n2029 ) | ( n234 & ~n2029 ) ;
  assign n2031 = n2029 | n2030 ;
  assign n2032 = n146 | n331 ;
  assign n2033 = n642 | n775 ;
  assign n2034 = ( ~n2031 & n2032 ) | ( ~n2031 & n2033 ) | ( n2032 & n2033 ) ;
  assign n2035 = n2031 | n2034 ;
  assign n2036 = ( n1950 & n2028 ) | ( n1950 & ~n2035 ) | ( n2028 & ~n2035 ) ;
  assign n2037 = n2026 | n2036 ;
  assign n2038 = n2024 | n2037 ;
  assign n2039 = ( n576 & n1068 ) | ( n576 & ~n1993 ) | ( n1068 & ~n1993 ) ;
  assign n2040 = n1993 | n2039 ;
  assign n2041 = ( n2035 & ~n2038 ) | ( n2035 & n2040 ) | ( ~n2038 & n2040 ) ;
  assign n2042 = n2038 | n2041 ;
  assign n2043 = ( n41 & n44 ) | ( n41 & n66 ) | ( n44 & n66 ) ;
  assign n2044 = ( n534 & n590 ) | ( n534 & ~n2043 ) | ( n590 & ~n2043 ) ;
  assign n2045 = n2043 | n2044 ;
  assign n2046 = n537 | n613 ;
  assign n2047 = n824 | n2046 ;
  assign n2048 = n1389 | n2047 ;
  assign n2049 = n171 | n186 ;
  assign n2050 = ( n455 & n952 ) | ( n455 & ~n2049 ) | ( n952 & ~n2049 ) ;
  assign n2051 = n2049 | n2050 ;
  assign n2052 = n922 | n1366 ;
  assign n2053 = n394 | n985 ;
  assign n2054 = ( ~n2051 & n2052 ) | ( ~n2051 & n2053 ) | ( n2052 & n2053 ) ;
  assign n2055 = n2051 | n2054 ;
  assign n2056 = ( ~n2045 & n2048 ) | ( ~n2045 & n2055 ) | ( n2048 & n2055 ) ;
  assign n2057 = n2045 | n2056 ;
  assign n2058 = n177 | n581 ;
  assign n2059 = n67 | n536 ;
  assign n2060 = n161 | n2059 ;
  assign n2061 = ( n1489 & n1793 ) | ( n1489 & ~n2060 ) | ( n1793 & ~n2060 ) ;
  assign n2062 = n2060 | n2061 ;
  assign n2063 = ( n302 & ~n2058 ) | ( n302 & n2062 ) | ( ~n2058 & n2062 ) ;
  assign n2064 = n2058 | n2063 ;
  assign n2065 = ( ~n2042 & n2057 ) | ( ~n2042 & n2064 ) | ( n2057 & n2064 ) ;
  assign n2066 = n960 | n1595 ;
  assign n2067 = n144 | n762 ;
  assign n2068 = ( n1700 & ~n2066 ) | ( n1700 & n2067 ) | ( ~n2066 & n2067 ) ;
  assign n2069 = n2066 | n2068 ;
  assign n2070 = n448 | n487 ;
  assign n2071 = n895 | n1225 ;
  assign n2072 = n977 | n1376 ;
  assign n2073 = n120 | n185 ;
  assign n2074 = ( ~n494 & n2072 ) | ( ~n494 & n2073 ) | ( n2072 & n2073 ) ;
  assign n2075 = ( n494 & ~n2071 ) | ( n494 & n2074 ) | ( ~n2071 & n2074 ) ;
  assign n2076 = n2071 | n2075 ;
  assign n2077 = n258 | n433 ;
  assign n2078 = n272 | n806 ;
  assign n2079 = n1792 | n2078 ;
  assign n2080 = n208 | n567 ;
  assign n2081 = n150 | n1027 ;
  assign n2082 = n2080 | n2081 ;
  assign n2083 = n2079 | n2082 ;
  assign n2084 = n2077 | n2083 ;
  assign n2085 = n2076 | n2084 ;
  assign n2086 = n2070 | n2085 ;
  assign n2087 = ( ~n2064 & n2069 ) | ( ~n2064 & n2086 ) | ( n2069 & n2086 ) ;
  assign n2088 = ( ~n2042 & n2065 ) | ( ~n2042 & n2087 ) | ( n2065 & n2087 ) ;
  assign n2089 = n2042 | n2088 ;
  assign n2090 = n144 | n337 ;
  assign n2091 = ( n1171 & n1237 ) | ( n1171 & ~n2090 ) | ( n1237 & ~n2090 ) ;
  assign n2092 = n2090 | n2091 ;
  assign n2093 = n536 | n1169 ;
  assign n2094 = n440 | n567 ;
  assign n2095 = ( n215 & n505 ) | ( n215 & ~n2094 ) | ( n505 & ~n2094 ) ;
  assign n2096 = n2094 | n2095 ;
  assign n2097 = ( ~n2092 & n2093 ) | ( ~n2092 & n2096 ) | ( n2093 & n2096 ) ;
  assign n2098 = n2092 | n2097 ;
  assign n2099 = n60 | n544 ;
  assign n2100 = n662 | n806 ;
  assign n2101 = ( n356 & ~n2099 ) | ( n356 & n2100 ) | ( ~n2099 & n2100 ) ;
  assign n2102 = n2099 | n2101 ;
  assign n2103 = ( n1588 & n1600 ) | ( n1588 & ~n2102 ) | ( n1600 & ~n2102 ) ;
  assign n2104 = n2102 | n2103 ;
  assign n2105 = ( n44 & n97 ) | ( n44 & n152 ) | ( n97 & n152 ) ;
  assign n2106 = n1560 | n1762 ;
  assign n2107 = n171 | n504 ;
  assign n2108 = n661 | n2107 ;
  assign n2109 = ( ~n54 & n152 ) | ( ~n54 & n166 ) | ( n152 & n166 ) ;
  assign n2110 = ( n301 & n529 ) | ( n301 & ~n2109 ) | ( n529 & ~n2109 ) ;
  assign n2111 = n2109 | n2110 ;
  assign n2112 = ( ~n2106 & n2108 ) | ( ~n2106 & n2111 ) | ( n2108 & n2111 ) ;
  assign n2113 = ( ~n2105 & n2106 ) | ( ~n2105 & n2112 ) | ( n2106 & n2112 ) ;
  assign n2114 = n2105 | n2113 ;
  assign n2115 = ( ~n2098 & n2104 ) | ( ~n2098 & n2114 ) | ( n2104 & n2114 ) ;
  assign n2116 = n2098 | n2115 ;
  assign n2117 = n130 | n444 ;
  assign n2118 = ( n73 & n83 ) | ( n73 & n145 ) | ( n83 & n145 ) ;
  assign n2119 = n101 | n2118 ;
  assign n2120 = ( n582 & n2117 ) | ( n582 & ~n2119 ) | ( n2117 & ~n2119 ) ;
  assign n2121 = ( n361 & n719 ) | ( n361 & ~n947 ) | ( n719 & ~n947 ) ;
  assign n2122 = n947 | n2121 ;
  assign n2123 = ( n2119 & ~n2120 ) | ( n2119 & n2122 ) | ( ~n2120 & n2122 ) ;
  assign n2124 = n2120 | n2123 ;
  assign n2125 = n1688 | n1838 ;
  assign n2126 = n45 | n762 ;
  assign n2127 = n51 | n227 ;
  assign n2128 = n545 | n2127 ;
  assign n2129 = ( ~n259 & n550 ) | ( ~n259 & n679 ) | ( n550 & n679 ) ;
  assign n2130 = n259 | n2129 ;
  assign n2131 = ( n66 & n102 ) | ( n66 & n160 ) | ( n102 & n160 ) ;
  assign n2132 = ( n581 & n764 ) | ( n581 & ~n2131 ) | ( n764 & ~n2131 ) ;
  assign n2133 = n2131 | n2132 ;
  assign n2134 = ( ~n2128 & n2130 ) | ( ~n2128 & n2133 ) | ( n2130 & n2133 ) ;
  assign n2135 = n2128 | n2134 ;
  assign n2136 = ( ~n2125 & n2126 ) | ( ~n2125 & n2135 ) | ( n2126 & n2135 ) ;
  assign n2137 = n2125 | n2136 ;
  assign n2138 = n383 | n1024 ;
  assign n2139 = ( n1625 & n1680 ) | ( n1625 & ~n2138 ) | ( n1680 & ~n2138 ) ;
  assign n2140 = n2138 | n2139 ;
  assign n2141 = ( ~n2124 & n2137 ) | ( ~n2124 & n2140 ) | ( n2137 & n2140 ) ;
  assign n2142 = n2124 | n2141 ;
  assign n2143 = n154 | n600 ;
  assign n2144 = n111 | n120 ;
  assign n2145 = n382 | n2144 ;
  assign n2146 = n234 | n479 ;
  assign n2147 = n261 | n992 ;
  assign n2148 = ( n775 & n890 ) | ( n775 & ~n2147 ) | ( n890 & ~n2147 ) ;
  assign n2149 = n2147 | n2148 ;
  assign n2150 = ( ~n2145 & n2146 ) | ( ~n2145 & n2149 ) | ( n2146 & n2149 ) ;
  assign n2151 = n2145 | n2150 ;
  assign n2152 = n360 | n447 ;
  assign n2153 = ( n492 & n642 ) | ( n492 & ~n2152 ) | ( n642 & ~n2152 ) ;
  assign n2154 = n2152 | n2153 ;
  assign n2155 = ( ~n2143 & n2151 ) | ( ~n2143 & n2154 ) | ( n2151 & n2154 ) ;
  assign n2156 = n2143 | n2155 ;
  assign n2157 = ( ~n2116 & n2142 ) | ( ~n2116 & n2156 ) | ( n2142 & n2156 ) ;
  assign n2158 = n732 | n1048 ;
  assign n2159 = n203 | n2158 ;
  assign n2160 = ( n1057 & n1510 ) | ( n1057 & ~n2159 ) | ( n1510 & ~n2159 ) ;
  assign n2161 = n2159 | n2160 ;
  assign n2162 = n1145 | n1914 ;
  assign n2163 = n488 | n517 ;
  assign n2164 = n331 | n666 ;
  assign n2165 = ( n865 & n1027 ) | ( n865 & ~n2164 ) | ( n1027 & ~n2164 ) ;
  assign n2166 = n2164 | n2165 ;
  assign n2167 = n132 | n483 ;
  assign n2168 = ( n118 & ~n2166 ) | ( n118 & n2167 ) | ( ~n2166 & n2167 ) ;
  assign n2169 = n2166 | n2168 ;
  assign n2170 = ( ~n2162 & n2163 ) | ( ~n2162 & n2169 ) | ( n2163 & n2169 ) ;
  assign n2171 = n2162 | n2170 ;
  assign n2172 = ( ~n2156 & n2161 ) | ( ~n2156 & n2171 ) | ( n2161 & n2171 ) ;
  assign n2173 = ( ~n2116 & n2157 ) | ( ~n2116 & n2172 ) | ( n2157 & n2172 ) ;
  assign n2174 = n2116 | n2173 ;
  assign n2175 = n981 | n1711 ;
  assign n2176 = n104 | n273 ;
  assign n2177 = ( n165 & n1074 ) | ( n165 & ~n2176 ) | ( n1074 & ~n2176 ) ;
  assign n2178 = n2176 | n2177 ;
  assign n2179 = ( n781 & ~n2175 ) | ( n781 & n2178 ) | ( ~n2175 & n2178 ) ;
  assign n2180 = n2175 | n2179 ;
  assign n2181 = n338 | n1376 ;
  assign n2182 = n1171 | n2181 ;
  assign n2183 = n479 | n544 ;
  assign n2184 = ( n168 & n933 ) | ( n168 & ~n2183 ) | ( n933 & ~n2183 ) ;
  assign n2185 = n2183 | n2184 ;
  assign n2186 = n2182 | n2185 ;
  assign n2187 = ( n360 & ~n566 ) | ( n360 & n1082 ) | ( ~n566 & n1082 ) ;
  assign n2188 = n566 | n2187 ;
  assign n2189 = ( ~n231 & n551 ) | ( ~n231 & n599 ) | ( n551 & n599 ) ;
  assign n2190 = n231 | n2189 ;
  assign n2191 = ( ~n2186 & n2188 ) | ( ~n2186 & n2190 ) | ( n2188 & n2190 ) ;
  assign n2192 = n2186 | n2191 ;
  assign n2193 = ( n2069 & ~n2180 ) | ( n2069 & n2192 ) | ( ~n2180 & n2192 ) ;
  assign n2194 = n2180 | n2193 ;
  assign n2195 = n777 | n977 ;
  assign n2196 = ( n367 & n655 ) | ( n367 & ~n1237 ) | ( n655 & ~n1237 ) ;
  assign n2197 = n1237 | n2196 ;
  assign n2198 = n536 | n691 ;
  assign n2199 = ( ~n2195 & n2197 ) | ( ~n2195 & n2198 ) | ( n2197 & n2198 ) ;
  assign n2200 = n2195 | n2199 ;
  assign n2201 = n211 | n1366 ;
  assign n2202 = ( n1346 & n1961 ) | ( n1346 & ~n2201 ) | ( n1961 & ~n2201 ) ;
  assign n2203 = n2201 | n2202 ;
  assign n2204 = n294 | n890 ;
  assign n2205 = ( n98 & n100 ) | ( n98 & n116 ) | ( n100 & n116 ) ;
  assign n2206 = n2204 | n2205 ;
  assign n2207 = n465 | n759 ;
  assign n2208 = n233 | n582 ;
  assign n2209 = n2207 | n2208 ;
  assign n2210 = ( ~n185 & n205 ) | ( ~n185 & n545 ) | ( n205 & n545 ) ;
  assign n2211 = n185 | n2210 ;
  assign n2212 = ( ~n2206 & n2209 ) | ( ~n2206 & n2211 ) | ( n2209 & n2211 ) ;
  assign n2213 = n2206 | n2212 ;
  assign n2214 = n259 | n661 ;
  assign n2215 = n591 | n992 ;
  assign n2216 = ( n1694 & ~n2214 ) | ( n1694 & n2215 ) | ( ~n2214 & n2215 ) ;
  assign n2217 = n2214 | n2216 ;
  assign n2218 = ( ~n2203 & n2213 ) | ( ~n2203 & n2217 ) | ( n2213 & n2217 ) ;
  assign n2219 = ( ~n2200 & n2203 ) | ( ~n2200 & n2218 ) | ( n2203 & n2218 ) ;
  assign n2220 = ( n66 & n102 ) | ( n66 & n216 ) | ( n102 & n216 ) ;
  assign n2221 = ( n41 & n44 ) | ( n41 & n122 ) | ( n44 & n122 ) ;
  assign n2222 = n2220 | n2221 ;
  assign n2223 = n2200 | n2222 ;
  assign n2224 = n449 | n1510 ;
  assign n2225 = n112 | n348 ;
  assign n2226 = ( n131 & n137 ) | ( n131 & ~n2225 ) | ( n137 & ~n2225 ) ;
  assign n2227 = n2225 | n2226 ;
  assign n2228 = ( ~n2222 & n2224 ) | ( ~n2222 & n2227 ) | ( n2224 & n2227 ) ;
  assign n2229 = ( ~n2219 & n2223 ) | ( ~n2219 & n2228 ) | ( n2223 & n2228 ) ;
  assign n2230 = n2219 | n2229 ;
  assign n2231 = n2194 | n2230 ;
  assign n2232 = n489 | n856 ;
  assign n2233 = n1758 | n2232 ;
  assign n2234 = ( n73 & n97 ) | ( n73 & n166 ) | ( n97 & n166 ) ;
  assign n2235 = n613 | n747 ;
  assign n2236 = n638 | n2235 ;
  assign n2237 = n1048 | n1059 ;
  assign n2238 = n123 | n2237 ;
  assign n2239 = n337 | n732 ;
  assign n2240 = ( n153 & n286 ) | ( n153 & ~n2239 ) | ( n286 & ~n2239 ) ;
  assign n2241 = n2239 | n2240 ;
  assign n2242 = ( ~n2236 & n2238 ) | ( ~n2236 & n2241 ) | ( n2238 & n2241 ) ;
  assign n2243 = n2236 | n2242 ;
  assign n2244 = ( ~n2233 & n2234 ) | ( ~n2233 & n2243 ) | ( n2234 & n2243 ) ;
  assign n2245 = n2233 | n2244 ;
  assign n2246 = n229 | n654 ;
  assign n2247 = n2033 | n2246 ;
  assign n2248 = n395 | n1870 ;
  assign n2249 = ( n266 & ~n395 ) | ( n266 & n630 ) | ( ~n395 & n630 ) ;
  assign n2250 = ( n55 & n696 ) | ( n55 & ~n956 ) | ( n696 & ~n956 ) ;
  assign n2251 = n956 | n2250 ;
  assign n2252 = ( ~n208 & n2249 ) | ( ~n208 & n2251 ) | ( n2249 & n2251 ) ;
  assign n2253 = ( n208 & ~n2248 ) | ( n208 & n2252 ) | ( ~n2248 & n2252 ) ;
  assign n2254 = ( ~n715 & n2248 ) | ( ~n715 & n2253 ) | ( n2248 & n2253 ) ;
  assign n2255 = n715 | n2254 ;
  assign n2256 = n662 | n666 ;
  assign n2257 = ( n383 & ~n1077 ) | ( n383 & n2256 ) | ( ~n1077 & n2256 ) ;
  assign n2258 = n1077 | n2257 ;
  assign n2259 = ( ~n2246 & n2255 ) | ( ~n2246 & n2258 ) | ( n2255 & n2258 ) ;
  assign n2260 = n217 | n299 ;
  assign n2261 = ( n44 & n145 ) | ( n44 & n152 ) | ( n145 & n152 ) ;
  assign n2262 = n316 | n2261 ;
  assign n2263 = n290 | n838 ;
  assign n2264 = n783 | n2263 ;
  assign n2265 = ( ~n2260 & n2262 ) | ( ~n2260 & n2264 ) | ( n2262 & n2264 ) ;
  assign n2266 = n2260 | n2265 ;
  assign n2267 = ( ~n2247 & n2259 ) | ( ~n2247 & n2266 ) | ( n2259 & n2266 ) ;
  assign n2268 = n2247 | n2267 ;
  assign n2269 = ( ~n2231 & n2245 ) | ( ~n2231 & n2268 ) | ( n2245 & n2268 ) ;
  assign n2270 = n2231 | n2269 ;
  assign n2271 = n446 | n1722 ;
  assign n2272 = n75 & n717 ;
  assign n2273 = ( n317 & ~n977 ) | ( n317 & n1477 ) | ( ~n977 & n1477 ) ;
  assign n2274 = n977 | n2273 ;
  assign n2275 = ( ~n2271 & n2272 ) | ( ~n2271 & n2274 ) | ( n2272 & n2274 ) ;
  assign n2276 = n2271 | n2275 ;
  assign n2277 = n204 | n921 ;
  assign n2278 = n193 | n1626 ;
  assign n2279 = n2277 | n2278 ;
  assign n2280 = n507 | n1556 ;
  assign n2281 = n753 | n2280 ;
  assign n2282 = n171 | n189 ;
  assign n2283 = ( n777 & n795 ) | ( n777 & ~n2282 ) | ( n795 & ~n2282 ) ;
  assign n2284 = n2282 | n2283 ;
  assign n2285 = n67 | n1001 ;
  assign n2286 = ( n254 & n2122 ) | ( n254 & ~n2285 ) | ( n2122 & ~n2285 ) ;
  assign n2287 = n2285 | n2286 ;
  assign n2288 = ( ~n2281 & n2284 ) | ( ~n2281 & n2287 ) | ( n2284 & n2287 ) ;
  assign n2289 = n2281 | n2288 ;
  assign n2290 = n45 | n483 ;
  assign n2291 = ( n1050 & n1912 ) | ( n1050 & ~n2290 ) | ( n1912 & ~n2290 ) ;
  assign n2292 = n2290 | n2291 ;
  assign n2293 = ( ~n2279 & n2289 ) | ( ~n2279 & n2292 ) | ( n2289 & n2292 ) ;
  assign n2294 = n2279 | n2293 ;
  assign n2295 = ( n1937 & ~n2276 ) | ( n1937 & n2294 ) | ( ~n2276 & n2294 ) ;
  assign n2296 = n2276 | n2295 ;
  assign n2297 = ( n673 & n2194 ) | ( n673 & n2296 ) | ( n2194 & n2296 ) ;
  assign n2298 = n673 & ~n2297 ;
  assign n2299 = n224 | n295 ;
  assign n2300 = n549 | n2299 ;
  assign n2301 = ( n48 & n66 ) | ( n48 & n160 ) | ( n66 & n160 ) ;
  assign n2302 = n312 | n2301 ;
  assign n2303 = n146 | n239 ;
  assign n2304 = ( ~n2300 & n2302 ) | ( ~n2300 & n2303 ) | ( n2302 & n2303 ) ;
  assign n2305 = n2300 | n2304 ;
  assign n2306 = n193 | n873 ;
  assign n2307 = n111 | n2306 ;
  assign n2308 = n211 | n972 ;
  assign n2309 = n177 | n2308 ;
  assign n2310 = n485 | n713 ;
  assign n2311 = ( n59 & n73 ) | ( n59 & n83 ) | ( n73 & n83 ) ;
  assign n2312 = n195 | n1225 ;
  assign n2313 = ( n2181 & ~n2311 ) | ( n2181 & n2312 ) | ( ~n2311 & n2312 ) ;
  assign n2314 = n2311 | n2313 ;
  assign n2315 = ( ~n2309 & n2310 ) | ( ~n2309 & n2314 ) | ( n2310 & n2314 ) ;
  assign n2316 = n2309 | n2315 ;
  assign n2317 = ( n66 & n84 ) | ( n66 & n109 ) | ( n84 & n109 ) ;
  assign n2318 = ( n142 & n150 ) | ( n142 & ~n2317 ) | ( n150 & ~n2317 ) ;
  assign n2319 = n2317 | n2318 ;
  assign n2320 = ( n2307 & ~n2316 ) | ( n2307 & n2319 ) | ( ~n2316 & n2319 ) ;
  assign n2321 = n492 | n545 ;
  assign n2322 = n2011 | n2321 ;
  assign n2323 = ( n44 & n84 ) | ( n44 & n1450 ) | ( n84 & n1450 ) ;
  assign n2324 = n995 | n1001 ;
  assign n2325 = n196 | n876 ;
  assign n2326 = n2324 | n2325 ;
  assign n2327 = n2323 | n2326 ;
  assign n2328 = n316 | n581 ;
  assign n2329 = ( ~n2322 & n2327 ) | ( ~n2322 & n2328 ) | ( n2327 & n2328 ) ;
  assign n2330 = n2322 | n2329 ;
  assign n2331 = ( n2316 & ~n2320 ) | ( n2316 & n2330 ) | ( ~n2320 & n2330 ) ;
  assign n2332 = ( ~n774 & n2320 ) | ( ~n774 & n2331 ) | ( n2320 & n2331 ) ;
  assign n2333 = ( n774 & ~n2305 ) | ( n774 & n2332 ) | ( ~n2305 & n2332 ) ;
  assign n2334 = n2305 | n2333 ;
  assign n2335 = n772 | n2334 ;
  assign n2336 = n686 | n991 ;
  assign n2337 = n61 | n396 ;
  assign n2338 = n1980 | n2008 ;
  assign n2339 = n268 | n540 ;
  assign n2340 = n115 | n2339 ;
  assign n2341 = n2338 | n2340 ;
  assign n2342 = ( ~n2336 & n2337 ) | ( ~n2336 & n2341 ) | ( n2337 & n2341 ) ;
  assign n2343 = n2336 | n2342 ;
  assign n2344 = ( n72 & n109 ) | ( n72 & n166 ) | ( n109 & n166 ) ;
  assign n2345 = n445 | n2344 ;
  assign n2346 = n331 | n917 ;
  assign n2347 = n1494 | n2346 ;
  assign n2348 = n691 | n1660 ;
  assign n2349 = n227 | n2348 ;
  assign n2350 = ( n2345 & ~n2347 ) | ( n2345 & n2349 ) | ( ~n2347 & n2349 ) ;
  assign n2351 = ( n1700 & n2347 ) | ( n1700 & ~n2350 ) | ( n2347 & ~n2350 ) ;
  assign n2352 = n2350 | n2351 ;
  assign n2353 = n171 | n851 ;
  assign n2354 = n1031 | n1436 ;
  assign n2355 = n2353 | n2354 ;
  assign n2356 = n435 | n444 ;
  assign n2357 = n1096 | n1346 ;
  assign n2358 = ( n1600 & ~n2356 ) | ( n1600 & n2357 ) | ( ~n2356 & n2357 ) ;
  assign n2359 = n2356 | n2358 ;
  assign n2360 = n913 | n2232 ;
  assign n2361 = n240 | n352 ;
  assign n2362 = n586 | n591 ;
  assign n2363 = n144 | n888 ;
  assign n2364 = ( ~n2361 & n2362 ) | ( ~n2361 & n2363 ) | ( n2362 & n2363 ) ;
  assign n2365 = n2361 | n2364 ;
  assign n2366 = n85 | n347 ;
  assign n2367 = n228 | n2366 ;
  assign n2368 = ( ~n2360 & n2365 ) | ( ~n2360 & n2367 ) | ( n2365 & n2367 ) ;
  assign n2369 = n2360 | n2368 ;
  assign n2370 = ( ~n2355 & n2359 ) | ( ~n2355 & n2369 ) | ( n2359 & n2369 ) ;
  assign n2371 = n2355 | n2370 ;
  assign n2372 = ( ~n2343 & n2352 ) | ( ~n2343 & n2371 ) | ( n2352 & n2371 ) ;
  assign n2373 = n2343 | n2372 ;
  assign n2374 = n74 | n104 ;
  assign n2375 = ( n507 & n947 ) | ( n507 & ~n2374 ) | ( n947 & ~n2374 ) ;
  assign n2376 = n2374 | n2375 ;
  assign n2377 = n587 | n807 ;
  assign n2378 = ( n626 & ~n2376 ) | ( n626 & n2377 ) | ( ~n2376 & n2377 ) ;
  assign n2379 = n2376 | n2378 ;
  assign n2380 = n101 | n1068 ;
  assign n2381 = ( n993 & ~n1163 ) | ( n993 & n2380 ) | ( ~n1163 & n2380 ) ;
  assign n2382 = ( ~n327 & n1163 ) | ( ~n327 & n2381 ) | ( n1163 & n2381 ) ;
  assign n2383 = ( n327 & n1969 ) | ( n327 & ~n2382 ) | ( n1969 & ~n2382 ) ;
  assign n2384 = n2382 | n2383 ;
  assign n2385 = n290 | n402 ;
  assign n2386 = n163 | n285 ;
  assign n2387 = ( n255 & n2385 ) | ( n255 & ~n2386 ) | ( n2385 & ~n2386 ) ;
  assign n2388 = n67 | n696 ;
  assign n2389 = ( n238 & n514 ) | ( n238 & ~n2388 ) | ( n514 & ~n2388 ) ;
  assign n2390 = n2388 | n2389 ;
  assign n2391 = ( n2386 & ~n2387 ) | ( n2386 & n2390 ) | ( ~n2387 & n2390 ) ;
  assign n2392 = n2387 | n2391 ;
  assign n2393 = ( ~n2379 & n2384 ) | ( ~n2379 & n2392 ) | ( n2384 & n2392 ) ;
  assign n2394 = n2379 | n2393 ;
  assign n2395 = ( ~n2335 & n2373 ) | ( ~n2335 & n2394 ) | ( n2373 & n2394 ) ;
  assign n2396 = n2335 | n2395 ;
  assign n2397 = n2033 | n2181 ;
  assign n2398 = n238 | n732 ;
  assign n2399 = n225 | n348 ;
  assign n2400 = ( n807 & ~n2398 ) | ( n807 & n2399 ) | ( ~n2398 & n2399 ) ;
  assign n2401 = n2398 | n2400 ;
  assign n2402 = n76 | n441 ;
  assign n2403 = n582 | n2402 ;
  assign n2404 = ( ~n2397 & n2401 ) | ( ~n2397 & n2403 ) | ( n2401 & n2403 ) ;
  assign n2405 = n2397 | n2404 ;
  assign n2406 = ( n48 & n50 ) | ( n48 & n66 ) | ( n50 & n66 ) ;
  assign n2407 = n1313 | n2406 ;
  assign n2408 = n1160 | n2407 ;
  assign n2409 = n592 | n1122 ;
  assign n2410 = n2408 | n2409 ;
  assign n2411 = ( n2197 & n2405 ) | ( n2197 & ~n2410 ) | ( n2405 & ~n2410 ) ;
  assign n2412 = n295 | n613 ;
  assign n2413 = n2214 | n2412 ;
  assign n2414 = n266 | n890 ;
  assign n2415 = ( n192 & n517 ) | ( n192 & ~n791 ) | ( n517 & ~n791 ) ;
  assign n2416 = n791 | n2415 ;
  assign n2417 = ( n317 & n528 ) | ( n317 & ~n865 ) | ( n528 & ~n865 ) ;
  assign n2418 = n865 | n2417 ;
  assign n2419 = ( n2284 & ~n2416 ) | ( n2284 & n2418 ) | ( ~n2416 & n2418 ) ;
  assign n2420 = n2416 | n2419 ;
  assign n2421 = ( ~n2413 & n2414 ) | ( ~n2413 & n2420 ) | ( n2414 & n2420 ) ;
  assign n2422 = n2413 | n2421 ;
  assign n2423 = ( n2410 & ~n2411 ) | ( n2410 & n2422 ) | ( ~n2411 & n2422 ) ;
  assign n2424 = n2411 | n2423 ;
  assign n2425 = ( n512 & n1595 ) | ( n512 & ~n2424 ) | ( n1595 & ~n2424 ) ;
  assign n2426 = n2424 | n2425 ;
  assign n2427 = n362 | n500 ;
  assign n2428 = n277 | n2427 ;
  assign n2429 = n176 | n489 ;
  assign n2430 = n193 | n2429 ;
  assign n2431 = n239 | n992 ;
  assign n2432 = n232 | n2431 ;
  assign n2433 = n147 | n941 ;
  assign n2434 = n981 | n1626 ;
  assign n2435 = ( n567 & ~n2433 ) | ( n567 & n2434 ) | ( ~n2433 & n2434 ) ;
  assign n2436 = n2433 | n2435 ;
  assign n2437 = ( n610 & ~n2432 ) | ( n610 & n2436 ) | ( ~n2432 & n2436 ) ;
  assign n2438 = n2432 | n2437 ;
  assign n2439 = n218 & ~n1225 ;
  assign n2440 = ( n164 & n261 ) | ( n164 & n2439 ) | ( n261 & n2439 ) ;
  assign n2441 = n2439 & ~n2440 ;
  assign n2442 = n267 | n1068 ;
  assign n2443 = n917 | n1526 ;
  assign n2444 = n45 | n1692 ;
  assign n2445 = ( ~n2442 & n2443 ) | ( ~n2442 & n2444 ) | ( n2443 & n2444 ) ;
  assign n2446 = n2442 | n2445 ;
  assign n2447 = ( n1945 & ~n2438 ) | ( n1945 & n2446 ) | ( ~n2438 & n2446 ) ;
  assign n2448 = ( n2438 & n2441 ) | ( n2438 & ~n2447 ) | ( n2441 & ~n2447 ) ;
  assign n2449 = ( n2430 & ~n2438 ) | ( n2430 & n2448 ) | ( ~n2438 & n2448 ) ;
  assign n2450 = ( n2428 & ~n2430 ) | ( n2428 & n2449 ) | ( ~n2430 & n2449 ) ;
  assign n2451 = ~n2428 & n2450 ;
  assign n2452 = n290 | n759 ;
  assign n2453 = ( n545 & n562 ) | ( n545 & ~n2452 ) | ( n562 & ~n2452 ) ;
  assign n2454 = n2452 | n2453 ;
  assign n2455 = n435 | n1031 ;
  assign n2456 = ( n255 & n273 ) | ( n255 & ~n2455 ) | ( n273 & ~n2455 ) ;
  assign n2457 = n2455 | n2456 ;
  assign n2458 = n203 | n540 ;
  assign n2459 = n873 | n2458 ;
  assign n2460 = ( ~n2454 & n2457 ) | ( ~n2454 & n2459 ) | ( n2457 & n2459 ) ;
  assign n2461 = n2454 | n2460 ;
  assign n2462 = ( n2426 & n2451 ) | ( n2426 & ~n2461 ) | ( n2451 & ~n2461 ) ;
  assign n2463 = n690 | n1646 ;
  assign n2464 = n137 | n952 ;
  assign n2465 = ( n653 & n1059 ) | ( n653 & ~n2464 ) | ( n1059 & ~n2464 ) ;
  assign n2466 = n2464 | n2465 ;
  assign n2467 = n115 | n534 ;
  assign n2468 = ( n1608 & n1929 ) | ( n1608 & ~n2467 ) | ( n1929 & ~n2467 ) ;
  assign n2469 = n2467 | n2468 ;
  assign n2470 = ( n48 & n72 ) | ( n48 & n216 ) | ( n72 & n216 ) ;
  assign n2471 = ( n55 & n523 ) | ( n55 & ~n2470 ) | ( n523 & ~n2470 ) ;
  assign n2472 = n2470 | n2471 ;
  assign n2473 = ( ~n2466 & n2469 ) | ( ~n2466 & n2472 ) | ( n2469 & n2472 ) ;
  assign n2474 = n2466 | n2473 ;
  assign n2475 = ( n300 & n482 ) | ( n300 & ~n1494 ) | ( n482 & ~n1494 ) ;
  assign n2476 = n1494 | n2475 ;
  assign n2477 = ( ~n2463 & n2474 ) | ( ~n2463 & n2476 ) | ( n2474 & n2476 ) ;
  assign n2478 = n2463 | n2477 ;
  assign n2479 = ( n124 & n433 ) | ( n124 & ~n1027 ) | ( n433 & ~n1027 ) ;
  assign n2480 = n1027 | n2479 ;
  assign n2481 = ( n123 & n360 ) | ( n123 & ~n698 ) | ( n360 & ~n698 ) ;
  assign n2482 = n698 | n2481 ;
  assign n2483 = n331 | n2482 ;
  assign n2484 = n132 | n329 ;
  assign n2485 = ( n253 & ~n885 ) | ( n253 & n2484 ) | ( ~n885 & n2484 ) ;
  assign n2486 = ( ~n331 & n885 ) | ( ~n331 & n2485 ) | ( n885 & n2485 ) ;
  assign n2487 = ( ~n2480 & n2483 ) | ( ~n2480 & n2486 ) | ( n2483 & n2486 ) ;
  assign n2488 = n2480 | n2487 ;
  assign n2489 = ( ~n2461 & n2478 ) | ( ~n2461 & n2488 ) | ( n2478 & n2488 ) ;
  assign n2490 = ( n2426 & n2462 ) | ( n2426 & ~n2489 ) | ( n2462 & ~n2489 ) ;
  assign n2491 = ~n2426 & n2490 ;
  assign n2492 = ( n97 & n98 ) | ( n97 & n119 ) | ( n98 & n119 ) ;
  assign n2493 = n642 | n2492 ;
  assign n2494 = n379 | n549 ;
  assign n2495 = n876 | n2494 ;
  assign n2496 = n328 | n985 ;
  assign n2497 = n445 | n1341 ;
  assign n2498 = n492 | n582 ;
  assign n2499 = ( ~n1173 & n2497 ) | ( ~n1173 & n2498 ) | ( n2497 & n2498 ) ;
  assign n2500 = ( n1173 & ~n2496 ) | ( n1173 & n2499 ) | ( ~n2496 & n2499 ) ;
  assign n2501 = n2496 | n2500 ;
  assign n2502 = ( n69 & ~n2495 ) | ( n69 & n2501 ) | ( ~n2495 & n2501 ) ;
  assign n2503 = ( ~n2493 & n2495 ) | ( ~n2493 & n2502 ) | ( n2495 & n2502 ) ;
  assign n2504 = ( n44 & n57 ) | ( n44 & n216 ) | ( n57 & n216 ) ;
  assign n2505 = ( n136 & n149 ) | ( n136 & n166 ) | ( n149 & n166 ) ;
  assign n2506 = n895 | n2505 ;
  assign n2507 = ( n488 & n1450 ) | ( n488 & ~n1689 ) | ( n1450 & ~n1689 ) ;
  assign n2508 = n1689 | n2507 ;
  assign n2509 = ( n2504 & ~n2506 ) | ( n2504 & n2508 ) | ( ~n2506 & n2508 ) ;
  assign n2510 = ( n2446 & n2506 ) | ( n2446 & ~n2509 ) | ( n2506 & ~n2509 ) ;
  assign n2511 = n2509 | n2510 ;
  assign n2512 = n2493 | n2511 ;
  assign n2513 = ( n337 & n921 ) | ( n337 & ~n2032 ) | ( n921 & ~n2032 ) ;
  assign n2514 = n2032 | n2513 ;
  assign n2515 = ( n233 & n1096 ) | ( n233 & ~n1237 ) | ( n1096 & ~n1237 ) ;
  assign n2516 = n1237 | n2515 ;
  assign n2517 = ( n612 & ~n2514 ) | ( n612 & n2516 ) | ( ~n2514 & n2516 ) ;
  assign n2518 = n2514 | n2517 ;
  assign n2519 = ( ~n2503 & n2512 ) | ( ~n2503 & n2518 ) | ( n2512 & n2518 ) ;
  assign n2520 = n2503 | n2519 ;
  assign n2521 = n517 | n1056 ;
  assign n2522 = n215 | n912 ;
  assign n2523 = n995 | n2522 ;
  assign n2524 = n2521 | n2523 ;
  assign n2525 = ( n163 & n873 ) | ( n163 & ~n1620 ) | ( n873 & ~n1620 ) ;
  assign n2526 = n1620 | n2525 ;
  assign n2527 = n1346 | n1376 ;
  assign n2528 = n217 | n609 ;
  assign n2529 = ( n942 & ~n2431 ) | ( n942 & n2528 ) | ( ~n2431 & n2528 ) ;
  assign n2530 = ( n2431 & ~n2527 ) | ( n2431 & n2529 ) | ( ~n2527 & n2529 ) ;
  assign n2531 = n2527 | n2530 ;
  assign n2532 = ( ~n2524 & n2526 ) | ( ~n2524 & n2531 ) | ( n2526 & n2531 ) ;
  assign n2533 = n2524 | n2532 ;
  assign n2534 = ( ~n805 & n2520 ) | ( ~n805 & n2533 ) | ( n2520 & n2533 ) ;
  assign n2535 = ( n75 & n80 ) | ( n75 & n116 ) | ( n80 & n116 ) ;
  assign n2536 = ( n666 & n928 ) | ( n666 & ~n2535 ) | ( n928 & ~n2535 ) ;
  assign n2537 = n2535 | n2536 ;
  assign n2538 = n1678 | n2167 ;
  assign n2539 = n51 | n81 ;
  assign n2540 = ( n259 & n613 ) | ( n259 & ~n2539 ) | ( n613 & ~n2539 ) ;
  assign n2541 = n2539 | n2540 ;
  assign n2542 = ( ~n2537 & n2538 ) | ( ~n2537 & n2541 ) | ( n2538 & n2541 ) ;
  assign n2543 = n2537 | n2542 ;
  assign n2544 = n285 | n444 ;
  assign n2545 = ( n151 & ~n1132 ) | ( n151 & n2544 ) | ( ~n1132 & n2544 ) ;
  assign n2546 = n1132 | n2545 ;
  assign n2547 = ( n312 & n466 ) | ( n312 & ~n2546 ) | ( n466 & ~n2546 ) ;
  assign n2548 = n2546 | n2547 ;
  assign n2549 = n1907 | n2548 ;
  assign n2550 = ( ~n2533 & n2543 ) | ( ~n2533 & n2549 ) | ( n2543 & n2549 ) ;
  assign n2551 = ( ~n805 & n2534 ) | ( ~n805 & n2550 ) | ( n2534 & n2550 ) ;
  assign n2552 = n805 | n2551 ;
  assign n2553 = n81 | n207 ;
  assign n2554 = n104 | n888 ;
  assign n2555 = ( n847 & ~n2553 ) | ( n847 & n2554 ) | ( ~n2553 & n2554 ) ;
  assign n2556 = n2553 | n2555 ;
  assign n2557 = n148 | n662 ;
  assign n2558 = n638 | n1237 ;
  assign n2559 = ( n64 & n145 ) | ( n64 & n152 ) | ( n145 & n152 ) ;
  assign n2560 = ( n536 & n865 ) | ( n536 & ~n2559 ) | ( n865 & ~n2559 ) ;
  assign n2561 = n2559 | n2560 ;
  assign n2562 = ( ~n2557 & n2558 ) | ( ~n2557 & n2561 ) | ( n2558 & n2561 ) ;
  assign n2563 = ( n1680 & n2557 ) | ( n1680 & ~n2562 ) | ( n2557 & ~n2562 ) ;
  assign n2564 = n2562 | n2563 ;
  assign n2565 = n2556 | n2564 ;
  assign n2566 = ( n57 & n64 ) | ( n57 & n149 ) | ( n64 & n149 ) ;
  assign n2567 = n91 | n2566 ;
  assign n2568 = ( n444 & n655 ) | ( n444 & ~n2567 ) | ( n655 & ~n2567 ) ;
  assign n2569 = n2567 | n2568 ;
  assign n2570 = ( n72 & n160 ) | ( n72 & n216 ) | ( n160 & n216 ) ;
  assign n2571 = n132 | n2570 ;
  assign n2572 = n79 | n587 ;
  assign n2573 = ( n187 & ~n2571 ) | ( n187 & n2572 ) | ( ~n2571 & n2572 ) ;
  assign n2574 = n2571 | n2573 ;
  assign n2575 = n567 | n775 ;
  assign n2576 = n873 | n1068 ;
  assign n2577 = n661 | n990 ;
  assign n2578 = ( n1770 & ~n2576 ) | ( n1770 & n2577 ) | ( ~n2576 & n2577 ) ;
  assign n2579 = n2576 | n2578 ;
  assign n2580 = ( ~n2574 & n2575 ) | ( ~n2574 & n2579 ) | ( n2575 & n2579 ) ;
  assign n2581 = n2574 | n2580 ;
  assign n2582 = ( ~n2565 & n2569 ) | ( ~n2565 & n2581 ) | ( n2569 & n2581 ) ;
  assign n2583 = n2565 | n2582 ;
  assign n2584 = ( n57 & n80 ) | ( n57 & n160 ) | ( n80 & n160 ) ;
  assign n2585 = n299 | n2584 ;
  assign n2586 = n2416 | n2585 ;
  assign n2587 = n1512 | n1543 ;
  assign n2588 = ( n866 & n2011 ) | ( n866 & ~n2587 ) | ( n2011 & ~n2587 ) ;
  assign n2589 = n2587 | n2588 ;
  assign n2590 = ( n50 & n64 ) | ( n50 & n109 ) | ( n64 & n109 ) ;
  assign n2591 = ( n85 & n1048 ) | ( n85 & ~n2590 ) | ( n1048 & ~n2590 ) ;
  assign n2592 = n2590 | n2591 ;
  assign n2593 = ( n379 & n959 ) | ( n379 & ~n2592 ) | ( n959 & ~n2592 ) ;
  assign n2594 = n2592 | n2593 ;
  assign n2595 = ( n2586 & n2589 ) | ( n2586 & ~n2594 ) | ( n2589 & ~n2594 ) ;
  assign n2596 = ( ~n161 & n204 ) | ( ~n161 & n434 ) | ( n204 & n434 ) ;
  assign n2597 = n161 | n2596 ;
  assign n2598 = n298 | n1940 ;
  assign n2599 = n435 | n2598 ;
  assign n2600 = ( ~n227 & n231 ) | ( ~n227 & n1700 ) | ( n231 & n1700 ) ;
  assign n2601 = ( n227 & ~n435 ) | ( n227 & n2600 ) | ( ~n435 & n2600 ) ;
  assign n2602 = ( ~n2597 & n2599 ) | ( ~n2597 & n2601 ) | ( n2599 & n2601 ) ;
  assign n2603 = n2597 | n2602 ;
  assign n2604 = ( n2594 & ~n2595 ) | ( n2594 & n2603 ) | ( ~n2595 & n2603 ) ;
  assign n2605 = n2595 | n2604 ;
  assign n2606 = n67 | n653 ;
  assign n2607 = n163 | n239 ;
  assign n2608 = n171 | n295 ;
  assign n2609 = ( ~n2606 & n2607 ) | ( ~n2606 & n2608 ) | ( n2607 & n2608 ) ;
  assign n2610 = n2606 | n2609 ;
  assign n2611 = n523 | n1082 ;
  assign n2612 = n719 | n746 ;
  assign n2613 = n2611 | n2612 ;
  assign n2614 = ( ~n54 & n129 ) | ( ~n54 & n136 ) | ( n129 & n136 ) ;
  assign n2615 = n347 | n995 ;
  assign n2616 = ( n1356 & ~n2614 ) | ( n1356 & n2615 ) | ( ~n2614 & n2615 ) ;
  assign n2617 = n2614 | n2616 ;
  assign n2618 = ( n80 & n100 ) | ( n80 & n145 ) | ( n100 & n145 ) ;
  assign n2619 = n396 | n2618 ;
  assign n2620 = n786 | n1044 ;
  assign n2621 = ( n123 & n215 ) | ( n123 & ~n2620 ) | ( n215 & ~n2620 ) ;
  assign n2622 = n2620 | n2621 ;
  assign n2623 = ( n2010 & ~n2619 ) | ( n2010 & n2622 ) | ( ~n2619 & n2622 ) ;
  assign n2624 = ( ~n2617 & n2619 ) | ( ~n2617 & n2623 ) | ( n2619 & n2623 ) ;
  assign n2625 = n2617 | n2624 ;
  assign n2626 = ( n904 & ~n2613 ) | ( n904 & n2625 ) | ( ~n2613 & n2625 ) ;
  assign n2627 = n2613 | n2626 ;
  assign n2628 = n455 | n1096 ;
  assign n2629 = ( ~n260 & n658 ) | ( ~n260 & n1793 ) | ( n658 & n1793 ) ;
  assign n2630 = ( n260 & ~n2628 ) | ( n260 & n2629 ) | ( ~n2628 & n2629 ) ;
  assign n2631 = n2628 | n2630 ;
  assign n2632 = ( ~n2610 & n2627 ) | ( ~n2610 & n2631 ) | ( n2627 & n2631 ) ;
  assign n2633 = n2610 | n2632 ;
  assign n2634 = ( ~n2583 & n2605 ) | ( ~n2583 & n2633 ) | ( n2605 & n2633 ) ;
  assign n2635 = n2583 | n2634 ;
  assign n2636 = n197 | n856 ;
  assign n2637 = n2321 | n2636 ;
  assign n2638 = n225 | n1116 ;
  assign n2639 = n195 | n448 ;
  assign n2640 = n203 | n712 ;
  assign n2641 = ( n48 & n57 ) | ( n48 & n166 ) | ( n57 & n166 ) ;
  assign n2642 = ( ~n2639 & n2640 ) | ( ~n2639 & n2641 ) | ( n2640 & n2641 ) ;
  assign n2643 = n2639 | n2642 ;
  assign n2644 = ( n2637 & n2638 ) | ( n2637 & ~n2643 ) | ( n2638 & ~n2643 ) ;
  assign n2645 = ( n103 & n1483 ) | ( n103 & ~n2052 ) | ( n1483 & ~n2052 ) ;
  assign n2646 = n2052 | n2645 ;
  assign n2647 = ( n44 & n50 ) | ( n44 & n59 ) | ( n50 & n59 ) ;
  assign n2648 = n435 | n2647 ;
  assign n2649 = n1948 | n2648 ;
  assign n2650 = ( n66 & n129 ) | ( n66 & n145 ) | ( n129 & n145 ) ;
  assign n2651 = ( n132 & n528 ) | ( n132 & ~n2650 ) | ( n528 & ~n2650 ) ;
  assign n2652 = n2650 | n2651 ;
  assign n2653 = ( n2523 & ~n2648 ) | ( n2523 & n2652 ) | ( ~n2648 & n2652 ) ;
  assign n2654 = n79 | n941 ;
  assign n2655 = n45 | n992 ;
  assign n2656 = ( n2067 & ~n2654 ) | ( n2067 & n2655 ) | ( ~n2654 & n2655 ) ;
  assign n2657 = n2654 | n2656 ;
  assign n2658 = ( ~n2649 & n2653 ) | ( ~n2649 & n2657 ) | ( n2653 & n2657 ) ;
  assign n2659 = n2649 | n2658 ;
  assign n2660 = ( ~n1444 & n2646 ) | ( ~n1444 & n2659 ) | ( n2646 & n2659 ) ;
  assign n2661 = n111 | n153 ;
  assign n2662 = ( n353 & n1526 ) | ( n353 & ~n2661 ) | ( n1526 & ~n2661 ) ;
  assign n2663 = n2661 | n2662 ;
  assign n2664 = n328 | n990 ;
  assign n2665 = n135 | n2664 ;
  assign n2666 = n85 | n262 ;
  assign n2667 = ( n218 & ~n1477 ) | ( n218 & n2666 ) | ( ~n1477 & n2666 ) ;
  assign n2668 = ~n2666 & n2667 ;
  assign n2669 = ( n2663 & ~n2665 ) | ( n2663 & n2668 ) | ( ~n2665 & n2668 ) ;
  assign n2670 = ~n2663 & n2669 ;
  assign n2671 = n517 | n1001 ;
  assign n2672 = ( n44 & n57 ) | ( n44 & n59 ) | ( n57 & n59 ) ;
  assign n2673 = ( n656 & ~n2671 ) | ( n656 & n2672 ) | ( ~n2671 & n2672 ) ;
  assign n2674 = n2671 | n2673 ;
  assign n2675 = ( n2646 & n2670 ) | ( n2646 & ~n2674 ) | ( n2670 & ~n2674 ) ;
  assign n2676 = ( n1444 & ~n2660 ) | ( n1444 & n2675 ) | ( ~n2660 & n2675 ) ;
  assign n2677 = ~n1444 & n2676 ;
  assign n2678 = ( ~n2643 & n2644 ) | ( ~n2643 & n2677 ) | ( n2644 & n2677 ) ;
  assign n2679 = ~n2644 & n2678 ;
  assign n2680 = n104 | n272 ;
  assign n2681 = n837 | n2680 ;
  assign n2682 = n540 | n1048 ;
  assign n2683 = n206 | n266 ;
  assign n2684 = n2682 | n2683 ;
  assign n2685 = ( n598 & ~n2680 ) | ( n598 & n2684 ) | ( ~n2680 & n2684 ) ;
  assign n2686 = n678 | n2685 ;
  assign n2687 = ( n171 & n544 ) | ( n171 & ~n2557 ) | ( n544 & ~n2557 ) ;
  assign n2688 = n2557 | n2687 ;
  assign n2689 = n301 | n1225 ;
  assign n2690 = ( n259 & n878 ) | ( n259 & ~n2689 ) | ( n878 & ~n2689 ) ;
  assign n2691 = n2689 | n2690 ;
  assign n2692 = ( n77 & n235 ) | ( n77 & ~n2691 ) | ( n235 & ~n2691 ) ;
  assign n2693 = n2691 | n2692 ;
  assign n2694 = ( n2482 & ~n2688 ) | ( n2482 & n2693 ) | ( ~n2688 & n2693 ) ;
  assign n2695 = n2688 | n2694 ;
  assign n2696 = ( ~n2681 & n2686 ) | ( ~n2681 & n2695 ) | ( n2686 & n2695 ) ;
  assign n2697 = n2681 | n2696 ;
  assign n2698 = n2679 & ~n2697 ;
  assign n2699 = n389 | n402 ;
  assign n2700 = ( n159 & n1892 ) | ( n159 & ~n2699 ) | ( n1892 & ~n2699 ) ;
  assign n2701 = n2699 | n2700 ;
  assign n2702 = n806 | n1254 ;
  assign n2703 = n848 | n2702 ;
  assign n2704 = n92 | n261 ;
  assign n2705 = n356 | n1059 ;
  assign n2706 = n838 | n1169 ;
  assign n2707 = ( ~n2704 & n2705 ) | ( ~n2704 & n2706 ) | ( n2705 & n2706 ) ;
  assign n2708 = n2704 | n2707 ;
  assign n2709 = n586 | n977 ;
  assign n2710 = n292 | n2709 ;
  assign n2711 = ( ~n2703 & n2708 ) | ( ~n2703 & n2710 ) | ( n2708 & n2710 ) ;
  assign n2712 = n2703 | n2711 ;
  assign n2713 = ( n80 & n102 ) | ( n80 & n160 ) | ( n102 & n160 ) ;
  assign n2714 = ( n212 & n493 ) | ( n212 & ~n2713 ) | ( n493 & ~n2713 ) ;
  assign n2715 = n2713 | n2714 ;
  assign n2716 = ( ~n2701 & n2712 ) | ( ~n2701 & n2715 ) | ( n2712 & n2715 ) ;
  assign n2717 = n2701 | n2716 ;
  assign n2718 = n755 | n888 ;
  assign n2719 = n302 | n529 ;
  assign n2720 = n193 | n500 ;
  assign n2721 = n298 | n2720 ;
  assign n2722 = ( ~n2718 & n2719 ) | ( ~n2718 & n2721 ) | ( n2719 & n2721 ) ;
  assign n2723 = n2718 | n2722 ;
  assign n2724 = ( n2698 & n2717 ) | ( n2698 & n2723 ) | ( n2717 & n2723 ) ;
  assign n2725 = n2698 & ~n2724 ;
  assign n2726 = n482 | n856 ;
  assign n2727 = n142 | n878 ;
  assign n2728 = n2726 | n2727 ;
  assign n2729 = n1547 | n2672 ;
  assign n2730 = n655 | n685 ;
  assign n2731 = n445 | n992 ;
  assign n2732 = n202 | n2731 ;
  assign n2733 = n224 | n348 ;
  assign n2734 = ( ~n2730 & n2732 ) | ( ~n2730 & n2733 ) | ( n2732 & n2733 ) ;
  assign n2735 = n2730 | n2734 ;
  assign n2736 = ( ~n2728 & n2729 ) | ( ~n2728 & n2735 ) | ( n2729 & n2735 ) ;
  assign n2737 = n2728 | n2736 ;
  assign n2738 = n193 | n266 ;
  assign n2739 = n288 | n1002 ;
  assign n2740 = ( n1023 & ~n2738 ) | ( n1023 & n2739 ) | ( ~n2738 & n2739 ) ;
  assign n2741 = n2738 | n2740 ;
  assign n2742 = n917 | n1313 ;
  assign n2743 = n931 | n1512 ;
  assign n2744 = n1079 | n2743 ;
  assign n2745 = n367 | n514 ;
  assign n2746 = ( n302 & n638 ) | ( n302 & ~n2745 ) | ( n638 & ~n2745 ) ;
  assign n2747 = n2745 | n2746 ;
  assign n2748 = ( n118 & n563 ) | ( n118 & ~n2747 ) | ( n563 & ~n2747 ) ;
  assign n2749 = n2747 | n2748 ;
  assign n2750 = ( ~n2741 & n2744 ) | ( ~n2741 & n2749 ) | ( n2744 & n2749 ) ;
  assign n2751 = n164 | n732 ;
  assign n2752 = ( ~n2742 & n2750 ) | ( ~n2742 & n2751 ) | ( n2750 & n2751 ) ;
  assign n2753 = n2742 | n2752 ;
  assign n2754 = ( ~n2737 & n2741 ) | ( ~n2737 & n2753 ) | ( n2741 & n2753 ) ;
  assign n2755 = n2737 | n2754 ;
  assign n2756 = ( n177 & n512 ) | ( n177 & ~n2755 ) | ( n512 & ~n2755 ) ;
  assign n2757 = n2755 | n2756 ;
  assign n2758 = n295 | n537 ;
  assign n2759 = n207 | n2758 ;
  assign n2760 = ( n238 & n267 ) | ( n238 & ~n1363 ) | ( n267 & ~n1363 ) ;
  assign n2761 = ( n130 & n1363 ) | ( n130 & ~n1608 ) | ( n1363 & ~n1608 ) ;
  assign n2762 = n1608 | n2761 ;
  assign n2763 = ( ~n2759 & n2760 ) | ( ~n2759 & n2762 ) | ( n2760 & n2762 ) ;
  assign n2764 = n2759 | n2763 ;
  assign n2765 = n519 | n1365 ;
  assign n2766 = n153 | n591 ;
  assign n2767 = n2765 | n2766 ;
  assign n2768 = ( n73 & n75 ) | ( n73 & n129 ) | ( n75 & n129 ) ;
  assign n2769 = n120 | n565 ;
  assign n2770 = ( n135 & ~n2768 ) | ( n135 & n2769 ) | ( ~n2768 & n2769 ) ;
  assign n2771 = n2768 | n2770 ;
  assign n2772 = ( ~n2098 & n2767 ) | ( ~n2098 & n2771 ) | ( n2767 & n2771 ) ;
  assign n2773 = ( n2098 & ~n2764 ) | ( n2098 & n2772 ) | ( ~n2764 & n2772 ) ;
  assign n2774 = ~n1006 & n1049 ;
  assign n2775 = ( ~n2764 & n2773 ) | ( ~n2764 & n2774 ) | ( n2773 & n2774 ) ;
  assign n2776 = ~n2773 & n2775 ;
  assign n2777 = n654 | n1144 ;
  assign n2778 = n1057 | n2777 ;
  assign n2779 = n137 | n696 ;
  assign n2780 = n205 | n361 ;
  assign n2781 = ( n2709 & ~n2779 ) | ( n2709 & n2780 ) | ( ~n2779 & n2780 ) ;
  assign n2782 = n2779 | n2781 ;
  assign n2783 = ( n1598 & ~n2778 ) | ( n1598 & n2782 ) | ( ~n2778 & n2782 ) ;
  assign n2784 = n2778 | n2783 ;
  assign n2785 = ( n2757 & n2776 ) | ( n2757 & ~n2784 ) | ( n2776 & ~n2784 ) ;
  assign n2786 = n192 | n490 ;
  assign n2787 = ( n44 & n75 ) | ( n44 & n80 ) | ( n75 & n80 ) ;
  assign n2788 = n2033 | n2705 ;
  assign n2789 = ( ~n490 & n2787 ) | ( ~n490 & n2788 ) | ( n2787 & n2788 ) ;
  assign n2790 = n146 | n228 ;
  assign n2791 = n641 | n1366 ;
  assign n2792 = n317 | n360 ;
  assign n2793 = ( ~n2790 & n2791 ) | ( ~n2790 & n2792 ) | ( n2791 & n2792 ) ;
  assign n2794 = n2790 | n2793 ;
  assign n2795 = ( ~n2786 & n2789 ) | ( ~n2786 & n2794 ) | ( n2789 & n2794 ) ;
  assign n2796 = n2786 | n2795 ;
  assign n2797 = n151 | n782 ;
  assign n2798 = n51 | n92 ;
  assign n2799 = n1660 | n2798 ;
  assign n2800 = n171 | n203 ;
  assign n2801 = ( n273 & n1526 ) | ( n273 & ~n1692 ) | ( n1526 & ~n1692 ) ;
  assign n2802 = n1692 | n2801 ;
  assign n2803 = n85 | n316 ;
  assign n2804 = ( ~n2800 & n2802 ) | ( ~n2800 & n2803 ) | ( n2802 & n2803 ) ;
  assign n2805 = n2800 | n2804 ;
  assign n2806 = ( ~n2797 & n2799 ) | ( ~n2797 & n2805 ) | ( n2799 & n2805 ) ;
  assign n2807 = n2797 | n2806 ;
  assign n2808 = ( ~n2784 & n2796 ) | ( ~n2784 & n2807 ) | ( n2796 & n2807 ) ;
  assign n2809 = ( n2757 & n2785 ) | ( n2757 & ~n2808 ) | ( n2785 & ~n2808 ) ;
  assign n2810 = ~n2757 & n2809 ;
  assign n2811 = n123 | n691 ;
  assign n2812 = n2399 | n2811 ;
  assign n2813 = ( n891 & ~n2362 ) | ( n891 & n2812 ) | ( ~n2362 & n2812 ) ;
  assign n2814 = ( n55 & n2362 ) | ( n55 & ~n2813 ) | ( n2362 & ~n2813 ) ;
  assign n2815 = n2813 | n2814 ;
  assign n2816 = n2276 | n2815 ;
  assign n2817 = ( n80 & n136 ) | ( n80 & n166 ) | ( n136 & n166 ) ;
  assign n2818 = n188 | n2817 ;
  assign n2819 = n112 | n153 ;
  assign n2820 = ( n85 & n299 ) | ( n85 & ~n2819 ) | ( n299 & ~n2819 ) ;
  assign n2821 = n2819 | n2820 ;
  assign n2822 = n367 | n489 ;
  assign n2823 = ( n895 & n2665 ) | ( n895 & ~n2822 ) | ( n2665 & ~n2822 ) ;
  assign n2824 = n2822 | n2823 ;
  assign n2825 = ( ~n2818 & n2821 ) | ( ~n2818 & n2824 ) | ( n2821 & n2824 ) ;
  assign n2826 = n2818 | n2825 ;
  assign n2827 = n148 | n1110 ;
  assign n2828 = n329 | n1277 ;
  assign n2829 = n2827 | n2828 ;
  assign n2830 = n286 | n482 ;
  assign n2831 = n331 | n985 ;
  assign n2832 = ( n653 & n1116 ) | ( n653 & ~n2831 ) | ( n1116 & ~n2831 ) ;
  assign n2833 = n2831 | n2832 ;
  assign n2834 = ( n912 & ~n2830 ) | ( n912 & n2833 ) | ( ~n2830 & n2833 ) ;
  assign n2835 = n2830 | n2834 ;
  assign n2836 = n260 | n1662 ;
  assign n2837 = ( ~n2829 & n2835 ) | ( ~n2829 & n2836 ) | ( n2835 & n2836 ) ;
  assign n2838 = ( n2528 & ~n2829 ) | ( n2528 & n2837 ) | ( ~n2829 & n2837 ) ;
  assign n2839 = n2829 | n2838 ;
  assign n2840 = ( ~n2816 & n2826 ) | ( ~n2816 & n2839 ) | ( n2826 & n2839 ) ;
  assign n2841 = n2816 | n2840 ;
  assign n2842 = ( n2116 & n2334 ) | ( n2116 & ~n2841 ) | ( n2334 & ~n2841 ) ;
  assign n2843 = n2841 | n2842 ;
  assign n2844 = ( n347 & n592 ) | ( n347 & ~n1024 ) | ( n592 & ~n1024 ) ;
  assign n2845 = n1024 | n2844 ;
  assign n2846 = n806 | n992 ;
  assign n2847 = n130 | n1314 ;
  assign n2848 = ( n1356 & n1860 ) | ( n1356 & ~n2847 ) | ( n1860 & ~n2847 ) ;
  assign n2849 = n2847 | n2848 ;
  assign n2850 = n318 | n956 ;
  assign n2851 = ( n41 & n84 ) | ( n41 & n145 ) | ( n84 & n145 ) ;
  assign n2852 = ( n148 & n549 ) | ( n148 & ~n2851 ) | ( n549 & ~n2851 ) ;
  assign n2853 = n2851 | n2852 ;
  assign n2854 = ( n661 & ~n2850 ) | ( n661 & n2853 ) | ( ~n2850 & n2853 ) ;
  assign n2855 = n2850 | n2854 ;
  assign n2856 = ( n2846 & ~n2849 ) | ( n2846 & n2855 ) | ( ~n2849 & n2855 ) ;
  assign n2857 = n163 | n562 ;
  assign n2858 = ( n2071 & ~n2849 ) | ( n2071 & n2857 ) | ( ~n2849 & n2857 ) ;
  assign n2859 = n2849 | n2858 ;
  assign n2860 = ( ~n2845 & n2856 ) | ( ~n2845 & n2859 ) | ( n2856 & n2859 ) ;
  assign n2861 = n2845 | n2860 ;
  assign n2862 = n485 | n885 ;
  assign n2863 = n300 | n465 ;
  assign n2864 = n675 | n985 ;
  assign n2865 = ( n64 & n75 ) | ( n64 & n149 ) | ( n75 & n149 ) ;
  assign n2866 = ( n783 & ~n2864 ) | ( n783 & n2865 ) | ( ~n2864 & n2865 ) ;
  assign n2867 = n2864 | n2866 ;
  assign n2868 = ( ~n2862 & n2863 ) | ( ~n2862 & n2867 ) | ( n2863 & n2867 ) ;
  assign n2869 = n2862 | n2868 ;
  assign n2870 = n648 | n1839 ;
  assign n2871 = n1340 | n2870 ;
  assign n2872 = n796 | n1940 ;
  assign n2873 = n922 | n2033 ;
  assign n2874 = n2872 | n2873 ;
  assign n2875 = ( n116 & n129 ) | ( n116 & n136 ) | ( n129 & n136 ) ;
  assign n2876 = ( n273 & ~n1340 ) | ( n273 & n2875 ) | ( ~n1340 & n2875 ) ;
  assign n2877 = ( ~n2871 & n2874 ) | ( ~n2871 & n2876 ) | ( n2874 & n2876 ) ;
  assign n2878 = n2871 | n2877 ;
  assign n2879 = ( ~n2861 & n2869 ) | ( ~n2861 & n2878 ) | ( n2869 & n2878 ) ;
  assign n2880 = n811 | n1396 ;
  assign n2881 = n67 | n331 ;
  assign n2882 = n185 | n2881 ;
  assign n2883 = n186 | n301 ;
  assign n2884 = ( n218 & ~n1600 ) | ( n218 & n2883 ) | ( ~n1600 & n2883 ) ;
  assign n2885 = ~n2883 & n2884 ;
  assign n2886 = ( n205 & n352 ) | ( n205 & ~n1611 ) | ( n352 & ~n1611 ) ;
  assign n2887 = n1611 | n2886 ;
  assign n2888 = n942 | n2620 ;
  assign n2889 = ( ~n791 & n2077 ) | ( ~n791 & n2888 ) | ( n2077 & n2888 ) ;
  assign n2890 = ( n791 & ~n1611 ) | ( n791 & n2889 ) | ( ~n1611 & n2889 ) ;
  assign n2891 = ( n2885 & n2887 ) | ( n2885 & n2890 ) | ( n2887 & n2890 ) ;
  assign n2892 = n2885 & ~n2891 ;
  assign n2893 = ( n1449 & ~n2882 ) | ( n1449 & n2892 ) | ( ~n2882 & n2892 ) ;
  assign n2894 = n111 | n440 ;
  assign n2895 = n746 | n2894 ;
  assign n2896 = n293 | n666 ;
  assign n2897 = n2163 | n2896 ;
  assign n2898 = n101 | n261 ;
  assign n2899 = n340 | n2126 ;
  assign n2900 = ( n59 & n64 ) | ( n59 & n102 ) | ( n64 & n102 ) ;
  assign n2901 = ( n1041 & ~n2899 ) | ( n1041 & n2900 ) | ( ~n2899 & n2900 ) ;
  assign n2902 = n2899 | n2901 ;
  assign n2903 = ( ~n2897 & n2898 ) | ( ~n2897 & n2902 ) | ( n2898 & n2902 ) ;
  assign n2904 = n2897 | n2903 ;
  assign n2905 = ( ~n2882 & n2895 ) | ( ~n2882 & n2904 ) | ( n2895 & n2904 ) ;
  assign n2906 = ( n1449 & n2893 ) | ( n1449 & ~n2905 ) | ( n2893 & ~n2905 ) ;
  assign n2907 = ~n1449 & n2906 ;
  assign n2908 = ( ~n2861 & n2880 ) | ( ~n2861 & n2907 ) | ( n2880 & n2907 ) ;
  assign n2909 = ( n2879 & ~n2880 ) | ( n2879 & n2908 ) | ( ~n2880 & n2908 ) ;
  assign n2910 = ~n2879 & n2909 ;
  assign n2911 = n295 | n587 ;
  assign n2912 = ( n445 & n1824 ) | ( n445 & ~n2911 ) | ( n1824 & ~n2911 ) ;
  assign n2913 = n2911 | n2912 ;
  assign n2914 = n207 | n1556 ;
  assign n2915 = n1460 | n1487 ;
  assign n2916 = ( n1588 & n2321 ) | ( n1588 & ~n2915 ) | ( n2321 & ~n2915 ) ;
  assign n2917 = n2915 | n2916 ;
  assign n2918 = n762 | n851 ;
  assign n2919 = n773 | n2654 ;
  assign n2920 = n2918 | n2919 ;
  assign n2921 = ( n2914 & n2917 ) | ( n2914 & ~n2920 ) | ( n2917 & ~n2920 ) ;
  assign n2922 = ( n2646 & n2920 ) | ( n2646 & ~n2921 ) | ( n2920 & ~n2921 ) ;
  assign n2923 = n2921 | n2922 ;
  assign n2924 = n265 | n507 ;
  assign n2925 = ( n167 & n947 ) | ( n167 & ~n2924 ) | ( n947 & ~n2924 ) ;
  assign n2926 = n2924 | n2925 ;
  assign n2927 = ( ~n2913 & n2923 ) | ( ~n2913 & n2926 ) | ( n2923 & n2926 ) ;
  assign n2928 = n2913 | n2927 ;
  assign n2929 = n489 | n885 ;
  assign n2930 = n124 | n775 ;
  assign n2931 = n2929 | n2930 ;
  assign n2932 = n1679 | n2818 ;
  assign n2933 = n839 | n878 ;
  assign n2934 = n45 | n262 ;
  assign n2935 = n117 | n2934 ;
  assign n2936 = ( ~n2932 & n2933 ) | ( ~n2932 & n2935 ) | ( n2933 & n2935 ) ;
  assign n2937 = n2932 | n2936 ;
  assign n2938 = n1928 | n2072 ;
  assign n2939 = ( ~n2931 & n2937 ) | ( ~n2931 & n2938 ) | ( n2937 & n2938 ) ;
  assign n2940 = n2931 | n2939 ;
  assign n2941 = n329 | n759 ;
  assign n2942 = ( n302 & n685 ) | ( n302 & ~n2941 ) | ( n685 & ~n2941 ) ;
  assign n2943 = n2941 | n2942 ;
  assign n2944 = n865 | n1450 ;
  assign n2945 = n395 | n734 ;
  assign n2946 = ( n224 & n361 ) | ( n224 & ~n2945 ) | ( n361 & ~n2945 ) ;
  assign n2947 = n2945 | n2946 ;
  assign n2948 = ( ~n2943 & n2944 ) | ( ~n2943 & n2947 ) | ( n2944 & n2947 ) ;
  assign n2949 = ( n172 & ~n2943 ) | ( n172 & n2948 ) | ( ~n2943 & n2948 ) ;
  assign n2950 = n2943 | n2949 ;
  assign n2951 = ( n218 & ~n383 ) | ( n218 & n1716 ) | ( ~n383 & n1716 ) ;
  assign n2952 = ~n1716 & n2951 ;
  assign n2953 = n312 | n1421 ;
  assign n2954 = ( n98 & n160 ) | ( n98 & n166 ) | ( n160 & n166 ) ;
  assign n2955 = ( n747 & ~n2953 ) | ( n747 & n2954 ) | ( ~n2953 & n2954 ) ;
  assign n2956 = n2953 | n2955 ;
  assign n2957 = ( n648 & n2768 ) | ( n648 & ~n2857 ) | ( n2768 & ~n2857 ) ;
  assign n2958 = n2857 | n2957 ;
  assign n2959 = ( ~n1350 & n2956 ) | ( ~n1350 & n2958 ) | ( n2956 & n2958 ) ;
  assign n2960 = ( n1350 & n2952 ) | ( n1350 & n2959 ) | ( n2952 & n2959 ) ;
  assign n2961 = n2952 & ~n2960 ;
  assign n2962 = ( n2940 & ~n2950 ) | ( n2940 & n2961 ) | ( ~n2950 & n2961 ) ;
  assign n2963 = ~n2940 & n2962 ;
  assign n2964 = ( ~n2605 & n2928 ) | ( ~n2605 & n2963 ) | ( n2928 & n2963 ) ;
  assign n2965 = ~n2928 & n2964 ;
  assign n2966 = n55 | n565 ;
  assign n2967 = n218 & ~n796 ;
  assign n2968 = ~n2966 & n2967 ;
  assign n2969 = n265 | n781 ;
  assign n2970 = ( n44 & n102 ) | ( n44 & n160 ) | ( n102 & n160 ) ;
  assign n2971 = n514 | n2970 ;
  assign n2972 = ( n961 & ~n2969 ) | ( n961 & n2971 ) | ( ~n2969 & n2971 ) ;
  assign n2973 = ( n1533 & n2969 ) | ( n1533 & ~n2972 ) | ( n2969 & ~n2972 ) ;
  assign n2974 = n2972 | n2973 ;
  assign n2975 = n360 | n777 ;
  assign n2976 = n2346 | n2975 ;
  assign n2977 = ( n2968 & n2974 ) | ( n2968 & n2976 ) | ( n2974 & n2976 ) ;
  assign n2978 = n2968 & ~n2977 ;
  assign n2979 = n1001 | n1421 ;
  assign n2980 = n2611 | n2664 ;
  assign n2981 = ( n44 & n66 ) | ( n44 & n92 ) | ( n66 & n92 ) ;
  assign n2982 = n186 | n337 ;
  assign n2983 = ( ~n2980 & n2981 ) | ( ~n2980 & n2982 ) | ( n2981 & n2982 ) ;
  assign n2984 = n2980 | n2983 ;
  assign n2985 = ( ~n1120 & n2355 ) | ( ~n1120 & n2984 ) | ( n2355 & n2984 ) ;
  assign n2986 = n1120 | n2985 ;
  assign n2987 = ( n445 & ~n2979 ) | ( n445 & n2986 ) | ( ~n2979 & n2986 ) ;
  assign n2988 = n2979 | n2987 ;
  assign n2989 = n349 | n384 ;
  assign n2990 = ( n866 & n1792 ) | ( n866 & ~n2989 ) | ( n1792 & ~n2989 ) ;
  assign n2991 = n2989 | n2990 ;
  assign n2992 = ( n2978 & n2988 ) | ( n2978 & n2991 ) | ( n2988 & n2991 ) ;
  assign n2993 = n2978 & ~n2992 ;
  assign n2994 = n1341 | n1692 ;
  assign n2995 = ( n66 & n80 ) | ( n66 & n109 ) | ( n80 & n109 ) ;
  assign n2996 = ( n301 & n697 ) | ( n301 & ~n2995 ) | ( n697 & ~n2995 ) ;
  assign n2997 = n2995 | n2996 ;
  assign n2998 = n1096 | n1110 ;
  assign n2999 = ( ~n2994 & n2997 ) | ( ~n2994 & n2998 ) | ( n2997 & n2998 ) ;
  assign n3000 = n2994 | n2999 ;
  assign n3001 = n1737 | n2093 ;
  assign n3002 = n1472 | n1487 ;
  assign n3003 = n85 | n361 ;
  assign n3004 = n891 | n2214 ;
  assign n3005 = n3003 | n3004 ;
  assign n3006 = ( ~n3001 & n3002 ) | ( ~n3001 & n3005 ) | ( n3002 & n3005 ) ;
  assign n3007 = ( n320 & n1507 ) | ( n320 & ~n3001 ) | ( n1507 & ~n3001 ) ;
  assign n3008 = n3001 | n3007 ;
  assign n3009 = n3006 | n3008 ;
  assign n3010 = ( n195 & n675 ) | ( n195 & ~n981 ) | ( n675 & ~n981 ) ;
  assign n3011 = n981 | n3010 ;
  assign n3012 = ( n2622 & ~n3008 ) | ( n2622 & n3011 ) | ( ~n3008 & n3011 ) ;
  assign n3013 = ( ~n3000 & n3009 ) | ( ~n3000 & n3012 ) | ( n3009 & n3012 ) ;
  assign n3014 = n3000 | n3013 ;
  assign n3015 = n165 | n2215 ;
  assign n3016 = ( n1377 & n1974 ) | ( n1377 & ~n3015 ) | ( n1974 & ~n3015 ) ;
  assign n3017 = n3015 | n3016 ;
  assign n3018 = n254 | n367 ;
  assign n3019 = ( n490 & n566 ) | ( n490 & ~n3018 ) | ( n566 & ~n3018 ) ;
  assign n3020 = n3018 | n3019 ;
  assign n3021 = ( n72 & n84 ) | ( n72 & n149 ) | ( n84 & n149 ) ;
  assign n3022 = n775 | n3021 ;
  assign n3023 = ( n347 & n686 ) | ( n347 & ~n3022 ) | ( n686 & ~n3022 ) ;
  assign n3024 = n3022 | n3023 ;
  assign n3025 = ( ~n3017 & n3020 ) | ( ~n3017 & n3024 ) | ( n3020 & n3024 ) ;
  assign n3026 = n130 | n174 ;
  assign n3027 = ( n2047 & ~n3025 ) | ( n2047 & n3026 ) | ( ~n3025 & n3026 ) ;
  assign n3028 = n3025 | n3027 ;
  assign n3029 = n3017 | n3028 ;
  assign n3030 = n203 | n662 ;
  assign n3031 = n1547 | n3030 ;
  assign n3032 = n255 | n655 ;
  assign n3033 = n112 | n838 ;
  assign n3034 = ( n66 & n73 ) | ( n66 & n84 ) | ( n73 & n84 ) ;
  assign n3035 = n197 | n3034 ;
  assign n3036 = ( ~n3032 & n3033 ) | ( ~n3032 & n3035 ) | ( n3033 & n3035 ) ;
  assign n3037 = n3032 | n3036 ;
  assign n3038 = ( n149 & n152 ) | ( n149 & n534 ) | ( n152 & n534 ) ;
  assign n3039 = ( ~n3031 & n3037 ) | ( ~n3031 & n3038 ) | ( n3037 & n3038 ) ;
  assign n3040 = n3031 | n3039 ;
  assign n3041 = n105 | n353 ;
  assign n3042 = n746 | n3041 ;
  assign n3043 = ( ~n3029 & n3040 ) | ( ~n3029 & n3042 ) | ( n3040 & n3042 ) ;
  assign n3044 = n3029 | n3043 ;
  assign n3045 = ( n2993 & n3014 ) | ( n2993 & n3044 ) | ( n3014 & n3044 ) ;
  assign n3046 = n2993 & ~n3045 ;
  assign n3047 = n164 | n1720 ;
  assign n3048 = ( n658 & n981 ) | ( n658 & ~n3047 ) | ( n981 & ~n3047 ) ;
  assign n3049 = n3047 | n3048 ;
  assign n3050 = n1134 | n2835 ;
  assign n3051 = n888 | n960 ;
  assign n3052 = n2431 | n3051 ;
  assign n3053 = n337 | n590 ;
  assign n3054 = ( n2327 & ~n3052 ) | ( n2327 & n3053 ) | ( ~n3052 & n3053 ) ;
  assign n3055 = n3052 | n3054 ;
  assign n3056 = ( ~n3049 & n3050 ) | ( ~n3049 & n3055 ) | ( n3050 & n3055 ) ;
  assign n3057 = n3049 | n3056 ;
  assign n3058 = n384 | n577 ;
  assign n3059 = n228 | n3058 ;
  assign n3060 = n1793 | n2362 ;
  assign n3061 = n272 | n928 ;
  assign n3062 = n352 | n796 ;
  assign n3063 = n177 | n3062 ;
  assign n3064 = ( n1593 & ~n3061 ) | ( n1593 & n3063 ) | ( ~n3061 & n3063 ) ;
  assign n3065 = n3061 | n3064 ;
  assign n3066 = ( n2654 & ~n3060 ) | ( n2654 & n3065 ) | ( ~n3060 & n3065 ) ;
  assign n3067 = n3060 | n3066 ;
  assign n3068 = n1856 | n1995 ;
  assign n3069 = ( n74 & n959 ) | ( n74 & ~n2821 ) | ( n959 & ~n2821 ) ;
  assign n3070 = n2821 | n3069 ;
  assign n3071 = ( n504 & n551 ) | ( n504 & ~n2256 ) | ( n551 & ~n2256 ) ;
  assign n3072 = n2256 | n3071 ;
  assign n3073 = ( ~n3068 & n3070 ) | ( ~n3068 & n3072 ) | ( n3070 & n3072 ) ;
  assign n3074 = ( ~n3067 & n3068 ) | ( ~n3067 & n3073 ) | ( n3068 & n3073 ) ;
  assign n3075 = ( ~n3059 & n3067 ) | ( ~n3059 & n3074 ) | ( n3067 & n3074 ) ;
  assign n3076 = n3059 | n3075 ;
  assign n3077 = ( n2426 & ~n3057 ) | ( n2426 & n3076 ) | ( ~n3057 & n3076 ) ;
  assign n3078 = n3057 | n3077 ;
  assign n3079 = n123 | n630 ;
  assign n3080 = ( n72 & n84 ) | ( n72 & n216 ) | ( n84 & n216 ) ;
  assign n3081 = n466 | n3080 ;
  assign n3082 = n3079 | n3081 ;
  assign n3083 = n567 | n762 ;
  assign n3084 = n1826 | n3083 ;
  assign n3085 = ( n1425 & ~n3082 ) | ( n1425 & n3084 ) | ( ~n3082 & n3084 ) ;
  assign n3086 = n3082 | n3085 ;
  assign n3087 = ( n448 & n689 ) | ( n448 & ~n3086 ) | ( n689 & ~n3086 ) ;
  assign n3088 = n3086 | n3087 ;
  assign n3089 = n1488 | n1887 ;
  assign n3090 = n720 | n2966 ;
  assign n3091 = ( n98 & n149 ) | ( n98 & n1116 ) | ( n149 & n1116 ) ;
  assign n3092 = ( n164 & n273 ) | ( n164 & ~n3091 ) | ( n273 & ~n3091 ) ;
  assign n3093 = n3091 | n3092 ;
  assign n3094 = ( n3089 & ~n3090 ) | ( n3089 & n3093 ) | ( ~n3090 & n3093 ) ;
  assign n3095 = ( n2200 & n3090 ) | ( n2200 & ~n3094 ) | ( n3090 & ~n3094 ) ;
  assign n3096 = n3094 | n3095 ;
  assign n3097 = ( n44 & n57 ) | ( n44 & n66 ) | ( n57 & n66 ) ;
  assign n3098 = n238 | n1366 ;
  assign n3099 = ( n1658 & ~n1998 ) | ( n1658 & n3098 ) | ( ~n1998 & n3098 ) ;
  assign n3100 = n1998 | n3099 ;
  assign n3101 = ( n2882 & ~n3097 ) | ( n2882 & n3100 ) | ( ~n3097 & n3100 ) ;
  assign n3102 = ( n1059 & n3097 ) | ( n1059 & ~n3101 ) | ( n3097 & ~n3101 ) ;
  assign n3103 = n3101 | n3102 ;
  assign n3104 = n189 | n233 ;
  assign n3105 = n362 | n3104 ;
  assign n3106 = ( n2702 & ~n3103 ) | ( n2702 & n3105 ) | ( ~n3103 & n3105 ) ;
  assign n3107 = n3103 | n3106 ;
  assign n3108 = n133 | n1613 ;
  assign n3109 = n174 | n586 ;
  assign n3110 = ( n2929 & ~n3108 ) | ( n2929 & n3109 ) | ( ~n3108 & n3109 ) ;
  assign n3111 = ( n41 & n80 ) | ( n41 & n119 ) | ( n80 & n119 ) ;
  assign n3112 = ( n338 & n540 ) | ( n338 & ~n3111 ) | ( n540 & ~n3111 ) ;
  assign n3113 = n3111 | n3112 ;
  assign n3114 = ( n153 & n205 ) | ( n153 & ~n928 ) | ( n205 & ~n928 ) ;
  assign n3115 = n928 | n3114 ;
  assign n3116 = ( ~n1963 & n3113 ) | ( ~n1963 & n3115 ) | ( n3113 & n3115 ) ;
  assign n3117 = n3110 | n3116 ;
  assign n3118 = n3108 | n3117 ;
  assign n3119 = n241 | n599 ;
  assign n3120 = ( n202 & n1027 ) | ( n202 & ~n3119 ) | ( n1027 & ~n3119 ) ;
  assign n3121 = n3119 | n3120 ;
  assign n3122 = ( n1963 & ~n3118 ) | ( n1963 & n3121 ) | ( ~n3118 & n3121 ) ;
  assign n3123 = n3118 | n3122 ;
  assign n3124 = ( ~n3096 & n3107 ) | ( ~n3096 & n3123 ) | ( n3107 & n3123 ) ;
  assign n3125 = n3096 | n3124 ;
  assign n3126 = n3088 | n3125 ;
  assign n3127 = ( ~n78 & n149 ) | ( ~n78 & n1313 ) | ( n149 & n1313 ) ;
  assign n3128 = n329 | n851 ;
  assign n3129 = ( n76 & n516 ) | ( n76 & ~n3128 ) | ( n516 & ~n3128 ) ;
  assign n3130 = n3128 | n3129 ;
  assign n3131 = n115 | n713 ;
  assign n3132 = ( n150 & ~n783 ) | ( n150 & n3131 ) | ( ~n783 & n3131 ) ;
  assign n3133 = ( ~n76 & n783 ) | ( ~n76 & n3132 ) | ( n783 & n3132 ) ;
  assign n3134 = ( ~n3127 & n3130 ) | ( ~n3127 & n3133 ) | ( n3130 & n3133 ) ;
  assign n3135 = n3127 | n3134 ;
  assign n3136 = n517 | n2726 ;
  assign n3137 = n316 | n3136 ;
  assign n3138 = ( n120 & n1277 ) | ( n120 & ~n3137 ) | ( n1277 & ~n3137 ) ;
  assign n3139 = n3137 | n3138 ;
  assign n3140 = n1652 | n1732 ;
  assign n3141 = ( n70 & n71 ) | ( n70 & n302 ) | ( n71 & n302 ) ;
  assign n3142 = ( n57 & n149 ) | ( n57 & n3141 ) | ( n149 & n3141 ) ;
  assign n3143 = ( n203 & ~n256 ) | ( n203 & n657 ) | ( ~n256 & n657 ) ;
  assign n3144 = n256 | n3143 ;
  assign n3145 = ( n3140 & ~n3142 ) | ( n3140 & n3144 ) | ( ~n3142 & n3144 ) ;
  assign n3146 = ( n1838 & n3142 ) | ( n1838 & ~n3145 ) | ( n3142 & ~n3145 ) ;
  assign n3147 = n3145 | n3146 ;
  assign n3148 = ( n2359 & ~n3139 ) | ( n2359 & n3147 ) | ( ~n3139 & n3147 ) ;
  assign n3149 = n3139 | n3148 ;
  assign n3150 = ( n426 & ~n3135 ) | ( n426 & n3149 ) | ( ~n3135 & n3149 ) ;
  assign n3151 = n3135 | n3150 ;
  assign n3152 = ( n1141 & ~n3126 ) | ( n1141 & n3151 ) | ( ~n3126 & n3151 ) ;
  assign n3153 = n3126 | n3152 ;
  assign n3154 = n447 | n941 ;
  assign n3155 = n208 | n563 ;
  assign n3156 = ( n1928 & ~n3154 ) | ( n1928 & n3155 ) | ( ~n3154 & n3155 ) ;
  assign n3157 = n3154 | n3156 ;
  assign n3158 = n528 | n895 ;
  assign n3159 = n493 | n519 ;
  assign n3160 = ( n1672 & ~n3158 ) | ( n1672 & n3159 ) | ( ~n3158 & n3159 ) ;
  assign n3161 = n3158 | n3160 ;
  assign n3162 = n445 | n455 ;
  assign n3163 = n686 | n2100 ;
  assign n3164 = ( n2672 & ~n3162 ) | ( n2672 & n3163 ) | ( ~n3162 & n3163 ) ;
  assign n3165 = n3162 | n3164 ;
  assign n3166 = ( ~n3157 & n3161 ) | ( ~n3157 & n3165 ) | ( n3161 & n3165 ) ;
  assign n3167 = n3157 | n3166 ;
  assign n3168 = n45 | n888 ;
  assign n3169 = n2607 | n3168 ;
  assign n3170 = n81 | n320 ;
  assign n3171 = ( n489 & n595 ) | ( n489 & ~n3170 ) | ( n595 & ~n3170 ) ;
  assign n3172 = n3170 | n3171 ;
  assign n3173 = n74 | n1032 ;
  assign n3174 = n1526 | n3173 ;
  assign n3175 = ( n293 & n1430 ) | ( n293 & ~n1526 ) | ( n1430 & ~n1526 ) ;
  assign n3176 = ( ~n3172 & n3174 ) | ( ~n3172 & n3175 ) | ( n3174 & n3175 ) ;
  assign n3177 = n3172 | n3176 ;
  assign n3178 = n235 | n1690 ;
  assign n3179 = ( ~n3169 & n3177 ) | ( ~n3169 & n3178 ) | ( n3177 & n3178 ) ;
  assign n3180 = n3169 | n3179 ;
  assign n3181 = n810 | n887 ;
  assign n3182 = n150 | n291 ;
  assign n3183 = n79 | n1001 ;
  assign n3184 = n960 | n3183 ;
  assign n3185 = n261 | n329 ;
  assign n3186 = ( ~n3182 & n3184 ) | ( ~n3182 & n3185 ) | ( n3184 & n3185 ) ;
  assign n3187 = n3182 | n3186 ;
  assign n3188 = ( n977 & ~n3181 ) | ( n977 & n3187 ) | ( ~n3181 & n3187 ) ;
  assign n3189 = n3181 | n3188 ;
  assign n3190 = ( ~n3167 & n3180 ) | ( ~n3167 & n3189 ) | ( n3180 & n3189 ) ;
  assign n3191 = n3167 | n3190 ;
  assign n3192 = ( n48 & ~n54 ) | ( n48 & n75 ) | ( ~n54 & n75 ) ;
  assign n3193 = ( n274 & n1450 ) | ( n274 & ~n3192 ) | ( n1450 & ~n3192 ) ;
  assign n3194 = n3192 | n3193 ;
  assign n3195 = ( n482 & ~n746 ) | ( n482 & n1377 ) | ( ~n746 & n1377 ) ;
  assign n3196 = n746 | n3195 ;
  assign n3197 = n85 | n638 ;
  assign n3198 = ( n1692 & n3196 ) | ( n1692 & ~n3197 ) | ( n3196 & ~n3197 ) ;
  assign n3199 = n931 | n1533 ;
  assign n3200 = ( ~n785 & n2105 ) | ( ~n785 & n3199 ) | ( n2105 & n3199 ) ;
  assign n3201 = ( n3197 & ~n3198 ) | ( n3197 & n3200 ) | ( ~n3198 & n3200 ) ;
  assign n3202 = n3198 | n3201 ;
  assign n3203 = ( n581 & ~n2188 ) | ( n581 & n2528 ) | ( ~n2188 & n2528 ) ;
  assign n3204 = n2188 | n3203 ;
  assign n3205 = ( n785 & n1978 ) | ( n785 & ~n3063 ) | ( n1978 & ~n3063 ) ;
  assign n3206 = n3063 | n3205 ;
  assign n3207 = ( n1125 & ~n3204 ) | ( n1125 & n3206 ) | ( ~n3204 & n3206 ) ;
  assign n3208 = ( ~n3202 & n3204 ) | ( ~n3202 & n3207 ) | ( n3204 & n3207 ) ;
  assign n3209 = ( ~n3194 & n3202 ) | ( ~n3194 & n3208 ) | ( n3202 & n3208 ) ;
  assign n3210 = n3194 | n3209 ;
  assign n3211 = ( n254 & n655 ) | ( n254 & ~n1110 ) | ( n655 & ~n1110 ) ;
  assign n3212 = n1110 | n3211 ;
  assign n3213 = ( n80 & n98 ) | ( n80 & n145 ) | ( n98 & n145 ) ;
  assign n3214 = n465 | n3213 ;
  assign n3215 = n241 | n328 ;
  assign n3216 = ( n173 & n839 ) | ( n173 & ~n3215 ) | ( n839 & ~n3215 ) ;
  assign n3217 = n3215 | n3216 ;
  assign n3218 = ( ~n3212 & n3214 ) | ( ~n3212 & n3217 ) | ( n3214 & n3217 ) ;
  assign n3219 = n3212 | n3218 ;
  assign n3220 = n170 | n338 ;
  assign n3221 = n231 | n661 ;
  assign n3222 = ( n83 & n109 ) | ( n83 & n145 ) | ( n109 & n145 ) ;
  assign n3223 = ( n1068 & ~n3221 ) | ( n1068 & n3222 ) | ( ~n3221 & n3222 ) ;
  assign n3224 = n3221 | n3223 ;
  assign n3225 = ( n2682 & ~n3220 ) | ( n2682 & n3224 ) | ( ~n3220 & n3224 ) ;
  assign n3226 = n3220 | n3225 ;
  assign n3227 = n1915 | n2033 ;
  assign n3228 = n516 | n625 ;
  assign n3229 = n185 | n786 ;
  assign n3230 = ( ~n657 & n876 ) | ( ~n657 & n1523 ) | ( n876 & n1523 ) ;
  assign n3231 = n657 | n3230 ;
  assign n3232 = ( n1365 & ~n3229 ) | ( n1365 & n3231 ) | ( ~n3229 & n3231 ) ;
  assign n3233 = n3229 | n3232 ;
  assign n3234 = ( ~n3227 & n3228 ) | ( ~n3227 & n3233 ) | ( n3228 & n3233 ) ;
  assign n3235 = n3227 | n3234 ;
  assign n3236 = ( ~n3219 & n3226 ) | ( ~n3219 & n3235 ) | ( n3226 & n3235 ) ;
  assign n3237 = n3219 | n3236 ;
  assign n3238 = ( ~n3191 & n3210 ) | ( ~n3191 & n3237 ) | ( n3210 & n3237 ) ;
  assign n3239 = n3191 | n3238 ;
  assign n3240 = n2928 | n3040 ;
  assign n3241 = n193 | n1346 ;
  assign n3242 = n891 | n3241 ;
  assign n3243 = ( n2237 & ~n2443 ) | ( n2237 & n3242 ) | ( ~n2443 & n3242 ) ;
  assign n3244 = ( ~n1741 & n2443 ) | ( ~n1741 & n3243 ) | ( n2443 & n3243 ) ;
  assign n3245 = n433 | n482 ;
  assign n3246 = ( n101 & n839 ) | ( n101 & ~n3245 ) | ( n839 & ~n3245 ) ;
  assign n3247 = n3245 | n3246 ;
  assign n3248 = n1172 | n1254 ;
  assign n3249 = n224 | n529 ;
  assign n3250 = ( n188 & n238 ) | ( n188 & ~n3249 ) | ( n238 & ~n3249 ) ;
  assign n3251 = n3249 | n3250 ;
  assign n3252 = ( ~n3247 & n3248 ) | ( ~n3247 & n3251 ) | ( n3248 & n3251 ) ;
  assign n3253 = n3247 | n3252 ;
  assign n3254 = ( n1741 & ~n3244 ) | ( n1741 & n3253 ) | ( ~n3244 & n3253 ) ;
  assign n3255 = n3244 | n3254 ;
  assign n3256 = n1144 | n2672 ;
  assign n3257 = n943 | n3256 ;
  assign n3258 = n567 | n928 ;
  assign n3259 = ( n971 & ~n3257 ) | ( n971 & n3258 ) | ( ~n3257 & n3258 ) ;
  assign n3260 = n3257 | n3259 ;
  assign n3261 = ( n441 & ~n447 ) | ( n441 & n550 ) | ( ~n447 & n550 ) ;
  assign n3262 = n447 | n3261 ;
  assign n3263 = ( ~n1047 & n1435 ) | ( ~n1047 & n1870 ) | ( n1435 & n1870 ) ;
  assign n3264 = n1047 | n3263 ;
  assign n3265 = n186 | n886 ;
  assign n3266 = ( n356 & n933 ) | ( n356 & ~n3265 ) | ( n933 & ~n3265 ) ;
  assign n3267 = n3265 | n3266 ;
  assign n3268 = ( ~n3262 & n3264 ) | ( ~n3262 & n3267 ) | ( n3264 & n3267 ) ;
  assign n3269 = n3262 | n3268 ;
  assign n3270 = ( ~n3255 & n3260 ) | ( ~n3255 & n3269 ) | ( n3260 & n3269 ) ;
  assign n3271 = ( ~n3240 & n3255 ) | ( ~n3240 & n3270 ) | ( n3255 & n3270 ) ;
  assign n3272 = n667 & ~n2324 ;
  assign n3273 = n137 | n329 ;
  assign n3274 = ( ~n52 & n512 ) | ( ~n52 & n952 ) | ( n512 & n952 ) ;
  assign n3275 = n52 | n3274 ;
  assign n3276 = ( n3272 & n3273 ) | ( n3272 & n3275 ) | ( n3273 & n3275 ) ;
  assign n3277 = n3272 & ~n3276 ;
  assign n3278 = n258 | n824 ;
  assign n3279 = ( n734 & n1297 ) | ( n734 & ~n3278 ) | ( n1297 & ~n3278 ) ;
  assign n3280 = n3278 | n3279 ;
  assign n3281 = n144 | n959 ;
  assign n3282 = ( n2188 & ~n3280 ) | ( n2188 & n3281 ) | ( ~n3280 & n3281 ) ;
  assign n3283 = n3280 | n3282 ;
  assign n3284 = n206 | n960 ;
  assign n3285 = ( n41 & n80 ) | ( n41 & n100 ) | ( n80 & n100 ) ;
  assign n3286 = n3284 | n3285 ;
  assign n3287 = n104 | n1376 ;
  assign n3288 = n293 | n641 ;
  assign n3289 = n489 | n1450 ;
  assign n3290 = ( ~n3287 & n3288 ) | ( ~n3287 & n3289 ) | ( n3288 & n3289 ) ;
  assign n3291 = n3287 | n3290 ;
  assign n3292 = ( n91 & n440 ) | ( n91 & ~n2362 ) | ( n440 & ~n2362 ) ;
  assign n3293 = n2362 | n3292 ;
  assign n3294 = ( ~n3286 & n3291 ) | ( ~n3286 & n3293 ) | ( n3291 & n3293 ) ;
  assign n3295 = n3286 | n3294 ;
  assign n3296 = ( n3277 & n3283 ) | ( n3277 & n3295 ) | ( n3283 & n3295 ) ;
  assign n3297 = n3277 & ~n3296 ;
  assign n3298 = ~n2521 & n3297 ;
  assign n3299 = ( ~n3240 & n3271 ) | ( ~n3240 & n3298 ) | ( n3271 & n3298 ) ;
  assign n3300 = ~n3271 & n3299 ;
  assign n3301 = ( n148 & n388 ) | ( n148 & ~n1699 ) | ( n388 & ~n1699 ) ;
  assign n3302 = n1699 | n3301 ;
  assign n3303 = ( n98 & n145 ) | ( n98 & n166 ) | ( n145 & n166 ) ;
  assign n3304 = n889 | n3303 ;
  assign n3305 = n3098 | n3304 ;
  assign n3306 = n142 | n921 ;
  assign n3307 = n261 | n956 ;
  assign n3308 = ( n100 & n102 ) | ( n100 & n145 ) | ( n102 & n145 ) ;
  assign n3309 = n172 | n3308 ;
  assign n3310 = ( n207 & ~n3307 ) | ( n207 & n3309 ) | ( ~n3307 & n3309 ) ;
  assign n3311 = n3307 | n3310 ;
  assign n3312 = ( ~n3305 & n3306 ) | ( ~n3305 & n3311 ) | ( n3306 & n3311 ) ;
  assign n3313 = n3305 | n3312 ;
  assign n3314 = n503 | n3313 ;
  assign n3315 = n272 | n320 ;
  assign n3316 = n167 | n3315 ;
  assign n3317 = n228 | n876 ;
  assign n3318 = ( n3080 & ~n3316 ) | ( n3080 & n3317 ) | ( ~n3316 & n3317 ) ;
  assign n3319 = n3316 | n3318 ;
  assign n3320 = ( n1726 & ~n3313 ) | ( n1726 & n3319 ) | ( ~n3313 & n3319 ) ;
  assign n3321 = ( ~n3302 & n3314 ) | ( ~n3302 & n3320 ) | ( n3314 & n3320 ) ;
  assign n3322 = n3302 | n3321 ;
  assign n3323 = n3297 & ~n3322 ;
  assign n3324 = n2846 | n2864 ;
  assign n3325 = n1145 | n1732 ;
  assign n3326 = n67 | n352 ;
  assign n3327 = ( n544 & n638 ) | ( n544 & ~n3326 ) | ( n638 & ~n3326 ) ;
  assign n3328 = n3326 | n3327 ;
  assign n3329 = n1078 | n2033 ;
  assign n3330 = ( n59 & ~n78 ) | ( n59 & n100 ) | ( ~n78 & n100 ) ;
  assign n3331 = ( n132 & n505 ) | ( n132 & ~n3330 ) | ( n505 & ~n3330 ) ;
  assign n3332 = n3330 | n3331 ;
  assign n3333 = ( n113 & n446 ) | ( n113 & ~n3332 ) | ( n446 & ~n3332 ) ;
  assign n3334 = n3332 | n3333 ;
  assign n3335 = ( ~n3328 & n3329 ) | ( ~n3328 & n3334 ) | ( n3329 & n3334 ) ;
  assign n3336 = n3328 | n3335 ;
  assign n3337 = ( ~n3324 & n3325 ) | ( ~n3324 & n3336 ) | ( n3325 & n3336 ) ;
  assign n3338 = n3324 | n3337 ;
  assign n3339 = ( n119 & n122 ) | ( n119 & n129 ) | ( n122 & n129 ) ;
  assign n3340 = n1625 | n3339 ;
  assign n3341 = ( n92 & n796 ) | ( n92 & ~n1430 ) | ( n796 & ~n1430 ) ;
  assign n3342 = n1430 | n3341 ;
  assign n3343 = ( ~n468 & n684 ) | ( ~n468 & n1363 ) | ( n684 & n1363 ) ;
  assign n3344 = n468 | n3343 ;
  assign n3345 = ( n41 & n64 ) | ( n41 & n119 ) | ( n64 & n119 ) ;
  assign n3346 = ( n448 & n912 ) | ( n448 & ~n3345 ) | ( n912 & ~n3345 ) ;
  assign n3347 = n3345 | n3346 ;
  assign n3348 = ( ~n3342 & n3344 ) | ( ~n3342 & n3347 ) | ( n3344 & n3347 ) ;
  assign n3349 = n3342 | n3348 ;
  assign n3350 = ( ~n2040 & n3340 ) | ( ~n2040 & n3349 ) | ( n3340 & n3349 ) ;
  assign n3351 = n192 | n947 ;
  assign n3352 = ( n2040 & ~n3350 ) | ( n2040 & n3351 ) | ( ~n3350 & n3351 ) ;
  assign n3353 = n3350 | n3352 ;
  assign n3354 = ( n3323 & n3338 ) | ( n3323 & n3353 ) | ( n3338 & n3353 ) ;
  assign n3355 = n3323 & ~n3354 ;
  assign n3356 = ( n44 & n84 ) | ( n44 & n129 ) | ( n84 & n129 ) ;
  assign n3357 = n577 | n3356 ;
  assign n3358 = n295 | n528 ;
  assign n3359 = n685 | n3358 ;
  assign n3360 = ( n3281 & ~n3356 ) | ( n3281 & n3359 ) | ( ~n3356 & n3359 ) ;
  assign n3361 = n85 | n394 ;
  assign n3362 = n202 | n824 ;
  assign n3363 = ( n692 & ~n3361 ) | ( n692 & n3362 ) | ( ~n3361 & n3362 ) ;
  assign n3364 = n3361 | n3363 ;
  assign n3365 = ( ~n3357 & n3360 ) | ( ~n3357 & n3364 ) | ( n3360 & n3364 ) ;
  assign n3366 = n3357 | n3365 ;
  assign n3367 = ( n393 & n440 ) | ( n393 & ~n592 ) | ( n440 & ~n592 ) ;
  assign n3368 = n592 | n3367 ;
  assign n3369 = n353 | n1044 ;
  assign n3370 = n82 | n3369 ;
  assign n3371 = n115 | n3370 ;
  assign n3372 = ( n72 & ~n78 ) | ( n72 & n122 ) | ( ~n78 & n122 ) ;
  assign n3373 = ( ~n3368 & n3371 ) | ( ~n3368 & n3372 ) | ( n3371 & n3372 ) ;
  assign n3374 = n3368 | n3373 ;
  assign n3375 = n117 | n233 ;
  assign n3376 = ( n783 & n1059 ) | ( n783 & ~n3375 ) | ( n1059 & ~n3375 ) ;
  assign n3377 = n3375 | n3376 ;
  assign n3378 = n104 | n1313 ;
  assign n3379 = n2126 | n3378 ;
  assign n3380 = ( n362 & n535 ) | ( n362 & ~n2126 ) | ( n535 & ~n2126 ) ;
  assign n3381 = ( ~n3377 & n3379 ) | ( ~n3377 & n3380 ) | ( n3379 & n3380 ) ;
  assign n3382 = ( ~n3374 & n3377 ) | ( ~n3374 & n3381 ) | ( n3377 & n3381 ) ;
  assign n3383 = n3374 | n3382 ;
  assign n3384 = n2431 | n2497 ;
  assign n3385 = n891 | n3384 ;
  assign n3386 = ( ~n3366 & n3383 ) | ( ~n3366 & n3385 ) | ( n3383 & n3385 ) ;
  assign n3387 = n3366 | n3386 ;
  assign n3388 = ( n673 & ~n1989 ) | ( n673 & n3387 ) | ( ~n1989 & n3387 ) ;
  assign n3389 = ~n3387 & n3388 ;
  assign n3390 = n74 | n732 ;
  assign n3391 = n587 | n691 ;
  assign n3392 = ( n66 & n152 ) | ( n66 & n216 ) | ( n152 & n216 ) ;
  assign n3393 = ( n565 & n995 ) | ( n565 & ~n3392 ) | ( n995 & ~n3392 ) ;
  assign n3394 = n3392 | n3393 ;
  assign n3395 = ( n3390 & ~n3391 ) | ( n3390 & n3394 ) | ( ~n3391 & n3394 ) ;
  assign n3396 = ( n961 & n3391 ) | ( n961 & ~n3395 ) | ( n3391 & ~n3395 ) ;
  assign n3397 = n3395 | n3396 ;
  assign n3398 = n2759 | n3397 ;
  assign n3399 = ( n83 & n129 ) | ( n83 & n160 ) | ( n129 & n160 ) ;
  assign n3400 = ( n262 & n265 ) | ( n262 & ~n3399 ) | ( n265 & ~n3399 ) ;
  assign n3401 = n3399 | n3400 ;
  assign n3402 = ( n103 & n796 ) | ( n103 & ~n1346 ) | ( n796 & ~n1346 ) ;
  assign n3403 = n1346 | n3402 ;
  assign n3404 = n101 | n1027 ;
  assign n3405 = n2576 | n3404 ;
  assign n3406 = n186 | n242 ;
  assign n3407 = n377 | n1235 ;
  assign n3408 = ( n1435 & n1887 ) | ( n1435 & ~n3407 ) | ( n1887 & ~n3407 ) ;
  assign n3409 = n3407 | n3408 ;
  assign n3410 = ( ~n3405 & n3406 ) | ( ~n3405 & n3409 ) | ( n3406 & n3409 ) ;
  assign n3411 = n3405 | n3410 ;
  assign n3412 = ( ~n3401 & n3403 ) | ( ~n3401 & n3411 ) | ( n3403 & n3411 ) ;
  assign n3413 = ( n3398 & n3401 ) | ( n3398 & ~n3412 ) | ( n3401 & ~n3412 ) ;
  assign n3414 = ( n161 & n592 ) | ( n161 & ~n1626 ) | ( n592 & ~n1626 ) ;
  assign n3415 = n1626 | n3414 ;
  assign n3416 = n1116 | n2896 ;
  assign n3417 = n131 | n352 ;
  assign n3418 = n689 | n760 ;
  assign n3419 = ( n3416 & ~n3417 ) | ( n3416 & n3418 ) | ( ~n3417 & n3418 ) ;
  assign n3420 = n337 | n886 ;
  assign n3421 = ( n3417 & ~n3419 ) | ( n3417 & n3420 ) | ( ~n3419 & n3420 ) ;
  assign n3422 = n3419 | n3421 ;
  assign n3423 = n563 | n2163 ;
  assign n3424 = n3168 | n3423 ;
  assign n3425 = ( ~n3415 & n3422 ) | ( ~n3415 & n3424 ) | ( n3422 & n3424 ) ;
  assign n3426 = n3415 | n3425 ;
  assign n3427 = ( n3412 & ~n3413 ) | ( n3412 & n3426 ) | ( ~n3413 & n3426 ) ;
  assign n3428 = n3413 | n3427 ;
  assign n3429 = n383 | n449 ;
  assign n3430 = ( n241 & n810 ) | ( n241 & ~n2498 ) | ( n810 & ~n2498 ) ;
  assign n3431 = n2498 | n3430 ;
  assign n3432 = n59 | n84 ;
  assign n3433 = ( n98 & n116 ) | ( n98 & n3432 ) | ( n116 & n3432 ) ;
  assign n3434 = ( n172 & n416 ) | ( n172 & ~n3433 ) | ( n416 & ~n3433 ) ;
  assign n3435 = n3433 | n3434 ;
  assign n3436 = ( n64 & n102 ) | ( n64 & n216 ) | ( n102 & n216 ) ;
  assign n3437 = ( n528 & n1001 ) | ( n528 & ~n3436 ) | ( n1001 & ~n3436 ) ;
  assign n3438 = n3436 | n3437 ;
  assign n3439 = ( ~n3431 & n3435 ) | ( ~n3431 & n3438 ) | ( n3435 & n3438 ) ;
  assign n3440 = n3431 | n3439 ;
  assign n3441 = ( n2544 & ~n3429 ) | ( n2544 & n3440 ) | ( ~n3429 & n3440 ) ;
  assign n3442 = n3429 | n3441 ;
  assign n3443 = ( n151 & n317 ) | ( n151 & ~n1005 ) | ( n317 & ~n1005 ) ;
  assign n3444 = n1005 | n3443 ;
  assign n3445 = n76 | n124 ;
  assign n3446 = ( n41 & n50 ) | ( n41 & n109 ) | ( n50 & n109 ) ;
  assign n3447 = ( n775 & ~n3445 ) | ( n775 & n3446 ) | ( ~n3445 & n3446 ) ;
  assign n3448 = n3445 | n3447 ;
  assign n3449 = ( n1493 & n2522 ) | ( n1493 & ~n3448 ) | ( n2522 & ~n3448 ) ;
  assign n3450 = n3448 | n3449 ;
  assign n3451 = ( n3442 & n3444 ) | ( n3442 & ~n3450 ) | ( n3444 & ~n3450 ) ;
  assign n3452 = n865 | n2598 ;
  assign n3453 = ( n117 & n294 ) | ( n117 & ~n3303 ) | ( n294 & ~n3303 ) ;
  assign n3454 = n3303 | n3453 ;
  assign n3455 = n1174 | n1976 ;
  assign n3456 = ( n2067 & n2680 ) | ( n2067 & ~n3455 ) | ( n2680 & ~n3455 ) ;
  assign n3457 = n3455 | n3456 ;
  assign n3458 = ( ~n3452 & n3454 ) | ( ~n3452 & n3457 ) | ( n3454 & n3457 ) ;
  assign n3459 = n3452 | n3458 ;
  assign n3460 = ( n59 & n66 ) | ( n59 & n80 ) | ( n66 & n80 ) ;
  assign n3461 = ( ~n2474 & n2727 ) | ( ~n2474 & n3460 ) | ( n2727 & n3460 ) ;
  assign n3462 = n2474 | n3461 ;
  assign n3463 = ( n167 & n291 ) | ( n167 & ~n731 ) | ( n291 & ~n731 ) ;
  assign n3464 = n731 | n3463 ;
  assign n3465 = ( ~n3459 & n3462 ) | ( ~n3459 & n3464 ) | ( n3462 & n3464 ) ;
  assign n3466 = n3459 | n3465 ;
  assign n3467 = ( n3450 & ~n3451 ) | ( n3450 & n3466 ) | ( ~n3451 & n3466 ) ;
  assign n3468 = n3451 | n3467 ;
  assign n3469 = ( n188 & n440 ) | ( n188 & ~n1879 ) | ( n440 & ~n1879 ) ;
  assign n3470 = n1879 | n3469 ;
  assign n3471 = ( n66 & ~n78 ) | ( n66 & n116 ) | ( ~n78 & n116 ) ;
  assign n3472 = n713 | n3471 ;
  assign n3473 = n657 | n824 ;
  assign n3474 = n123 | n3162 ;
  assign n3475 = n3473 | n3474 ;
  assign n3476 = ( ~n3470 & n3472 ) | ( ~n3470 & n3475 ) | ( n3472 & n3475 ) ;
  assign n3477 = n3470 | n3476 ;
  assign n3478 = ( ~n3428 & n3468 ) | ( ~n3428 & n3477 ) | ( n3468 & n3477 ) ;
  assign n3479 = n3428 | n3478 ;
  assign n3480 = ( n64 & n119 ) | ( n64 & n136 ) | ( n119 & n136 ) ;
  assign n3481 = n103 | n3480 ;
  assign n3482 = n349 | n1235 ;
  assign n3483 = n3481 | n3482 ;
  assign n3484 = n85 | n1556 ;
  assign n3485 = n131 | n3484 ;
  assign n3486 = ( n2441 & n3483 ) | ( n2441 & ~n3485 ) | ( n3483 & ~n3485 ) ;
  assign n3487 = ~n3483 & n3486 ;
  assign n3488 = n75 | n122 ;
  assign n3489 = ( n44 & n83 ) | ( n44 & n3488 ) | ( n83 & n3488 ) ;
  assign n3490 = ( n419 & n2262 ) | ( n419 & ~n3489 ) | ( n2262 & ~n3489 ) ;
  assign n3491 = n3489 | n3490 ;
  assign n3492 = n3226 | n3491 ;
  assign n3493 = n383 | n1172 ;
  assign n3494 = ( n159 & n1594 ) | ( n159 & ~n3493 ) | ( n1594 & ~n3493 ) ;
  assign n3495 = n3493 | n3494 ;
  assign n3496 = ( n3487 & n3492 ) | ( n3487 & n3495 ) | ( n3492 & n3495 ) ;
  assign n3497 = n3487 & ~n3496 ;
  assign n3498 = ( n102 & n136 ) | ( n102 & n145 ) | ( n136 & n145 ) ;
  assign n3499 = n394 | n3498 ;
  assign n3500 = n359 | n3204 ;
  assign n3501 = n193 | n512 ;
  assign n3502 = ( ~n208 & n648 ) | ( ~n208 & n1658 ) | ( n648 & n1658 ) ;
  assign n3503 = ( n208 & ~n3501 ) | ( n208 & n3502 ) | ( ~n3501 & n3502 ) ;
  assign n3504 = n3501 | n3503 ;
  assign n3505 = n60 | n312 ;
  assign n3506 = ( n795 & n2791 ) | ( n795 & ~n3505 ) | ( n2791 & ~n3505 ) ;
  assign n3507 = n3505 | n3506 ;
  assign n3508 = ( ~n3500 & n3504 ) | ( ~n3500 & n3507 ) | ( n3504 & n3507 ) ;
  assign n3509 = n3500 | n3508 ;
  assign n3510 = n3499 | n3509 ;
  assign n3511 = n295 | n1220 ;
  assign n3512 = n242 | n485 ;
  assign n3513 = ( n302 & n666 ) | ( n302 & ~n3512 ) | ( n666 & ~n3512 ) ;
  assign n3514 = n3512 | n3513 ;
  assign n3515 = ( n505 & ~n3511 ) | ( n505 & n3514 ) | ( ~n3511 & n3514 ) ;
  assign n3516 = n3511 | n3515 ;
  assign n3517 = n101 | n549 ;
  assign n3518 = ( n488 & n536 ) | ( n488 & ~n3517 ) | ( n536 & ~n3517 ) ;
  assign n3519 = n3517 | n3518 ;
  assign n3520 = n266 | n519 ;
  assign n3521 = n889 | n3520 ;
  assign n3522 = n254 | n977 ;
  assign n3523 = n74 | n921 ;
  assign n3524 = ( ~n3521 & n3522 ) | ( ~n3521 & n3523 ) | ( n3522 & n3523 ) ;
  assign n3525 = n3521 | n3524 ;
  assign n3526 = ( n482 & n1237 ) | ( n482 & ~n2607 ) | ( n1237 & ~n2607 ) ;
  assign n3527 = n2607 | n3526 ;
  assign n3528 = ( ~n3519 & n3525 ) | ( ~n3519 & n3527 ) | ( n3525 & n3527 ) ;
  assign n3529 = n3519 | n3528 ;
  assign n3530 = ( ~n3510 & n3516 ) | ( ~n3510 & n3529 ) | ( n3516 & n3529 ) ;
  assign n3531 = n3510 | n3530 ;
  assign n3532 = ( n3466 & n3497 ) | ( n3466 & n3531 ) | ( n3497 & n3531 ) ;
  assign n3533 = n3497 & ~n3532 ;
  assign n3534 = ~n3479 & n3533 ;
  assign n3535 = n301 | n420 ;
  assign n3536 = n273 | n952 ;
  assign n3537 = ( n1780 & ~n3535 ) | ( n1780 & n3536 ) | ( ~n3535 & n3536 ) ;
  assign n3538 = n3535 | n3537 ;
  assign n3539 = n807 | n2929 ;
  assign n3540 = n130 | n1589 ;
  assign n3541 = ( n1380 & n1782 ) | ( n1380 & ~n1915 ) | ( n1782 & ~n1915 ) ;
  assign n3542 = n1915 | n3541 ;
  assign n3543 = ( n177 & ~n1024 ) | ( n177 & n1116 ) | ( ~n1024 & n1116 ) ;
  assign n3544 = n1024 | n3543 ;
  assign n3545 = ( ~n3540 & n3542 ) | ( ~n3540 & n3544 ) | ( n3542 & n3544 ) ;
  assign n3546 = n3540 | n3545 ;
  assign n3547 = ( n850 & ~n3539 ) | ( n850 & n3546 ) | ( ~n3539 & n3546 ) ;
  assign n3548 = n3539 | n3547 ;
  assign n3549 = ( n581 & n1169 ) | ( n581 & ~n1237 ) | ( n1169 & ~n1237 ) ;
  assign n3550 = n1237 | n3549 ;
  assign n3551 = n51 | n290 ;
  assign n3552 = n685 | n696 ;
  assign n3553 = ( ~n3550 & n3551 ) | ( ~n3550 & n3552 ) | ( n3551 & n3552 ) ;
  assign n3554 = n3550 | n3553 ;
  assign n3555 = ( ~n3538 & n3548 ) | ( ~n3538 & n3554 ) | ( n3548 & n3554 ) ;
  assign n3556 = n3538 | n3555 ;
  assign n3557 = n368 | n1660 ;
  assign n3558 = ( n434 & n1314 ) | ( n434 & ~n3557 ) | ( n1314 & ~n3557 ) ;
  assign n3559 = n3557 | n3558 ;
  assign n3560 = n146 | n591 ;
  assign n3561 = ( n195 & n734 ) | ( n195 & ~n3560 ) | ( n734 & ~n3560 ) ;
  assign n3562 = n3560 | n3561 ;
  assign n3563 = n105 | n170 ;
  assign n3564 = n285 | n3563 ;
  assign n3565 = ( n3559 & ~n3562 ) | ( n3559 & n3564 ) | ( ~n3562 & n3564 ) ;
  assign n3566 = n256 | n2727 ;
  assign n3567 = n1929 | n2636 ;
  assign n3568 = n218 & ~n956 ;
  assign n3569 = n300 | n493 ;
  assign n3570 = n3568 & ~n3569 ;
  assign n3571 = ( n66 & n116 ) | ( n66 & n136 ) | ( n116 & n136 ) ;
  assign n3572 = n3570 & ~n3571 ;
  assign n3573 = ( n3566 & ~n3567 ) | ( n3566 & n3572 ) | ( ~n3567 & n3572 ) ;
  assign n3574 = ~n3566 & n3573 ;
  assign n3575 = ( ~n3562 & n3565 ) | ( ~n3562 & n3574 ) | ( n3565 & n3574 ) ;
  assign n3576 = ( n1017 & ~n3565 ) | ( n1017 & n3575 ) | ( ~n3565 & n3575 ) ;
  assign n3577 = ~n1017 & n3576 ;
  assign n3578 = n2941 | n2981 ;
  assign n3579 = n675 | n796 ;
  assign n3580 = ( n1712 & n2105 ) | ( n1712 & ~n3579 ) | ( n2105 & ~n3579 ) ;
  assign n3581 = n3579 | n3580 ;
  assign n3582 = n791 | n2576 ;
  assign n3583 = ( ~n3578 & n3581 ) | ( ~n3578 & n3582 ) | ( n3581 & n3582 ) ;
  assign n3584 = n3578 | n3583 ;
  assign n3585 = ( n3556 & n3577 ) | ( n3556 & ~n3584 ) | ( n3577 & ~n3584 ) ;
  assign n3586 = ~n3556 & n3585 ;
  assign n3587 = ( n3479 & ~n3534 ) | ( n3479 & n3586 ) | ( ~n3534 & n3586 ) ;
  assign n3588 = ( ~n3389 & n3533 ) | ( ~n3389 & n3587 ) | ( n3533 & n3587 ) ;
  assign n3589 = ( n3389 & ~n3479 ) | ( n3389 & n3588 ) | ( ~n3479 & n3588 ) ;
  assign n3590 = ( n3355 & n3389 ) | ( n3355 & n3589 ) | ( n3389 & n3589 ) ;
  assign n3591 = ( n3300 & n3355 ) | ( n3300 & n3590 ) | ( n3355 & n3590 ) ;
  assign n3592 = ( ~n3239 & n3300 ) | ( ~n3239 & n3591 ) | ( n3300 & n3591 ) ;
  assign n3593 = ( n3153 & n3239 ) | ( n3153 & ~n3592 ) | ( n3239 & ~n3592 ) ;
  assign n3594 = ( n3078 & n3153 ) | ( n3078 & n3593 ) | ( n3153 & n3593 ) ;
  assign n3595 = ( ~n3046 & n3078 ) | ( ~n3046 & n3594 ) | ( n3078 & n3594 ) ;
  assign n3596 = ( n2965 & n3046 ) | ( n2965 & ~n3595 ) | ( n3046 & ~n3595 ) ;
  assign n3597 = ( n2910 & n2965 ) | ( n2910 & n3596 ) | ( n2965 & n3596 ) ;
  assign n3598 = ( ~n2843 & n2910 ) | ( ~n2843 & n3597 ) | ( n2910 & n3597 ) ;
  assign n3599 = ( n2810 & ~n2843 ) | ( n2810 & n3598 ) | ( ~n2843 & n3598 ) ;
  assign n3600 = ( n2725 & n2810 ) | ( n2725 & n3599 ) | ( n2810 & n3599 ) ;
  assign n3601 = ( ~n2635 & n2725 ) | ( ~n2635 & n3600 ) | ( n2725 & n3600 ) ;
  assign n3602 = ( n2552 & n2635 ) | ( n2552 & ~n3601 ) | ( n2635 & ~n3601 ) ;
  assign n3603 = ( ~n2491 & n2552 ) | ( ~n2491 & n3602 ) | ( n2552 & n3602 ) ;
  assign n3604 = ( n2396 & ~n2491 ) | ( n2396 & n3603 ) | ( ~n2491 & n3603 ) ;
  assign n3605 = ( ~n2298 & n2396 ) | ( ~n2298 & n3604 ) | ( n2396 & n3604 ) ;
  assign n3606 = ( n2270 & ~n2298 ) | ( n2270 & n3605 ) | ( ~n2298 & n3605 ) ;
  assign n3607 = ( n2174 & n2270 ) | ( n2174 & n3606 ) | ( n2270 & n3606 ) ;
  assign n3608 = ( n2089 & n2174 ) | ( n2089 & n3607 ) | ( n2174 & n3607 ) ;
  assign n3609 = ( ~n2023 & n2089 ) | ( ~n2023 & n3608 ) | ( n2089 & n3608 ) ;
  assign n3610 = ( n1926 & ~n2023 ) | ( n1926 & n3609 ) | ( ~n2023 & n3609 ) ;
  assign n3611 = ( n1852 & n1926 ) | ( n1852 & n3610 ) | ( n1926 & n3610 ) ;
  assign n3612 = ( ~n1750 & n1852 ) | ( ~n1750 & n3611 ) | ( n1852 & n3611 ) ;
  assign n3613 = ( n1669 & n1750 ) | ( n1669 & ~n3612 ) | ( n1750 & ~n3612 ) ;
  assign n3614 = ( ~n1576 & n1669 ) | ( ~n1576 & n3613 ) | ( n1669 & n3613 ) ;
  assign n3615 = ( n1458 & n1576 ) | ( n1458 & ~n3614 ) | ( n1576 & ~n3614 ) ;
  assign n3616 = ( ~n1338 & n1458 ) | ( ~n1338 & n3615 ) | ( n1458 & n3615 ) ;
  assign n3617 = ( n1267 & ~n1338 ) | ( n1267 & n3616 ) | ( ~n1338 & n3616 ) ;
  assign n3618 = ( ~n1246 & n1267 ) | ( ~n1246 & n3617 ) | ( n1267 & n3617 ) ;
  assign n3619 = ( n1246 & n1290 ) | ( n1246 & ~n3618 ) | ( n1290 & ~n3618 ) ;
  assign n3620 = ( n1246 & n1290 ) | ( n1246 & ~n3619 ) | ( n1290 & ~n3619 ) ;
  assign n3621 = ( n3618 & n3619 ) | ( n3618 & ~n3620 ) | ( n3619 & ~n3620 ) ;
  assign n3622 = n1248 & n3621 ;
  assign n3623 = n1292 | n3622 ;
  assign n3624 = ( n1040 & n1157 ) | ( n1040 & ~n3623 ) | ( n1157 & ~n3623 ) ;
  assign n3625 = ( n744 & n1040 ) | ( n744 & ~n3624 ) | ( n1040 & ~n3624 ) ;
  assign n3626 = ( n1040 & n1157 ) | ( n1040 & n3623 ) | ( n1157 & n3623 ) ;
  assign n3627 = ( n744 & n1157 ) | ( n744 & ~n3626 ) | ( n1157 & ~n3626 ) ;
  assign n3628 = ( ~n744 & n3625 ) | ( ~n744 & n3627 ) | ( n3625 & n3627 ) ;
  assign n3629 = n607 & ~n1246 ;
  assign n3630 = ( ~n41 & n54 ) | ( ~n41 & n78 ) | ( n54 & n78 ) ;
  assign n3631 = ( n463 & ~n1363 ) | ( n463 & n1595 ) | ( ~n1363 & n1595 ) ;
  assign n3632 = n1363 | n3631 ;
  assign n3633 = n1835 | n1870 ;
  assign n3634 = ( n3630 & ~n3632 ) | ( n3630 & n3633 ) | ( ~n3632 & n3633 ) ;
  assign n3635 = ( n63 & n70 ) | ( n63 & n261 ) | ( n70 & n261 ) ;
  assign n3636 = ( ~n54 & n166 ) | ( ~n54 & n3635 ) | ( n166 & n3635 ) ;
  assign n3637 = ( n57 & ~n78 ) | ( n57 & n145 ) | ( ~n78 & n145 ) ;
  assign n3638 = ( n1326 & ~n3636 ) | ( n1326 & n3637 ) | ( ~n3636 & n3637 ) ;
  assign n3639 = n3636 | n3638 ;
  assign n3640 = ( n3633 & n3634 ) | ( n3633 & n3639 ) | ( n3634 & n3639 ) ;
  assign n3641 = n3634 & ~n3640 ;
  assign n3642 = n267 | n455 ;
  assign n3643 = n217 | n641 ;
  assign n3644 = n747 | n1940 ;
  assign n3645 = ( n41 & n152 ) | ( n41 & n216 ) | ( n152 & n216 ) ;
  assign n3646 = n138 | n1122 ;
  assign n3647 = ( n66 & n72 ) | ( n66 & n122 ) | ( n72 & n122 ) ;
  assign n3648 = ( ~n3645 & n3646 ) | ( ~n3645 & n3647 ) | ( n3646 & n3647 ) ;
  assign n3649 = n3645 | n3648 ;
  assign n3650 = ( ~n3643 & n3644 ) | ( ~n3643 & n3649 ) | ( n3644 & n3649 ) ;
  assign n3651 = n3643 | n3650 ;
  assign n3652 = n428 | n3651 ;
  assign n3653 = ( n75 & n102 ) | ( n75 & n136 ) | ( n102 & n136 ) ;
  assign n3654 = ( ~n3088 & n3652 ) | ( ~n3088 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3655 = n3088 | n3654 ;
  assign n3656 = n408 | n3655 ;
  assign n3657 = ( n3641 & n3642 ) | ( n3641 & n3656 ) | ( n3642 & n3656 ) ;
  assign n3658 = n3641 & ~n3657 ;
  assign n3659 = n606 & ~n3658 ;
  assign n3660 = n3629 | n3659 ;
  assign n3661 = n1250 | n1290 ;
  assign n3662 = ( ~n1290 & n3660 ) | ( ~n1290 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3663 = ( n1290 & n3619 ) | ( n1290 & n3658 ) | ( n3619 & n3658 ) ;
  assign n3664 = ( n1290 & ~n3619 ) | ( n1290 & n3658 ) | ( ~n3619 & n3658 ) ;
  assign n3665 = ( n3619 & ~n3663 ) | ( n3619 & n3664 ) | ( ~n3663 & n3664 ) ;
  assign n3666 = n1248 & ~n3665 ;
  assign n3667 = n3662 | n3666 ;
  assign n3668 = n253 | n1254 ;
  assign n3669 = ( n41 & n44 ) | ( n41 & n72 ) | ( n44 & n72 ) ;
  assign n3670 = n591 | n3669 ;
  assign n3671 = ( ~n450 & n1032 ) | ( ~n450 & n3097 ) | ( n1032 & n3097 ) ;
  assign n3672 = n450 | n3671 ;
  assign n3673 = ( ~n3668 & n3670 ) | ( ~n3668 & n3672 ) | ( n3670 & n3672 ) ;
  assign n3674 = n3668 | n3673 ;
  assign n3675 = n84 | n952 ;
  assign n3676 = ( n152 & n160 ) | ( n152 & n3675 ) | ( n160 & n3675 ) ;
  assign n3677 = ( n41 & n50 ) | ( n41 & n160 ) | ( n50 & n160 ) ;
  assign n3678 = ( n2954 & ~n3676 ) | ( n2954 & n3677 ) | ( ~n3676 & n3677 ) ;
  assign n3679 = n3676 | n3678 ;
  assign n3680 = n147 | n441 ;
  assign n3681 = n1202 | n2787 ;
  assign n3682 = ( n75 & ~n78 ) | ( n75 & n160 ) | ( ~n78 & n160 ) ;
  assign n3683 = n3357 | n3682 ;
  assign n3684 = n3681 | n3683 ;
  assign n3685 = n3680 | n3684 ;
  assign n3686 = ( ~n3674 & n3679 ) | ( ~n3674 & n3685 ) | ( n3679 & n3685 ) ;
  assign n3687 = n3674 | n3686 ;
  assign n3688 = n254 | n3687 ;
  assign n3689 = n413 | n3688 ;
  assign n3690 = ( n3657 & ~n3663 ) | ( n3657 & n3689 ) | ( ~n3663 & n3689 ) ;
  assign n3691 = n3658 & ~n3690 ;
  assign n3692 = n3641 & ~n3689 ;
  assign n3693 = n3691 & ~n3692 ;
  assign n3694 = x28 | x29 ;
  assign n3695 = x26 | x27 ;
  assign n3696 = ( x26 & x27 ) | ( x26 & ~n3695 ) | ( x27 & ~n3695 ) ;
  assign n3697 = n3695 & ~n3696 ;
  assign n3698 = ( ~n46 & n53 ) | ( ~n46 & n3697 ) | ( n53 & n3697 ) ;
  assign n3699 = ( x28 & x29 ) | ( x28 & n3698 ) | ( x29 & n3698 ) ;
  assign n3700 = n3694 & ~n3699 ;
  assign n3701 = n3693 & n3700 ;
  assign n3702 = ( ~x29 & n3667 ) | ( ~x29 & n3701 ) | ( n3667 & n3701 ) ;
  assign n3703 = ( n3667 & n3701 ) | ( n3667 & ~n3702 ) | ( n3701 & ~n3702 ) ;
  assign n3704 = ( x29 & n3702 ) | ( x29 & ~n3703 ) | ( n3702 & ~n3703 ) ;
  assign n3705 = n3628 & n3704 ;
  assign n3706 = ~n3628 & n3704 ;
  assign n3707 = ( n3628 & ~n3705 ) | ( n3628 & n3706 ) | ( ~n3705 & n3706 ) ;
  assign n3708 = n1173 | n3637 ;
  assign n3709 = n337 | n465 ;
  assign n3710 = n1341 | n3709 ;
  assign n3711 = ( ~n54 & n80 ) | ( ~n54 & n102 ) | ( n80 & n102 ) ;
  assign n3712 = ( n734 & n1526 ) | ( n734 & ~n2224 ) | ( n1526 & ~n2224 ) ;
  assign n3713 = n2224 | n3712 ;
  assign n3714 = ( ~n3710 & n3711 ) | ( ~n3710 & n3713 ) | ( n3711 & n3713 ) ;
  assign n3715 = n3710 | n3714 ;
  assign n3716 = ( ~n2672 & n3708 ) | ( ~n2672 & n3715 ) | ( n3708 & n3715 ) ;
  assign n3717 = ( ~n923 & n2672 ) | ( ~n923 & n3716 ) | ( n2672 & n3716 ) ;
  assign n3718 = n992 | n1031 ;
  assign n3719 = ( n167 & n746 ) | ( n167 & ~n3718 ) | ( n746 & ~n3718 ) ;
  assign n3720 = n3718 | n3719 ;
  assign n3721 = ( n151 & n2362 ) | ( n151 & ~n2528 ) | ( n2362 & ~n2528 ) ;
  assign n3722 = ( n382 & n577 ) | ( n382 & ~n2528 ) | ( n577 & ~n2528 ) ;
  assign n3723 = n2528 | n3722 ;
  assign n3724 = ( ~n3720 & n3721 ) | ( ~n3720 & n3723 ) | ( n3721 & n3723 ) ;
  assign n3725 = n3720 | n3724 ;
  assign n3726 = ( n59 & n75 ) | ( n59 & n102 ) | ( n75 & n102 ) ;
  assign n3727 = n1225 | n3726 ;
  assign n3728 = ( n1772 & ~n3725 ) | ( n1772 & n3727 ) | ( ~n3725 & n3727 ) ;
  assign n3729 = n3725 | n3728 ;
  assign n3730 = n211 | n1280 ;
  assign n3731 = n348 | n764 ;
  assign n3732 = ( n1110 & ~n3730 ) | ( n1110 & n3731 ) | ( ~n3730 & n3731 ) ;
  assign n3733 = n3730 | n3732 ;
  assign n3734 = n272 | n500 ;
  assign n3735 = ( n316 & n517 ) | ( n316 & ~n3361 ) | ( n517 & ~n3361 ) ;
  assign n3736 = n3361 | n3735 ;
  assign n3737 = ( n780 & ~n3734 ) | ( n780 & n3736 ) | ( ~n3734 & n3736 ) ;
  assign n3738 = ( ~n3733 & n3734 ) | ( ~n3733 & n3737 ) | ( n3734 & n3737 ) ;
  assign n3739 = n3733 | n3738 ;
  assign n3740 = n176 | n360 ;
  assign n3741 = n254 | n3740 ;
  assign n3742 = n356 | n873 ;
  assign n3743 = n64 | n109 ;
  assign n3744 = ( n72 & n116 ) | ( n72 & n3743 ) | ( n116 & n3743 ) ;
  assign n3745 = ( n1133 & n3742 ) | ( n1133 & ~n3744 ) | ( n3742 & ~n3744 ) ;
  assign n3746 = n230 | n485 ;
  assign n3747 = n188 | n3746 ;
  assign n3748 = ( n3744 & ~n3745 ) | ( n3744 & n3747 ) | ( ~n3745 & n3747 ) ;
  assign n3749 = n3745 | n3748 ;
  assign n3750 = n137 | n290 ;
  assign n3751 = n885 | n3750 ;
  assign n3752 = ( n466 & n1136 ) | ( n466 & ~n3751 ) | ( n1136 & ~n3751 ) ;
  assign n3753 = n3751 | n3752 ;
  assign n3754 = ( ~n3741 & n3749 ) | ( ~n3741 & n3753 ) | ( n3749 & n3753 ) ;
  assign n3755 = n3741 | n3754 ;
  assign n3756 = ( ~n3729 & n3739 ) | ( ~n3729 & n3755 ) | ( n3739 & n3755 ) ;
  assign n3757 = n3729 | n3756 ;
  assign n3758 = n377 | n416 ;
  assign n3759 = n479 | n689 ;
  assign n3760 = n696 | n806 ;
  assign n3761 = n713 | n3760 ;
  assign n3762 = ( n528 & ~n3759 ) | ( n528 & n3761 ) | ( ~n3759 & n3761 ) ;
  assign n3763 = n3759 | n3762 ;
  assign n3764 = n123 | n144 ;
  assign n3765 = ( n228 & n1044 ) | ( n228 & ~n3764 ) | ( n1044 & ~n3764 ) ;
  assign n3766 = n3764 | n3765 ;
  assign n3767 = ( ~n377 & n3763 ) | ( ~n377 & n3766 ) | ( n3763 & n3766 ) ;
  assign n3768 = ( ~n1922 & n3758 ) | ( ~n1922 & n3767 ) | ( n3758 & n3767 ) ;
  assign n3769 = n1922 | n3768 ;
  assign n3770 = n923 | n3769 ;
  assign n3771 = ( ~n3717 & n3757 ) | ( ~n3717 & n3770 ) | ( n3757 & n3770 ) ;
  assign n3772 = n3717 | n3771 ;
  assign n3773 = ~n607 & n1458 ;
  assign n3774 = n1250 & ~n1338 ;
  assign n3775 = ( n1458 & ~n3773 ) | ( n1458 & n3774 ) | ( ~n3773 & n3774 ) ;
  assign n3776 = n606 & ~n1267 ;
  assign n3777 = ( n606 & n3775 ) | ( n606 & ~n3776 ) | ( n3775 & ~n3776 ) ;
  assign n3778 = ( n1267 & n1338 ) | ( n1267 & n3616 ) | ( n1338 & n3616 ) ;
  assign n3779 = ( n1338 & n3617 ) | ( n1338 & ~n3778 ) | ( n3617 & ~n3778 ) ;
  assign n3780 = n1248 & ~n3779 ;
  assign n3781 = n3777 | n3780 ;
  assign n3782 = ( ~n902 & n3772 ) | ( ~n902 & n3781 ) | ( n3772 & n3781 ) ;
  assign n3783 = ( n902 & n1039 ) | ( n902 & ~n1040 ) | ( n1039 & ~n1040 ) ;
  assign n3784 = ( x26 & n1040 ) | ( x26 & ~n3783 ) | ( n1040 & ~n3783 ) ;
  assign n3785 = n606 & ~n1246 ;
  assign n3786 = n607 & ~n1338 ;
  assign n3787 = n3785 | n3786 ;
  assign n3788 = ~n1250 & n1267 ;
  assign n3789 = ( n1267 & n3787 ) | ( n1267 & ~n3788 ) | ( n3787 & ~n3788 ) ;
  assign n3790 = ( n1246 & ~n1267 ) | ( n1246 & n3617 ) | ( ~n1267 & n3617 ) ;
  assign n3791 = ( ~n3617 & n3618 ) | ( ~n3617 & n3790 ) | ( n3618 & n3790 ) ;
  assign n3792 = n1248 & ~n3791 ;
  assign n3793 = n3789 | n3792 ;
  assign n3794 = ( n3782 & ~n3784 ) | ( n3782 & n3793 ) | ( ~n3784 & n3793 ) ;
  assign n3795 = ( n3623 & n3624 ) | ( n3623 & ~n3626 ) | ( n3624 & ~n3626 ) ;
  assign n3796 = ~n3690 & n3692 ;
  assign n3797 = ( n3692 & n3693 ) | ( n3692 & ~n3796 ) | ( n3693 & ~n3796 ) ;
  assign n3798 = ( x29 & ~n3694 ) | ( x29 & n3697 ) | ( ~n3694 & n3697 ) ;
  assign n3799 = ( x28 & ~n3694 ) | ( x28 & n3798 ) | ( ~n3694 & n3798 ) ;
  assign n3800 = n3697 & ~n3799 ;
  assign n3801 = n3797 & n3800 ;
  assign n3802 = ( n43 & n108 ) | ( n43 & ~n3697 ) | ( n108 & ~n3697 ) ;
  assign n3803 = ~n3692 & n3802 ;
  assign n3804 = ( n3658 & n3694 ) | ( n3658 & n3699 ) | ( n3694 & n3699 ) ;
  assign n3805 = ( n3694 & n3803 ) | ( n3694 & ~n3804 ) | ( n3803 & ~n3804 ) ;
  assign n3806 = ( ~x29 & n3801 ) | ( ~x29 & n3805 ) | ( n3801 & n3805 ) ;
  assign n3807 = ( n3801 & n3805 ) | ( n3801 & ~n3806 ) | ( n3805 & ~n3806 ) ;
  assign n3808 = ( x29 & n3806 ) | ( x29 & ~n3807 ) | ( n3806 & ~n3807 ) ;
  assign n3809 = ( n3794 & n3795 ) | ( n3794 & n3808 ) | ( n3795 & n3808 ) ;
  assign n3810 = n293 | n465 ;
  assign n3811 = ( n186 & n675 ) | ( n186 & ~n1692 ) | ( n675 & ~n1692 ) ;
  assign n3812 = n1692 | n3811 ;
  assign n3813 = ( n3221 & ~n3810 ) | ( n3221 & n3812 ) | ( ~n3810 & n3812 ) ;
  assign n3814 = n3810 | n3813 ;
  assign n3815 = n2316 | n3281 ;
  assign n3816 = ( n505 & n810 ) | ( n505 & ~n2443 ) | ( n810 & ~n2443 ) ;
  assign n3817 = n2443 | n3816 ;
  assign n3818 = n103 | n450 ;
  assign n3819 = n101 | n732 ;
  assign n3820 = ( n298 & n1082 ) | ( n298 & ~n3819 ) | ( n1082 & ~n3819 ) ;
  assign n3821 = n3819 | n3820 ;
  assign n3822 = ( n167 & ~n3818 ) | ( n167 & n3821 ) | ( ~n3818 & n3821 ) ;
  assign n3823 = n3818 | n3822 ;
  assign n3824 = ( ~n3815 & n3817 ) | ( ~n3815 & n3823 ) | ( n3817 & n3823 ) ;
  assign n3825 = n3815 | n3824 ;
  assign n3826 = n690 | n723 ;
  assign n3827 = n205 | n242 ;
  assign n3828 = n433 | n795 ;
  assign n3829 = ( n1556 & ~n3827 ) | ( n1556 & n3828 ) | ( ~n3827 & n3828 ) ;
  assign n3830 = n3827 | n3829 ;
  assign n3831 = ( n2846 & ~n3826 ) | ( n2846 & n3830 ) | ( ~n3826 & n3830 ) ;
  assign n3832 = n3826 | n3831 ;
  assign n3833 = ( n3814 & n3825 ) | ( n3814 & ~n3832 ) | ( n3825 & ~n3832 ) ;
  assign n3834 = n761 | n1522 ;
  assign n3835 = n188 | n273 ;
  assign n3836 = ( n57 & n73 ) | ( n57 & n84 ) | ( n73 & n84 ) ;
  assign n3837 = ( n545 & n1116 ) | ( n545 & ~n3836 ) | ( n1116 & ~n3836 ) ;
  assign n3838 = n3836 | n3837 ;
  assign n3839 = ( ~n3834 & n3835 ) | ( ~n3834 & n3838 ) | ( n3835 & n3838 ) ;
  assign n3840 = n3834 | n3839 ;
  assign n3841 = n142 | n582 ;
  assign n3842 = n1608 | n3841 ;
  assign n3843 = ( n57 & n100 ) | ( n57 & n109 ) | ( n100 & n109 ) ;
  assign n3844 = ( n41 & n48 ) | ( n41 & n129 ) | ( n48 & n129 ) ;
  assign n3845 = n990 | n3844 ;
  assign n3846 = ( n1405 & ~n3843 ) | ( n1405 & n3845 ) | ( ~n3843 & n3845 ) ;
  assign n3847 = n3843 | n3846 ;
  assign n3848 = ( n3038 & ~n3842 ) | ( n3038 & n3847 ) | ( ~n3842 & n3847 ) ;
  assign n3849 = n3842 | n3848 ;
  assign n3850 = ( n1509 & n2459 ) | ( n1509 & ~n3849 ) | ( n2459 & ~n3849 ) ;
  assign n3851 = n3849 | n3850 ;
  assign n3852 = n295 | n782 ;
  assign n3853 = n856 | n3852 ;
  assign n3854 = n92 | n550 ;
  assign n3855 = n1690 | n2766 ;
  assign n3856 = n3854 | n3855 ;
  assign n3857 = n507 | n642 ;
  assign n3858 = ( ~n3853 & n3856 ) | ( ~n3853 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3859 = n3853 | n3858 ;
  assign n3860 = n445 | n945 ;
  assign n3861 = ( n50 & ~n78 ) | ( n50 & n149 ) | ( ~n78 & n149 ) ;
  assign n3862 = n74 | n466 ;
  assign n3863 = n272 | n3862 ;
  assign n3864 = ( ~n3860 & n3861 ) | ( ~n3860 & n3863 ) | ( n3861 & n3863 ) ;
  assign n3865 = n3860 | n3864 ;
  assign n3866 = ( n3450 & ~n3859 ) | ( n3450 & n3865 ) | ( ~n3859 & n3865 ) ;
  assign n3867 = n3859 | n3866 ;
  assign n3868 = ( ~n3840 & n3851 ) | ( ~n3840 & n3867 ) | ( n3851 & n3867 ) ;
  assign n3869 = n3840 | n3868 ;
  assign n3870 = ( n3832 & ~n3833 ) | ( n3832 & n3869 ) | ( ~n3833 & n3869 ) ;
  assign n3871 = n3833 | n3870 ;
  assign n3872 = n703 | n1132 ;
  assign n3873 = n137 | n1450 ;
  assign n3874 = n144 | n225 ;
  assign n3875 = ( n132 & n301 ) | ( n132 & ~n3874 ) | ( n301 & ~n3874 ) ;
  assign n3876 = n3874 | n3875 ;
  assign n3877 = ( ~n3872 & n3873 ) | ( ~n3872 & n3876 ) | ( n3873 & n3876 ) ;
  assign n3878 = n3872 | n3877 ;
  assign n3879 = n262 | n642 ;
  assign n3880 = n2258 | n3879 ;
  assign n3881 = ( ~n657 & n685 ) | ( ~n657 & n1689 ) | ( n685 & n1689 ) ;
  assign n3882 = n657 | n3881 ;
  assign n3883 = n960 | n1171 ;
  assign n3884 = ( n185 & n534 ) | ( n185 & ~n3883 ) | ( n534 & ~n3883 ) ;
  assign n3885 = n3883 | n3884 ;
  assign n3886 = ( n73 & ~n78 ) | ( n73 & n84 ) | ( ~n78 & n84 ) ;
  assign n3887 = ( n72 & n75 ) | ( n72 & n136 ) | ( n75 & n136 ) ;
  assign n3888 = n3886 | n3887 ;
  assign n3889 = ( n239 & ~n609 ) | ( n239 & n3888 ) | ( ~n609 & n3888 ) ;
  assign n3890 = ( n517 & n609 ) | ( n517 & ~n3889 ) | ( n609 & ~n3889 ) ;
  assign n3891 = n3889 | n3890 ;
  assign n3892 = ( n727 & ~n3885 ) | ( n727 & n3891 ) | ( ~n3885 & n3891 ) ;
  assign n3893 = n3885 | n3892 ;
  assign n3894 = ( ~n3880 & n3882 ) | ( ~n3880 & n3893 ) | ( n3882 & n3893 ) ;
  assign n3895 = n3880 | n3894 ;
  assign n3896 = n377 | n1048 ;
  assign n3897 = n168 | n599 ;
  assign n3898 = ( n3391 & ~n3896 ) | ( n3391 & n3897 ) | ( ~n3896 & n3897 ) ;
  assign n3899 = n3896 | n3898 ;
  assign n3900 = n266 | n273 ;
  assign n3901 = ( n1376 & n1593 ) | ( n1376 & ~n3900 ) | ( n1593 & ~n3900 ) ;
  assign n3902 = n3900 | n3901 ;
  assign n3903 = ( ~n256 & n530 ) | ( ~n256 & n1056 ) | ( n530 & n1056 ) ;
  assign n3904 = n256 | n3903 ;
  assign n3905 = ( ~n3899 & n3902 ) | ( ~n3899 & n3904 ) | ( n3902 & n3904 ) ;
  assign n3906 = n3899 | n3905 ;
  assign n3907 = ( n3878 & n3895 ) | ( n3878 & ~n3906 ) | ( n3895 & ~n3906 ) ;
  assign n3908 = n292 | n1976 ;
  assign n3909 = n2518 | n3908 ;
  assign n3910 = ( ~n302 & n479 ) | ( ~n302 & n732 ) | ( n479 & n732 ) ;
  assign n3911 = n302 | n3910 ;
  assign n3912 = ( n163 & n211 ) | ( n163 & ~n1731 ) | ( n211 & ~n1731 ) ;
  assign n3913 = n1731 | n3912 ;
  assign n3914 = ( ~n3908 & n3911 ) | ( ~n3908 & n3913 ) | ( n3911 & n3913 ) ;
  assign n3915 = n330 | n361 ;
  assign n3916 = n590 | n3915 ;
  assign n3917 = ( n1660 & n2204 ) | ( n1660 & ~n3916 ) | ( n2204 & ~n3916 ) ;
  assign n3918 = n3916 | n3917 ;
  assign n3919 = n991 | n1145 ;
  assign n3920 = n904 | n2929 ;
  assign n3921 = ( n1655 & ~n3919 ) | ( n1655 & n3920 ) | ( ~n3919 & n3920 ) ;
  assign n3922 = n3919 | n3921 ;
  assign n3923 = ( n1035 & ~n3918 ) | ( n1035 & n3922 ) | ( ~n3918 & n3922 ) ;
  assign n3924 = n3918 | n3923 ;
  assign n3925 = ( n3909 & n3914 ) | ( n3909 & ~n3924 ) | ( n3914 & ~n3924 ) ;
  assign n3926 = n105 | n234 ;
  assign n3927 = ( n783 & n822 ) | ( n783 & ~n3926 ) | ( n822 & ~n3926 ) ;
  assign n3928 = n3926 | n3927 ;
  assign n3929 = n288 | n1008 ;
  assign n3930 = n507 | n638 ;
  assign n3931 = n74 | n91 ;
  assign n3932 = ( ~n654 & n1998 ) | ( ~n654 & n3931 ) | ( n1998 & n3931 ) ;
  assign n3933 = ( n654 & ~n3930 ) | ( n654 & n3932 ) | ( ~n3930 & n3932 ) ;
  assign n3934 = n3930 | n3933 ;
  assign n3935 = n161 | n857 ;
  assign n3936 = ( n3929 & n3934 ) | ( n3929 & ~n3935 ) | ( n3934 & ~n3935 ) ;
  assign n3937 = ( n1350 & n3935 ) | ( n1350 & ~n3936 ) | ( n3935 & ~n3936 ) ;
  assign n3938 = n3936 | n3937 ;
  assign n3939 = ( ~n78 & n84 ) | ( ~n78 & n216 ) | ( n84 & n216 ) ;
  assign n3940 = ( n992 & n1556 ) | ( n992 & ~n3939 ) | ( n1556 & ~n3939 ) ;
  assign n3941 = n3939 | n3940 ;
  assign n3942 = ( ~n3928 & n3938 ) | ( ~n3928 & n3941 ) | ( n3938 & n3941 ) ;
  assign n3943 = n3928 | n3942 ;
  assign n3944 = ( n3924 & ~n3925 ) | ( n3924 & n3943 ) | ( ~n3925 & n3943 ) ;
  assign n3945 = n3925 | n3944 ;
  assign n3946 = ( n3906 & ~n3907 ) | ( n3906 & n3945 ) | ( ~n3907 & n3945 ) ;
  assign n3947 = n3907 | n3946 ;
  assign n3948 = ( ~x23 & n3871 ) | ( ~x23 & n3947 ) | ( n3871 & n3947 ) ;
  assign n3949 = n606 | n1338 ;
  assign n3950 = n1250 & n1458 ;
  assign n3951 = ( ~n1338 & n3949 ) | ( ~n1338 & n3950 ) | ( n3949 & n3950 ) ;
  assign n3952 = n607 & ~n1576 ;
  assign n3953 = ( n607 & n3951 ) | ( n607 & ~n3952 ) | ( n3951 & ~n3952 ) ;
  assign n3954 = ( n1338 & n1458 ) | ( n1338 & ~n3615 ) | ( n1458 & ~n3615 ) ;
  assign n3955 = ( ~n1458 & n3616 ) | ( ~n1458 & n3954 ) | ( n3616 & n3954 ) ;
  assign n3956 = n1248 & ~n3955 ;
  assign n3957 = n3953 | n3956 ;
  assign n3958 = ( ~n902 & n3948 ) | ( ~n902 & n3957 ) | ( n3948 & n3957 ) ;
  assign n3959 = n489 | n1007 ;
  assign n3960 = ( n116 & n160 ) | ( n116 & n166 ) | ( n160 & n166 ) ;
  assign n3961 = n173 | n685 ;
  assign n3962 = n218 & ~n361 ;
  assign n3963 = ( n978 & ~n2399 ) | ( n978 & n3962 ) | ( ~n2399 & n3962 ) ;
  assign n3964 = ( ~n978 & n3961 ) | ( ~n978 & n3963 ) | ( n3961 & n3963 ) ;
  assign n3965 = ~n3961 & n3964 ;
  assign n3966 = ( n3959 & ~n3960 ) | ( n3959 & n3965 ) | ( ~n3960 & n3965 ) ;
  assign n3967 = ~n3959 & n3966 ;
  assign n3968 = n395 | n1174 ;
  assign n3969 = n212 | n888 ;
  assign n3970 = n3968 | n3969 ;
  assign n3971 = n505 | n544 ;
  assign n3972 = ( n57 & n72 ) | ( n57 & n116 ) | ( n72 & n116 ) ;
  assign n3973 = ( n2306 & n3971 ) | ( n2306 & ~n3972 ) | ( n3971 & ~n3972 ) ;
  assign n3974 = ( n104 & n205 ) | ( n104 & ~n1059 ) | ( n205 & ~n1059 ) ;
  assign n3975 = n1059 | n3974 ;
  assign n3976 = ( n3972 & ~n3973 ) | ( n3972 & n3975 ) | ( ~n3973 & n3975 ) ;
  assign n3977 = n3973 | n3976 ;
  assign n3978 = ( n3967 & n3970 ) | ( n3967 & ~n3977 ) | ( n3970 & ~n3977 ) ;
  assign n3979 = ( n1775 & n3970 ) | ( n1775 & n3978 ) | ( n3970 & n3978 ) ;
  assign n3980 = n3978 & ~n3979 ;
  assign n3981 = n2057 | n3210 ;
  assign n3982 = n1116 | n2575 ;
  assign n3983 = n231 | n657 ;
  assign n3984 = n688 | n3983 ;
  assign n3985 = ( n974 & ~n3982 ) | ( n974 & n3984 ) | ( ~n3982 & n3984 ) ;
  assign n3986 = n3982 | n3985 ;
  assign n3987 = ( n124 & n536 ) | ( n124 & ~n928 ) | ( n536 & ~n928 ) ;
  assign n3988 = n928 | n3987 ;
  assign n3989 = ( n80 & n83 ) | ( n80 & n97 ) | ( n83 & n97 ) ;
  assign n3990 = ( n189 & ~n3988 ) | ( n189 & n3989 ) | ( ~n3988 & n3989 ) ;
  assign n3991 = n3988 | n3990 ;
  assign n3992 = n1185 | n1253 ;
  assign n3993 = ( n2799 & n3991 ) | ( n2799 & ~n3992 ) | ( n3991 & ~n3992 ) ;
  assign n3994 = ( n75 & n97 ) | ( n75 & n119 ) | ( n97 & n119 ) ;
  assign n3995 = ( n3992 & ~n3993 ) | ( n3992 & n3994 ) | ( ~n3993 & n3994 ) ;
  assign n3996 = n3993 | n3995 ;
  assign n3997 = n753 | n1365 ;
  assign n3998 = n551 | n913 ;
  assign n3999 = n3997 | n3998 ;
  assign n4000 = ( ~n3986 & n3996 ) | ( ~n3986 & n3999 ) | ( n3996 & n3999 ) ;
  assign n4001 = n3986 | n4000 ;
  assign n4002 = ( n3980 & n3981 ) | ( n3980 & n4001 ) | ( n3981 & n4001 ) ;
  assign n4003 = n3980 & ~n4002 ;
  assign n4004 = n291 | n455 ;
  assign n4005 = n212 | n4004 ;
  assign n4006 = n723 | n3051 ;
  assign n4007 = n115 | n224 ;
  assign n4008 = n1515 | n4007 ;
  assign n4009 = n4006 | n4008 ;
  assign n4010 = ( n1148 & ~n4005 ) | ( n1148 & n4009 ) | ( ~n4005 & n4009 ) ;
  assign n4011 = n4005 | n4010 ;
  assign n4012 = n815 | n2726 ;
  assign n4013 = n259 | n1096 ;
  assign n4014 = ( n48 & n84 ) | ( n48 & n100 ) | ( n84 & n100 ) ;
  assign n4015 = n416 | n4014 ;
  assign n4016 = ( n41 & n145 ) | ( n41 & n933 ) | ( n145 & n933 ) ;
  assign n4017 = ( ~n4013 & n4015 ) | ( ~n4013 & n4016 ) | ( n4015 & n4016 ) ;
  assign n4018 = n4013 | n4017 ;
  assign n4019 = ( n3975 & n4012 ) | ( n3975 & ~n4018 ) | ( n4012 & ~n4018 ) ;
  assign n4020 = n1220 | n1751 ;
  assign n4021 = ( n4018 & ~n4019 ) | ( n4018 & n4020 ) | ( ~n4019 & n4020 ) ;
  assign n4022 = n4019 | n4021 ;
  assign n4023 = ( n2815 & ~n4011 ) | ( n2815 & n4022 ) | ( ~n4011 & n4022 ) ;
  assign n4024 = n4011 | n4023 ;
  assign n4025 = n2511 | n4024 ;
  assign n4026 = ( n476 & n2307 ) | ( n476 & ~n3514 ) | ( n2307 & ~n3514 ) ;
  assign n4027 = n3514 | n4026 ;
  assign n4028 = n231 | n3173 ;
  assign n4029 = n293 | n941 ;
  assign n4030 = n388 | n582 ;
  assign n4031 = ( n1129 & ~n4029 ) | ( n1129 & n4030 ) | ( ~n4029 & n4030 ) ;
  assign n4032 = n4029 | n4031 ;
  assign n4033 = n4028 | n4032 ;
  assign n4034 = n824 | n2798 ;
  assign n4035 = n286 | n690 ;
  assign n4036 = n4034 | n4035 ;
  assign n4037 = n124 | n165 ;
  assign n4038 = n347 | n1314 ;
  assign n4039 = n4037 | n4038 ;
  assign n4040 = n4036 | n4039 ;
  assign n4041 = ( ~n4027 & n4033 ) | ( ~n4027 & n4040 ) | ( n4033 & n4040 ) ;
  assign n4042 = n4027 | n4041 ;
  assign n4043 = n789 | n1720 ;
  assign n4044 = n137 | n186 ;
  assign n4045 = ( n239 & n599 ) | ( n239 & ~n4044 ) | ( n599 & ~n4044 ) ;
  assign n4046 = n4044 | n4045 ;
  assign n4047 = n178 | n3539 ;
  assign n4048 = n1839 | n2029 ;
  assign n4049 = n1533 | n1891 ;
  assign n4050 = n4048 | n4049 ;
  assign n4051 = n4047 | n4050 ;
  assign n4052 = ( ~n4043 & n4046 ) | ( ~n4043 & n4051 ) | ( n4046 & n4051 ) ;
  assign n4053 = n4043 | n4052 ;
  assign n4054 = ( n1278 & n2266 ) | ( n1278 & ~n4053 ) | ( n2266 & ~n4053 ) ;
  assign n4055 = n4053 | n4054 ;
  assign n4056 = ( ~n4025 & n4042 ) | ( ~n4025 & n4055 ) | ( n4042 & n4055 ) ;
  assign n4057 = n4025 | n4056 ;
  assign n4058 = ( n1526 & n1556 ) | ( n1526 & ~n3879 ) | ( n1556 & ~n3879 ) ;
  assign n4059 = n3879 | n4058 ;
  assign n4060 = n1174 | n1320 ;
  assign n4061 = n394 | n1870 ;
  assign n4062 = n153 | n4061 ;
  assign n4063 = ( ~n4059 & n4060 ) | ( ~n4059 & n4062 ) | ( n4060 & n4062 ) ;
  assign n4064 = n4059 | n4063 ;
  assign n4065 = n238 | n753 ;
  assign n4066 = n978 | n1720 ;
  assign n4067 = ( n2181 & n2214 ) | ( n2181 & ~n4066 ) | ( n2214 & ~n4066 ) ;
  assign n4068 = n4066 | n4067 ;
  assign n4069 = n164 | n493 ;
  assign n4070 = n3168 | n4069 ;
  assign n4071 = ( n4065 & n4068 ) | ( n4065 & ~n4070 ) | ( n4068 & ~n4070 ) ;
  assign n4072 = n123 | n506 ;
  assign n4073 = ( n4070 & ~n4071 ) | ( n4070 & n4072 ) | ( ~n4071 & n4072 ) ;
  assign n4074 = n4071 | n4073 ;
  assign n4075 = n54 & ~n83 ;
  assign n4076 = ( n50 & n119 ) | ( n50 & ~n4075 ) | ( n119 & ~n4075 ) ;
  assign n4077 = ( n2073 & ~n3571 ) | ( n2073 & n4076 ) | ( ~n3571 & n4076 ) ;
  assign n4078 = n3571 | n4077 ;
  assign n4079 = ( ~n4064 & n4074 ) | ( ~n4064 & n4078 ) | ( n4074 & n4078 ) ;
  assign n4080 = n4064 | n4079 ;
  assign n4081 = n1356 | n1522 ;
  assign n4082 = ( n866 & n1078 ) | ( n866 & ~n4081 ) | ( n1078 & ~n4081 ) ;
  assign n4083 = n4081 | n4082 ;
  assign n4084 = ( n1311 & ~n3212 ) | ( n1311 & n4083 ) | ( ~n3212 & n4083 ) ;
  assign n4085 = n60 | n448 ;
  assign n4086 = ( n291 & n928 ) | ( n291 & ~n4085 ) | ( n928 & ~n4085 ) ;
  assign n4087 = n4085 | n4086 ;
  assign n4088 = ( n3212 & ~n4084 ) | ( n3212 & n4087 ) | ( ~n4084 & n4087 ) ;
  assign n4089 = n4084 | n4088 ;
  assign n4090 = n538 | n1838 ;
  assign n4091 = n1199 | n1363 ;
  assign n4092 = n599 | n990 ;
  assign n4093 = n294 | n361 ;
  assign n4094 = ( ~n132 & n549 ) | ( ~n132 & n689 ) | ( n549 & n689 ) ;
  assign n4095 = n132 | n4094 ;
  assign n4096 = ( ~n4092 & n4093 ) | ( ~n4092 & n4095 ) | ( n4093 & n4095 ) ;
  assign n4097 = n4092 | n4096 ;
  assign n4098 = ( ~n4090 & n4091 ) | ( ~n4090 & n4097 ) | ( n4091 & n4097 ) ;
  assign n4099 = n4090 | n4098 ;
  assign n4100 = n1009 | n1237 ;
  assign n4101 = n1647 | n4100 ;
  assign n4102 = ( n41 & ~n54 ) | ( n41 & n152 ) | ( ~n54 & n152 ) ;
  assign n4103 = ( n73 & n80 ) | ( n73 & n352 ) | ( n80 & n352 ) ;
  assign n4104 = n4102 | n4103 ;
  assign n4105 = n479 | n1225 ;
  assign n4106 = n203 | n4105 ;
  assign n4107 = ( n686 & n2011 ) | ( n686 & ~n4106 ) | ( n2011 & ~n4106 ) ;
  assign n4108 = n4106 | n4107 ;
  assign n4109 = ( ~n4101 & n4104 ) | ( ~n4101 & n4108 ) | ( n4104 & n4108 ) ;
  assign n4110 = n4101 | n4109 ;
  assign n4111 = ( n2548 & ~n4099 ) | ( n2548 & n4110 ) | ( ~n4099 & n4110 ) ;
  assign n4112 = n4099 | n4111 ;
  assign n4113 = n419 | n3339 ;
  assign n4114 = n171 | n856 ;
  assign n4115 = n202 | n500 ;
  assign n4116 = ( n941 & n992 ) | ( n941 & ~n1341 ) | ( n992 & ~n1341 ) ;
  assign n4117 = n1341 | n4116 ;
  assign n4118 = ( n135 & ~n4115 ) | ( n135 & n4117 ) | ( ~n4115 & n4117 ) ;
  assign n4119 = n4115 | n4118 ;
  assign n4120 = ( ~n4113 & n4114 ) | ( ~n4113 & n4119 ) | ( n4114 & n4119 ) ;
  assign n4121 = n4113 | n4120 ;
  assign n4122 = ( ~n4089 & n4112 ) | ( ~n4089 & n4121 ) | ( n4112 & n4121 ) ;
  assign n4123 = n4089 | n4122 ;
  assign n4124 = ( n102 & n116 ) | ( n102 & n129 ) | ( n116 & n129 ) ;
  assign n4125 = n1365 | n4124 ;
  assign n4126 = ( n98 & n102 ) | ( n98 & n122 ) | ( n102 & n122 ) ;
  assign n4127 = ( n48 & n50 ) | ( n48 & n83 ) | ( n50 & n83 ) ;
  assign n4128 = n4126 | n4127 ;
  assign n4129 = ( n145 & n261 ) | ( n145 & n3635 ) | ( n261 & n3635 ) ;
  assign n4130 = ( n241 & n353 ) | ( n241 & ~n4129 ) | ( n353 & ~n4129 ) ;
  assign n4131 = n4129 | n4130 ;
  assign n4132 = ( n4125 & ~n4128 ) | ( n4125 & n4131 ) | ( ~n4128 & n4131 ) ;
  assign n4133 = n878 | n1059 ;
  assign n4134 = n386 | n4133 ;
  assign n4135 = ( n4128 & ~n4132 ) | ( n4128 & n4134 ) | ( ~n4132 & n4134 ) ;
  assign n4136 = n4132 | n4135 ;
  assign n4137 = ( ~n4080 & n4123 ) | ( ~n4080 & n4136 ) | ( n4123 & n4136 ) ;
  assign n4138 = n4080 | n4137 ;
  assign n4139 = ( ~x20 & n4057 ) | ( ~x20 & n4138 ) | ( n4057 & n4138 ) ;
  assign n4140 = ~n607 & n1852 ;
  assign n4141 = n1250 & ~n1750 ;
  assign n4142 = ( n1852 & ~n4140 ) | ( n1852 & n4141 ) | ( ~n4140 & n4141 ) ;
  assign n4143 = n606 & n1669 ;
  assign n4144 = ( n606 & n4142 ) | ( n606 & ~n4143 ) | ( n4142 & ~n4143 ) ;
  assign n4145 = ( n1669 & n1750 ) | ( n1669 & ~n3613 ) | ( n1750 & ~n3613 ) ;
  assign n4146 = ( n3612 & n3613 ) | ( n3612 & ~n4145 ) | ( n3613 & ~n4145 ) ;
  assign n4147 = n1248 & n4146 ;
  assign n4148 = n4144 | n4147 ;
  assign n4149 = ( n4003 & n4139 ) | ( n4003 & n4148 ) | ( n4139 & n4148 ) ;
  assign n4150 = ( n3871 & n4003 ) | ( n3871 & ~n4149 ) | ( n4003 & ~n4149 ) ;
  assign n4151 = ( n3871 & n3947 ) | ( n3871 & ~n3948 ) | ( n3947 & ~n3948 ) ;
  assign n4152 = ( x23 & n3948 ) | ( x23 & ~n4151 ) | ( n3948 & ~n4151 ) ;
  assign n4153 = ~n606 & n1458 ;
  assign n4154 = n607 & ~n1669 ;
  assign n4155 = ( n1458 & ~n4153 ) | ( n1458 & n4154 ) | ( ~n4153 & n4154 ) ;
  assign n4156 = ~n1250 & n1576 ;
  assign n4157 = ( n1576 & n4155 ) | ( n1576 & ~n4156 ) | ( n4155 & ~n4156 ) ;
  assign n4158 = ( n1458 & n1576 ) | ( n1458 & ~n3615 ) | ( n1576 & ~n3615 ) ;
  assign n4159 = ( n3614 & n3615 ) | ( n3614 & ~n4158 ) | ( n3615 & ~n4158 ) ;
  assign n4160 = n1248 & ~n4159 ;
  assign n4161 = n4157 | n4160 ;
  assign n4162 = ( n4150 & n4152 ) | ( n4150 & ~n4161 ) | ( n4152 & ~n4161 ) ;
  assign n4163 = ( n902 & ~n3948 ) | ( n902 & n3957 ) | ( ~n3948 & n3957 ) ;
  assign n4164 = ( ~n3957 & n3958 ) | ( ~n3957 & n4163 ) | ( n3958 & n4163 ) ;
  assign n4165 = n3621 & n3800 ;
  assign n4166 = ~n1290 & n3799 ;
  assign n4167 = ~n1246 & n3802 ;
  assign n4168 = ( ~n1267 & n3694 ) | ( ~n1267 & n3699 ) | ( n3694 & n3699 ) ;
  assign n4169 = ( n3694 & n4167 ) | ( n3694 & ~n4168 ) | ( n4167 & ~n4168 ) ;
  assign n4170 = ( ~n4165 & n4166 ) | ( ~n4165 & n4169 ) | ( n4166 & n4169 ) ;
  assign n4171 = ( ~x29 & n4165 ) | ( ~x29 & n4170 ) | ( n4165 & n4170 ) ;
  assign n4172 = ( n4165 & n4170 ) | ( n4165 & ~n4171 ) | ( n4170 & ~n4171 ) ;
  assign n4173 = ( x29 & n4171 ) | ( x29 & ~n4172 ) | ( n4171 & ~n4172 ) ;
  assign n4174 = ( n4162 & n4164 ) | ( n4162 & ~n4173 ) | ( n4164 & ~n4173 ) ;
  assign n4175 = ( n3772 & n3781 ) | ( n3772 & ~n3782 ) | ( n3781 & ~n3782 ) ;
  assign n4176 = ( n902 & n3782 ) | ( n902 & ~n4175 ) | ( n3782 & ~n4175 ) ;
  assign n4177 = ( ~n3958 & n4174 ) | ( ~n3958 & n4176 ) | ( n4174 & n4176 ) ;
  assign n4178 = ( ~n3782 & n3784 ) | ( ~n3782 & n3793 ) | ( n3784 & n3793 ) ;
  assign n4179 = ( ~n3793 & n3794 ) | ( ~n3793 & n4178 ) | ( n3794 & n4178 ) ;
  assign n4180 = ( n3658 & n3663 ) | ( n3658 & ~n3692 ) | ( n3663 & ~n3692 ) ;
  assign n4181 = ( n3658 & n3663 ) | ( n3658 & ~n4180 ) | ( n3663 & ~n4180 ) ;
  assign n4182 = ( n3692 & n4180 ) | ( n3692 & ~n4181 ) | ( n4180 & ~n4181 ) ;
  assign n4183 = n3800 & ~n4182 ;
  assign n4184 = ~n1290 & n3700 ;
  assign n4185 = n3692 & n3799 ;
  assign n4186 = ~n3658 & n3802 ;
  assign n4187 = ( n3799 & ~n4185 ) | ( n3799 & n4186 ) | ( ~n4185 & n4186 ) ;
  assign n4188 = ( ~n4183 & n4184 ) | ( ~n4183 & n4187 ) | ( n4184 & n4187 ) ;
  assign n4189 = ( ~x29 & n4183 ) | ( ~x29 & n4188 ) | ( n4183 & n4188 ) ;
  assign n4190 = ( n4183 & n4188 ) | ( n4183 & ~n4189 ) | ( n4188 & ~n4189 ) ;
  assign n4191 = ( x29 & n4189 ) | ( x29 & ~n4190 ) | ( n4189 & ~n4190 ) ;
  assign n4192 = ( n4177 & n4179 ) | ( n4177 & ~n4191 ) | ( n4179 & ~n4191 ) ;
  assign n4193 = x23 | x24 ;
  assign n4194 = ( x23 & x24 ) | ( x23 & ~n4193 ) | ( x24 & ~n4193 ) ;
  assign n4195 = n4193 & ~n4194 ;
  assign n4196 = ( ~n39 & n56 ) | ( ~n39 & n4195 ) | ( n56 & n4195 ) ;
  assign n4197 = x25 | x26 ;
  assign n4198 = x25 & x26 ;
  assign n4199 = n4197 & ~n4198 ;
  assign n4200 = ~n4196 & n4199 ;
  assign n4201 = ( n4195 & ~n4197 ) | ( n4195 & n4198 ) | ( ~n4197 & n4198 ) ;
  assign n4202 = n4195 & ~n4201 ;
  assign n4203 = ~n3691 & n4202 ;
  assign n4204 = ( ~n3692 & n4200 ) | ( ~n3692 & n4203 ) | ( n4200 & n4203 ) ;
  assign n4205 = x26 | n4204 ;
  assign n4206 = ( x26 & n4204 ) | ( x26 & ~n4205 ) | ( n4204 & ~n4205 ) ;
  assign n4207 = n4205 & ~n4206 ;
  assign n4208 = ~n3665 & n3800 ;
  assign n4209 = ~n1290 & n3802 ;
  assign n4210 = n1246 & n3700 ;
  assign n4211 = ~n3658 & n3799 ;
  assign n4212 = ( n3700 & ~n4210 ) | ( n3700 & n4211 ) | ( ~n4210 & n4211 ) ;
  assign n4213 = ( ~n4208 & n4209 ) | ( ~n4208 & n4212 ) | ( n4209 & n4212 ) ;
  assign n4214 = ( ~x29 & n4208 ) | ( ~x29 & n4213 ) | ( n4208 & n4213 ) ;
  assign n4215 = ( n4208 & n4213 ) | ( n4208 & ~n4214 ) | ( n4213 & ~n4214 ) ;
  assign n4216 = ( x29 & n4214 ) | ( x29 & ~n4215 ) | ( n4214 & ~n4215 ) ;
  assign n4217 = ( n4174 & n4176 ) | ( n4174 & ~n4177 ) | ( n4176 & ~n4177 ) ;
  assign n4218 = ( n3958 & n4177 ) | ( n3958 & ~n4217 ) | ( n4177 & ~n4217 ) ;
  assign n4219 = ( n4207 & n4216 ) | ( n4207 & n4218 ) | ( n4216 & n4218 ) ;
  assign n4220 = ( n59 & n97 ) | ( n59 & n129 ) | ( n97 & n129 ) ;
  assign n4221 = n111 | n796 ;
  assign n4222 = n4220 | n4221 ;
  assign n4223 = n317 | n1341 ;
  assign n4224 = n512 | n4223 ;
  assign n4225 = n1964 | n4224 ;
  assign n4226 = n4222 | n4225 ;
  assign n4227 = n528 | n1173 ;
  assign n4228 = n211 | n576 ;
  assign n4229 = ( n745 & n4227 ) | ( n745 & ~n4228 ) | ( n4227 & ~n4228 ) ;
  assign n4230 = n115 | n144 ;
  assign n4231 = n960 | n992 ;
  assign n4232 = ( n148 & n895 ) | ( n148 & ~n4231 ) | ( n895 & ~n4231 ) ;
  assign n4233 = n4231 | n4232 ;
  assign n4234 = ( n172 & ~n4230 ) | ( n172 & n4233 ) | ( ~n4230 & n4233 ) ;
  assign n4235 = n4230 | n4234 ;
  assign n4236 = ( n4228 & ~n4229 ) | ( n4228 & n4235 ) | ( ~n4229 & n4235 ) ;
  assign n4237 = n4229 | n4236 ;
  assign n4238 = n1793 | n2011 ;
  assign n4239 = n2024 | n4238 ;
  assign n4240 = ( n1055 & n1558 ) | ( n1055 & ~n4239 ) | ( n1558 & ~n4239 ) ;
  assign n4241 = n4239 | n4240 ;
  assign n4242 = ( ~n4226 & n4237 ) | ( ~n4226 & n4241 ) | ( n4237 & n4241 ) ;
  assign n4243 = n4226 | n4242 ;
  assign n4244 = n2093 | n2256 ;
  assign n4245 = ( n689 & ~n981 ) | ( n689 & n2214 ) | ( ~n981 & n2214 ) ;
  assign n4246 = n981 | n4245 ;
  assign n4247 = n226 | n1739 ;
  assign n4248 = ( ~n4244 & n4246 ) | ( ~n4244 & n4247 ) | ( n4246 & n4247 ) ;
  assign n4249 = n4244 | n4248 ;
  assign n4250 = n140 | n1634 ;
  assign n4251 = n189 | n205 ;
  assign n4252 = ( n534 & n1365 ) | ( n534 & ~n4251 ) | ( n1365 & ~n4251 ) ;
  assign n4253 = n4251 | n4252 ;
  assign n4254 = n691 | n851 ;
  assign n4255 = n104 | n240 ;
  assign n4256 = n261 | n4255 ;
  assign n4257 = n753 | n3523 ;
  assign n4258 = n4256 | n4257 ;
  assign n4259 = ( n150 & ~n4254 ) | ( n150 & n4258 ) | ( ~n4254 & n4258 ) ;
  assign n4260 = n4254 | n4259 ;
  assign n4261 = ( ~n4250 & n4253 ) | ( ~n4250 & n4260 ) | ( n4253 & n4260 ) ;
  assign n4262 = ( ~n637 & n933 ) | ( ~n637 & n1835 ) | ( n933 & n1835 ) ;
  assign n4263 = n637 | n4262 ;
  assign n4264 = ( n4250 & ~n4261 ) | ( n4250 & n4263 ) | ( ~n4261 & n4263 ) ;
  assign n4265 = n4261 | n4264 ;
  assign n4266 = ( n394 & n1044 ) | ( n394 & ~n2430 ) | ( n1044 & ~n2430 ) ;
  assign n4267 = n2430 | n4266 ;
  assign n4268 = ( ~n4249 & n4265 ) | ( ~n4249 & n4267 ) | ( n4265 & n4267 ) ;
  assign n4269 = n4249 | n4268 ;
  assign n4270 = n4243 | n4269 ;
  assign n4271 = n207 | n337 ;
  assign n4272 = n117 | n4271 ;
  assign n4273 = n320 | n978 ;
  assign n4274 = ( n2204 & n3841 ) | ( n2204 & ~n4273 ) | ( n3841 & ~n4273 ) ;
  assign n4275 = ( n356 & n1510 ) | ( n356 & ~n4273 ) | ( n1510 & ~n4273 ) ;
  assign n4276 = n4273 | n4275 ;
  assign n4277 = ( ~n4272 & n4274 ) | ( ~n4272 & n4276 ) | ( n4274 & n4276 ) ;
  assign n4278 = n4272 | n4277 ;
  assign n4279 = n1833 | n3103 ;
  assign n4280 = ~n2070 & n2885 ;
  assign n4281 = ( n4278 & ~n4279 ) | ( n4278 & n4280 ) | ( ~n4279 & n4280 ) ;
  assign n4282 = ( n4270 & ~n4278 ) | ( n4270 & n4281 ) | ( ~n4278 & n4281 ) ;
  assign n4283 = ~n4270 & n4282 ;
  assign n4284 = n607 | n2023 ;
  assign n4285 = n1250 & n1926 ;
  assign n4286 = ( ~n2023 & n4284 ) | ( ~n2023 & n4285 ) | ( n4284 & n4285 ) ;
  assign n4287 = n606 & ~n1852 ;
  assign n4288 = ( n606 & n4286 ) | ( n606 & ~n4287 ) | ( n4286 & ~n4287 ) ;
  assign n4289 = ( n1852 & ~n1926 ) | ( n1852 & n3610 ) | ( ~n1926 & n3610 ) ;
  assign n4290 = ( n1926 & ~n3611 ) | ( n1926 & n4289 ) | ( ~n3611 & n4289 ) ;
  assign n4291 = n1248 & n4290 ;
  assign n4292 = n4288 | n4291 ;
  assign n4293 = ( n4057 & n4283 ) | ( n4057 & ~n4292 ) | ( n4283 & ~n4292 ) ;
  assign n4294 = ( n4057 & n4138 ) | ( n4057 & ~n4139 ) | ( n4138 & ~n4139 ) ;
  assign n4295 = ( x20 & n4139 ) | ( x20 & ~n4294 ) | ( n4139 & ~n4294 ) ;
  assign n4296 = n1250 & n1852 ;
  assign n4297 = n607 & n1926 ;
  assign n4298 = n4296 | n4297 ;
  assign n4299 = n606 & n1750 ;
  assign n4300 = ( n606 & n4298 ) | ( n606 & ~n4299 ) | ( n4298 & ~n4299 ) ;
  assign n4301 = ( n1750 & ~n1852 ) | ( n1750 & n3611 ) | ( ~n1852 & n3611 ) ;
  assign n4302 = ( ~n3611 & n3612 ) | ( ~n3611 & n4301 ) | ( n3612 & n4301 ) ;
  assign n4303 = n1248 & ~n4302 ;
  assign n4304 = n4300 | n4303 ;
  assign n4305 = ( n4293 & n4295 ) | ( n4293 & ~n4304 ) | ( n4295 & ~n4304 ) ;
  assign n4306 = ( n4003 & ~n4139 ) | ( n4003 & n4148 ) | ( ~n4139 & n4148 ) ;
  assign n4307 = ( n4139 & ~n4149 ) | ( n4139 & n4306 ) | ( ~n4149 & n4306 ) ;
  assign n4308 = n3800 & ~n3955 ;
  assign n4309 = ~n1338 & n3799 ;
  assign n4310 = n1458 & n3802 ;
  assign n4311 = ( ~n1576 & n3694 ) | ( ~n1576 & n3699 ) | ( n3694 & n3699 ) ;
  assign n4312 = ( n3694 & n4310 ) | ( n3694 & ~n4311 ) | ( n4310 & ~n4311 ) ;
  assign n4313 = ( ~n4308 & n4309 ) | ( ~n4308 & n4312 ) | ( n4309 & n4312 ) ;
  assign n4314 = ( ~x29 & n4308 ) | ( ~x29 & n4313 ) | ( n4308 & n4313 ) ;
  assign n4315 = ( n4308 & n4313 ) | ( n4308 & ~n4314 ) | ( n4313 & ~n4314 ) ;
  assign n4316 = ( x29 & n4314 ) | ( x29 & ~n4315 ) | ( n4314 & ~n4315 ) ;
  assign n4317 = ( ~n4305 & n4307 ) | ( ~n4305 & n4316 ) | ( n4307 & n4316 ) ;
  assign n4318 = ( n3871 & n4148 ) | ( n3871 & ~n4306 ) | ( n4148 & ~n4306 ) ;
  assign n4319 = ( ~n3871 & n4150 ) | ( ~n3871 & n4318 ) | ( n4150 & n4318 ) ;
  assign n4320 = n607 | n1750 ;
  assign n4321 = n1250 & ~n1669 ;
  assign n4322 = ( ~n1750 & n4320 ) | ( ~n1750 & n4321 ) | ( n4320 & n4321 ) ;
  assign n4323 = n606 & ~n1576 ;
  assign n4324 = ( n606 & n4322 ) | ( n606 & ~n4323 ) | ( n4322 & ~n4323 ) ;
  assign n4325 = ( n1576 & n1669 ) | ( n1576 & ~n3613 ) | ( n1669 & ~n3613 ) ;
  assign n4326 = ( ~n1669 & n3614 ) | ( ~n1669 & n4325 ) | ( n3614 & n4325 ) ;
  assign n4327 = n1248 & n4326 ;
  assign n4328 = n4324 | n4327 ;
  assign n4329 = ( n4317 & n4319 ) | ( n4317 & n4328 ) | ( n4319 & n4328 ) ;
  assign n4330 = ( n4150 & ~n4152 ) | ( n4150 & n4161 ) | ( ~n4152 & n4161 ) ;
  assign n4331 = ( ~n4150 & n4162 ) | ( ~n4150 & n4330 ) | ( n4162 & n4330 ) ;
  assign n4332 = ~n3791 & n3800 ;
  assign n4333 = n1267 & n3802 ;
  assign n4334 = ~n1246 & n3799 ;
  assign n4335 = ( n1338 & n3694 ) | ( n1338 & n3699 ) | ( n3694 & n3699 ) ;
  assign n4336 = ( n3694 & n4334 ) | ( n3694 & ~n4335 ) | ( n4334 & ~n4335 ) ;
  assign n4337 = ( ~n4332 & n4333 ) | ( ~n4332 & n4336 ) | ( n4333 & n4336 ) ;
  assign n4338 = ( ~x29 & n4332 ) | ( ~x29 & n4337 ) | ( n4332 & n4337 ) ;
  assign n4339 = ( n4332 & n4337 ) | ( n4332 & ~n4338 ) | ( n4337 & ~n4338 ) ;
  assign n4340 = ( x29 & n4338 ) | ( x29 & ~n4339 ) | ( n4338 & ~n4339 ) ;
  assign n4341 = ( n4329 & n4331 ) | ( n4329 & n4340 ) | ( n4331 & n4340 ) ;
  assign n4342 = ( n4162 & ~n4164 ) | ( n4162 & n4173 ) | ( ~n4164 & n4173 ) ;
  assign n4343 = ( ~n4162 & n4174 ) | ( ~n4162 & n4342 ) | ( n4174 & n4342 ) ;
  assign n4344 = n3797 & n4202 ;
  assign n4345 = ( n65 & n70 ) | ( n65 & ~n4195 ) | ( n70 & ~n4195 ) ;
  assign n4346 = ~n3692 & n4345 ;
  assign n4347 = ~n3658 & n4200 ;
  assign n4348 = n4346 | n4347 ;
  assign n4349 = ( ~x26 & n4344 ) | ( ~x26 & n4348 ) | ( n4344 & n4348 ) ;
  assign n4350 = ( n4344 & n4348 ) | ( n4344 & ~n4349 ) | ( n4348 & ~n4349 ) ;
  assign n4351 = ( x26 & n4349 ) | ( x26 & ~n4350 ) | ( n4349 & ~n4350 ) ;
  assign n4352 = ( n4341 & n4343 ) | ( n4341 & n4351 ) | ( n4343 & n4351 ) ;
  assign n4353 = ~n3779 & n3800 ;
  assign n4354 = n1267 & n3799 ;
  assign n4355 = n1458 & ~n3700 ;
  assign n4356 = ~n1338 & n3802 ;
  assign n4357 = ( n1458 & ~n4355 ) | ( n1458 & n4356 ) | ( ~n4355 & n4356 ) ;
  assign n4358 = ( ~n4353 & n4354 ) | ( ~n4353 & n4357 ) | ( n4354 & n4357 ) ;
  assign n4359 = ( ~x29 & n4353 ) | ( ~x29 & n4358 ) | ( n4353 & n4358 ) ;
  assign n4360 = ( n4353 & n4358 ) | ( n4353 & ~n4359 ) | ( n4358 & ~n4359 ) ;
  assign n4361 = ( x29 & n4359 ) | ( x29 & ~n4360 ) | ( n4359 & ~n4360 ) ;
  assign n4362 = ( ~n4317 & n4319 ) | ( ~n4317 & n4328 ) | ( n4319 & n4328 ) ;
  assign n4363 = ( n4317 & ~n4329 ) | ( n4317 & n4362 ) | ( ~n4329 & n4362 ) ;
  assign n4364 = ~n3665 & n4202 ;
  assign n4365 = ~n1290 & n4345 ;
  assign n4366 = n1246 & n4200 ;
  assign n4367 = ~n3658 & n4201 ;
  assign n4368 = ( n4200 & ~n4366 ) | ( n4200 & n4367 ) | ( ~n4366 & n4367 ) ;
  assign n4369 = ( ~n4364 & n4365 ) | ( ~n4364 & n4368 ) | ( n4365 & n4368 ) ;
  assign n4370 = ( ~x26 & n4364 ) | ( ~x26 & n4369 ) | ( n4364 & n4369 ) ;
  assign n4371 = ( n4364 & n4369 ) | ( n4364 & ~n4370 ) | ( n4369 & ~n4370 ) ;
  assign n4372 = ( x26 & n4370 ) | ( x26 & ~n4371 ) | ( n4370 & ~n4371 ) ;
  assign n4373 = ( n4361 & n4363 ) | ( n4361 & n4372 ) | ( n4363 & n4372 ) ;
  assign n4374 = ~n4182 & n4202 ;
  assign n4375 = ~n1290 & n4200 ;
  assign n4376 = ~n3692 & n4201 ;
  assign n4377 = ~n3658 & n4345 ;
  assign n4378 = n4376 | n4377 ;
  assign n4379 = ( ~n4374 & n4375 ) | ( ~n4374 & n4378 ) | ( n4375 & n4378 ) ;
  assign n4380 = ( ~x26 & n4374 ) | ( ~x26 & n4379 ) | ( n4374 & n4379 ) ;
  assign n4381 = ( n4374 & n4379 ) | ( n4374 & ~n4380 ) | ( n4379 & ~n4380 ) ;
  assign n4382 = ( x26 & n4380 ) | ( x26 & ~n4381 ) | ( n4380 & ~n4381 ) ;
  assign n4383 = ( n4329 & ~n4331 ) | ( n4329 & n4340 ) | ( ~n4331 & n4340 ) ;
  assign n4384 = ( n4331 & ~n4341 ) | ( n4331 & n4383 ) | ( ~n4341 & n4383 ) ;
  assign n4385 = ( n4373 & n4382 ) | ( n4373 & n4384 ) | ( n4382 & n4384 ) ;
  assign n4386 = n1009 | n2071 ;
  assign n4387 = n263 | n1695 ;
  assign n4388 = n81 | n338 ;
  assign n4389 = n259 | n1068 ;
  assign n4390 = ( n66 & n97 ) | ( n66 & n119 ) | ( n97 & n119 ) ;
  assign n4391 = n4389 | n4390 ;
  assign n4392 = ( n389 & ~n4388 ) | ( n389 & n4391 ) | ( ~n4388 & n4391 ) ;
  assign n4393 = n4388 | n4392 ;
  assign n4394 = ( ~n4386 & n4387 ) | ( ~n4386 & n4393 ) | ( n4387 & n4393 ) ;
  assign n4395 = n4386 | n4394 ;
  assign n4396 = n1623 | n3135 ;
  assign n4397 = n320 | n922 ;
  assign n4398 = ( ~n648 & n1131 ) | ( ~n648 & n2612 ) | ( n1131 & n2612 ) ;
  assign n4399 = ( n648 & ~n4397 ) | ( n648 & n4398 ) | ( ~n4397 & n4398 ) ;
  assign n4400 = n4397 | n4399 ;
  assign n4401 = ( ~n4395 & n4396 ) | ( ~n4395 & n4400 ) | ( n4396 & n4400 ) ;
  assign n4402 = n4395 | n4401 ;
  assign n4403 = n250 & ~n1188 ;
  assign n4404 = ( ~n3338 & n4402 ) | ( ~n3338 & n4403 ) | ( n4402 & n4403 ) ;
  assign n4405 = ~n4402 & n4404 ;
  assign n4406 = n117 | n523 ;
  assign n4407 = ( n299 & n1068 ) | ( n299 & ~n4406 ) | ( n1068 & ~n4406 ) ;
  assign n4408 = n4406 | n4407 ;
  assign n4409 = n262 | n293 ;
  assign n4410 = n2765 | n4409 ;
  assign n4411 = ( n41 & n44 ) | ( n41 & n98 ) | ( n44 & n98 ) ;
  assign n4412 = n963 | n4411 ;
  assign n4413 = n1700 | n4412 ;
  assign n4414 = ( ~n4408 & n4410 ) | ( ~n4408 & n4413 ) | ( n4410 & n4413 ) ;
  assign n4415 = n4408 | n4414 ;
  assign n4416 = n1974 | n2355 ;
  assign n4417 = n2671 | n4223 ;
  assign n4418 = n746 | n878 ;
  assign n4419 = n395 | n2181 ;
  assign n4420 = n4034 | n4419 ;
  assign n4421 = ( ~n4417 & n4418 ) | ( ~n4417 & n4420 ) | ( n4418 & n4420 ) ;
  assign n4422 = n4417 | n4421 ;
  assign n4423 = n144 | n444 ;
  assign n4424 = ( n230 & n890 ) | ( n230 & ~n4423 ) | ( n890 & ~n4423 ) ;
  assign n4425 = n4423 | n4424 ;
  assign n4426 = n435 | n922 ;
  assign n4427 = ( n2205 & ~n4425 ) | ( n2205 & n4426 ) | ( ~n4425 & n4426 ) ;
  assign n4428 = n4425 | n4427 ;
  assign n4429 = ( ~n4416 & n4422 ) | ( ~n4416 & n4428 ) | ( n4422 & n4428 ) ;
  assign n4430 = n4416 | n4429 ;
  assign n4431 = ( n320 & n529 ) | ( n320 & ~n551 ) | ( n529 & ~n551 ) ;
  assign n4432 = n551 | n4431 ;
  assign n4433 = ( n194 & n1315 ) | ( n194 & ~n4432 ) | ( n1315 & ~n4432 ) ;
  assign n4434 = n4432 | n4433 ;
  assign n4435 = n204 | n290 ;
  assign n4436 = n661 | n4435 ;
  assign n4437 = ( n4430 & ~n4434 ) | ( n4430 & n4436 ) | ( ~n4434 & n4436 ) ;
  assign n4438 = ( n154 & n4434 ) | ( n154 & ~n4437 ) | ( n4434 & ~n4437 ) ;
  assign n4439 = n4437 | n4438 ;
  assign n4440 = n1506 | n4439 ;
  assign n4441 = n778 | n2553 ;
  assign n4442 = n1057 | n1595 ;
  assign n4443 = ( n2256 & n2429 ) | ( n2256 & ~n4442 ) | ( n2429 & ~n4442 ) ;
  assign n4444 = n4442 | n4443 ;
  assign n4445 = ( ~n107 & n4441 ) | ( ~n107 & n4444 ) | ( n4441 & n4444 ) ;
  assign n4446 = ( n107 & n3162 ) | ( n107 & ~n4445 ) | ( n3162 & ~n4445 ) ;
  assign n4447 = n4445 | n4446 ;
  assign n4448 = ( ~n4415 & n4440 ) | ( ~n4415 & n4447 ) | ( n4440 & n4447 ) ;
  assign n4449 = n4415 | n4448 ;
  assign n4450 = ( x17 & n4405 ) | ( x17 & ~n4449 ) | ( n4405 & ~n4449 ) ;
  assign n4451 = n1250 & ~n2023 ;
  assign n4452 = n607 & n2089 ;
  assign n4453 = n4451 | n4452 ;
  assign n4454 = n606 & ~n1926 ;
  assign n4455 = ( n606 & n4453 ) | ( n606 & ~n4454 ) | ( n4453 & ~n4454 ) ;
  assign n4456 = ( ~n1926 & n2023 ) | ( ~n1926 & n3609 ) | ( n2023 & n3609 ) ;
  assign n4457 = ( ~n3609 & n3610 ) | ( ~n3609 & n4456 ) | ( n3610 & n4456 ) ;
  assign n4458 = n1248 & ~n4457 ;
  assign n4459 = n4455 | n4458 ;
  assign n4460 = ( n4057 & n4450 ) | ( n4057 & ~n4459 ) | ( n4450 & ~n4459 ) ;
  assign n4461 = ( n196 & n595 ) | ( n196 & ~n1695 ) | ( n595 & ~n1695 ) ;
  assign n4462 = n1695 | n4461 ;
  assign n4463 = ( n98 & n100 ) | ( n98 & n109 ) | ( n100 & n109 ) ;
  assign n4464 = ( n1060 & ~n4462 ) | ( n1060 & n4463 ) | ( ~n4462 & n4463 ) ;
  assign n4465 = n4462 | n4464 ;
  assign n4466 = n163 | n176 ;
  assign n4467 = n1865 | n2146 ;
  assign n4468 = n4466 | n4467 ;
  assign n4469 = n807 | n2256 ;
  assign n4470 = n3552 | n4469 ;
  assign n4471 = ( ~n4465 & n4468 ) | ( ~n4465 & n4470 ) | ( n4468 & n4470 ) ;
  assign n4472 = n4465 | n4471 ;
  assign n4473 = ( n961 & n2001 ) | ( n961 & ~n2163 ) | ( n2001 & ~n2163 ) ;
  assign n4474 = n2163 | n4473 ;
  assign n4475 = n91 | n1430 ;
  assign n4476 = ( n3302 & ~n4474 ) | ( n3302 & n4475 ) | ( ~n4474 & n4475 ) ;
  assign n4477 = n4474 | n4476 ;
  assign n4478 = n195 | n865 ;
  assign n4479 = ( n144 & n193 ) | ( n144 & ~n1314 ) | ( n193 & ~n1314 ) ;
  assign n4480 = n1314 | n4479 ;
  assign n4481 = ( n653 & ~n4478 ) | ( n653 & n4480 ) | ( ~n4478 & n4480 ) ;
  assign n4482 = n4478 | n4481 ;
  assign n4483 = ( n2895 & n3485 ) | ( n2895 & ~n4482 ) | ( n3485 & ~n4482 ) ;
  assign n4484 = n4482 | n4483 ;
  assign n4485 = ( ~n4472 & n4477 ) | ( ~n4472 & n4484 ) | ( n4477 & n4484 ) ;
  assign n4486 = n4472 | n4485 ;
  assign n4487 = ( ~n301 & n534 ) | ( ~n301 & n591 ) | ( n534 & n591 ) ;
  assign n4488 = n301 | n4487 ;
  assign n4489 = n105 | n3162 ;
  assign n4490 = n188 | n876 ;
  assign n4491 = n753 | n4490 ;
  assign n4492 = ( ~n4488 & n4489 ) | ( ~n4488 & n4491 ) | ( n4489 & n4491 ) ;
  assign n4493 = n4488 | n4492 ;
  assign n4494 = n192 | n285 ;
  assign n4495 = n356 | n895 ;
  assign n4496 = ( ~n159 & n4028 ) | ( ~n159 & n4495 ) | ( n4028 & n4495 ) ;
  assign n4497 = ( n159 & ~n4494 ) | ( n159 & n4496 ) | ( ~n4494 & n4496 ) ;
  assign n4498 = n4494 | n4497 ;
  assign n4499 = n101 | n435 ;
  assign n4500 = ( n1169 & n1365 ) | ( n1169 & ~n4499 ) | ( n1365 & ~n4499 ) ;
  assign n4501 = n4499 | n4500 ;
  assign n4502 = ( n83 & n97 ) | ( n83 & n145 ) | ( n97 & n145 ) ;
  assign n4503 = n1477 | n4502 ;
  assign n4504 = n3063 | n4503 ;
  assign n4505 = ( n376 & n1315 ) | ( n376 & ~n4503 ) | ( n1315 & ~n4503 ) ;
  assign n4506 = ( ~n4501 & n4504 ) | ( ~n4501 & n4505 ) | ( n4504 & n4505 ) ;
  assign n4507 = n4501 | n4506 ;
  assign n4508 = ( n4493 & ~n4498 ) | ( n4493 & n4507 ) | ( ~n4498 & n4507 ) ;
  assign n4509 = n67 | n786 ;
  assign n4510 = n550 | n4509 ;
  assign n4511 = n1143 | n4510 ;
  assign n4512 = ( n75 & ~n78 ) | ( n75 & n116 ) | ( ~n78 & n116 ) ;
  assign n4513 = ( n242 & n600 ) | ( n242 & ~n4512 ) | ( n600 & ~n4512 ) ;
  assign n4514 = n4512 | n4513 ;
  assign n4515 = n1044 | n1171 ;
  assign n4516 = ( ~n545 & n1008 ) | ( ~n545 & n4515 ) | ( n1008 & n4515 ) ;
  assign n4517 = ( n317 & n545 ) | ( n317 & ~n4516 ) | ( n545 & ~n4516 ) ;
  assign n4518 = n4516 | n4517 ;
  assign n4519 = ( ~n1573 & n3464 ) | ( ~n1573 & n4518 ) | ( n3464 & n4518 ) ;
  assign n4520 = ( n1573 & ~n4514 ) | ( n1573 & n4519 ) | ( ~n4514 & n4519 ) ;
  assign n4521 = n4514 | n4520 ;
  assign n4522 = ( n55 & n1225 ) | ( n55 & ~n2323 ) | ( n1225 & ~n2323 ) ;
  assign n4523 = n2323 | n4522 ;
  assign n4524 = ( ~n4511 & n4521 ) | ( ~n4511 & n4523 ) | ( n4521 & n4523 ) ;
  assign n4525 = n4511 | n4524 ;
  assign n4526 = n1418 | n1489 ;
  assign n4527 = n112 | n261 ;
  assign n4528 = ( n168 & n642 ) | ( n168 & ~n4527 ) | ( n642 & ~n4527 ) ;
  assign n4529 = n4527 | n4528 ;
  assign n4530 = n212 | n1231 ;
  assign n4531 = ( n100 & n152 ) | ( n100 & n240 ) | ( n152 & n240 ) ;
  assign n4532 = ( n174 & n523 ) | ( n174 & ~n4531 ) | ( n523 & ~n4531 ) ;
  assign n4533 = n4531 | n4532 ;
  assign n4534 = ( ~n4529 & n4530 ) | ( ~n4529 & n4533 ) | ( n4530 & n4533 ) ;
  assign n4535 = n4529 | n4534 ;
  assign n4536 = ( n2576 & ~n4526 ) | ( n2576 & n4535 ) | ( ~n4526 & n4535 ) ;
  assign n4537 = n4526 | n4536 ;
  assign n4538 = ( ~n4498 & n4525 ) | ( ~n4498 & n4537 ) | ( n4525 & n4537 ) ;
  assign n4539 = n4498 | n4538 ;
  assign n4540 = ( ~n4486 & n4508 ) | ( ~n4486 & n4539 ) | ( n4508 & n4539 ) ;
  assign n4541 = n4486 | n4540 ;
  assign n4542 = n512 | n638 ;
  assign n4543 = n104 | n233 ;
  assign n4544 = ( ~n188 & n254 ) | ( ~n188 & n320 ) | ( n254 & n320 ) ;
  assign n4545 = n188 | n4544 ;
  assign n4546 = ( ~n4542 & n4543 ) | ( ~n4542 & n4545 ) | ( n4543 & n4545 ) ;
  assign n4547 = n4542 | n4546 ;
  assign n4548 = n523 | n1122 ;
  assign n4549 = ( n1878 & ~n4235 ) | ( n1878 & n4548 ) | ( ~n4235 & n4548 ) ;
  assign n4550 = n4235 | n4549 ;
  assign n4551 = n550 | n1110 ;
  assign n4552 = n773 | n1928 ;
  assign n4553 = n4551 | n4552 ;
  assign n4554 = ( n83 & n129 ) | ( n83 & n149 ) | ( n129 & n149 ) ;
  assign n4555 = ( n3194 & ~n4553 ) | ( n3194 & n4554 ) | ( ~n4553 & n4554 ) ;
  assign n4556 = n4553 | n4555 ;
  assign n4557 = ( ~n4547 & n4550 ) | ( ~n4547 & n4556 ) | ( n4550 & n4556 ) ;
  assign n4558 = n4547 | n4557 ;
  assign n4559 = n3128 | n3569 ;
  assign n4560 = ( n75 & n97 ) | ( n75 & n102 ) | ( n97 & n102 ) ;
  assign n4561 = n337 | n4560 ;
  assign n4562 = ( n1421 & n2073 ) | ( n1421 & ~n4561 ) | ( n2073 & ~n4561 ) ;
  assign n4563 = n4561 | n4562 ;
  assign n4564 = ( n4412 & ~n4559 ) | ( n4412 & n4563 ) | ( ~n4559 & n4563 ) ;
  assign n4565 = ( n957 & n4559 ) | ( n957 & ~n4564 ) | ( n4559 & ~n4564 ) ;
  assign n4566 = n4564 | n4565 ;
  assign n4567 = ( n60 & n299 ) | ( n60 & ~n789 ) | ( n299 & ~n789 ) ;
  assign n4568 = n789 | n4567 ;
  assign n4569 = ( n72 & n97 ) | ( n72 & n145 ) | ( n97 & n145 ) ;
  assign n4570 = ( n1132 & n2361 ) | ( n1132 & ~n4569 ) | ( n2361 & ~n4569 ) ;
  assign n4571 = n4569 | n4570 ;
  assign n4572 = n137 | n267 ;
  assign n4573 = ( n195 & n215 ) | ( n195 & ~n4572 ) | ( n215 & ~n4572 ) ;
  assign n4574 = n4572 | n4573 ;
  assign n4575 = ( ~n4568 & n4571 ) | ( ~n4568 & n4574 ) | ( n4571 & n4574 ) ;
  assign n4576 = ( n64 & n145 ) | ( n64 & n234 ) | ( n145 & n234 ) ;
  assign n4577 = n3351 | n4576 ;
  assign n4578 = ( n1304 & ~n4568 ) | ( n1304 & n4577 ) | ( ~n4568 & n4577 ) ;
  assign n4579 = n4568 | n4578 ;
  assign n4580 = ( ~n4566 & n4575 ) | ( ~n4566 & n4579 ) | ( n4575 & n4579 ) ;
  assign n4581 = n4566 | n4580 ;
  assign n4582 = n1220 | n1400 ;
  assign n4583 = n913 | n4582 ;
  assign n4584 = n2787 | n2954 ;
  assign n4585 = n189 | n537 ;
  assign n4586 = n117 | n4585 ;
  assign n4587 = ( ~n4582 & n4584 ) | ( ~n4582 & n4586 ) | ( n4584 & n4586 ) ;
  assign n4588 = n292 | n2380 ;
  assign n4589 = ( n134 & ~n2128 ) | ( n134 & n4588 ) | ( ~n2128 & n4588 ) ;
  assign n4590 = n2128 | n4589 ;
  assign n4591 = ( ~n4583 & n4587 ) | ( ~n4583 & n4590 ) | ( n4587 & n4590 ) ;
  assign n4592 = n4583 | n4591 ;
  assign n4593 = ( ~n4558 & n4581 ) | ( ~n4558 & n4592 ) | ( n4581 & n4592 ) ;
  assign n4594 = ( n59 & n84 ) | ( n59 & n149 ) | ( n84 & n149 ) ;
  assign n4595 = n888 | n4594 ;
  assign n4596 = ( n1864 & n2648 ) | ( n1864 & ~n4595 ) | ( n2648 & ~n4595 ) ;
  assign n4597 = n4595 | n4596 ;
  assign n4598 = n316 | n609 ;
  assign n4599 = ( n2053 & ~n2185 ) | ( n2053 & n4598 ) | ( ~n2185 & n4598 ) ;
  assign n4600 = n3214 | n4599 ;
  assign n4601 = n239 | n1031 ;
  assign n4602 = ~n1057 & n3962 ;
  assign n4603 = ~n4601 & n4602 ;
  assign n4604 = ( ~n2185 & n4600 ) | ( ~n2185 & n4603 ) | ( n4600 & n4603 ) ;
  assign n4605 = ~n4600 & n4604 ;
  assign n4606 = ( n4592 & ~n4597 ) | ( n4592 & n4605 ) | ( ~n4597 & n4605 ) ;
  assign n4607 = ( n4558 & ~n4593 ) | ( n4558 & n4606 ) | ( ~n4593 & n4606 ) ;
  assign n4608 = ~n4558 & n4607 ;
  assign n4609 = ( x14 & ~n4541 ) | ( x14 & n4608 ) | ( ~n4541 & n4608 ) ;
  assign n4610 = n215 | n519 ;
  assign n4611 = n186 | n4610 ;
  assign n4612 = ( n48 & n66 ) | ( n48 & n75 ) | ( n66 & n75 ) ;
  assign n4613 = n933 | n4612 ;
  assign n4614 = n2310 | n4613 ;
  assign n4615 = n4611 | n4614 ;
  assign n4616 = n1837 | n3233 ;
  assign n4617 = n731 | n4616 ;
  assign n4618 = n523 | n613 ;
  assign n4619 = n2798 | n3104 ;
  assign n4620 = ( n889 & ~n4618 ) | ( n889 & n4619 ) | ( ~n4618 & n4619 ) ;
  assign n4621 = n4618 | n4620 ;
  assign n4622 = ( n3491 & ~n4616 ) | ( n3491 & n4621 ) | ( ~n4616 & n4621 ) ;
  assign n4623 = ( ~n4615 & n4617 ) | ( ~n4615 & n4622 ) | ( n4617 & n4622 ) ;
  assign n4624 = n4615 | n4623 ;
  assign n4625 = n1155 | n4624 ;
  assign n4626 = n55 | n512 ;
  assign n4627 = ( n356 & n795 ) | ( n356 & ~n4626 ) | ( n795 & ~n4626 ) ;
  assign n4628 = n4626 | n4627 ;
  assign n4629 = n529 | n642 ;
  assign n4630 = ( n131 & n173 ) | ( n131 & ~n4629 ) | ( n173 & ~n4629 ) ;
  assign n4631 = n4629 | n4630 ;
  assign n4632 = ( n4577 & n4628 ) | ( n4577 & ~n4631 ) | ( n4628 & ~n4631 ) ;
  assign n4633 = n656 | n959 ;
  assign n4634 = n376 | n3637 ;
  assign n4635 = ( n2956 & ~n4633 ) | ( n2956 & n4634 ) | ( ~n4633 & n4634 ) ;
  assign n4636 = n4633 | n4635 ;
  assign n4637 = ( n4631 & ~n4632 ) | ( n4631 & n4636 ) | ( ~n4632 & n4636 ) ;
  assign n4638 = n4632 | n4637 ;
  assign n4639 = ( n4477 & ~n4625 ) | ( n4477 & n4638 ) | ( ~n4625 & n4638 ) ;
  assign n4640 = n4625 | n4639 ;
  assign n4641 = n607 | n2298 ;
  assign n4642 = n1250 & n2270 ;
  assign n4643 = ( ~n2298 & n4641 ) | ( ~n2298 & n4642 ) | ( n4641 & n4642 ) ;
  assign n4644 = n606 & ~n2174 ;
  assign n4645 = ( n606 & n4643 ) | ( n606 & ~n4644 ) | ( n4643 & ~n4644 ) ;
  assign n4646 = ( n2174 & ~n2270 ) | ( n2174 & n3606 ) | ( ~n2270 & n3606 ) ;
  assign n4647 = ( n2270 & ~n3607 ) | ( n2270 & n4646 ) | ( ~n3607 & n4646 ) ;
  assign n4648 = n1248 & n4647 ;
  assign n4649 = n4645 | n4648 ;
  assign n4650 = ( n4609 & n4640 ) | ( n4609 & n4649 ) | ( n4640 & n4649 ) ;
  assign n4651 = ( n4405 & ~n4609 ) | ( n4405 & n4650 ) | ( ~n4609 & n4650 ) ;
  assign n4652 = ( x17 & ~n4405 ) | ( x17 & n4449 ) | ( ~n4405 & n4449 ) ;
  assign n4653 = ( ~x17 & n4450 ) | ( ~x17 & n4652 ) | ( n4450 & n4652 ) ;
  assign n4654 = ~n607 & n2174 ;
  assign n4655 = n1250 & n2089 ;
  assign n4656 = ( n2174 & ~n4654 ) | ( n2174 & n4655 ) | ( ~n4654 & n4655 ) ;
  assign n4657 = n606 & n2023 ;
  assign n4658 = ( n606 & n4656 ) | ( n606 & ~n4657 ) | ( n4656 & ~n4657 ) ;
  assign n4659 = ( n2023 & ~n2089 ) | ( n2023 & n3608 ) | ( ~n2089 & n3608 ) ;
  assign n4660 = ( ~n3608 & n3609 ) | ( ~n3608 & n4659 ) | ( n3609 & n4659 ) ;
  assign n4661 = n1248 & ~n4660 ;
  assign n4662 = n4658 | n4661 ;
  assign n4663 = ( n4651 & n4653 ) | ( n4651 & n4662 ) | ( n4653 & n4662 ) ;
  assign n4664 = ( n4057 & n4450 ) | ( n4057 & n4459 ) | ( n4450 & n4459 ) ;
  assign n4665 = ( n4459 & n4460 ) | ( n4459 & ~n4664 ) | ( n4460 & ~n4664 ) ;
  assign n4666 = n3800 & n4146 ;
  assign n4667 = ~n1669 & n3799 ;
  assign n4668 = n1852 & ~n3700 ;
  assign n4669 = ~n1750 & n3802 ;
  assign n4670 = ( n1852 & ~n4668 ) | ( n1852 & n4669 ) | ( ~n4668 & n4669 ) ;
  assign n4671 = ( ~n4666 & n4667 ) | ( ~n4666 & n4670 ) | ( n4667 & n4670 ) ;
  assign n4672 = ( ~x29 & n4666 ) | ( ~x29 & n4671 ) | ( n4666 & n4671 ) ;
  assign n4673 = ( n4666 & n4671 ) | ( n4666 & ~n4672 ) | ( n4671 & ~n4672 ) ;
  assign n4674 = ( x29 & n4672 ) | ( x29 & ~n4673 ) | ( n4672 & ~n4673 ) ;
  assign n4675 = ( n4663 & n4665 ) | ( n4663 & n4674 ) | ( n4665 & n4674 ) ;
  assign n4676 = ( n4057 & ~n4283 ) | ( n4057 & n4292 ) | ( ~n4283 & n4292 ) ;
  assign n4677 = ( ~n4057 & n4293 ) | ( ~n4057 & n4676 ) | ( n4293 & n4676 ) ;
  assign n4678 = ( ~n4460 & n4675 ) | ( ~n4460 & n4677 ) | ( n4675 & n4677 ) ;
  assign n4679 = n3800 & ~n4159 ;
  assign n4680 = n1458 & n3799 ;
  assign n4681 = ~n1669 & n3700 ;
  assign n4682 = n1576 & n3802 ;
  assign n4683 = n4681 | n4682 ;
  assign n4684 = ( ~n4679 & n4680 ) | ( ~n4679 & n4683 ) | ( n4680 & n4683 ) ;
  assign n4685 = ( ~x29 & n4679 ) | ( ~x29 & n4684 ) | ( n4679 & n4684 ) ;
  assign n4686 = ( n4679 & n4684 ) | ( n4679 & ~n4685 ) | ( n4684 & ~n4685 ) ;
  assign n4687 = ( x29 & n4685 ) | ( x29 & ~n4686 ) | ( n4685 & ~n4686 ) ;
  assign n4688 = ( n4293 & ~n4295 ) | ( n4293 & n4304 ) | ( ~n4295 & n4304 ) ;
  assign n4689 = ( ~n4293 & n4305 ) | ( ~n4293 & n4688 ) | ( n4305 & n4688 ) ;
  assign n4690 = ( n4678 & n4687 ) | ( n4678 & n4689 ) | ( n4687 & n4689 ) ;
  assign n4691 = ( n4307 & n4316 ) | ( n4307 & ~n4317 ) | ( n4316 & ~n4317 ) ;
  assign n4692 = ( n4305 & n4317 ) | ( n4305 & ~n4691 ) | ( n4317 & ~n4691 ) ;
  assign n4693 = n3621 & n4202 ;
  assign n4694 = ~n1290 & n4201 ;
  assign n4695 = ~n1246 & n4345 ;
  assign n4696 = n1267 & n4200 ;
  assign n4697 = n4695 | n4696 ;
  assign n4698 = ( ~n4693 & n4694 ) | ( ~n4693 & n4697 ) | ( n4694 & n4697 ) ;
  assign n4699 = ( ~x26 & n4693 ) | ( ~x26 & n4698 ) | ( n4693 & n4698 ) ;
  assign n4700 = ( n4693 & n4698 ) | ( n4693 & ~n4699 ) | ( n4698 & ~n4699 ) ;
  assign n4701 = ( x26 & n4699 ) | ( x26 & ~n4700 ) | ( n4699 & ~n4700 ) ;
  assign n4702 = ( n4690 & ~n4692 ) | ( n4690 & n4701 ) | ( ~n4692 & n4701 ) ;
  assign n4703 = x20 | x21 ;
  assign n4704 = x21 & x22 ;
  assign n4705 = x22 | x23 ;
  assign n4706 = x22 & x23 ;
  assign n4707 = n4705 & ~n4706 ;
  assign n4708 = ( x20 & ~x22 ) | ( x20 & n4707 ) | ( ~x22 & n4707 ) ;
  assign n4709 = ( ~n4703 & n4704 ) | ( ~n4703 & n4708 ) | ( n4704 & n4708 ) ;
  assign n4710 = x20 & x21 ;
  assign n4711 = n4703 & ~n4710 ;
  assign n4712 = ( ~n4705 & n4706 ) | ( ~n4705 & n4711 ) | ( n4706 & n4711 ) ;
  assign n4713 = n4711 & ~n4712 ;
  assign n4714 = ~n3691 & n4713 ;
  assign n4715 = ( ~n3692 & n4709 ) | ( ~n3692 & n4714 ) | ( n4709 & n4714 ) ;
  assign n4716 = x23 | n4715 ;
  assign n4717 = ( x23 & n4715 ) | ( x23 & ~n4716 ) | ( n4715 & ~n4716 ) ;
  assign n4718 = n4716 & ~n4717 ;
  assign n4719 = ( n4361 & ~n4363 ) | ( n4361 & n4372 ) | ( ~n4363 & n4372 ) ;
  assign n4720 = ( n4363 & ~n4373 ) | ( n4363 & n4719 ) | ( ~n4373 & n4719 ) ;
  assign n4721 = ( n4702 & n4718 ) | ( n4702 & n4720 ) | ( n4718 & n4720 ) ;
  assign n4722 = ( n4405 & n4650 ) | ( n4405 & ~n4651 ) | ( n4650 & ~n4651 ) ;
  assign n4723 = ( n4609 & n4651 ) | ( n4609 & ~n4722 ) | ( n4651 & ~n4722 ) ;
  assign n4724 = ~n607 & n2270 ;
  assign n4725 = n1250 & n2174 ;
  assign n4726 = ( n2270 & ~n4724 ) | ( n2270 & n4725 ) | ( ~n4724 & n4725 ) ;
  assign n4727 = n606 & ~n2089 ;
  assign n4728 = ( n606 & n4726 ) | ( n606 & ~n4727 ) | ( n4726 & ~n4727 ) ;
  assign n4729 = ( n2089 & ~n2174 ) | ( n2089 & n3607 ) | ( ~n2174 & n3607 ) ;
  assign n4730 = ( n2174 & ~n3608 ) | ( n2174 & n4729 ) | ( ~n3608 & n4729 ) ;
  assign n4731 = n1248 & n4730 ;
  assign n4732 = n4728 | n4731 ;
  assign n4733 = n3800 & n4290 ;
  assign n4734 = n1852 & n3799 ;
  assign n4735 = ~n2023 & n3700 ;
  assign n4736 = n1926 & n3802 ;
  assign n4737 = n4735 | n4736 ;
  assign n4738 = ( ~n4733 & n4734 ) | ( ~n4733 & n4737 ) | ( n4734 & n4737 ) ;
  assign n4739 = ( ~x29 & n4733 ) | ( ~x29 & n4738 ) | ( n4733 & n4738 ) ;
  assign n4740 = ( n4733 & n4738 ) | ( n4733 & ~n4739 ) | ( n4738 & ~n4739 ) ;
  assign n4741 = ( x29 & n4739 ) | ( x29 & ~n4740 ) | ( n4739 & ~n4740 ) ;
  assign n4742 = ( ~n4723 & n4732 ) | ( ~n4723 & n4741 ) | ( n4732 & n4741 ) ;
  assign n4743 = ( n4651 & ~n4653 ) | ( n4651 & n4662 ) | ( ~n4653 & n4662 ) ;
  assign n4744 = ( n4653 & ~n4663 ) | ( n4653 & n4743 ) | ( ~n4663 & n4743 ) ;
  assign n4745 = n3800 & ~n4302 ;
  assign n4746 = ~n1750 & n3799 ;
  assign n4747 = n1852 & n3802 ;
  assign n4748 = ( ~n1926 & n3694 ) | ( ~n1926 & n3699 ) | ( n3694 & n3699 ) ;
  assign n4749 = ( n3694 & n4747 ) | ( n3694 & ~n4748 ) | ( n4747 & ~n4748 ) ;
  assign n4750 = ( ~n4745 & n4746 ) | ( ~n4745 & n4749 ) | ( n4746 & n4749 ) ;
  assign n4751 = ( ~x29 & n4745 ) | ( ~x29 & n4750 ) | ( n4745 & n4750 ) ;
  assign n4752 = ( n4745 & n4750 ) | ( n4745 & ~n4751 ) | ( n4750 & ~n4751 ) ;
  assign n4753 = ( x29 & n4751 ) | ( x29 & ~n4752 ) | ( n4751 & ~n4752 ) ;
  assign n4754 = ( n4742 & n4744 ) | ( n4742 & n4753 ) | ( n4744 & n4753 ) ;
  assign n4755 = ( n4663 & ~n4665 ) | ( n4663 & n4674 ) | ( ~n4665 & n4674 ) ;
  assign n4756 = ( n4665 & ~n4675 ) | ( n4665 & n4755 ) | ( ~n4675 & n4755 ) ;
  assign n4757 = ~n3955 & n4202 ;
  assign n4758 = ~n1338 & n4201 ;
  assign n4759 = n1458 & n4345 ;
  assign n4760 = n1576 & n4200 ;
  assign n4761 = n4759 | n4760 ;
  assign n4762 = ( ~n4757 & n4758 ) | ( ~n4757 & n4761 ) | ( n4758 & n4761 ) ;
  assign n4763 = ( ~x26 & n4757 ) | ( ~x26 & n4762 ) | ( n4757 & n4762 ) ;
  assign n4764 = ( n4757 & n4762 ) | ( n4757 & ~n4763 ) | ( n4762 & ~n4763 ) ;
  assign n4765 = ( x26 & n4763 ) | ( x26 & ~n4764 ) | ( n4763 & ~n4764 ) ;
  assign n4766 = ( n4754 & n4756 ) | ( n4754 & n4765 ) | ( n4756 & n4765 ) ;
  assign n4767 = ( n4675 & n4677 ) | ( n4675 & ~n4678 ) | ( n4677 & ~n4678 ) ;
  assign n4768 = ( n4460 & n4678 ) | ( n4460 & ~n4767 ) | ( n4678 & ~n4767 ) ;
  assign n4769 = n3800 & n4326 ;
  assign n4770 = n1576 & n3799 ;
  assign n4771 = n1750 | n3700 ;
  assign n4772 = ~n1669 & n3802 ;
  assign n4773 = ( ~n1750 & n4771 ) | ( ~n1750 & n4772 ) | ( n4771 & n4772 ) ;
  assign n4774 = ( ~n4769 & n4770 ) | ( ~n4769 & n4773 ) | ( n4770 & n4773 ) ;
  assign n4775 = ( ~x29 & n4769 ) | ( ~x29 & n4774 ) | ( n4769 & n4774 ) ;
  assign n4776 = ( n4769 & n4774 ) | ( n4769 & ~n4775 ) | ( n4774 & ~n4775 ) ;
  assign n4777 = ( x29 & n4775 ) | ( x29 & ~n4776 ) | ( n4775 & ~n4776 ) ;
  assign n4778 = ~n3779 & n4202 ;
  assign n4779 = n1267 & n4201 ;
  assign n4780 = n1458 & ~n4200 ;
  assign n4781 = ~n1338 & n4345 ;
  assign n4782 = ( n1458 & ~n4780 ) | ( n1458 & n4781 ) | ( ~n4780 & n4781 ) ;
  assign n4783 = ( ~n4778 & n4779 ) | ( ~n4778 & n4782 ) | ( n4779 & n4782 ) ;
  assign n4784 = ( ~x26 & n4778 ) | ( ~x26 & n4783 ) | ( n4778 & n4783 ) ;
  assign n4785 = ( n4778 & n4783 ) | ( n4778 & ~n4784 ) | ( n4783 & ~n4784 ) ;
  assign n4786 = ( x26 & n4784 ) | ( x26 & ~n4785 ) | ( n4784 & ~n4785 ) ;
  assign n4787 = ( ~n4768 & n4777 ) | ( ~n4768 & n4786 ) | ( n4777 & n4786 ) ;
  assign n4788 = ( n4777 & n4786 ) | ( n4777 & ~n4787 ) | ( n4786 & ~n4787 ) ;
  assign n4789 = ( n4768 & n4787 ) | ( n4768 & ~n4788 ) | ( n4787 & ~n4788 ) ;
  assign n4790 = ~n3665 & n4713 ;
  assign n4791 = ~x20 & x22 ;
  assign n4792 = ( ~n4704 & n4710 ) | ( ~n4704 & n4791 ) | ( n4710 & n4791 ) ;
  assign n4793 = ~n1290 & n4792 ;
  assign n4794 = ~n1246 & n4709 ;
  assign n4795 = ~n3658 & n4712 ;
  assign n4796 = n4794 | n4795 ;
  assign n4797 = ( ~n4790 & n4793 ) | ( ~n4790 & n4796 ) | ( n4793 & n4796 ) ;
  assign n4798 = ( ~x23 & n4790 ) | ( ~x23 & n4797 ) | ( n4790 & n4797 ) ;
  assign n4799 = ( n4790 & n4797 ) | ( n4790 & ~n4798 ) | ( n4797 & ~n4798 ) ;
  assign n4800 = ( x23 & n4798 ) | ( x23 & ~n4799 ) | ( n4798 & ~n4799 ) ;
  assign n4801 = ( n4766 & ~n4789 ) | ( n4766 & n4800 ) | ( ~n4789 & n4800 ) ;
  assign n4802 = n3692 & n4712 ;
  assign n4803 = ~n3658 & n4792 ;
  assign n4804 = ( n4712 & ~n4802 ) | ( n4712 & n4803 ) | ( ~n4802 & n4803 ) ;
  assign n4805 = ~n1290 & n4709 ;
  assign n4806 = n4804 | n4805 ;
  assign n4807 = ~n4182 & n4713 ;
  assign n4808 = ( x23 & n4806 ) | ( x23 & ~n4807 ) | ( n4806 & ~n4807 ) ;
  assign n4809 = ( ~x23 & n4806 ) | ( ~x23 & n4807 ) | ( n4806 & n4807 ) ;
  assign n4810 = ( ~n4806 & n4808 ) | ( ~n4806 & n4809 ) | ( n4808 & n4809 ) ;
  assign n4811 = ( ~n4678 & n4687 ) | ( ~n4678 & n4689 ) | ( n4687 & n4689 ) ;
  assign n4812 = ( n4678 & ~n4690 ) | ( n4678 & n4811 ) | ( ~n4690 & n4811 ) ;
  assign n4813 = ~n3791 & n4202 ;
  assign n4814 = n1267 & n4345 ;
  assign n4815 = ~n1246 & n4201 ;
  assign n4816 = ~n1338 & n4200 ;
  assign n4817 = n4815 | n4816 ;
  assign n4818 = ( ~n4813 & n4814 ) | ( ~n4813 & n4817 ) | ( n4814 & n4817 ) ;
  assign n4819 = ( ~x26 & n4813 ) | ( ~x26 & n4818 ) | ( n4813 & n4818 ) ;
  assign n4820 = ( n4813 & n4818 ) | ( n4813 & ~n4819 ) | ( n4818 & ~n4819 ) ;
  assign n4821 = ( x26 & n4819 ) | ( x26 & ~n4820 ) | ( n4819 & ~n4820 ) ;
  assign n4822 = ( n4787 & n4812 ) | ( n4787 & n4821 ) | ( n4812 & n4821 ) ;
  assign n4823 = ( ~n4787 & n4812 ) | ( ~n4787 & n4821 ) | ( n4812 & n4821 ) ;
  assign n4824 = ( n4787 & ~n4822 ) | ( n4787 & n4823 ) | ( ~n4822 & n4823 ) ;
  assign n4825 = ( n4801 & n4810 ) | ( n4801 & n4824 ) | ( n4810 & n4824 ) ;
  assign n4826 = n887 | n2077 ;
  assign n4827 = n45 | n1235 ;
  assign n4828 = n519 | n1171 ;
  assign n4829 = n1492 | n4828 ;
  assign n4830 = ( n465 & ~n4827 ) | ( n465 & n4829 ) | ( ~n4827 & n4829 ) ;
  assign n4831 = n4827 | n4830 ;
  assign n4832 = n204 | n382 ;
  assign n4833 = ( ~n4826 & n4831 ) | ( ~n4826 & n4832 ) | ( n4831 & n4832 ) ;
  assign n4834 = n4826 | n4833 ;
  assign n4835 = n2726 | n3841 ;
  assign n4836 = n91 | n362 ;
  assign n4837 = n1718 | n4836 ;
  assign n4838 = ( ~n1714 & n4835 ) | ( ~n1714 & n4837 ) | ( n4835 & n4837 ) ;
  assign n4839 = ( n1714 & ~n4834 ) | ( n1714 & n4838 ) | ( ~n4834 & n4838 ) ;
  assign n4840 = n103 | n719 ;
  assign n4841 = n4397 | n4840 ;
  assign n4842 = ( n4834 & ~n4839 ) | ( n4834 & n4841 ) | ( ~n4839 & n4841 ) ;
  assign n4843 = n4839 | n4842 ;
  assign n4844 = n1022 | n1613 ;
  assign n4845 = n4043 | n4844 ;
  assign n4846 = ( n895 & ~n957 ) | ( n895 & n1254 ) | ( ~n957 & n1254 ) ;
  assign n4847 = n957 | n4846 ;
  assign n4848 = n479 | n921 ;
  assign n4849 = n261 | n661 ;
  assign n4850 = ( n884 & ~n4848 ) | ( n884 & n4849 ) | ( ~n4848 & n4849 ) ;
  assign n4851 = n4848 | n4850 ;
  assign n4852 = ( n1159 & n2067 ) | ( n1159 & ~n4851 ) | ( n2067 & ~n4851 ) ;
  assign n4853 = n4851 | n4852 ;
  assign n4854 = n124 | n267 ;
  assign n4855 = ( n566 & n586 ) | ( n566 & ~n4854 ) | ( n586 & ~n4854 ) ;
  assign n4856 = n4854 | n4855 ;
  assign n4857 = ( ~n4847 & n4853 ) | ( ~n4847 & n4856 ) | ( n4853 & n4856 ) ;
  assign n4858 = n4847 | n4857 ;
  assign n4859 = ( n3749 & ~n4845 ) | ( n3749 & n4858 ) | ( ~n4845 & n4858 ) ;
  assign n4860 = n4845 | n4859 ;
  assign n4861 = n137 | n272 ;
  assign n4862 = ( n912 & n1449 ) | ( n912 & ~n4861 ) | ( n1449 & ~n4861 ) ;
  assign n4863 = n4861 | n4862 ;
  assign n4864 = ( n197 & n294 ) | ( n197 & ~n1512 ) | ( n294 & ~n1512 ) ;
  assign n4865 = n1512 | n4864 ;
  assign n4866 = n240 | n455 ;
  assign n4867 = ( n227 & n488 ) | ( n227 & ~n4866 ) | ( n488 & ~n4866 ) ;
  assign n4868 = n4866 | n4867 ;
  assign n4869 = ( n1979 & n3994 ) | ( n1979 & ~n4868 ) | ( n3994 & ~n4868 ) ;
  assign n4870 = n4868 | n4869 ;
  assign n4871 = ( n4863 & n4865 ) | ( n4863 & ~n4870 ) | ( n4865 & ~n4870 ) ;
  assign n4872 = n255 | n331 ;
  assign n4873 = n79 | n1110 ;
  assign n4874 = n4872 | n4873 ;
  assign n4875 = ( n4870 & ~n4871 ) | ( n4870 & n4874 ) | ( ~n4871 & n4874 ) ;
  assign n4876 = n4871 | n4875 ;
  assign n4877 = n4860 | n4876 ;
  assign n4878 = n1793 | n3339 ;
  assign n4879 = ( n2845 & ~n4874 ) | ( n2845 & n4878 ) | ( ~n4874 & n4878 ) ;
  assign n4880 = n77 | n1510 ;
  assign n4881 = n3391 | n4880 ;
  assign n4882 = n697 | n1237 ;
  assign n4883 = n224 | n576 ;
  assign n4884 = ( n3499 & ~n4882 ) | ( n3499 & n4883 ) | ( ~n4882 & n4883 ) ;
  assign n4885 = n4882 | n4884 ;
  assign n4886 = n170 | n562 ;
  assign n4887 = ( n1169 & n3241 ) | ( n1169 & ~n4886 ) | ( n3241 & ~n4886 ) ;
  assign n4888 = n4886 | n4887 ;
  assign n4889 = ( ~n4881 & n4885 ) | ( ~n4881 & n4888 ) | ( n4885 & n4888 ) ;
  assign n4890 = n4881 | n4889 ;
  assign n4891 = ( ~n4876 & n4879 ) | ( ~n4876 & n4890 ) | ( n4879 & n4890 ) ;
  assign n4892 = ( ~n4843 & n4877 ) | ( ~n4843 & n4891 ) | ( n4877 & n4891 ) ;
  assign n4893 = n4843 | n4892 ;
  assign n4894 = n606 & ~n2298 ;
  assign n4895 = n607 & ~n2491 ;
  assign n4896 = n4894 | n4895 ;
  assign n4897 = ~n1250 & n2396 ;
  assign n4898 = ( n2396 & n4896 ) | ( n2396 & ~n4897 ) | ( n4896 & ~n4897 ) ;
  assign n4899 = ( n2298 & ~n2396 ) | ( n2298 & n3604 ) | ( ~n2396 & n3604 ) ;
  assign n4900 = ( ~n3604 & n3605 ) | ( ~n3604 & n4899 ) | ( n3605 & n4899 ) ;
  assign n4901 = n1248 & ~n4900 ;
  assign n4902 = n4898 | n4901 ;
  assign n4903 = ( ~n4541 & n4893 ) | ( ~n4541 & n4902 ) | ( n4893 & n4902 ) ;
  assign n4904 = ( ~x14 & n4541 ) | ( ~x14 & n4608 ) | ( n4541 & n4608 ) ;
  assign n4905 = ( ~n4608 & n4609 ) | ( ~n4608 & n4904 ) | ( n4609 & n4904 ) ;
  assign n4906 = n1250 | n2298 ;
  assign n4907 = n606 & n2270 ;
  assign n4908 = ( ~n2298 & n4906 ) | ( ~n2298 & n4907 ) | ( n4906 & n4907 ) ;
  assign n4909 = n607 & ~n2396 ;
  assign n4910 = ( n607 & n4908 ) | ( n607 & ~n4909 ) | ( n4908 & ~n4909 ) ;
  assign n4911 = ( ~n2270 & n2298 ) | ( ~n2270 & n3605 ) | ( n2298 & n3605 ) ;
  assign n4912 = ( ~n3605 & n3606 ) | ( ~n3605 & n4911 ) | ( n3606 & n4911 ) ;
  assign n4913 = n1248 & ~n4912 ;
  assign n4914 = n4910 | n4913 ;
  assign n4915 = ( n4903 & n4905 ) | ( n4903 & n4914 ) | ( n4905 & n4914 ) ;
  assign n4916 = ( ~n4609 & n4640 ) | ( ~n4609 & n4649 ) | ( n4640 & n4649 ) ;
  assign n4917 = ( n4609 & ~n4650 ) | ( n4609 & n4916 ) | ( ~n4650 & n4916 ) ;
  assign n4918 = n3800 & ~n4457 ;
  assign n4919 = n1926 & n3799 ;
  assign n4920 = ~n2023 & n3802 ;
  assign n4921 = ( ~n2089 & n3694 ) | ( ~n2089 & n3699 ) | ( n3694 & n3699 ) ;
  assign n4922 = ( n3694 & n4920 ) | ( n3694 & ~n4921 ) | ( n4920 & ~n4921 ) ;
  assign n4923 = ( ~n4918 & n4919 ) | ( ~n4918 & n4922 ) | ( n4919 & n4922 ) ;
  assign n4924 = ( ~x29 & n4918 ) | ( ~x29 & n4923 ) | ( n4918 & n4923 ) ;
  assign n4925 = ( n4918 & n4923 ) | ( n4918 & ~n4924 ) | ( n4923 & ~n4924 ) ;
  assign n4926 = ( x29 & n4924 ) | ( x29 & ~n4925 ) | ( n4924 & ~n4925 ) ;
  assign n4927 = ( n4915 & n4917 ) | ( n4915 & n4926 ) | ( n4917 & n4926 ) ;
  assign n4928 = ( n4732 & n4741 ) | ( n4732 & ~n4742 ) | ( n4741 & ~n4742 ) ;
  assign n4929 = ( n4723 & n4742 ) | ( n4723 & ~n4928 ) | ( n4742 & ~n4928 ) ;
  assign n4930 = n4202 & n4326 ;
  assign n4931 = n1576 & n4201 ;
  assign n4932 = n1750 | n4200 ;
  assign n4933 = ~n1669 & n4345 ;
  assign n4934 = ( ~n1750 & n4932 ) | ( ~n1750 & n4933 ) | ( n4932 & n4933 ) ;
  assign n4935 = ( ~n4930 & n4931 ) | ( ~n4930 & n4934 ) | ( n4931 & n4934 ) ;
  assign n4936 = ( ~x26 & n4930 ) | ( ~x26 & n4935 ) | ( n4930 & n4935 ) ;
  assign n4937 = ( n4930 & n4935 ) | ( n4930 & ~n4936 ) | ( n4935 & ~n4936 ) ;
  assign n4938 = ( x26 & n4936 ) | ( x26 & ~n4937 ) | ( n4936 & ~n4937 ) ;
  assign n4939 = ( n4927 & ~n4929 ) | ( n4927 & n4938 ) | ( ~n4929 & n4938 ) ;
  assign n4940 = ( n4742 & ~n4744 ) | ( n4742 & n4753 ) | ( ~n4744 & n4753 ) ;
  assign n4941 = ( n4744 & ~n4754 ) | ( n4744 & n4940 ) | ( ~n4754 & n4940 ) ;
  assign n4942 = ~n4159 & n4202 ;
  assign n4943 = n1458 & n4201 ;
  assign n4944 = ~n1669 & n4200 ;
  assign n4945 = n1576 & n4345 ;
  assign n4946 = n4944 | n4945 ;
  assign n4947 = ( ~n4942 & n4943 ) | ( ~n4942 & n4946 ) | ( n4943 & n4946 ) ;
  assign n4948 = ( ~x26 & n4942 ) | ( ~x26 & n4947 ) | ( n4942 & n4947 ) ;
  assign n4949 = ( n4942 & n4947 ) | ( n4942 & ~n4948 ) | ( n4947 & ~n4948 ) ;
  assign n4950 = ( x26 & n4948 ) | ( x26 & ~n4949 ) | ( n4948 & ~n4949 ) ;
  assign n4951 = ( n4939 & n4941 ) | ( n4939 & n4950 ) | ( n4941 & n4950 ) ;
  assign n4952 = ( ~n4754 & n4756 ) | ( ~n4754 & n4765 ) | ( n4756 & n4765 ) ;
  assign n4953 = ( n4754 & ~n4766 ) | ( n4754 & n4952 ) | ( ~n4766 & n4952 ) ;
  assign n4954 = n3621 & n4713 ;
  assign n4955 = ~n1290 & n4712 ;
  assign n4956 = ~n1246 & n4792 ;
  assign n4957 = n1267 & n4709 ;
  assign n4958 = n4956 | n4957 ;
  assign n4959 = ( ~n4954 & n4955 ) | ( ~n4954 & n4958 ) | ( n4955 & n4958 ) ;
  assign n4960 = ( ~x23 & n4954 ) | ( ~x23 & n4959 ) | ( n4954 & n4959 ) ;
  assign n4961 = ( n4954 & n4959 ) | ( n4954 & ~n4960 ) | ( n4959 & ~n4960 ) ;
  assign n4962 = ( x23 & n4960 ) | ( x23 & ~n4961 ) | ( n4960 & ~n4961 ) ;
  assign n4963 = ( n4951 & n4953 ) | ( n4951 & n4962 ) | ( n4953 & n4962 ) ;
  assign n4964 = x19 | x20 ;
  assign n4965 = x19 & x20 ;
  assign n4966 = n4964 & ~n4965 ;
  assign n4967 = x17 & x18 ;
  assign n4968 = x17 | x18 ;
  assign n4969 = ( n4966 & n4967 ) | ( n4966 & ~n4968 ) | ( n4967 & ~n4968 ) ;
  assign n4970 = x18 | x19 ;
  assign n4971 = x17 & ~x19 ;
  assign n4972 = ( ~n4968 & n4970 ) | ( ~n4968 & n4971 ) | ( n4970 & n4971 ) ;
  assign n4973 = n4969 & ~n4972 ;
  assign n4974 = n4966 & ~n4969 ;
  assign n4975 = ~n3691 & n4974 ;
  assign n4976 = ( ~n3692 & n4973 ) | ( ~n3692 & n4975 ) | ( n4973 & n4975 ) ;
  assign n4977 = x20 | n4976 ;
  assign n4978 = ( x20 & n4976 ) | ( x20 & ~n4977 ) | ( n4976 & ~n4977 ) ;
  assign n4979 = n4977 & ~n4978 ;
  assign n4980 = ( ~n4766 & n4789 ) | ( ~n4766 & n4800 ) | ( n4789 & n4800 ) ;
  assign n4981 = ( ~n4800 & n4801 ) | ( ~n4800 & n4980 ) | ( n4801 & n4980 ) ;
  assign n4982 = ( n4963 & n4979 ) | ( n4963 & ~n4981 ) | ( n4979 & ~n4981 ) ;
  assign n4983 = n51 | n1096 ;
  assign n4984 = n500 | n4983 ;
  assign n4985 = n774 | n4984 ;
  assign n4986 = n3879 | n4985 ;
  assign n4987 = n67 | n290 ;
  assign n4988 = n489 | n528 ;
  assign n4989 = n1445 | n4988 ;
  assign n4990 = ( n2802 & ~n4985 ) | ( n2802 & n4989 ) | ( ~n4985 & n4989 ) ;
  assign n4991 = n4987 | n4990 ;
  assign n4992 = n1708 | n2636 ;
  assign n4993 = ( n83 & n136 ) | ( n83 & n166 ) | ( n136 & n166 ) ;
  assign n4994 = ( n2924 & ~n4992 ) | ( n2924 & n4993 ) | ( ~n4992 & n4993 ) ;
  assign n4995 = n4992 | n4994 ;
  assign n4996 = ( n224 & n240 ) | ( n224 & ~n1976 ) | ( n240 & ~n1976 ) ;
  assign n4997 = n1976 | n4996 ;
  assign n4998 = ( ~n4987 & n4995 ) | ( ~n4987 & n4997 ) | ( n4995 & n4997 ) ;
  assign n4999 = ( ~n4986 & n4991 ) | ( ~n4986 & n4998 ) | ( n4991 & n4998 ) ;
  assign n5000 = n4986 | n4999 ;
  assign n5001 = n1323 | n3362 ;
  assign n5002 = n348 | n488 ;
  assign n5003 = n368 | n447 ;
  assign n5004 = ( n45 & ~n234 ) | ( n45 & n696 ) | ( ~n234 & n696 ) ;
  assign n5005 = n234 | n5004 ;
  assign n5006 = ( n885 & ~n5003 ) | ( n885 & n5005 ) | ( ~n5003 & n5005 ) ;
  assign n5007 = n5003 | n5006 ;
  assign n5008 = n287 | n4601 ;
  assign n5009 = ( n2377 & ~n5007 ) | ( n2377 & n5008 ) | ( ~n5007 & n5008 ) ;
  assign n5010 = n5007 | n5009 ;
  assign n5011 = ( ~n5001 & n5002 ) | ( ~n5001 & n5010 ) | ( n5002 & n5010 ) ;
  assign n5012 = n5001 | n5011 ;
  assign n5013 = n2564 | n4493 ;
  assign n5014 = ( n383 & n675 ) | ( n383 & ~n943 ) | ( n675 & ~n943 ) ;
  assign n5015 = n943 | n5014 ;
  assign n5016 = n120 | n171 ;
  assign n5017 = n485 | n5016 ;
  assign n5018 = ( ~n54 & n57 ) | ( ~n54 & n97 ) | ( n57 & n97 ) ;
  assign n5019 = n786 | n5018 ;
  assign n5020 = ( n299 & n395 ) | ( n299 & ~n1974 ) | ( n395 & ~n1974 ) ;
  assign n5021 = n1974 | n5020 ;
  assign n5022 = ( n702 & ~n4133 ) | ( n702 & n5021 ) | ( ~n4133 & n5021 ) ;
  assign n5023 = ( n4133 & ~n5019 ) | ( n4133 & n5022 ) | ( ~n5019 & n5022 ) ;
  assign n5024 = ( ~n5017 & n5019 ) | ( ~n5017 & n5023 ) | ( n5019 & n5023 ) ;
  assign n5025 = n5017 | n5024 ;
  assign n5026 = ( ~n5013 & n5015 ) | ( ~n5013 & n5025 ) | ( n5015 & n5025 ) ;
  assign n5027 = n5013 | n5026 ;
  assign n5028 = ( ~n1667 & n5012 ) | ( ~n1667 & n5027 ) | ( n5012 & n5027 ) ;
  assign n5029 = ( n1667 & ~n5000 ) | ( n1667 & n5028 ) | ( ~n5000 & n5028 ) ;
  assign n5030 = n5000 | n5029 ;
  assign n5031 = n3851 | n4011 ;
  assign n5032 = n163 | n719 ;
  assign n5033 = n360 | n655 ;
  assign n5034 = ( n144 & n1477 ) | ( n144 & ~n5033 ) | ( n1477 & ~n5033 ) ;
  assign n5035 = n5033 | n5034 ;
  assign n5036 = ( n653 & ~n5032 ) | ( n653 & n5035 ) | ( ~n5032 & n5035 ) ;
  assign n5037 = n5032 | n5036 ;
  assign n5038 = n718 | n2236 ;
  assign n5039 = n1929 | n2093 ;
  assign n5040 = n1593 | n1976 ;
  assign n5041 = n518 | n577 ;
  assign n5042 = ( n133 & n1024 ) | ( n133 & ~n5041 ) | ( n1024 & ~n5041 ) ;
  assign n5043 = n5041 | n5042 ;
  assign n5044 = ( ~n5039 & n5040 ) | ( ~n5039 & n5043 ) | ( n5040 & n5043 ) ;
  assign n5045 = n5039 | n5044 ;
  assign n5046 = ( ~n5037 & n5038 ) | ( ~n5037 & n5045 ) | ( n5038 & n5045 ) ;
  assign n5047 = n5037 | n5046 ;
  assign n5048 = ( ~n5012 & n5031 ) | ( ~n5012 & n5047 ) | ( n5031 & n5047 ) ;
  assign n5049 = n689 | n783 ;
  assign n5050 = n1863 | n5049 ;
  assign n5051 = n1057 | n2353 ;
  assign n5052 = ( n83 & n109 ) | ( n83 & n119 ) | ( n109 & n119 ) ;
  assign n5053 = n732 | n5052 ;
  assign n5054 = ( n384 & n2672 ) | ( n384 & ~n5053 ) | ( n2672 & ~n5053 ) ;
  assign n5055 = n5053 | n5054 ;
  assign n5056 = n103 | n227 ;
  assign n5057 = ( n293 & n537 ) | ( n293 & ~n5056 ) | ( n537 & ~n5056 ) ;
  assign n5058 = n5056 | n5057 ;
  assign n5059 = ( ~n5051 & n5055 ) | ( ~n5051 & n5058 ) | ( n5055 & n5058 ) ;
  assign n5060 = n5051 | n5059 ;
  assign n5061 = n230 | n448 ;
  assign n5062 = n918 | n2654 ;
  assign n5063 = n5061 | n5062 ;
  assign n5064 = ( n5050 & ~n5060 ) | ( n5050 & n5063 ) | ( ~n5060 & n5063 ) ;
  assign n5065 = n188 | n2248 ;
  assign n5066 = ( ~n540 & n581 ) | ( ~n540 & n5065 ) | ( n581 & n5065 ) ;
  assign n5067 = n661 | n838 ;
  assign n5068 = ( ~n176 & n3406 ) | ( ~n176 & n5067 ) | ( n3406 & n5067 ) ;
  assign n5069 = n176 | n3994 ;
  assign n5070 = n5068 | n5069 ;
  assign n5071 = ( n3329 & ~n5066 ) | ( n3329 & n5070 ) | ( ~n5066 & n5070 ) ;
  assign n5072 = n5066 | n5071 ;
  assign n5073 = ( n5060 & ~n5064 ) | ( n5060 & n5072 ) | ( ~n5064 & n5072 ) ;
  assign n5074 = n5064 | n5073 ;
  assign n5075 = ( n5012 & ~n5048 ) | ( n5012 & n5074 ) | ( ~n5048 & n5074 ) ;
  assign n5076 = n5048 | n5075 ;
  assign n5077 = ( ~x11 & n5030 ) | ( ~x11 & n5076 ) | ( n5030 & n5076 ) ;
  assign n5078 = n1250 & ~n2491 ;
  assign n5079 = n607 & n2552 ;
  assign n5080 = n5078 | n5079 ;
  assign n5081 = n606 & ~n2396 ;
  assign n5082 = ( n606 & n5080 ) | ( n606 & ~n5081 ) | ( n5080 & ~n5081 ) ;
  assign n5083 = ( n2396 & n2491 ) | ( n2396 & n3603 ) | ( n2491 & n3603 ) ;
  assign n5084 = ( n2491 & n3604 ) | ( n2491 & ~n5083 ) | ( n3604 & ~n5083 ) ;
  assign n5085 = n1248 & ~n5084 ;
  assign n5086 = n5082 | n5085 ;
  assign n5087 = ( ~n4541 & n5077 ) | ( ~n4541 & n5086 ) | ( n5077 & n5086 ) ;
  assign n5088 = n444 | n1313 ;
  assign n5089 = n174 | n433 ;
  assign n5090 = ( n3144 & ~n5088 ) | ( n3144 & n5089 ) | ( ~n5088 & n5089 ) ;
  assign n5091 = n5088 | n5090 ;
  assign n5092 = n384 | n1711 ;
  assign n5093 = ( n3306 & n3501 ) | ( n3306 & ~n3879 ) | ( n3501 & ~n3879 ) ;
  assign n5094 = n3879 | n5093 ;
  assign n5095 = ( ~n4048 & n5092 ) | ( ~n4048 & n5094 ) | ( n5092 & n5094 ) ;
  assign n5096 = ( n4048 & n4597 ) | ( n4048 & ~n5095 ) | ( n4597 & ~n5095 ) ;
  assign n5097 = n5095 | n5096 ;
  assign n5098 = ( n85 & n455 ) | ( n85 & ~n981 ) | ( n455 & ~n981 ) ;
  assign n5099 = n981 | n5098 ;
  assign n5100 = ( ~n5091 & n5097 ) | ( ~n5091 & n5099 ) | ( n5097 & n5099 ) ;
  assign n5101 = n5091 | n5100 ;
  assign n5102 = n523 | n1031 ;
  assign n5103 = ( n519 & n638 ) | ( n519 & ~n5102 ) | ( n638 & ~n5102 ) ;
  assign n5104 = n5102 | n5103 ;
  assign n5105 = n115 | n947 ;
  assign n5106 = ( n3121 & ~n5104 ) | ( n3121 & n5105 ) | ( ~n5104 & n5105 ) ;
  assign n5107 = n5104 | n5106 ;
  assign n5108 = n132 | n277 ;
  assign n5109 = n445 | n567 ;
  assign n5110 = ( n238 & n582 ) | ( n238 & ~n5109 ) | ( n582 & ~n5109 ) ;
  assign n5111 = n5109 | n5110 ;
  assign n5112 = ( n777 & ~n5108 ) | ( n777 & n5111 ) | ( ~n5108 & n5111 ) ;
  assign n5113 = n5108 | n5112 ;
  assign n5114 = ( n2102 & ~n2188 ) | ( n2102 & n4530 ) | ( ~n2188 & n4530 ) ;
  assign n5115 = n2188 | n5114 ;
  assign n5116 = n323 | n746 ;
  assign n5117 = n1511 | n1526 ;
  assign n5118 = n5116 | n5117 ;
  assign n5119 = ( ~n5113 & n5115 ) | ( ~n5113 & n5118 ) | ( n5115 & n5118 ) ;
  assign n5120 = n5113 | n5119 ;
  assign n5121 = ~n92 & n218 ;
  assign n5122 = ( n83 & n102 ) | ( n83 & n116 ) | ( n102 & n116 ) ;
  assign n5123 = n514 | n5122 ;
  assign n5124 = n272 | n312 ;
  assign n5125 = ( n207 & n1692 ) | ( n207 & ~n5124 ) | ( n1692 & ~n5124 ) ;
  assign n5126 = n5124 | n5125 ;
  assign n5127 = ( n5121 & n5123 ) | ( n5121 & ~n5126 ) | ( n5123 & ~n5126 ) ;
  assign n5128 = ( n3931 & n5123 ) | ( n3931 & n5127 ) | ( n5123 & n5127 ) ;
  assign n5129 = n5127 & ~n5128 ;
  assign n5130 = ( n5107 & ~n5120 ) | ( n5107 & n5129 ) | ( ~n5120 & n5129 ) ;
  assign n5131 = ~n5107 & n5130 ;
  assign n5132 = n716 | n2215 ;
  assign n5133 = n1012 | n5132 ;
  assign n5134 = n760 | n3079 ;
  assign n5135 = ( n886 & n1225 ) | ( n886 & ~n5134 ) | ( n1225 & ~n5134 ) ;
  assign n5136 = n5134 | n5135 ;
  assign n5137 = ( n253 & ~n5133 ) | ( n253 & n5136 ) | ( ~n5133 & n5136 ) ;
  assign n5138 = n5133 | n5137 ;
  assign n5139 = n317 | n448 ;
  assign n5140 = n111 | n394 ;
  assign n5141 = ( n349 & n676 ) | ( n349 & ~n5140 ) | ( n676 & ~n5140 ) ;
  assign n5142 = n5140 | n5141 ;
  assign n5143 = ( n609 & ~n5139 ) | ( n609 & n5142 ) | ( ~n5139 & n5142 ) ;
  assign n5144 = n5139 | n5143 ;
  assign n5145 = n299 | n952 ;
  assign n5146 = n933 | n1913 ;
  assign n5147 = n5145 | n5146 ;
  assign n5148 = ( ~n5138 & n5144 ) | ( ~n5138 & n5147 ) | ( n5144 & n5147 ) ;
  assign n5149 = n2782 | n5053 ;
  assign n5150 = n5138 | n5149 ;
  assign n5151 = n81 | n1237 ;
  assign n5152 = n941 | n4840 ;
  assign n5153 = ( n3284 & ~n5151 ) | ( n3284 & n5152 ) | ( ~n5151 & n5152 ) ;
  assign n5154 = n5151 | n5153 ;
  assign n5155 = n878 | n928 ;
  assign n5156 = n492 | n517 ;
  assign n5157 = ( n2311 & ~n5155 ) | ( n2311 & n5156 ) | ( ~n5155 & n5156 ) ;
  assign n5158 = n5155 | n5157 ;
  assign n5159 = ( ~n5149 & n5154 ) | ( ~n5149 & n5158 ) | ( n5154 & n5158 ) ;
  assign n5160 = ( ~n5148 & n5150 ) | ( ~n5148 & n5159 ) | ( n5150 & n5159 ) ;
  assign n5161 = n5148 | n5160 ;
  assign n5162 = ( n5101 & n5131 ) | ( n5101 & ~n5161 ) | ( n5131 & ~n5161 ) ;
  assign n5163 = ~n5101 & n5162 ;
  assign n5164 = ( n83 & n84 ) | ( n83 & n145 ) | ( n84 & n145 ) ;
  assign n5165 = ( n517 & n537 ) | ( n517 & ~n5164 ) | ( n537 & ~n5164 ) ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = ( n434 & ~n3472 ) | ( n434 & n5166 ) | ( ~n3472 & n5166 ) ;
  assign n5168 = ( n396 & ~n3472 ) | ( n396 & n5167 ) | ( ~n3472 & n5167 ) ;
  assign n5169 = n243 | n2232 ;
  assign n5170 = n2558 | n5169 ;
  assign n5171 = ( n72 & n119 ) | ( n72 & n129 ) | ( n119 & n129 ) ;
  assign n5172 = n529 | n5171 ;
  assign n5173 = ( ~n230 & n285 ) | ( ~n230 & n5172 ) | ( n285 & n5172 ) ;
  assign n5174 = ( n230 & n1870 ) | ( n230 & ~n5173 ) | ( n1870 & ~n5173 ) ;
  assign n5175 = n5173 | n5174 ;
  assign n5176 = ( n919 & ~n5170 ) | ( n919 & n5175 ) | ( ~n5170 & n5175 ) ;
  assign n5177 = n5170 | n5176 ;
  assign n5178 = ( n3472 & ~n5168 ) | ( n3472 & n5177 ) | ( ~n5168 & n5177 ) ;
  assign n5179 = n5168 | n5178 ;
  assign n5180 = n836 | n3551 ;
  assign n5181 = n1312 | n1515 ;
  assign n5182 = ( n4263 & ~n5180 ) | ( n4263 & n5181 ) | ( ~n5180 & n5181 ) ;
  assign n5183 = n5180 | n5182 ;
  assign n5184 = n347 | n4551 ;
  assign n5185 = n45 | n653 ;
  assign n5186 = ( n123 & n136 ) | ( n123 & n469 ) | ( n136 & n469 ) ;
  assign n5187 = ( n240 & n1171 ) | ( n240 & ~n5186 ) | ( n1171 & ~n5186 ) ;
  assign n5188 = n5186 | n5187 ;
  assign n5189 = ( ~n5184 & n5185 ) | ( ~n5184 & n5188 ) | ( n5185 & n5188 ) ;
  assign n5190 = n5184 | n5189 ;
  assign n5191 = ( n5179 & ~n5183 ) | ( n5179 & n5190 ) | ( ~n5183 & n5190 ) ;
  assign n5192 = n4243 | n5191 ;
  assign n5193 = n1253 | n1487 ;
  assign n5194 = n91 | n331 ;
  assign n5195 = n3285 | n4554 ;
  assign n5196 = n5194 | n5195 ;
  assign n5197 = n124 | n131 ;
  assign n5198 = ( n265 & n746 ) | ( n265 & ~n5197 ) | ( n746 & ~n5197 ) ;
  assign n5199 = n5197 | n5198 ;
  assign n5200 = ( ~n5193 & n5196 ) | ( ~n5193 & n5199 ) | ( n5196 & n5199 ) ;
  assign n5201 = n5193 | n5200 ;
  assign n5202 = n487 | n5201 ;
  assign n5203 = n500 | n642 ;
  assign n5204 = ( n239 & n734 ) | ( n239 & ~n5203 ) | ( n734 & ~n5203 ) ;
  assign n5205 = n5203 | n5204 ;
  assign n5206 = ( n1032 & ~n3356 ) | ( n1032 & n5205 ) | ( ~n3356 & n5205 ) ;
  assign n5207 = n3356 | n5206 ;
  assign n5208 = n120 | n1808 ;
  assign n5209 = ( n208 & n666 ) | ( n208 & ~n1365 ) | ( n666 & ~n1365 ) ;
  assign n5210 = n1365 | n5209 ;
  assign n5211 = ( n1020 & n1589 ) | ( n1020 & ~n5210 ) | ( n1589 & ~n5210 ) ;
  assign n5212 = n5210 | n5211 ;
  assign n5213 = n161 | n1511 ;
  assign n5214 = ( n1078 & n2628 ) | ( n1078 & ~n5213 ) | ( n2628 & ~n5213 ) ;
  assign n5215 = n5213 | n5214 ;
  assign n5216 = ( ~n5208 & n5212 ) | ( ~n5208 & n5215 ) | ( n5212 & n5215 ) ;
  assign n5217 = ( ~n4246 & n5208 ) | ( ~n4246 & n5216 ) | ( n5208 & n5216 ) ;
  assign n5218 = n4246 | n5217 ;
  assign n5219 = ( ~n5202 & n5207 ) | ( ~n5202 & n5218 ) | ( n5207 & n5218 ) ;
  assign n5220 = n5202 | n5219 ;
  assign n5221 = ( n5183 & ~n5192 ) | ( n5183 & n5220 ) | ( ~n5192 & n5220 ) ;
  assign n5222 = n5192 | n5221 ;
  assign n5223 = ( x8 & n5163 ) | ( x8 & ~n5222 ) | ( n5163 & ~n5222 ) ;
  assign n5224 = n1250 & ~n2725 ;
  assign n5225 = n606 & n2635 ;
  assign n5226 = n5224 | n5225 ;
  assign n5227 = n607 & n2810 ;
  assign n5228 = ( n607 & n5226 ) | ( n607 & ~n5227 ) | ( n5226 & ~n5227 ) ;
  assign n5229 = ( ~n2810 & n2843 ) | ( ~n2810 & n3598 ) | ( n2843 & n3598 ) ;
  assign n5230 = ( n2725 & ~n2843 ) | ( n2725 & n5229 ) | ( ~n2843 & n5229 ) ;
  assign n5231 = ( n2635 & n3599 ) | ( n2635 & ~n5230 ) | ( n3599 & ~n5230 ) ;
  assign n5232 = ( ~n3600 & n3601 ) | ( ~n3600 & n5231 ) | ( n3601 & n5231 ) ;
  assign n5233 = n1248 & n5232 ;
  assign n5234 = n5228 | n5233 ;
  assign n5235 = ( n5030 & n5223 ) | ( n5030 & ~n5234 ) | ( n5223 & ~n5234 ) ;
  assign n5236 = n2021 | n2583 ;
  assign n5237 = n675 | n1031 ;
  assign n5238 = ( n493 & n2045 ) | ( n493 & ~n5237 ) | ( n2045 & ~n5237 ) ;
  assign n5239 = n5237 | n5238 ;
  assign n5240 = ( n50 & n59 ) | ( n50 & n129 ) | ( n59 & n129 ) ;
  assign n5241 = n745 | n5240 ;
  assign n5242 = ( n262 & n465 ) | ( n262 & ~n773 ) | ( n465 & ~n773 ) ;
  assign n5243 = n773 | n5242 ;
  assign n5244 = n5241 | n5243 ;
  assign n5245 = n2846 | n3303 ;
  assign n5246 = n131 | n1376 ;
  assign n5247 = n233 | n1171 ;
  assign n5248 = ( n648 & ~n5246 ) | ( n648 & n5247 ) | ( ~n5246 & n5247 ) ;
  assign n5249 = n5246 | n5248 ;
  assign n5250 = n224 | n352 ;
  assign n5251 = ( n51 & n1346 ) | ( n51 & ~n5250 ) | ( n1346 & ~n5250 ) ;
  assign n5252 = n5250 | n5251 ;
  assign n5253 = ( ~n5245 & n5249 ) | ( ~n5245 & n5252 ) | ( n5249 & n5252 ) ;
  assign n5254 = n5245 | n5253 ;
  assign n5255 = ( ~n5239 & n5244 ) | ( ~n5239 & n5254 ) | ( n5244 & n5254 ) ;
  assign n5256 = n5239 | n5255 ;
  assign n5257 = ( ~n2583 & n3865 ) | ( ~n2583 & n5256 ) | ( n3865 & n5256 ) ;
  assign n5258 = ( ~n2603 & n5236 ) | ( ~n2603 & n5257 ) | ( n5236 & n5257 ) ;
  assign n5259 = n2603 | n5258 ;
  assign n5260 = ( n5030 & n5235 ) | ( n5030 & ~n5259 ) | ( n5235 & ~n5259 ) ;
  assign n5261 = ( n5030 & n5076 ) | ( n5030 & ~n5077 ) | ( n5076 & ~n5077 ) ;
  assign n5262 = ( x11 & n5077 ) | ( x11 & ~n5261 ) | ( n5077 & ~n5261 ) ;
  assign n5263 = n606 & ~n2491 ;
  assign n5264 = n607 & n2635 ;
  assign n5265 = n5263 | n5264 ;
  assign n5266 = ~n1250 & n2552 ;
  assign n5267 = ( n2552 & n5265 ) | ( n2552 & ~n5266 ) | ( n5265 & ~n5266 ) ;
  assign n5268 = ( ~n2552 & n2725 ) | ( ~n2552 & n5231 ) | ( n2725 & n5231 ) ;
  assign n5269 = ( n2491 & n3601 ) | ( n2491 & ~n5268 ) | ( n3601 & ~n5268 ) ;
  assign n5270 = ( ~n2552 & n3603 ) | ( ~n2552 & n5269 ) | ( n3603 & n5269 ) ;
  assign n5271 = n1248 & ~n5270 ;
  assign n5272 = n5267 | n5271 ;
  assign n5273 = ( n5260 & n5262 ) | ( n5260 & ~n5272 ) | ( n5262 & ~n5272 ) ;
  assign n5274 = ( n4541 & ~n5077 ) | ( n4541 & n5086 ) | ( ~n5077 & n5086 ) ;
  assign n5275 = ( ~n5086 & n5087 ) | ( ~n5086 & n5274 ) | ( n5087 & n5274 ) ;
  assign n5276 = n3800 & n4647 ;
  assign n5277 = n2174 & n3799 ;
  assign n5278 = n2298 | n3700 ;
  assign n5279 = n2270 & n3802 ;
  assign n5280 = ( ~n2298 & n5278 ) | ( ~n2298 & n5279 ) | ( n5278 & n5279 ) ;
  assign n5281 = ( ~n5276 & n5277 ) | ( ~n5276 & n5280 ) | ( n5277 & n5280 ) ;
  assign n5282 = ( ~x29 & n5276 ) | ( ~x29 & n5281 ) | ( n5276 & n5281 ) ;
  assign n5283 = ( n5276 & n5281 ) | ( n5276 & ~n5282 ) | ( n5281 & ~n5282 ) ;
  assign n5284 = ( x29 & n5282 ) | ( x29 & ~n5283 ) | ( n5282 & ~n5283 ) ;
  assign n5285 = ( n5273 & n5275 ) | ( n5273 & ~n5284 ) | ( n5275 & ~n5284 ) ;
  assign n5286 = ( n4893 & n4902 ) | ( n4893 & ~n4903 ) | ( n4902 & ~n4903 ) ;
  assign n5287 = ( n4541 & n4903 ) | ( n4541 & ~n5286 ) | ( n4903 & ~n5286 ) ;
  assign n5288 = ( ~n5087 & n5285 ) | ( ~n5087 & n5287 ) | ( n5285 & n5287 ) ;
  assign n5289 = n3800 & ~n4660 ;
  assign n5290 = ~n2023 & n3799 ;
  assign n5291 = n2174 & n3700 ;
  assign n5292 = n2089 & n3802 ;
  assign n5293 = n5291 | n5292 ;
  assign n5294 = ( ~n5289 & n5290 ) | ( ~n5289 & n5293 ) | ( n5290 & n5293 ) ;
  assign n5295 = ( ~x29 & n5289 ) | ( ~x29 & n5294 ) | ( n5289 & n5294 ) ;
  assign n5296 = ( n5289 & n5294 ) | ( n5289 & ~n5295 ) | ( n5294 & ~n5295 ) ;
  assign n5297 = ( x29 & n5295 ) | ( x29 & ~n5296 ) | ( n5295 & ~n5296 ) ;
  assign n5298 = ( n4903 & ~n4905 ) | ( n4903 & n4914 ) | ( ~n4905 & n4914 ) ;
  assign n5299 = ( n4905 & ~n4915 ) | ( n4905 & n5298 ) | ( ~n4915 & n5298 ) ;
  assign n5300 = ( ~n5288 & n5297 ) | ( ~n5288 & n5299 ) | ( n5297 & n5299 ) ;
  assign n5301 = ( n4915 & ~n4917 ) | ( n4915 & n4926 ) | ( ~n4917 & n4926 ) ;
  assign n5302 = ( n4917 & ~n4927 ) | ( n4917 & n5301 ) | ( ~n4927 & n5301 ) ;
  assign n5303 = n4146 & n4202 ;
  assign n5304 = ~n1669 & n4201 ;
  assign n5305 = n1852 & ~n4200 ;
  assign n5306 = ~n1750 & n4345 ;
  assign n5307 = ( n1852 & ~n5305 ) | ( n1852 & n5306 ) | ( ~n5305 & n5306 ) ;
  assign n5308 = ( ~n5303 & n5304 ) | ( ~n5303 & n5307 ) | ( n5304 & n5307 ) ;
  assign n5309 = ( ~x26 & n5303 ) | ( ~x26 & n5308 ) | ( n5303 & n5308 ) ;
  assign n5310 = ( n5303 & n5308 ) | ( n5303 & ~n5309 ) | ( n5308 & ~n5309 ) ;
  assign n5311 = ( x26 & n5309 ) | ( x26 & ~n5310 ) | ( n5309 & ~n5310 ) ;
  assign n5312 = ( n5300 & n5302 ) | ( n5300 & n5311 ) | ( n5302 & n5311 ) ;
  assign n5313 = ( ~n4927 & n4929 ) | ( ~n4927 & n4938 ) | ( n4929 & n4938 ) ;
  assign n5314 = ( ~n4938 & n4939 ) | ( ~n4938 & n5313 ) | ( n4939 & n5313 ) ;
  assign n5315 = ~n3779 & n4713 ;
  assign n5316 = n1267 & n4712 ;
  assign n5317 = n1458 & ~n4709 ;
  assign n5318 = ~n1338 & n4792 ;
  assign n5319 = ( n1458 & ~n5317 ) | ( n1458 & n5318 ) | ( ~n5317 & n5318 ) ;
  assign n5320 = ( ~n5315 & n5316 ) | ( ~n5315 & n5319 ) | ( n5316 & n5319 ) ;
  assign n5321 = ( ~x23 & n5315 ) | ( ~x23 & n5320 ) | ( n5315 & n5320 ) ;
  assign n5322 = ( n5315 & n5320 ) | ( n5315 & ~n5321 ) | ( n5320 & ~n5321 ) ;
  assign n5323 = ( x23 & n5321 ) | ( x23 & ~n5322 ) | ( n5321 & ~n5322 ) ;
  assign n5324 = ( n5312 & ~n5314 ) | ( n5312 & n5323 ) | ( ~n5314 & n5323 ) ;
  assign n5325 = ~n3791 & n4713 ;
  assign n5326 = n1267 & n4792 ;
  assign n5327 = ~n1246 & n4712 ;
  assign n5328 = ~n1338 & n4709 ;
  assign n5329 = n5327 | n5328 ;
  assign n5330 = ( ~n5325 & n5326 ) | ( ~n5325 & n5329 ) | ( n5326 & n5329 ) ;
  assign n5331 = ( ~x23 & n5325 ) | ( ~x23 & n5330 ) | ( n5325 & n5330 ) ;
  assign n5332 = ( n5325 & n5330 ) | ( n5325 & ~n5331 ) | ( n5330 & ~n5331 ) ;
  assign n5333 = ( x23 & n5331 ) | ( x23 & ~n5332 ) | ( n5331 & ~n5332 ) ;
  assign n5334 = ( ~n4939 & n4941 ) | ( ~n4939 & n4950 ) | ( n4941 & n4950 ) ;
  assign n5335 = ( n4939 & ~n4951 ) | ( n4939 & n5334 ) | ( ~n4951 & n5334 ) ;
  assign n5336 = ( n5324 & n5333 ) | ( n5324 & n5335 ) | ( n5333 & n5335 ) ;
  assign n5337 = ( ~n4951 & n4953 ) | ( ~n4951 & n4962 ) | ( n4953 & n4962 ) ;
  assign n5338 = ( n4951 & ~n4963 ) | ( n4951 & n5337 ) | ( ~n4963 & n5337 ) ;
  assign n5339 = n3797 & n4974 ;
  assign n5340 = ~n3692 & n4972 ;
  assign n5341 = ~n3658 & n4973 ;
  assign n5342 = n5340 | n5341 ;
  assign n5343 = ( ~x20 & n5339 ) | ( ~x20 & n5342 ) | ( n5339 & n5342 ) ;
  assign n5344 = ( n5339 & n5342 ) | ( n5339 & ~n5343 ) | ( n5342 & ~n5343 ) ;
  assign n5345 = ( x20 & n5343 ) | ( x20 & ~n5344 ) | ( n5343 & ~n5344 ) ;
  assign n5346 = ( n5336 & n5338 ) | ( n5336 & n5345 ) | ( n5338 & n5345 ) ;
  assign n5347 = ( n5285 & n5287 ) | ( n5285 & ~n5288 ) | ( n5287 & ~n5288 ) ;
  assign n5348 = ( n5087 & n5288 ) | ( n5087 & ~n5347 ) | ( n5288 & ~n5347 ) ;
  assign n5349 = n3800 & n4730 ;
  assign n5350 = n2089 & n3799 ;
  assign n5351 = n2270 & n3700 ;
  assign n5352 = n2174 & n3802 ;
  assign n5353 = n5351 | n5352 ;
  assign n5354 = ( ~n5349 & n5350 ) | ( ~n5349 & n5353 ) | ( n5350 & n5353 ) ;
  assign n5355 = ( ~x29 & n5349 ) | ( ~x29 & n5354 ) | ( n5349 & n5354 ) ;
  assign n5356 = ( n5349 & n5354 ) | ( n5349 & ~n5355 ) | ( n5354 & ~n5355 ) ;
  assign n5357 = ( x29 & n5355 ) | ( x29 & ~n5356 ) | ( n5355 & ~n5356 ) ;
  assign n5358 = n4202 & n4290 ;
  assign n5359 = n1852 & n4201 ;
  assign n5360 = ~n2023 & n4200 ;
  assign n5361 = n1926 & n4345 ;
  assign n5362 = n5360 | n5361 ;
  assign n5363 = ( ~n5358 & n5359 ) | ( ~n5358 & n5362 ) | ( n5359 & n5362 ) ;
  assign n5364 = ( ~x26 & n5358 ) | ( ~x26 & n5363 ) | ( n5358 & n5363 ) ;
  assign n5365 = ( n5358 & n5363 ) | ( n5358 & ~n5364 ) | ( n5363 & ~n5364 ) ;
  assign n5366 = ( x26 & n5364 ) | ( x26 & ~n5365 ) | ( n5364 & ~n5365 ) ;
  assign n5367 = ( n5348 & n5357 ) | ( n5348 & n5366 ) | ( n5357 & n5366 ) ;
  assign n5368 = ( n5297 & n5299 ) | ( n5297 & ~n5300 ) | ( n5299 & ~n5300 ) ;
  assign n5369 = ( n5288 & n5300 ) | ( n5288 & ~n5368 ) | ( n5300 & ~n5368 ) ;
  assign n5370 = n4202 & ~n4302 ;
  assign n5371 = ~n1750 & n4201 ;
  assign n5372 = n1852 & n4345 ;
  assign n5373 = n1926 & n4200 ;
  assign n5374 = n5372 | n5373 ;
  assign n5375 = ( ~n5370 & n5371 ) | ( ~n5370 & n5374 ) | ( n5371 & n5374 ) ;
  assign n5376 = ( ~x26 & n5370 ) | ( ~x26 & n5375 ) | ( n5370 & n5375 ) ;
  assign n5377 = ( n5370 & n5375 ) | ( n5370 & ~n5376 ) | ( n5375 & ~n5376 ) ;
  assign n5378 = ( x26 & n5376 ) | ( x26 & ~n5377 ) | ( n5376 & ~n5377 ) ;
  assign n5379 = ( n5367 & ~n5369 ) | ( n5367 & n5378 ) | ( ~n5369 & n5378 ) ;
  assign n5380 = ( n5300 & ~n5302 ) | ( n5300 & n5311 ) | ( ~n5302 & n5311 ) ;
  assign n5381 = ( n5302 & ~n5312 ) | ( n5302 & n5380 ) | ( ~n5312 & n5380 ) ;
  assign n5382 = ~n3955 & n4713 ;
  assign n5383 = ~n1338 & n4712 ;
  assign n5384 = n1458 & n4792 ;
  assign n5385 = n1576 & n4709 ;
  assign n5386 = n5384 | n5385 ;
  assign n5387 = ( ~n5382 & n5383 ) | ( ~n5382 & n5386 ) | ( n5383 & n5386 ) ;
  assign n5388 = ( ~x23 & n5382 ) | ( ~x23 & n5387 ) | ( n5382 & n5387 ) ;
  assign n5389 = ( n5382 & n5387 ) | ( n5382 & ~n5388 ) | ( n5387 & ~n5388 ) ;
  assign n5390 = ( x23 & n5388 ) | ( x23 & ~n5389 ) | ( n5388 & ~n5389 ) ;
  assign n5391 = ( n5379 & n5381 ) | ( n5379 & n5390 ) | ( n5381 & n5390 ) ;
  assign n5392 = ( ~n5312 & n5314 ) | ( ~n5312 & n5323 ) | ( n5314 & n5323 ) ;
  assign n5393 = ( ~n5323 & n5324 ) | ( ~n5323 & n5392 ) | ( n5324 & n5392 ) ;
  assign n5394 = ~n3665 & n4974 ;
  assign n5395 = ~n1290 & n4972 ;
  assign n5396 = ~n1246 & n4973 ;
  assign n5397 = ~n4967 & n4968 ;
  assign n5398 = ( ~n4964 & n4965 ) | ( ~n4964 & n5397 ) | ( n4965 & n5397 ) ;
  assign n5399 = ~n3658 & n5398 ;
  assign n5400 = n5396 | n5399 ;
  assign n5401 = ( ~n5394 & n5395 ) | ( ~n5394 & n5400 ) | ( n5395 & n5400 ) ;
  assign n5402 = ( ~x20 & n5394 ) | ( ~x20 & n5401 ) | ( n5394 & n5401 ) ;
  assign n5403 = ( n5394 & n5401 ) | ( n5394 & ~n5402 ) | ( n5401 & ~n5402 ) ;
  assign n5404 = ( x20 & n5402 ) | ( x20 & ~n5403 ) | ( n5402 & ~n5403 ) ;
  assign n5405 = ( n5391 & ~n5393 ) | ( n5391 & n5404 ) | ( ~n5393 & n5404 ) ;
  assign n5406 = n3692 & n5398 ;
  assign n5407 = ~n3658 & n4972 ;
  assign n5408 = ( n5398 & ~n5406 ) | ( n5398 & n5407 ) | ( ~n5406 & n5407 ) ;
  assign n5409 = ~n1290 & n4973 ;
  assign n5410 = n5408 | n5409 ;
  assign n5411 = ~n4182 & n4974 ;
  assign n5412 = ( x20 & n5410 ) | ( x20 & ~n5411 ) | ( n5410 & ~n5411 ) ;
  assign n5413 = ( ~x20 & n5410 ) | ( ~x20 & n5411 ) | ( n5410 & n5411 ) ;
  assign n5414 = ( ~n5410 & n5412 ) | ( ~n5410 & n5413 ) | ( n5412 & n5413 ) ;
  assign n5415 = ( ~n5324 & n5333 ) | ( ~n5324 & n5335 ) | ( n5333 & n5335 ) ;
  assign n5416 = ( n5324 & ~n5336 ) | ( n5324 & n5415 ) | ( ~n5336 & n5415 ) ;
  assign n5417 = ( n5405 & n5414 ) | ( n5405 & n5416 ) | ( n5414 & n5416 ) ;
  assign n5418 = ( n5030 & n5235 ) | ( n5030 & n5259 ) | ( n5235 & n5259 ) ;
  assign n5419 = ( n5259 & n5260 ) | ( n5259 & ~n5418 ) | ( n5260 & ~n5418 ) ;
  assign n5420 = n607 | n2725 ;
  assign n5421 = n1250 & n2635 ;
  assign n5422 = ( ~n2725 & n5420 ) | ( ~n2725 & n5421 ) | ( n5420 & n5421 ) ;
  assign n5423 = n606 & ~n2552 ;
  assign n5424 = ( n606 & n5422 ) | ( n606 & ~n5423 ) | ( n5422 & ~n5423 ) ;
  assign n5425 = ( ~n2635 & n3602 ) | ( ~n2635 & n5268 ) | ( n3602 & n5268 ) ;
  assign n5426 = n1248 & ~n5425 ;
  assign n5427 = n5424 | n5426 ;
  assign n5428 = n3800 & ~n4900 ;
  assign n5429 = n2396 & n3802 ;
  assign n5430 = ~n2298 & n3799 ;
  assign n5431 = ( n2491 & n3694 ) | ( n2491 & n3699 ) | ( n3694 & n3699 ) ;
  assign n5432 = ( n3694 & n5430 ) | ( n3694 & ~n5431 ) | ( n5430 & ~n5431 ) ;
  assign n5433 = ( ~n5428 & n5429 ) | ( ~n5428 & n5432 ) | ( n5429 & n5432 ) ;
  assign n5434 = ( ~x29 & n5428 ) | ( ~x29 & n5433 ) | ( n5428 & n5433 ) ;
  assign n5435 = ( n5428 & n5433 ) | ( n5428 & ~n5434 ) | ( n5433 & ~n5434 ) ;
  assign n5436 = ( x29 & n5434 ) | ( x29 & ~n5435 ) | ( n5434 & ~n5435 ) ;
  assign n5437 = ( n5419 & n5427 ) | ( n5419 & n5436 ) | ( n5427 & n5436 ) ;
  assign n5438 = ( n5260 & ~n5262 ) | ( n5260 & n5272 ) | ( ~n5262 & n5272 ) ;
  assign n5439 = ( ~n5260 & n5273 ) | ( ~n5260 & n5438 ) | ( n5273 & n5438 ) ;
  assign n5440 = n3800 & ~n4912 ;
  assign n5441 = n2396 & n3700 ;
  assign n5442 = n2298 | n3802 ;
  assign n5443 = n2270 & n3799 ;
  assign n5444 = ( ~n2298 & n5442 ) | ( ~n2298 & n5443 ) | ( n5442 & n5443 ) ;
  assign n5445 = ( ~n5440 & n5441 ) | ( ~n5440 & n5444 ) | ( n5441 & n5444 ) ;
  assign n5446 = ( ~x29 & n5440 ) | ( ~x29 & n5445 ) | ( n5440 & n5445 ) ;
  assign n5447 = ( n5440 & n5445 ) | ( n5440 & ~n5446 ) | ( n5445 & ~n5446 ) ;
  assign n5448 = ( x29 & n5446 ) | ( x29 & ~n5447 ) | ( n5446 & ~n5447 ) ;
  assign n5449 = ( n5437 & n5439 ) | ( n5437 & n5448 ) | ( n5439 & n5448 ) ;
  assign n5450 = ( n5273 & ~n5275 ) | ( n5273 & n5284 ) | ( ~n5275 & n5284 ) ;
  assign n5451 = ( ~n5273 & n5285 ) | ( ~n5273 & n5450 ) | ( n5285 & n5450 ) ;
  assign n5452 = n4202 & ~n4457 ;
  assign n5453 = n1926 & n4201 ;
  assign n5454 = ~n2023 & n4345 ;
  assign n5455 = n2089 & n4200 ;
  assign n5456 = n5454 | n5455 ;
  assign n5457 = ( ~n5452 & n5453 ) | ( ~n5452 & n5456 ) | ( n5453 & n5456 ) ;
  assign n5458 = ( ~x26 & n5452 ) | ( ~x26 & n5457 ) | ( n5452 & n5457 ) ;
  assign n5459 = ( n5452 & n5457 ) | ( n5452 & ~n5458 ) | ( n5457 & ~n5458 ) ;
  assign n5460 = ( x26 & n5458 ) | ( x26 & ~n5459 ) | ( n5458 & ~n5459 ) ;
  assign n5461 = ( n5449 & n5451 ) | ( n5449 & n5460 ) | ( n5451 & n5460 ) ;
  assign n5462 = ( n5348 & ~n5357 ) | ( n5348 & n5366 ) | ( ~n5357 & n5366 ) ;
  assign n5463 = ( n5357 & ~n5367 ) | ( n5357 & n5462 ) | ( ~n5367 & n5462 ) ;
  assign n5464 = n4326 & n4713 ;
  assign n5465 = n1576 & n4712 ;
  assign n5466 = n1750 | n4709 ;
  assign n5467 = ~n1669 & n4792 ;
  assign n5468 = ( ~n1750 & n5466 ) | ( ~n1750 & n5467 ) | ( n5466 & n5467 ) ;
  assign n5469 = ( ~n5464 & n5465 ) | ( ~n5464 & n5468 ) | ( n5465 & n5468 ) ;
  assign n5470 = ( ~x23 & n5464 ) | ( ~x23 & n5469 ) | ( n5464 & n5469 ) ;
  assign n5471 = ( n5464 & n5469 ) | ( n5464 & ~n5470 ) | ( n5469 & ~n5470 ) ;
  assign n5472 = ( x23 & n5470 ) | ( x23 & ~n5471 ) | ( n5470 & ~n5471 ) ;
  assign n5473 = ( n5461 & n5463 ) | ( n5461 & n5472 ) | ( n5463 & n5472 ) ;
  assign n5474 = ~n4159 & n4713 ;
  assign n5475 = n1458 & n4712 ;
  assign n5476 = ~n1669 & n4709 ;
  assign n5477 = n1576 & n4792 ;
  assign n5478 = n5476 | n5477 ;
  assign n5479 = ( ~n5474 & n5475 ) | ( ~n5474 & n5478 ) | ( n5475 & n5478 ) ;
  assign n5480 = ( ~x23 & n5474 ) | ( ~x23 & n5479 ) | ( n5474 & n5479 ) ;
  assign n5481 = ( n5474 & n5479 ) | ( n5474 & ~n5480 ) | ( n5479 & ~n5480 ) ;
  assign n5482 = ( x23 & n5480 ) | ( x23 & ~n5481 ) | ( n5480 & ~n5481 ) ;
  assign n5483 = ( ~n5367 & n5369 ) | ( ~n5367 & n5378 ) | ( n5369 & n5378 ) ;
  assign n5484 = ( ~n5378 & n5379 ) | ( ~n5378 & n5483 ) | ( n5379 & n5483 ) ;
  assign n5485 = ( n5473 & n5482 ) | ( n5473 & ~n5484 ) | ( n5482 & ~n5484 ) ;
  assign n5486 = ( n5379 & ~n5381 ) | ( n5379 & n5390 ) | ( ~n5381 & n5390 ) ;
  assign n5487 = ( n5381 & ~n5391 ) | ( n5381 & n5486 ) | ( ~n5391 & n5486 ) ;
  assign n5488 = n3621 & n4974 ;
  assign n5489 = ~n1290 & n5398 ;
  assign n5490 = n1267 & ~n4973 ;
  assign n5491 = ~n1246 & n4972 ;
  assign n5492 = ( n1267 & ~n5490 ) | ( n1267 & n5491 ) | ( ~n5490 & n5491 ) ;
  assign n5493 = ( ~n5488 & n5489 ) | ( ~n5488 & n5492 ) | ( n5489 & n5492 ) ;
  assign n5494 = ( ~x20 & n5488 ) | ( ~x20 & n5493 ) | ( n5488 & n5493 ) ;
  assign n5495 = ( n5488 & n5493 ) | ( n5488 & ~n5494 ) | ( n5493 & ~n5494 ) ;
  assign n5496 = ( x20 & n5494 ) | ( x20 & ~n5495 ) | ( n5494 & ~n5495 ) ;
  assign n5497 = ( n5485 & n5487 ) | ( n5485 & n5496 ) | ( n5487 & n5496 ) ;
  assign n5498 = x14 | x15 ;
  assign n5499 = x15 & x16 ;
  assign n5500 = x16 | x17 ;
  assign n5501 = x16 & x17 ;
  assign n5502 = n5500 & ~n5501 ;
  assign n5503 = ( x14 & ~x16 ) | ( x14 & n5502 ) | ( ~x16 & n5502 ) ;
  assign n5504 = ( ~n5498 & n5499 ) | ( ~n5498 & n5503 ) | ( n5499 & n5503 ) ;
  assign n5505 = x14 & x15 ;
  assign n5506 = n5498 & ~n5505 ;
  assign n5507 = ( ~n5500 & n5501 ) | ( ~n5500 & n5506 ) | ( n5501 & n5506 ) ;
  assign n5508 = n5506 & ~n5507 ;
  assign n5509 = ~n3691 & n5508 ;
  assign n5510 = ( ~n3692 & n5504 ) | ( ~n3692 & n5509 ) | ( n5504 & n5509 ) ;
  assign n5511 = x17 | n5510 ;
  assign n5512 = ( x17 & n5510 ) | ( x17 & ~n5511 ) | ( n5510 & ~n5511 ) ;
  assign n5513 = n5511 & ~n5512 ;
  assign n5514 = ( ~n5391 & n5393 ) | ( ~n5391 & n5404 ) | ( n5393 & n5404 ) ;
  assign n5515 = ( ~n5404 & n5405 ) | ( ~n5404 & n5514 ) | ( n5405 & n5514 ) ;
  assign n5516 = ( n5497 & n5513 ) | ( n5497 & ~n5515 ) | ( n5513 & ~n5515 ) ;
  assign n5517 = n242 | n258 ;
  assign n5518 = ( n1544 & n2496 ) | ( n1544 & ~n2527 ) | ( n2496 & ~n2527 ) ;
  assign n5519 = n2527 | n5518 ;
  assign n5520 = ( n933 & ~n5517 ) | ( n933 & n5519 ) | ( ~n5517 & n5519 ) ;
  assign n5521 = n5517 | n5520 ;
  assign n5522 = ( n846 & n1641 ) | ( n846 & ~n4581 ) | ( n1641 & ~n4581 ) ;
  assign n5523 = n4581 | n5522 ;
  assign n5524 = n1002 | n2158 ;
  assign n5525 = ( n697 & n1005 ) | ( n697 & ~n5524 ) | ( n1005 & ~n5524 ) ;
  assign n5526 = n5524 | n5525 ;
  assign n5527 = ( n59 & n64 ) | ( n59 & n72 ) | ( n64 & n72 ) ;
  assign n5528 = n2790 | n3258 ;
  assign n5529 = ( n1592 & ~n5527 ) | ( n1592 & n5528 ) | ( ~n5527 & n5528 ) ;
  assign n5530 = ( n1879 & n3727 ) | ( n1879 & ~n5527 ) | ( n3727 & ~n5527 ) ;
  assign n5531 = n5527 | n5530 ;
  assign n5532 = ( ~n5526 & n5529 ) | ( ~n5526 & n5531 ) | ( n5529 & n5531 ) ;
  assign n5533 = n5526 | n5532 ;
  assign n5534 = ( ~n5521 & n5523 ) | ( ~n5521 & n5533 ) | ( n5523 & n5533 ) ;
  assign n5535 = n5521 | n5534 ;
  assign n5536 = ( x2 & x5 ) | ( x2 & ~n5535 ) | ( x5 & ~n5535 ) ;
  assign n5537 = n607 & ~n2965 ;
  assign n5538 = n606 & n2843 ;
  assign n5539 = n5537 | n5538 ;
  assign n5540 = n1250 | n2910 ;
  assign n5541 = ( ~n2910 & n5539 ) | ( ~n2910 & n5540 ) | ( n5539 & n5540 ) ;
  assign n5542 = ( n2843 & n2910 ) | ( n2843 & n3597 ) | ( n2910 & n3597 ) ;
  assign n5543 = ( n2843 & n3598 ) | ( n2843 & ~n5542 ) | ( n3598 & ~n5542 ) ;
  assign n5544 = n1248 & n5543 ;
  assign n5545 = n5541 | n5544 ;
  assign n5546 = ( n5163 & ~n5536 ) | ( n5163 & n5545 ) | ( ~n5536 & n5545 ) ;
  assign n5547 = n189 | n1174 ;
  assign n5548 = n254 | n582 ;
  assign n5549 = ( n131 & n912 ) | ( n131 & ~n5548 ) | ( n912 & ~n5548 ) ;
  assign n5550 = n5548 | n5549 ;
  assign n5551 = ( n657 & ~n5547 ) | ( n657 & n5550 ) | ( ~n5547 & n5550 ) ;
  assign n5552 = n5547 | n5551 ;
  assign n5553 = ( n48 & n84 ) | ( n48 & n149 ) | ( n84 & n149 ) ;
  assign n5554 = n265 | n5553 ;
  assign n5555 = n5144 | n5554 ;
  assign n5556 = n1860 | n4389 ;
  assign n5557 = n1510 | n1737 ;
  assign n5558 = ( n5212 & ~n5556 ) | ( n5212 & n5557 ) | ( ~n5556 & n5557 ) ;
  assign n5559 = n5556 | n5558 ;
  assign n5560 = ( ~n5552 & n5555 ) | ( ~n5552 & n5559 ) | ( n5555 & n5559 ) ;
  assign n5561 = n5552 | n5560 ;
  assign n5562 = n1987 | n4112 ;
  assign n5563 = n1452 | n3817 ;
  assign n5564 = n5194 | n5563 ;
  assign n5565 = ( ~n1452 & n2163 ) | ( ~n1452 & n2414 ) | ( n2163 & n2414 ) ;
  assign n5566 = n92 | n293 ;
  assign n5567 = ( n586 & n1346 ) | ( n586 & ~n5566 ) | ( n1346 & ~n5566 ) ;
  assign n5568 = n5566 | n5567 ;
  assign n5569 = ( ~n5563 & n5565 ) | ( ~n5563 & n5568 ) | ( n5565 & n5568 ) ;
  assign n5570 = ( n2628 & n4069 ) | ( n2628 & ~n5569 ) | ( n4069 & ~n5569 ) ;
  assign n5571 = n5569 | n5570 ;
  assign n5572 = ( n267 & ~n1547 ) | ( n267 & n1660 ) | ( ~n1547 & n1660 ) ;
  assign n5573 = n1547 | n5572 ;
  assign n5574 = ( ~n5564 & n5571 ) | ( ~n5564 & n5573 ) | ( n5571 & n5573 ) ;
  assign n5575 = n5564 | n5574 ;
  assign n5576 = ( ~n5561 & n5562 ) | ( ~n5561 & n5575 ) | ( n5562 & n5575 ) ;
  assign n5577 = n5561 | n5576 ;
  assign n5578 = ( n5163 & n5546 ) | ( n5163 & n5577 ) | ( n5546 & n5577 ) ;
  assign n5579 = ( x8 & ~n5163 ) | ( x8 & n5222 ) | ( ~n5163 & n5222 ) ;
  assign n5580 = ( ~x8 & n5223 ) | ( ~x8 & n5579 ) | ( n5223 & n5579 ) ;
  assign n5581 = ~n607 & n2843 ;
  assign n5582 = n1250 & ~n2810 ;
  assign n5583 = ( n2843 & ~n5581 ) | ( n2843 & n5582 ) | ( ~n5581 & n5582 ) ;
  assign n5584 = n606 & n2725 ;
  assign n5585 = ( n606 & n5583 ) | ( n606 & ~n5584 ) | ( n5583 & ~n5584 ) ;
  assign n5586 = ( n2810 & ~n3600 ) | ( n2810 & n5230 ) | ( ~n3600 & n5230 ) ;
  assign n5587 = n1248 & ~n5586 ;
  assign n5588 = n5585 | n5587 ;
  assign n5589 = ( n5578 & n5580 ) | ( n5578 & n5588 ) | ( n5580 & n5588 ) ;
  assign n5590 = ( n5030 & n5223 ) | ( n5030 & n5234 ) | ( n5223 & n5234 ) ;
  assign n5591 = ( n5234 & n5235 ) | ( n5234 & ~n5590 ) | ( n5235 & ~n5590 ) ;
  assign n5592 = n3800 & ~n5084 ;
  assign n5593 = n2396 & n3799 ;
  assign n5594 = ~n2491 & n3802 ;
  assign n5595 = ( ~n2552 & n3694 ) | ( ~n2552 & n3699 ) | ( n3694 & n3699 ) ;
  assign n5596 = ( n3694 & n5594 ) | ( n3694 & ~n5595 ) | ( n5594 & ~n5595 ) ;
  assign n5597 = ( ~n5592 & n5593 ) | ( ~n5592 & n5596 ) | ( n5593 & n5596 ) ;
  assign n5598 = ( ~x29 & n5592 ) | ( ~x29 & n5597 ) | ( n5592 & n5597 ) ;
  assign n5599 = ( n5592 & n5597 ) | ( n5592 & ~n5598 ) | ( n5597 & ~n5598 ) ;
  assign n5600 = ( x29 & n5598 ) | ( x29 & ~n5599 ) | ( n5598 & ~n5599 ) ;
  assign n5601 = ( n5589 & n5591 ) | ( n5589 & n5600 ) | ( n5591 & n5600 ) ;
  assign n5602 = ( n5419 & ~n5427 ) | ( n5419 & n5436 ) | ( ~n5427 & n5436 ) ;
  assign n5603 = ( n5427 & ~n5437 ) | ( n5427 & n5602 ) | ( ~n5437 & n5602 ) ;
  assign n5604 = n4202 & n4730 ;
  assign n5605 = n2089 & n4201 ;
  assign n5606 = n2270 & n4200 ;
  assign n5607 = n2174 & n4345 ;
  assign n5608 = n5606 | n5607 ;
  assign n5609 = ( ~n5604 & n5605 ) | ( ~n5604 & n5608 ) | ( n5605 & n5608 ) ;
  assign n5610 = ( ~x26 & n5604 ) | ( ~x26 & n5609 ) | ( n5604 & n5609 ) ;
  assign n5611 = ( n5604 & n5609 ) | ( n5604 & ~n5610 ) | ( n5609 & ~n5610 ) ;
  assign n5612 = ( x26 & n5610 ) | ( x26 & ~n5611 ) | ( n5610 & ~n5611 ) ;
  assign n5613 = ( n5601 & n5603 ) | ( n5601 & n5612 ) | ( n5603 & n5612 ) ;
  assign n5614 = ( n5437 & ~n5439 ) | ( n5437 & n5448 ) | ( ~n5439 & n5448 ) ;
  assign n5615 = ( n5439 & ~n5449 ) | ( n5439 & n5614 ) | ( ~n5449 & n5614 ) ;
  assign n5616 = n4202 & ~n4660 ;
  assign n5617 = ~n2023 & n4201 ;
  assign n5618 = n2174 & n4200 ;
  assign n5619 = n2089 & n4345 ;
  assign n5620 = n5618 | n5619 ;
  assign n5621 = ( ~n5616 & n5617 ) | ( ~n5616 & n5620 ) | ( n5617 & n5620 ) ;
  assign n5622 = ( ~x26 & n5616 ) | ( ~x26 & n5621 ) | ( n5616 & n5621 ) ;
  assign n5623 = ( n5616 & n5621 ) | ( n5616 & ~n5622 ) | ( n5621 & ~n5622 ) ;
  assign n5624 = ( x26 & n5622 ) | ( x26 & ~n5623 ) | ( n5622 & ~n5623 ) ;
  assign n5625 = ( n5613 & n5615 ) | ( n5613 & n5624 ) | ( n5615 & n5624 ) ;
  assign n5626 = ( ~n5449 & n5451 ) | ( ~n5449 & n5460 ) | ( n5451 & n5460 ) ;
  assign n5627 = ( n5449 & ~n5461 ) | ( n5449 & n5626 ) | ( ~n5461 & n5626 ) ;
  assign n5628 = n4146 & n4713 ;
  assign n5629 = ~n1669 & n4712 ;
  assign n5630 = n1852 & ~n4709 ;
  assign n5631 = ~n1750 & n4792 ;
  assign n5632 = ( n1852 & ~n5630 ) | ( n1852 & n5631 ) | ( ~n5630 & n5631 ) ;
  assign n5633 = ( ~n5628 & n5629 ) | ( ~n5628 & n5632 ) | ( n5629 & n5632 ) ;
  assign n5634 = ( ~x23 & n5628 ) | ( ~x23 & n5633 ) | ( n5628 & n5633 ) ;
  assign n5635 = ( n5628 & n5633 ) | ( n5628 & ~n5634 ) | ( n5633 & ~n5634 ) ;
  assign n5636 = ( x23 & n5634 ) | ( x23 & ~n5635 ) | ( n5634 & ~n5635 ) ;
  assign n5637 = ( n5625 & n5627 ) | ( n5625 & n5636 ) | ( n5627 & n5636 ) ;
  assign n5638 = ( ~n5461 & n5463 ) | ( ~n5461 & n5472 ) | ( n5463 & n5472 ) ;
  assign n5639 = ( n5461 & ~n5473 ) | ( n5461 & n5638 ) | ( ~n5473 & n5638 ) ;
  assign n5640 = ~n3779 & n4974 ;
  assign n5641 = n1267 & n5398 ;
  assign n5642 = n1458 & ~n4973 ;
  assign n5643 = ~n1338 & n4972 ;
  assign n5644 = ( n1458 & ~n5642 ) | ( n1458 & n5643 ) | ( ~n5642 & n5643 ) ;
  assign n5645 = ( ~n5640 & n5641 ) | ( ~n5640 & n5644 ) | ( n5641 & n5644 ) ;
  assign n5646 = ( ~x20 & n5640 ) | ( ~x20 & n5645 ) | ( n5640 & n5645 ) ;
  assign n5647 = ( n5640 & n5645 ) | ( n5640 & ~n5646 ) | ( n5645 & ~n5646 ) ;
  assign n5648 = ( x20 & n5646 ) | ( x20 & ~n5647 ) | ( n5646 & ~n5647 ) ;
  assign n5649 = ( n5637 & n5639 ) | ( n5637 & n5648 ) | ( n5639 & n5648 ) ;
  assign n5650 = ( n5473 & ~n5482 ) | ( n5473 & n5484 ) | ( ~n5482 & n5484 ) ;
  assign n5651 = ( ~n5473 & n5485 ) | ( ~n5473 & n5650 ) | ( n5485 & n5650 ) ;
  assign n5652 = ~n3791 & n4974 ;
  assign n5653 = n1267 & n4972 ;
  assign n5654 = n1338 | n4973 ;
  assign n5655 = ~n1246 & n5398 ;
  assign n5656 = ( ~n1338 & n5654 ) | ( ~n1338 & n5655 ) | ( n5654 & n5655 ) ;
  assign n5657 = ( ~n5652 & n5653 ) | ( ~n5652 & n5656 ) | ( n5653 & n5656 ) ;
  assign n5658 = ( ~x20 & n5652 ) | ( ~x20 & n5657 ) | ( n5652 & n5657 ) ;
  assign n5659 = ( n5652 & n5657 ) | ( n5652 & ~n5658 ) | ( n5657 & ~n5658 ) ;
  assign n5660 = ( x20 & n5658 ) | ( x20 & ~n5659 ) | ( n5658 & ~n5659 ) ;
  assign n5661 = ( n5649 & ~n5651 ) | ( n5649 & n5660 ) | ( ~n5651 & n5660 ) ;
  assign n5662 = ( n5485 & ~n5487 ) | ( n5485 & n5496 ) | ( ~n5487 & n5496 ) ;
  assign n5663 = ( n5487 & ~n5497 ) | ( n5487 & n5662 ) | ( ~n5497 & n5662 ) ;
  assign n5664 = n3797 & n5508 ;
  assign n5665 = ~x14 & x16 ;
  assign n5666 = ( ~n5499 & n5505 ) | ( ~n5499 & n5665 ) | ( n5505 & n5665 ) ;
  assign n5667 = ~n3692 & n5666 ;
  assign n5668 = ~n3658 & n5504 ;
  assign n5669 = n5667 | n5668 ;
  assign n5670 = ( ~x17 & n5664 ) | ( ~x17 & n5669 ) | ( n5664 & n5669 ) ;
  assign n5671 = ( n5664 & n5669 ) | ( n5664 & ~n5670 ) | ( n5669 & ~n5670 ) ;
  assign n5672 = ( x17 & n5670 ) | ( x17 & ~n5671 ) | ( n5670 & ~n5671 ) ;
  assign n5673 = ( n5661 & n5663 ) | ( n5661 & n5672 ) | ( n5663 & n5672 ) ;
  assign n5674 = n167 | n402 ;
  assign n5675 = ( n66 & n152 ) | ( n66 & n160 ) | ( n152 & n160 ) ;
  assign n5676 = n675 | n5675 ;
  assign n5677 = ( n1526 & ~n5674 ) | ( n1526 & n5676 ) | ( ~n5674 & n5676 ) ;
  assign n5678 = n5674 | n5677 ;
  assign n5679 = n884 | n958 ;
  assign n5680 = ( n4463 & n4828 ) | ( n4463 & ~n5679 ) | ( n4828 & ~n5679 ) ;
  assign n5681 = n5679 | n5680 ;
  assign n5682 = n775 | n1718 ;
  assign n5683 = n299 | n5682 ;
  assign n5684 = ( n3104 & n3569 ) | ( n3104 & ~n5683 ) | ( n3569 & ~n5683 ) ;
  assign n5685 = n5683 | n5684 ;
  assign n5686 = ( ~n5678 & n5681 ) | ( ~n5678 & n5685 ) | ( n5681 & n5685 ) ;
  assign n5687 = n5678 | n5686 ;
  assign n5688 = ( ~n910 & n989 ) | ( ~n910 & n2373 ) | ( n989 & n2373 ) ;
  assign n5689 = n910 | n5688 ;
  assign n5690 = n1560 | n3416 ;
  assign n5691 = n260 | n383 ;
  assign n5692 = ( n923 & n2399 ) | ( n923 & ~n5691 ) | ( n2399 & ~n5691 ) ;
  assign n5693 = n5691 | n5692 ;
  assign n5694 = n1799 | n5154 ;
  assign n5695 = n231 | n1059 ;
  assign n5696 = ( n142 & n806 ) | ( n142 & ~n5695 ) | ( n806 & ~n5695 ) ;
  assign n5697 = n5695 | n5696 ;
  assign n5698 = ( ~n5693 & n5694 ) | ( ~n5693 & n5697 ) | ( n5694 & n5697 ) ;
  assign n5699 = n5693 | n5698 ;
  assign n5700 = ( n5241 & ~n5690 ) | ( n5241 & n5699 ) | ( ~n5690 & n5699 ) ;
  assign n5701 = n5690 | n5700 ;
  assign n5702 = ( ~n5687 & n5689 ) | ( ~n5687 & n5701 ) | ( n5689 & n5701 ) ;
  assign n5703 = n5687 | n5702 ;
  assign n5704 = n606 & n3078 ;
  assign n5705 = n607 & n3239 ;
  assign n5706 = n5704 | n5705 ;
  assign n5707 = ~n1250 & n3153 ;
  assign n5708 = ( n3153 & n5706 ) | ( n3153 & ~n5707 ) | ( n5706 & ~n5707 ) ;
  assign n5709 = ( n3078 & n3153 ) | ( n3078 & ~n3593 ) | ( n3153 & ~n3593 ) ;
  assign n5710 = ( n3593 & ~n3594 ) | ( n3593 & n5709 ) | ( ~n3594 & n5709 ) ;
  assign n5711 = n1248 & n5710 ;
  assign n5712 = n5708 | n5711 ;
  assign n5713 = ( x2 & n5703 ) | ( x2 & n5712 ) | ( n5703 & n5712 ) ;
  assign n5714 = n1687 | n3428 ;
  assign n5715 = n91 | n641 ;
  assign n5716 = ( n545 & n697 ) | ( n545 & ~n5715 ) | ( n697 & ~n5715 ) ;
  assign n5717 = n5715 | n5716 ;
  assign n5718 = n1380 | n1595 ;
  assign n5719 = n441 | n4238 ;
  assign n5720 = n5718 | n5719 ;
  assign n5721 = n5717 | n5720 ;
  assign n5722 = ( n1277 & n1891 ) | ( n1277 & ~n3841 ) | ( n1891 & ~n3841 ) ;
  assign n5723 = n3841 | n5722 ;
  assign n5724 = n2431 | n4872 ;
  assign n5725 = n261 | n519 ;
  assign n5726 = ( n1655 & ~n5724 ) | ( n1655 & n5725 ) | ( ~n5724 & n5725 ) ;
  assign n5727 = n5724 | n5726 ;
  assign n5728 = ( n4465 & ~n5723 ) | ( n4465 & n5727 ) | ( ~n5723 & n5727 ) ;
  assign n5729 = n5723 | n5728 ;
  assign n5730 = ( ~n1687 & n5721 ) | ( ~n1687 & n5729 ) | ( n5721 & n5729 ) ;
  assign n5731 = ( ~n861 & n5714 ) | ( ~n861 & n5730 ) | ( n5714 & n5730 ) ;
  assign n5732 = n861 | n5731 ;
  assign n5733 = ( x2 & n5713 ) | ( x2 & n5732 ) | ( n5713 & n5732 ) ;
  assign n5734 = n5066 | n5243 ;
  assign n5735 = n549 | n1225 ;
  assign n5736 = n535 | n3523 ;
  assign n5737 = ( n420 & ~n1441 ) | ( n420 & n5736 ) | ( ~n1441 & n5736 ) ;
  assign n5738 = n1441 | n5737 ;
  assign n5739 = ( n856 & ~n5735 ) | ( n856 & n5738 ) | ( ~n5735 & n5738 ) ;
  assign n5740 = n5735 | n5739 ;
  assign n5741 = n286 | n760 ;
  assign n5742 = ( n1277 & n1560 ) | ( n1277 & ~n5741 ) | ( n1560 & ~n5741 ) ;
  assign n5743 = n5741 | n5742 ;
  assign n5744 = ( ~n5734 & n5740 ) | ( ~n5734 & n5743 ) | ( n5740 & n5743 ) ;
  assign n5745 = n5734 | n5744 ;
  assign n5746 = n638 | n1027 ;
  assign n5747 = ( n57 & n84 ) | ( n57 & n149 ) | ( n84 & n149 ) ;
  assign n5748 = n488 | n5747 ;
  assign n5749 = ( n3030 & ~n5746 ) | ( n3030 & n5748 ) | ( ~n5746 & n5748 ) ;
  assign n5750 = n5746 | n5749 ;
  assign n5751 = n884 | n3734 ;
  assign n5752 = n4495 | n5751 ;
  assign n5753 = ( n5745 & ~n5750 ) | ( n5745 & n5752 ) | ( ~n5750 & n5752 ) ;
  assign n5754 = ( n2203 & n5750 ) | ( n2203 & ~n5753 ) | ( n5750 & ~n5753 ) ;
  assign n5755 = n5753 | n5754 ;
  assign n5756 = ( n3014 & n3297 ) | ( n3014 & n5755 ) | ( n3297 & n5755 ) ;
  assign n5757 = ( ~n1434 & n3297 ) | ( ~n1434 & n5756 ) | ( n3297 & n5756 ) ;
  assign n5758 = ~n5756 & n5757 ;
  assign n5759 = ( x2 & n5733 ) | ( x2 & ~n5758 ) | ( n5733 & ~n5758 ) ;
  assign n5760 = ( x2 & ~x5 ) | ( x2 & n5535 ) | ( ~x5 & n5535 ) ;
  assign n5761 = ( ~x2 & n5536 ) | ( ~x2 & n5760 ) | ( n5536 & n5760 ) ;
  assign n5762 = n607 | n3046 ;
  assign n5763 = n1250 & ~n2965 ;
  assign n5764 = ( ~n3046 & n5762 ) | ( ~n3046 & n5763 ) | ( n5762 & n5763 ) ;
  assign n5765 = n606 & n2910 ;
  assign n5766 = ( n606 & n5764 ) | ( n606 & ~n5765 ) | ( n5764 & ~n5765 ) ;
  assign n5767 = ( n2910 & n2965 ) | ( n2910 & ~n3596 ) | ( n2965 & ~n3596 ) ;
  assign n5768 = ( n3596 & ~n3597 ) | ( n3596 & n5767 ) | ( ~n3597 & n5767 ) ;
  assign n5769 = n1248 & ~n5768 ;
  assign n5770 = n5766 | n5769 ;
  assign n5771 = ( n5759 & n5761 ) | ( n5759 & n5770 ) | ( n5761 & n5770 ) ;
  assign n5772 = ( n5163 & n5545 ) | ( n5163 & ~n5546 ) | ( n5545 & ~n5546 ) ;
  assign n5773 = ( n5536 & n5546 ) | ( n5536 & ~n5772 ) | ( n5546 & ~n5772 ) ;
  assign n5774 = n3800 & n5232 ;
  assign n5775 = ~n2810 & n3700 ;
  assign n5776 = n2725 | n3802 ;
  assign n5777 = n2635 & n3799 ;
  assign n5778 = ( ~n2725 & n5776 ) | ( ~n2725 & n5777 ) | ( n5776 & n5777 ) ;
  assign n5779 = ( ~n5774 & n5775 ) | ( ~n5774 & n5778 ) | ( n5775 & n5778 ) ;
  assign n5780 = ( ~x29 & n5774 ) | ( ~x29 & n5779 ) | ( n5774 & n5779 ) ;
  assign n5781 = ( n5774 & n5779 ) | ( n5774 & ~n5780 ) | ( n5779 & ~n5780 ) ;
  assign n5782 = ( x29 & n5780 ) | ( x29 & ~n5781 ) | ( n5780 & ~n5781 ) ;
  assign n5783 = ( n5771 & ~n5773 ) | ( n5771 & n5782 ) | ( ~n5773 & n5782 ) ;
  assign n5784 = ( ~n5163 & n5546 ) | ( ~n5163 & n5577 ) | ( n5546 & n5577 ) ;
  assign n5785 = ( n5163 & ~n5578 ) | ( n5163 & n5784 ) | ( ~n5578 & n5784 ) ;
  assign n5786 = n607 | n2910 ;
  assign n5787 = n1250 & n2843 ;
  assign n5788 = ( ~n2910 & n5786 ) | ( ~n2910 & n5787 ) | ( n5786 & n5787 ) ;
  assign n5789 = n606 & n2810 ;
  assign n5790 = ( n606 & n5788 ) | ( n606 & ~n5789 ) | ( n5788 & ~n5789 ) ;
  assign n5791 = ( ~n3598 & n3599 ) | ( ~n3598 & n5229 ) | ( n3599 & n5229 ) ;
  assign n5792 = n1248 & n5791 ;
  assign n5793 = n5790 | n5792 ;
  assign n5794 = ( n5783 & n5785 ) | ( n5783 & n5793 ) | ( n5785 & n5793 ) ;
  assign n5795 = n3800 & ~n5270 ;
  assign n5796 = n2552 & n3802 ;
  assign n5797 = ~n2491 & n3799 ;
  assign n5798 = ( ~n2635 & n3694 ) | ( ~n2635 & n3699 ) | ( n3694 & n3699 ) ;
  assign n5799 = ( n3694 & n5797 ) | ( n3694 & ~n5798 ) | ( n5797 & ~n5798 ) ;
  assign n5800 = ( ~n5795 & n5796 ) | ( ~n5795 & n5799 ) | ( n5796 & n5799 ) ;
  assign n5801 = ( ~x29 & n5795 ) | ( ~x29 & n5800 ) | ( n5795 & n5800 ) ;
  assign n5802 = ( n5795 & n5800 ) | ( n5795 & ~n5801 ) | ( n5800 & ~n5801 ) ;
  assign n5803 = ( x29 & n5801 ) | ( x29 & ~n5802 ) | ( n5801 & ~n5802 ) ;
  assign n5804 = ( n5578 & ~n5580 ) | ( n5578 & n5588 ) | ( ~n5580 & n5588 ) ;
  assign n5805 = ( n5580 & ~n5589 ) | ( n5580 & n5804 ) | ( ~n5589 & n5804 ) ;
  assign n5806 = ( n5794 & n5803 ) | ( n5794 & n5805 ) | ( n5803 & n5805 ) ;
  assign n5807 = ( n5589 & ~n5591 ) | ( n5589 & n5600 ) | ( ~n5591 & n5600 ) ;
  assign n5808 = ( n5591 & ~n5601 ) | ( n5591 & n5807 ) | ( ~n5601 & n5807 ) ;
  assign n5809 = n4202 & n4647 ;
  assign n5810 = n2174 & n4201 ;
  assign n5811 = n2298 | n4200 ;
  assign n5812 = n2270 & n4345 ;
  assign n5813 = ( ~n2298 & n5811 ) | ( ~n2298 & n5812 ) | ( n5811 & n5812 ) ;
  assign n5814 = ( ~n5809 & n5810 ) | ( ~n5809 & n5813 ) | ( n5810 & n5813 ) ;
  assign n5815 = ( ~x26 & n5809 ) | ( ~x26 & n5814 ) | ( n5809 & n5814 ) ;
  assign n5816 = ( n5809 & n5814 ) | ( n5809 & ~n5815 ) | ( n5814 & ~n5815 ) ;
  assign n5817 = ( x26 & n5815 ) | ( x26 & ~n5816 ) | ( n5815 & ~n5816 ) ;
  assign n5818 = ( n5806 & n5808 ) | ( n5806 & n5817 ) | ( n5808 & n5817 ) ;
  assign n5819 = ( n5601 & ~n5603 ) | ( n5601 & n5612 ) | ( ~n5603 & n5612 ) ;
  assign n5820 = ( n5603 & ~n5613 ) | ( n5603 & n5819 ) | ( ~n5613 & n5819 ) ;
  assign n5821 = n4290 & n4713 ;
  assign n5822 = n1852 & n4712 ;
  assign n5823 = ~n2023 & n4709 ;
  assign n5824 = n1926 & n4792 ;
  assign n5825 = n5823 | n5824 ;
  assign n5826 = ( ~n5821 & n5822 ) | ( ~n5821 & n5825 ) | ( n5822 & n5825 ) ;
  assign n5827 = ( ~x23 & n5821 ) | ( ~x23 & n5826 ) | ( n5821 & n5826 ) ;
  assign n5828 = ( n5821 & n5826 ) | ( n5821 & ~n5827 ) | ( n5826 & ~n5827 ) ;
  assign n5829 = ( x23 & n5827 ) | ( x23 & ~n5828 ) | ( n5827 & ~n5828 ) ;
  assign n5830 = ( n5818 & n5820 ) | ( n5818 & n5829 ) | ( n5820 & n5829 ) ;
  assign n5831 = ~n4302 & n4713 ;
  assign n5832 = ~n1750 & n4712 ;
  assign n5833 = n1852 & n4792 ;
  assign n5834 = n1926 & n4709 ;
  assign n5835 = n5833 | n5834 ;
  assign n5836 = ( ~n5831 & n5832 ) | ( ~n5831 & n5835 ) | ( n5832 & n5835 ) ;
  assign n5837 = ( ~x23 & n5831 ) | ( ~x23 & n5836 ) | ( n5831 & n5836 ) ;
  assign n5838 = ( n5831 & n5836 ) | ( n5831 & ~n5837 ) | ( n5836 & ~n5837 ) ;
  assign n5839 = ( x23 & n5837 ) | ( x23 & ~n5838 ) | ( n5837 & ~n5838 ) ;
  assign n5840 = ( ~n5613 & n5615 ) | ( ~n5613 & n5624 ) | ( n5615 & n5624 ) ;
  assign n5841 = ( n5613 & ~n5625 ) | ( n5613 & n5840 ) | ( ~n5625 & n5840 ) ;
  assign n5842 = ( n5830 & n5839 ) | ( n5830 & n5841 ) | ( n5839 & n5841 ) ;
  assign n5843 = ( ~n5625 & n5627 ) | ( ~n5625 & n5636 ) | ( n5627 & n5636 ) ;
  assign n5844 = ( n5625 & ~n5637 ) | ( n5625 & n5843 ) | ( ~n5637 & n5843 ) ;
  assign n5845 = ~n3955 & n4974 ;
  assign n5846 = ~n1338 & n5398 ;
  assign n5847 = n1458 & n4972 ;
  assign n5848 = n1576 & n4973 ;
  assign n5849 = n5847 | n5848 ;
  assign n5850 = ( ~n5845 & n5846 ) | ( ~n5845 & n5849 ) | ( n5846 & n5849 ) ;
  assign n5851 = ( ~x20 & n5845 ) | ( ~x20 & n5850 ) | ( n5845 & n5850 ) ;
  assign n5852 = ( n5845 & n5850 ) | ( n5845 & ~n5851 ) | ( n5850 & ~n5851 ) ;
  assign n5853 = ( x20 & n5851 ) | ( x20 & ~n5852 ) | ( n5851 & ~n5852 ) ;
  assign n5854 = ( n5842 & n5844 ) | ( n5842 & n5853 ) | ( n5844 & n5853 ) ;
  assign n5855 = ( ~n5637 & n5639 ) | ( ~n5637 & n5648 ) | ( n5639 & n5648 ) ;
  assign n5856 = ( n5637 & ~n5649 ) | ( n5637 & n5855 ) | ( ~n5649 & n5855 ) ;
  assign n5857 = ~n3665 & n5508 ;
  assign n5858 = ~n1290 & n5666 ;
  assign n5859 = ~n1246 & n5504 ;
  assign n5860 = ~n3658 & n5507 ;
  assign n5861 = n5859 | n5860 ;
  assign n5862 = ( ~n5857 & n5858 ) | ( ~n5857 & n5861 ) | ( n5858 & n5861 ) ;
  assign n5863 = ( ~x17 & n5857 ) | ( ~x17 & n5862 ) | ( n5857 & n5862 ) ;
  assign n5864 = ( n5857 & n5862 ) | ( n5857 & ~n5863 ) | ( n5862 & ~n5863 ) ;
  assign n5865 = ( x17 & n5863 ) | ( x17 & ~n5864 ) | ( n5863 & ~n5864 ) ;
  assign n5866 = ( n5854 & n5856 ) | ( n5854 & n5865 ) | ( n5856 & n5865 ) ;
  assign n5867 = n3692 & n5507 ;
  assign n5868 = ~n3658 & n5666 ;
  assign n5869 = ( n5507 & ~n5867 ) | ( n5507 & n5868 ) | ( ~n5867 & n5868 ) ;
  assign n5870 = ~n1290 & n5504 ;
  assign n5871 = n5869 | n5870 ;
  assign n5872 = ~n4182 & n5508 ;
  assign n5873 = ( x17 & n5871 ) | ( x17 & ~n5872 ) | ( n5871 & ~n5872 ) ;
  assign n5874 = ( ~x17 & n5871 ) | ( ~x17 & n5872 ) | ( n5871 & n5872 ) ;
  assign n5875 = ( ~n5871 & n5873 ) | ( ~n5871 & n5874 ) | ( n5873 & n5874 ) ;
  assign n5876 = ( ~n5649 & n5651 ) | ( ~n5649 & n5660 ) | ( n5651 & n5660 ) ;
  assign n5877 = ( ~n5660 & n5661 ) | ( ~n5660 & n5876 ) | ( n5661 & n5876 ) ;
  assign n5878 = ( n5866 & n5875 ) | ( n5866 & ~n5877 ) | ( n5875 & ~n5877 ) ;
  assign n5879 = n3800 & ~n5425 ;
  assign n5880 = n2552 & n3799 ;
  assign n5881 = ~n2725 & n3700 ;
  assign n5882 = n2635 & n3802 ;
  assign n5883 = n5881 | n5882 ;
  assign n5884 = ( ~n5879 & n5880 ) | ( ~n5879 & n5883 ) | ( n5880 & n5883 ) ;
  assign n5885 = ( ~x29 & n5879 ) | ( ~x29 & n5884 ) | ( n5879 & n5884 ) ;
  assign n5886 = ( n5879 & n5884 ) | ( n5879 & ~n5885 ) | ( n5884 & ~n5885 ) ;
  assign n5887 = ( x29 & n5885 ) | ( x29 & ~n5886 ) | ( n5885 & ~n5886 ) ;
  assign n5888 = ( ~n5783 & n5785 ) | ( ~n5783 & n5793 ) | ( n5785 & n5793 ) ;
  assign n5889 = ( n5783 & ~n5794 ) | ( n5783 & n5888 ) | ( ~n5794 & n5888 ) ;
  assign n5890 = n4202 & ~n4900 ;
  assign n5891 = n2396 & n4345 ;
  assign n5892 = ~n2298 & n4201 ;
  assign n5893 = ~n2491 & n4200 ;
  assign n5894 = n5892 | n5893 ;
  assign n5895 = ( ~n5890 & n5891 ) | ( ~n5890 & n5894 ) | ( n5891 & n5894 ) ;
  assign n5896 = ( ~x26 & n5890 ) | ( ~x26 & n5895 ) | ( n5890 & n5895 ) ;
  assign n5897 = ( n5890 & n5895 ) | ( n5890 & ~n5896 ) | ( n5895 & ~n5896 ) ;
  assign n5898 = ( x26 & n5896 ) | ( x26 & ~n5897 ) | ( n5896 & ~n5897 ) ;
  assign n5899 = ( n5887 & n5889 ) | ( n5887 & n5898 ) | ( n5889 & n5898 ) ;
  assign n5900 = ( ~n5794 & n5803 ) | ( ~n5794 & n5805 ) | ( n5803 & n5805 ) ;
  assign n5901 = ( n5794 & ~n5806 ) | ( n5794 & n5900 ) | ( ~n5806 & n5900 ) ;
  assign n5902 = n4202 & ~n4912 ;
  assign n5903 = n2396 & n4200 ;
  assign n5904 = n2270 & ~n4201 ;
  assign n5905 = ~n2298 & n4345 ;
  assign n5906 = ( n2270 & ~n5904 ) | ( n2270 & n5905 ) | ( ~n5904 & n5905 ) ;
  assign n5907 = ( ~n5902 & n5903 ) | ( ~n5902 & n5906 ) | ( n5903 & n5906 ) ;
  assign n5908 = ( ~x26 & n5902 ) | ( ~x26 & n5907 ) | ( n5902 & n5907 ) ;
  assign n5909 = ( n5902 & n5907 ) | ( n5902 & ~n5908 ) | ( n5907 & ~n5908 ) ;
  assign n5910 = ( x26 & n5908 ) | ( x26 & ~n5909 ) | ( n5908 & ~n5909 ) ;
  assign n5911 = ( n5899 & n5901 ) | ( n5899 & n5910 ) | ( n5901 & n5910 ) ;
  assign n5912 = ( n5806 & ~n5808 ) | ( n5806 & n5817 ) | ( ~n5808 & n5817 ) ;
  assign n5913 = ( n5808 & ~n5818 ) | ( n5808 & n5912 ) | ( ~n5818 & n5912 ) ;
  assign n5914 = ~n4457 & n4713 ;
  assign n5915 = n1926 & n4712 ;
  assign n5916 = ~n2023 & n4792 ;
  assign n5917 = n2089 & n4709 ;
  assign n5918 = n5916 | n5917 ;
  assign n5919 = ( ~n5914 & n5915 ) | ( ~n5914 & n5918 ) | ( n5915 & n5918 ) ;
  assign n5920 = ( ~x23 & n5914 ) | ( ~x23 & n5919 ) | ( n5914 & n5919 ) ;
  assign n5921 = ( n5914 & n5919 ) | ( n5914 & ~n5920 ) | ( n5919 & ~n5920 ) ;
  assign n5922 = ( x23 & n5920 ) | ( x23 & ~n5921 ) | ( n5920 & ~n5921 ) ;
  assign n5923 = ( n5911 & n5913 ) | ( n5911 & n5922 ) | ( n5913 & n5922 ) ;
  assign n5924 = ( n5818 & ~n5820 ) | ( n5818 & n5829 ) | ( ~n5820 & n5829 ) ;
  assign n5925 = ( n5820 & ~n5830 ) | ( n5820 & n5924 ) | ( ~n5830 & n5924 ) ;
  assign n5926 = n4326 & n4974 ;
  assign n5927 = n1576 & n5398 ;
  assign n5928 = n1750 | n4973 ;
  assign n5929 = ~n1669 & n4972 ;
  assign n5930 = ( ~n1750 & n5928 ) | ( ~n1750 & n5929 ) | ( n5928 & n5929 ) ;
  assign n5931 = ( ~n5926 & n5927 ) | ( ~n5926 & n5930 ) | ( n5927 & n5930 ) ;
  assign n5932 = ( ~x20 & n5926 ) | ( ~x20 & n5931 ) | ( n5926 & n5931 ) ;
  assign n5933 = ( n5926 & n5931 ) | ( n5926 & ~n5932 ) | ( n5931 & ~n5932 ) ;
  assign n5934 = ( x20 & n5932 ) | ( x20 & ~n5933 ) | ( n5932 & ~n5933 ) ;
  assign n5935 = ( n5923 & n5925 ) | ( n5923 & n5934 ) | ( n5925 & n5934 ) ;
  assign n5936 = ( ~n5830 & n5839 ) | ( ~n5830 & n5841 ) | ( n5839 & n5841 ) ;
  assign n5937 = ( n5830 & ~n5842 ) | ( n5830 & n5936 ) | ( ~n5842 & n5936 ) ;
  assign n5938 = ~n4159 & n4974 ;
  assign n5939 = n1458 & n5398 ;
  assign n5940 = n1669 | n4973 ;
  assign n5941 = n1576 & n4972 ;
  assign n5942 = ( ~n1669 & n5940 ) | ( ~n1669 & n5941 ) | ( n5940 & n5941 ) ;
  assign n5943 = ( ~n5938 & n5939 ) | ( ~n5938 & n5942 ) | ( n5939 & n5942 ) ;
  assign n5944 = ( ~x20 & n5938 ) | ( ~x20 & n5943 ) | ( n5938 & n5943 ) ;
  assign n5945 = ( n5938 & n5943 ) | ( n5938 & ~n5944 ) | ( n5943 & ~n5944 ) ;
  assign n5946 = ( x20 & n5944 ) | ( x20 & ~n5945 ) | ( n5944 & ~n5945 ) ;
  assign n5947 = ( n5935 & n5937 ) | ( n5935 & n5946 ) | ( n5937 & n5946 ) ;
  assign n5948 = ( ~n5842 & n5844 ) | ( ~n5842 & n5853 ) | ( n5844 & n5853 ) ;
  assign n5949 = ( n5842 & ~n5854 ) | ( n5842 & n5948 ) | ( ~n5854 & n5948 ) ;
  assign n5950 = n3621 & n5508 ;
  assign n5951 = ~n1290 & n5507 ;
  assign n5952 = ~n1246 & n5666 ;
  assign n5953 = n1267 & n5504 ;
  assign n5954 = n5952 | n5953 ;
  assign n5955 = ( ~n5950 & n5951 ) | ( ~n5950 & n5954 ) | ( n5951 & n5954 ) ;
  assign n5956 = ( ~x17 & n5950 ) | ( ~x17 & n5955 ) | ( n5950 & n5955 ) ;
  assign n5957 = ( n5950 & n5955 ) | ( n5950 & ~n5956 ) | ( n5955 & ~n5956 ) ;
  assign n5958 = ( x17 & n5956 ) | ( x17 & ~n5957 ) | ( n5956 & ~n5957 ) ;
  assign n5959 = ( n5947 & n5949 ) | ( n5947 & n5958 ) | ( n5949 & n5958 ) ;
  assign n5960 = x13 | x14 ;
  assign n5961 = x13 & x14 ;
  assign n5962 = n5960 & ~n5961 ;
  assign n5963 = x11 & x12 ;
  assign n5964 = x11 | x12 ;
  assign n5965 = ( n5962 & n5963 ) | ( n5962 & ~n5964 ) | ( n5963 & ~n5964 ) ;
  assign n5966 = n5962 & ~n5965 ;
  assign n5967 = x12 | x13 ;
  assign n5968 = x11 & ~x13 ;
  assign n5969 = ( ~n5964 & n5967 ) | ( ~n5964 & n5968 ) | ( n5967 & n5968 ) ;
  assign n5970 = n5965 & ~n5969 ;
  assign n5971 = ~n3692 & n5970 ;
  assign n5972 = ( n3691 & n3692 ) | ( n3691 & n5966 ) | ( n3692 & n5966 ) ;
  assign n5973 = ( n5966 & n5971 ) | ( n5966 & ~n5972 ) | ( n5971 & ~n5972 ) ;
  assign n5974 = x14 | n5973 ;
  assign n5975 = ( x14 & n5973 ) | ( x14 & ~n5974 ) | ( n5973 & ~n5974 ) ;
  assign n5976 = n5974 & ~n5975 ;
  assign n5977 = ( n5854 & ~n5856 ) | ( n5854 & n5865 ) | ( ~n5856 & n5865 ) ;
  assign n5978 = ( n5856 & ~n5866 ) | ( n5856 & n5977 ) | ( ~n5866 & n5977 ) ;
  assign n5979 = ( n5959 & n5976 ) | ( n5959 & n5978 ) | ( n5976 & n5978 ) ;
  assign n5980 = n113 | n2303 ;
  assign n5981 = ( n102 & n145 ) | ( n102 & n216 ) | ( n145 & n216 ) ;
  assign n5982 = ( n41 & n48 ) | ( n41 & n132 ) | ( n48 & n132 ) ;
  assign n5983 = n5981 | n5982 ;
  assign n5984 = ( n3522 & ~n5980 ) | ( n3522 & n5983 ) | ( ~n5980 & n5983 ) ;
  assign n5985 = n5980 | n5984 ;
  assign n5986 = n684 | n1838 ;
  assign n5987 = n484 | n1543 ;
  assign n5988 = n1798 | n2078 ;
  assign n5989 = ( n5986 & ~n5987 ) | ( n5986 & n5988 ) | ( ~n5987 & n5988 ) ;
  assign n5990 = ( n59 & n152 ) | ( n59 & n839 ) | ( n152 & n839 ) ;
  assign n5991 = n3852 | n5990 ;
  assign n5992 = ( n5987 & ~n5989 ) | ( n5987 & n5991 ) | ( ~n5989 & n5991 ) ;
  assign n5993 = n5989 | n5992 ;
  assign n5994 = n920 | n3835 ;
  assign n5995 = n2654 | n3003 ;
  assign n5996 = n595 | n3035 ;
  assign n5997 = ( ~n5994 & n5995 ) | ( ~n5994 & n5996 ) | ( n5995 & n5996 ) ;
  assign n5998 = n5994 | n5997 ;
  assign n5999 = ( ~n5985 & n5993 ) | ( ~n5985 & n5998 ) | ( n5993 & n5998 ) ;
  assign n6000 = n5985 | n5999 ;
  assign n6001 = n2978 & ~n3943 ;
  assign n6002 = ( ~n4439 & n6000 ) | ( ~n4439 & n6001 ) | ( n6000 & n6001 ) ;
  assign n6003 = ~n6000 & n6002 ;
  assign n6004 = n1250 & ~n3533 ;
  assign n6005 = n607 & ~n3586 ;
  assign n6006 = n6004 | n6005 ;
  assign n6007 = n606 & ~n3479 ;
  assign n6008 = ( n606 & n6006 ) | ( n606 & ~n6007 ) | ( n6006 & ~n6007 ) ;
  assign n6009 = ~n3533 & n3586 ;
  assign n6010 = ( ~n1248 & n3479 ) | ( ~n1248 & n6009 ) | ( n3479 & n6009 ) ;
  assign n6011 = ( n3587 & n6008 ) | ( n3587 & ~n6010 ) | ( n6008 & ~n6010 ) ;
  assign n6012 = ~n6003 & n6011 ;
  assign n6013 = n1487 | n3460 ;
  assign n6014 = ( n57 & n75 ) | ( n57 & n122 ) | ( n75 & n122 ) ;
  assign n6015 = ( n146 & n211 ) | ( n146 & ~n6014 ) | ( n211 & ~n6014 ) ;
  assign n6016 = n6014 | n6015 ;
  assign n6017 = ( n1093 & ~n6013 ) | ( n1093 & n6016 ) | ( ~n6013 & n6016 ) ;
  assign n6018 = ( ~n2281 & n6013 ) | ( ~n2281 & n6017 ) | ( n6013 & n6017 ) ;
  assign n6019 = n2281 | n6018 ;
  assign n6020 = n489 | n523 ;
  assign n6021 = ( n113 & ~n489 ) | ( n113 & n3003 ) | ( ~n489 & n3003 ) ;
  assign n6022 = ( n185 & ~n6020 ) | ( n185 & n6021 ) | ( ~n6020 & n6021 ) ;
  assign n6023 = n6020 | n6022 ;
  assign n6024 = n2556 | n6023 ;
  assign n6025 = n838 | n1145 ;
  assign n6026 = n356 | n6025 ;
  assign n6027 = ( ~n6019 & n6024 ) | ( ~n6019 & n6026 ) | ( n6024 & n6026 ) ;
  assign n6028 = n6019 | n6027 ;
  assign n6029 = n2424 | n3477 ;
  assign n6030 = n287 | n1174 ;
  assign n6031 = n218 & ~n947 ;
  assign n6032 = n534 | n895 ;
  assign n6033 = ( n2571 & n6031 ) | ( n2571 & n6032 ) | ( n6031 & n6032 ) ;
  assign n6034 = n6031 & ~n6033 ;
  assign n6035 = ( ~n175 & n6030 ) | ( ~n175 & n6034 ) | ( n6030 & n6034 ) ;
  assign n6036 = ~n6030 & n6035 ;
  assign n6037 = n144 | n1870 ;
  assign n6038 = n1526 | n6037 ;
  assign n6039 = ( n782 & n837 ) | ( n782 & ~n6038 ) | ( n837 & ~n6038 ) ;
  assign n6040 = n6038 | n6039 ;
  assign n6041 = n566 | n2969 ;
  assign n6042 = n2029 | n3284 ;
  assign n6043 = n1079 | n2528 ;
  assign n6044 = ( n6041 & ~n6042 ) | ( n6041 & n6043 ) | ( ~n6042 & n6043 ) ;
  assign n6045 = ( n73 & n166 ) | ( n73 & n216 ) | ( n166 & n216 ) ;
  assign n6046 = ( n851 & n1001 ) | ( n851 & ~n6045 ) | ( n1001 & ~n6045 ) ;
  assign n6047 = n6045 | n6046 ;
  assign n6048 = ( n305 & ~n6040 ) | ( n305 & n6047 ) | ( ~n6040 & n6047 ) ;
  assign n6049 = ( n6042 & ~n6044 ) | ( n6042 & n6048 ) | ( ~n6044 & n6048 ) ;
  assign n6050 = n6044 | n6049 ;
  assign n6051 = ( n6036 & n6040 ) | ( n6036 & n6050 ) | ( n6040 & n6050 ) ;
  assign n6052 = n6036 & ~n6051 ;
  assign n6053 = ( n6028 & ~n6029 ) | ( n6028 & n6052 ) | ( ~n6029 & n6052 ) ;
  assign n6054 = ~n6028 & n6053 ;
  assign n6055 = n606 | n3389 ;
  assign n6056 = n607 & ~n3533 ;
  assign n6057 = ( ~n3389 & n6055 ) | ( ~n3389 & n6056 ) | ( n6055 & n6056 ) ;
  assign n6058 = ~n1250 & n3479 ;
  assign n6059 = ( n3479 & n6057 ) | ( n3479 & ~n6058 ) | ( n6057 & ~n6058 ) ;
  assign n6060 = ( ~n3479 & n3533 ) | ( ~n3479 & n3587 ) | ( n3533 & n3587 ) ;
  assign n6061 = ( n3588 & n3589 ) | ( n3588 & ~n6060 ) | ( n3589 & ~n6060 ) ;
  assign n6062 = n1248 & n6061 ;
  assign n6063 = n6059 | n6062 ;
  assign n6064 = ( n6012 & ~n6054 ) | ( n6012 & n6063 ) | ( ~n6054 & n6063 ) ;
  assign n6065 = n110 | n290 ;
  assign n6066 = n1477 | n6065 ;
  assign n6067 = n75 | n145 ;
  assign n6068 = ( n116 & n166 ) | ( n116 & n6067 ) | ( n166 & n6067 ) ;
  assign n6069 = n748 | n6068 ;
  assign n6070 = ( n1351 & n1715 ) | ( n1351 & ~n6069 ) | ( n1715 & ~n6069 ) ;
  assign n6071 = n6069 | n6070 ;
  assign n6072 = ( n4272 & ~n6066 ) | ( n4272 & n6071 ) | ( ~n6066 & n6071 ) ;
  assign n6073 = n6066 | n6072 ;
  assign n6074 = n996 | n4463 ;
  assign n6075 = n712 | n1113 ;
  assign n6076 = n679 | n782 ;
  assign n6077 = ( n416 & n551 ) | ( n416 & ~n6076 ) | ( n551 & ~n6076 ) ;
  assign n6078 = n6076 | n6077 ;
  assign n6079 = ( ~n6074 & n6075 ) | ( ~n6074 & n6078 ) | ( n6075 & n6078 ) ;
  assign n6080 = n6074 | n6079 ;
  assign n6081 = ( ~n3125 & n6073 ) | ( ~n3125 & n6080 ) | ( n6073 & n6080 ) ;
  assign n6082 = n170 | n567 ;
  assign n6083 = ( n173 & n544 ) | ( n173 & ~n6082 ) | ( n544 & ~n6082 ) ;
  assign n6084 = n6082 | n6083 ;
  assign n6085 = n2598 | n3941 ;
  assign n6086 = n217 | n441 ;
  assign n6087 = n148 | n6086 ;
  assign n6088 = ( ~n6084 & n6085 ) | ( ~n6084 & n6087 ) | ( n6085 & n6087 ) ;
  assign n6089 = n6084 | n6088 ;
  assign n6090 = ( ~n196 & n291 ) | ( ~n196 & n1001 ) | ( n291 & n1001 ) ;
  assign n6091 = n196 | n6090 ;
  assign n6092 = n448 | n795 ;
  assign n6093 = ( n1122 & ~n6091 ) | ( n1122 & n6092 ) | ( ~n6091 & n6092 ) ;
  assign n6094 = n6091 | n6093 ;
  assign n6095 = ( ~n6080 & n6089 ) | ( ~n6080 & n6094 ) | ( n6089 & n6094 ) ;
  assign n6096 = ( ~n3125 & n6081 ) | ( ~n3125 & n6095 ) | ( n6081 & n6095 ) ;
  assign n6097 = n3125 | n6096 ;
  assign n6098 = n606 & ~n3355 ;
  assign n6099 = n1250 & ~n3389 ;
  assign n6100 = n6098 | n6099 ;
  assign n6101 = n607 & ~n3479 ;
  assign n6102 = ( n607 & n6100 ) | ( n607 & ~n6101 ) | ( n6100 & ~n6101 ) ;
  assign n6103 = ( n3355 & ~n3389 ) | ( n3355 & n3589 ) | ( ~n3389 & n3589 ) ;
  assign n6104 = ( n3389 & ~n3590 ) | ( n3389 & n6103 ) | ( ~n3590 & n6103 ) ;
  assign n6105 = n1248 & ~n6104 ;
  assign n6106 = n6102 | n6105 ;
  assign n6107 = ( n6064 & n6097 ) | ( n6064 & n6106 ) | ( n6097 & n6106 ) ;
  assign n6108 = ( n455 & n587 ) | ( n455 & ~n3026 ) | ( n587 & ~n3026 ) ;
  assign n6109 = n3026 | n6108 ;
  assign n6110 = n144 | n203 ;
  assign n6111 = ( n2585 & n3245 ) | ( n2585 & ~n6110 ) | ( n3245 & ~n6110 ) ;
  assign n6112 = n6110 | n6111 ;
  assign n6113 = n172 | n1068 ;
  assign n6114 = n288 | n775 ;
  assign n6115 = ( n783 & n1059 ) | ( n783 & ~n6114 ) | ( n1059 & ~n6114 ) ;
  assign n6116 = n6114 | n6115 ;
  assign n6117 = n2577 | n2811 ;
  assign n6118 = n1589 | n2414 ;
  assign n6119 = ( n5249 & ~n6117 ) | ( n5249 & n6118 ) | ( ~n6117 & n6118 ) ;
  assign n6120 = n6117 | n6119 ;
  assign n6121 = ( ~n6113 & n6116 ) | ( ~n6113 & n6120 ) | ( n6116 & n6120 ) ;
  assign n6122 = ( ~n6112 & n6113 ) | ( ~n6112 & n6121 ) | ( n6113 & n6121 ) ;
  assign n6123 = ( ~n6109 & n6112 ) | ( ~n6109 & n6122 ) | ( n6112 & n6122 ) ;
  assign n6124 = n6109 | n6123 ;
  assign n6125 = n689 | n762 ;
  assign n6126 = ( n124 & n173 ) | ( n124 & ~n6125 ) | ( n173 & ~n6125 ) ;
  assign n6127 = n6125 | n6126 ;
  assign n6128 = n273 | n1048 ;
  assign n6129 = ( n2496 & n4983 ) | ( n2496 & ~n6128 ) | ( n4983 & ~n6128 ) ;
  assign n6130 = n6128 | n6129 ;
  assign n6131 = ( n81 & n911 ) | ( n81 & ~n3063 ) | ( n911 & ~n3063 ) ;
  assign n6132 = n3063 | n6131 ;
  assign n6133 = ( ~n6127 & n6130 ) | ( ~n6127 & n6132 ) | ( n6130 & n6132 ) ;
  assign n6134 = n6127 | n6133 ;
  assign n6135 = n478 | n3189 ;
  assign n6136 = n697 | n2047 ;
  assign n6137 = n164 | n225 ;
  assign n6138 = ( n963 & n1129 ) | ( n963 & ~n6137 ) | ( n1129 & ~n6137 ) ;
  assign n6139 = n6137 | n6138 ;
  assign n6140 = ( ~n836 & n856 ) | ( ~n836 & n1169 ) | ( n856 & n1169 ) ;
  assign n6141 = n836 | n6140 ;
  assign n6142 = ( ~n6136 & n6139 ) | ( ~n6136 & n6141 ) | ( n6139 & n6141 ) ;
  assign n6143 = n6136 | n6142 ;
  assign n6144 = ( ~n6134 & n6135 ) | ( ~n6134 & n6143 ) | ( n6135 & n6143 ) ;
  assign n6145 = n6134 | n6144 ;
  assign n6146 = ( n5131 & n6124 ) | ( n5131 & ~n6145 ) | ( n6124 & ~n6145 ) ;
  assign n6147 = ~n6124 & n6146 ;
  assign n6148 = n1250 & ~n3355 ;
  assign n6149 = n607 & ~n3389 ;
  assign n6150 = n6148 | n6149 ;
  assign n6151 = n606 & n3300 ;
  assign n6152 = ( n606 & n6150 ) | ( n606 & ~n6151 ) | ( n6150 & ~n6151 ) ;
  assign n6153 = ( n3300 & n3355 ) | ( n3300 & ~n3590 ) | ( n3355 & ~n3590 ) ;
  assign n6154 = ( n3590 & ~n3591 ) | ( n3590 & n6153 ) | ( ~n3591 & n6153 ) ;
  assign n6155 = n1248 & ~n6154 ;
  assign n6156 = n6152 | n6155 ;
  assign n6157 = ( n6107 & ~n6147 ) | ( n6107 & n6156 ) | ( ~n6147 & n6156 ) ;
  assign n6158 = n1083 | n1128 ;
  assign n6159 = n957 | n6158 ;
  assign n6160 = n2071 | n2671 ;
  assign n6161 = ( n2636 & n2683 ) | ( n2636 & ~n6160 ) | ( n2683 & ~n6160 ) ;
  assign n6162 = n6160 | n6161 ;
  assign n6163 = n1220 | n1793 ;
  assign n6164 = n331 | n2225 ;
  assign n6165 = n6163 | n6164 ;
  assign n6166 = ( ~n6158 & n6162 ) | ( ~n6158 & n6165 ) | ( n6162 & n6165 ) ;
  assign n6167 = ( ~n1707 & n6159 ) | ( ~n1707 & n6166 ) | ( n6159 & n6166 ) ;
  assign n6168 = n1707 | n6167 ;
  assign n6169 = n590 | n810 ;
  assign n6170 = n1254 | n1488 ;
  assign n6171 = ( n1790 & ~n6169 ) | ( n1790 & n6170 ) | ( ~n6169 & n6170 ) ;
  assign n6172 = n6169 | n6171 ;
  assign n6173 = n134 | n5072 ;
  assign n6174 = ( n228 & n734 ) | ( n228 & ~n981 ) | ( n734 & ~n981 ) ;
  assign n6175 = n981 | n6174 ;
  assign n6176 = ( ~n6172 & n6173 ) | ( ~n6172 & n6175 ) | ( n6173 & n6175 ) ;
  assign n6177 = n6172 | n6176 ;
  assign n6178 = ( n174 & ~n653 ) | ( n174 & n886 ) | ( ~n653 & n886 ) ;
  assign n6179 = n653 | n6178 ;
  assign n6180 = n59 | n72 ;
  assign n6181 = ( n64 & n109 ) | ( n64 & n6180 ) | ( n109 & n6180 ) ;
  assign n6182 = n482 | n2787 ;
  assign n6183 = n1110 | n6182 ;
  assign n6184 = ( ~n6179 & n6181 ) | ( ~n6179 & n6183 ) | ( n6181 & n6183 ) ;
  assign n6185 = ( n4984 & ~n6179 ) | ( n4984 & n6184 ) | ( ~n6179 & n6184 ) ;
  assign n6186 = n836 | n5247 ;
  assign n6187 = n1235 | n1543 ;
  assign n6188 = ( n4428 & ~n6186 ) | ( n4428 & n6187 ) | ( ~n6186 & n6187 ) ;
  assign n6189 = n6186 | n6188 ;
  assign n6190 = ( n6179 & ~n6185 ) | ( n6179 & n6189 ) | ( ~n6185 & n6189 ) ;
  assign n6191 = n6185 | n6190 ;
  assign n6192 = ( ~n6168 & n6177 ) | ( ~n6168 & n6191 ) | ( n6177 & n6191 ) ;
  assign n6193 = n6168 | n6192 ;
  assign n6194 = n607 & ~n3355 ;
  assign n6195 = n606 & n3239 ;
  assign n6196 = n6194 | n6195 ;
  assign n6197 = n1250 | n3300 ;
  assign n6198 = ( ~n3300 & n6196 ) | ( ~n3300 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6199 = ( n3239 & ~n3300 ) | ( n3239 & n3591 ) | ( ~n3300 & n3591 ) ;
  assign n6200 = ( ~n3591 & n3592 ) | ( ~n3591 & n6199 ) | ( n3592 & n6199 ) ;
  assign n6201 = n1248 & n6200 ;
  assign n6202 = n6198 | n6201 ;
  assign n6203 = ( n6157 & n6193 ) | ( n6157 & n6202 ) | ( n6193 & n6202 ) ;
  assign n6204 = n447 | n1001 ;
  assign n6205 = ( n529 & n549 ) | ( n529 & ~n6204 ) | ( n549 & ~n6204 ) ;
  assign n6206 = n6204 | n6205 ;
  assign n6207 = n1544 | n1893 ;
  assign n6208 = n762 | n1595 ;
  assign n6209 = n2011 | n2636 ;
  assign n6210 = ( n2819 & n3369 ) | ( n2819 & ~n6209 ) | ( n3369 & ~n6209 ) ;
  assign n6211 = n6209 | n6210 ;
  assign n6212 = ( ~n6207 & n6208 ) | ( ~n6207 & n6211 ) | ( n6208 & n6211 ) ;
  assign n6213 = n6207 | n6212 ;
  assign n6214 = ( n69 & n831 ) | ( n69 & ~n6213 ) | ( n831 & ~n6213 ) ;
  assign n6215 = n6213 | n6214 ;
  assign n6216 = n74 | n1632 ;
  assign n6217 = n5155 | n6216 ;
  assign n6218 = ( ~n6206 & n6215 ) | ( ~n6206 & n6217 ) | ( n6215 & n6217 ) ;
  assign n6219 = n6206 | n6218 ;
  assign n6220 = n4558 | n4566 ;
  assign n6221 = n2077 | n2181 ;
  assign n6222 = n133 | n1163 ;
  assign n6223 = n227 | n261 ;
  assign n6224 = ( ~n54 & n66 ) | ( ~n54 & n73 ) | ( n66 & n73 ) ;
  assign n6225 = n369 | n6224 ;
  assign n6226 = ( n483 & ~n6223 ) | ( n483 & n6225 ) | ( ~n6223 & n6225 ) ;
  assign n6227 = n6223 | n6226 ;
  assign n6228 = ( ~n6221 & n6222 ) | ( ~n6221 & n6227 ) | ( n6222 & n6227 ) ;
  assign n6229 = n6221 | n6228 ;
  assign n6230 = ( n2796 & ~n4468 ) | ( n2796 & n6229 ) | ( ~n4468 & n6229 ) ;
  assign n6231 = n3406 | n4601 ;
  assign n6232 = n4872 | n6231 ;
  assign n6233 = ( n4468 & ~n6230 ) | ( n4468 & n6232 ) | ( ~n6230 & n6232 ) ;
  assign n6234 = n6230 | n6233 ;
  assign n6235 = ( ~n6219 & n6220 ) | ( ~n6219 & n6234 ) | ( n6220 & n6234 ) ;
  assign n6236 = n6219 | n6235 ;
  assign n6237 = ~n1250 & n3239 ;
  assign n6238 = n606 & n3153 ;
  assign n6239 = ( n3239 & ~n6237 ) | ( n3239 & n6238 ) | ( ~n6237 & n6238 ) ;
  assign n6240 = n607 & n3300 ;
  assign n6241 = ( n607 & n6239 ) | ( n607 & ~n6240 ) | ( n6239 & ~n6240 ) ;
  assign n6242 = ( n3153 & n3239 ) | ( n3153 & ~n3593 ) | ( n3239 & ~n3593 ) ;
  assign n6243 = ( n3592 & n3593 ) | ( n3592 & ~n6242 ) | ( n3593 & ~n6242 ) ;
  assign n6244 = n1248 & ~n6243 ;
  assign n6245 = n6241 | n6244 ;
  assign n6246 = ( n6203 & n6236 ) | ( n6203 & n6245 ) | ( n6236 & n6245 ) ;
  assign n6247 = ( x2 & ~n5703 ) | ( x2 & n5712 ) | ( ~n5703 & n5712 ) ;
  assign n6248 = ( n5703 & ~n5713 ) | ( n5703 & n6247 ) | ( ~n5713 & n6247 ) ;
  assign n6249 = n3800 & ~n5768 ;
  assign n6250 = ~n2910 & n3799 ;
  assign n6251 = n3046 | n3700 ;
  assign n6252 = ~n2965 & n3802 ;
  assign n6253 = ( ~n3046 & n6251 ) | ( ~n3046 & n6252 ) | ( n6251 & n6252 ) ;
  assign n6254 = ( ~n6249 & n6250 ) | ( ~n6249 & n6253 ) | ( n6250 & n6253 ) ;
  assign n6255 = ( ~x29 & n6249 ) | ( ~x29 & n6254 ) | ( n6249 & n6254 ) ;
  assign n6256 = ( n6249 & n6254 ) | ( n6249 & ~n6255 ) | ( n6254 & ~n6255 ) ;
  assign n6257 = ( x29 & n6255 ) | ( x29 & ~n6256 ) | ( n6255 & ~n6256 ) ;
  assign n6258 = ( n6246 & n6248 ) | ( n6246 & n6257 ) | ( n6248 & n6257 ) ;
  assign n6259 = ( ~x2 & n5713 ) | ( ~x2 & n5732 ) | ( n5713 & n5732 ) ;
  assign n6260 = ( x2 & ~n5733 ) | ( x2 & n6259 ) | ( ~n5733 & n6259 ) ;
  assign n6261 = n1250 & n3078 ;
  assign n6262 = n606 & ~n3046 ;
  assign n6263 = n6261 | n6262 ;
  assign n6264 = n607 & ~n3153 ;
  assign n6265 = ( n607 & n6263 ) | ( n607 & ~n6264 ) | ( n6263 & ~n6264 ) ;
  assign n6266 = ( n3046 & ~n3078 ) | ( n3046 & n3594 ) | ( ~n3078 & n3594 ) ;
  assign n6267 = ( ~n3594 & n3595 ) | ( ~n3594 & n6266 ) | ( n3595 & n6266 ) ;
  assign n6268 = n1248 & ~n6267 ;
  assign n6269 = n6265 | n6268 ;
  assign n6270 = ( n6258 & n6260 ) | ( n6258 & n6269 ) | ( n6260 & n6269 ) ;
  assign n6271 = ( x2 & n5733 ) | ( x2 & n5758 ) | ( n5733 & n5758 ) ;
  assign n6272 = ( n5758 & n5759 ) | ( n5758 & ~n6271 ) | ( n5759 & ~n6271 ) ;
  assign n6273 = ~n607 & n3078 ;
  assign n6274 = n1250 & ~n3046 ;
  assign n6275 = ( n3078 & ~n6273 ) | ( n3078 & n6274 ) | ( ~n6273 & n6274 ) ;
  assign n6276 = n606 & n2965 ;
  assign n6277 = ( n606 & n6275 ) | ( n606 & ~n6276 ) | ( n6275 & ~n6276 ) ;
  assign n6278 = ( n2965 & n3046 ) | ( n2965 & ~n3596 ) | ( n3046 & ~n3596 ) ;
  assign n6279 = ( n3595 & n3596 ) | ( n3595 & ~n6278 ) | ( n3596 & ~n6278 ) ;
  assign n6280 = n1248 & n6279 ;
  assign n6281 = n6277 | n6280 ;
  assign n6282 = ( n6270 & ~n6272 ) | ( n6270 & n6281 ) | ( ~n6272 & n6281 ) ;
  assign n6283 = ( n5759 & ~n5761 ) | ( n5759 & n5770 ) | ( ~n5761 & n5770 ) ;
  assign n6284 = ( n5761 & ~n5771 ) | ( n5761 & n6283 ) | ( ~n5771 & n6283 ) ;
  assign n6285 = n3800 & ~n5586 ;
  assign n6286 = ~n2725 & n3799 ;
  assign n6287 = n2843 & n3700 ;
  assign n6288 = ~n2810 & n3802 ;
  assign n6289 = n6287 | n6288 ;
  assign n6290 = ( ~n6285 & n6286 ) | ( ~n6285 & n6289 ) | ( n6286 & n6289 ) ;
  assign n6291 = ( ~x29 & n6285 ) | ( ~x29 & n6290 ) | ( n6285 & n6290 ) ;
  assign n6292 = ( n6285 & n6290 ) | ( n6285 & ~n6291 ) | ( n6290 & ~n6291 ) ;
  assign n6293 = ( x29 & n6291 ) | ( x29 & ~n6292 ) | ( n6291 & ~n6292 ) ;
  assign n6294 = ( n6282 & n6284 ) | ( n6282 & n6293 ) | ( n6284 & n6293 ) ;
  assign n6295 = ( ~n5771 & n5773 ) | ( ~n5771 & n5782 ) | ( n5773 & n5782 ) ;
  assign n6296 = ( ~n5782 & n5783 ) | ( ~n5782 & n6295 ) | ( n5783 & n6295 ) ;
  assign n6297 = n4202 & ~n5084 ;
  assign n6298 = n2396 & n4201 ;
  assign n6299 = ~n2491 & n4345 ;
  assign n6300 = n2552 & n4200 ;
  assign n6301 = n6299 | n6300 ;
  assign n6302 = ( ~n6297 & n6298 ) | ( ~n6297 & n6301 ) | ( n6298 & n6301 ) ;
  assign n6303 = ( ~x26 & n6297 ) | ( ~x26 & n6302 ) | ( n6297 & n6302 ) ;
  assign n6304 = ( n6297 & n6302 ) | ( n6297 & ~n6303 ) | ( n6302 & ~n6303 ) ;
  assign n6305 = ( x26 & n6303 ) | ( x26 & ~n6304 ) | ( n6303 & ~n6304 ) ;
  assign n6306 = ( n6294 & ~n6296 ) | ( n6294 & n6305 ) | ( ~n6296 & n6305 ) ;
  assign n6307 = ( n5887 & ~n5889 ) | ( n5887 & n5898 ) | ( ~n5889 & n5898 ) ;
  assign n6308 = ( n5889 & ~n5899 ) | ( n5889 & n6307 ) | ( ~n5899 & n6307 ) ;
  assign n6309 = n4713 & n4730 ;
  assign n6310 = n2089 & n4712 ;
  assign n6311 = n2270 & n4709 ;
  assign n6312 = n2174 & n4792 ;
  assign n6313 = n6311 | n6312 ;
  assign n6314 = ( ~n6309 & n6310 ) | ( ~n6309 & n6313 ) | ( n6310 & n6313 ) ;
  assign n6315 = ( ~x23 & n6309 ) | ( ~x23 & n6314 ) | ( n6309 & n6314 ) ;
  assign n6316 = ( n6309 & n6314 ) | ( n6309 & ~n6315 ) | ( n6314 & ~n6315 ) ;
  assign n6317 = ( x23 & n6315 ) | ( x23 & ~n6316 ) | ( n6315 & ~n6316 ) ;
  assign n6318 = ( n6306 & n6308 ) | ( n6306 & n6317 ) | ( n6308 & n6317 ) ;
  assign n6319 = ~n4660 & n4713 ;
  assign n6320 = ~n2023 & n4712 ;
  assign n6321 = n2174 & n4709 ;
  assign n6322 = n2089 & n4792 ;
  assign n6323 = n6321 | n6322 ;
  assign n6324 = ( ~n6319 & n6320 ) | ( ~n6319 & n6323 ) | ( n6320 & n6323 ) ;
  assign n6325 = ( ~x23 & n6319 ) | ( ~x23 & n6324 ) | ( n6319 & n6324 ) ;
  assign n6326 = ( n6319 & n6324 ) | ( n6319 & ~n6325 ) | ( n6324 & ~n6325 ) ;
  assign n6327 = ( x23 & n6325 ) | ( x23 & ~n6326 ) | ( n6325 & ~n6326 ) ;
  assign n6328 = ( ~n5899 & n5901 ) | ( ~n5899 & n5910 ) | ( n5901 & n5910 ) ;
  assign n6329 = ( n5899 & ~n5911 ) | ( n5899 & n6328 ) | ( ~n5911 & n6328 ) ;
  assign n6330 = ( n6318 & n6327 ) | ( n6318 & n6329 ) | ( n6327 & n6329 ) ;
  assign n6331 = ( n5911 & ~n5913 ) | ( n5911 & n5922 ) | ( ~n5913 & n5922 ) ;
  assign n6332 = ( n5913 & ~n5923 ) | ( n5913 & n6331 ) | ( ~n5923 & n6331 ) ;
  assign n6333 = n4146 & n4974 ;
  assign n6334 = ~n1669 & n5398 ;
  assign n6335 = n1852 & ~n4973 ;
  assign n6336 = ~n1750 & n4972 ;
  assign n6337 = ( n1852 & ~n6335 ) | ( n1852 & n6336 ) | ( ~n6335 & n6336 ) ;
  assign n6338 = ( ~n6333 & n6334 ) | ( ~n6333 & n6337 ) | ( n6334 & n6337 ) ;
  assign n6339 = ( ~x20 & n6333 ) | ( ~x20 & n6338 ) | ( n6333 & n6338 ) ;
  assign n6340 = ( n6333 & n6338 ) | ( n6333 & ~n6339 ) | ( n6338 & ~n6339 ) ;
  assign n6341 = ( x20 & n6339 ) | ( x20 & ~n6340 ) | ( n6339 & ~n6340 ) ;
  assign n6342 = ( n6330 & n6332 ) | ( n6330 & n6341 ) | ( n6332 & n6341 ) ;
  assign n6343 = ( n5923 & ~n5925 ) | ( n5923 & n5934 ) | ( ~n5925 & n5934 ) ;
  assign n6344 = ( n5925 & ~n5935 ) | ( n5925 & n6343 ) | ( ~n5935 & n6343 ) ;
  assign n6345 = ~n3779 & n5508 ;
  assign n6346 = n1267 & n5507 ;
  assign n6347 = n1458 & ~n5504 ;
  assign n6348 = ~n1338 & n5666 ;
  assign n6349 = ( n1458 & ~n6347 ) | ( n1458 & n6348 ) | ( ~n6347 & n6348 ) ;
  assign n6350 = ( ~n6345 & n6346 ) | ( ~n6345 & n6349 ) | ( n6346 & n6349 ) ;
  assign n6351 = ( ~x17 & n6345 ) | ( ~x17 & n6350 ) | ( n6345 & n6350 ) ;
  assign n6352 = ( n6345 & n6350 ) | ( n6345 & ~n6351 ) | ( n6350 & ~n6351 ) ;
  assign n6353 = ( x17 & n6351 ) | ( x17 & ~n6352 ) | ( n6351 & ~n6352 ) ;
  assign n6354 = ( n6342 & n6344 ) | ( n6342 & n6353 ) | ( n6344 & n6353 ) ;
  assign n6355 = ~n3791 & n5508 ;
  assign n6356 = n1267 & n5666 ;
  assign n6357 = ~n1246 & n5507 ;
  assign n6358 = ~n1338 & n5504 ;
  assign n6359 = n6357 | n6358 ;
  assign n6360 = ( ~n6355 & n6356 ) | ( ~n6355 & n6359 ) | ( n6356 & n6359 ) ;
  assign n6361 = ( ~x17 & n6355 ) | ( ~x17 & n6360 ) | ( n6355 & n6360 ) ;
  assign n6362 = ( n6355 & n6360 ) | ( n6355 & ~n6361 ) | ( n6360 & ~n6361 ) ;
  assign n6363 = ( x17 & n6361 ) | ( x17 & ~n6362 ) | ( n6361 & ~n6362 ) ;
  assign n6364 = ( ~n5935 & n5937 ) | ( ~n5935 & n5946 ) | ( n5937 & n5946 ) ;
  assign n6365 = ( n5935 & ~n5947 ) | ( n5935 & n6364 ) | ( ~n5947 & n6364 ) ;
  assign n6366 = ( n6354 & n6363 ) | ( n6354 & n6365 ) | ( n6363 & n6365 ) ;
  assign n6367 = n3797 & n5966 ;
  assign n6368 = ~n3692 & n5969 ;
  assign n6369 = ~n3658 & n5970 ;
  assign n6370 = n6368 | n6369 ;
  assign n6371 = ( ~x14 & n6367 ) | ( ~x14 & n6370 ) | ( n6367 & n6370 ) ;
  assign n6372 = ( n6367 & n6370 ) | ( n6367 & ~n6371 ) | ( n6370 & ~n6371 ) ;
  assign n6373 = ( x14 & n6371 ) | ( x14 & ~n6372 ) | ( n6371 & ~n6372 ) ;
  assign n6374 = ( n5947 & ~n5949 ) | ( n5947 & n5958 ) | ( ~n5949 & n5958 ) ;
  assign n6375 = ( n5949 & ~n5959 ) | ( n5949 & n6374 ) | ( ~n5959 & n6374 ) ;
  assign n6376 = ( n6366 & n6373 ) | ( n6366 & n6375 ) | ( n6373 & n6375 ) ;
  assign n6377 = n3800 & n5791 ;
  assign n6378 = ~n2810 & n3799 ;
  assign n6379 = n2910 | n3700 ;
  assign n6380 = n2843 & n3802 ;
  assign n6381 = ( ~n2910 & n6379 ) | ( ~n2910 & n6380 ) | ( n6379 & n6380 ) ;
  assign n6382 = ( ~n6377 & n6378 ) | ( ~n6377 & n6381 ) | ( n6378 & n6381 ) ;
  assign n6383 = ( ~x29 & n6377 ) | ( ~x29 & n6382 ) | ( n6377 & n6382 ) ;
  assign n6384 = ( n6377 & n6382 ) | ( n6377 & ~n6383 ) | ( n6382 & ~n6383 ) ;
  assign n6385 = ( x29 & n6383 ) | ( x29 & ~n6384 ) | ( n6383 & ~n6384 ) ;
  assign n6386 = ( ~n6270 & n6272 ) | ( ~n6270 & n6281 ) | ( n6272 & n6281 ) ;
  assign n6387 = ( ~n6281 & n6282 ) | ( ~n6281 & n6386 ) | ( n6282 & n6386 ) ;
  assign n6388 = n4202 & ~n5425 ;
  assign n6389 = n2552 & n4201 ;
  assign n6390 = ~n2725 & n4200 ;
  assign n6391 = n2635 & n4345 ;
  assign n6392 = n6390 | n6391 ;
  assign n6393 = ( ~n6388 & n6389 ) | ( ~n6388 & n6392 ) | ( n6389 & n6392 ) ;
  assign n6394 = ( ~x26 & n6388 ) | ( ~x26 & n6393 ) | ( n6388 & n6393 ) ;
  assign n6395 = ( n6388 & n6393 ) | ( n6388 & ~n6394 ) | ( n6393 & ~n6394 ) ;
  assign n6396 = ( x26 & n6394 ) | ( x26 & ~n6395 ) | ( n6394 & ~n6395 ) ;
  assign n6397 = ( n6385 & ~n6387 ) | ( n6385 & n6396 ) | ( ~n6387 & n6396 ) ;
  assign n6398 = n4202 & ~n5270 ;
  assign n6399 = n2552 & n4345 ;
  assign n6400 = ~n2491 & n4201 ;
  assign n6401 = n2635 & n4200 ;
  assign n6402 = n6400 | n6401 ;
  assign n6403 = ( ~n6398 & n6399 ) | ( ~n6398 & n6402 ) | ( n6399 & n6402 ) ;
  assign n6404 = ( ~x26 & n6398 ) | ( ~x26 & n6403 ) | ( n6398 & n6403 ) ;
  assign n6405 = ( n6398 & n6403 ) | ( n6398 & ~n6404 ) | ( n6403 & ~n6404 ) ;
  assign n6406 = ( x26 & n6404 ) | ( x26 & ~n6405 ) | ( n6404 & ~n6405 ) ;
  assign n6407 = ( n6282 & ~n6284 ) | ( n6282 & n6293 ) | ( ~n6284 & n6293 ) ;
  assign n6408 = ( n6284 & ~n6294 ) | ( n6284 & n6407 ) | ( ~n6294 & n6407 ) ;
  assign n6409 = ( n6397 & n6406 ) | ( n6397 & n6408 ) | ( n6406 & n6408 ) ;
  assign n6410 = ( ~n6294 & n6296 ) | ( ~n6294 & n6305 ) | ( n6296 & n6305 ) ;
  assign n6411 = ( ~n6305 & n6306 ) | ( ~n6305 & n6410 ) | ( n6306 & n6410 ) ;
  assign n6412 = n4647 & n4713 ;
  assign n6413 = n2174 & n4712 ;
  assign n6414 = n2298 | n4709 ;
  assign n6415 = n2270 & n4792 ;
  assign n6416 = ( ~n2298 & n6414 ) | ( ~n2298 & n6415 ) | ( n6414 & n6415 ) ;
  assign n6417 = ( ~n6412 & n6413 ) | ( ~n6412 & n6416 ) | ( n6413 & n6416 ) ;
  assign n6418 = ( ~x23 & n6412 ) | ( ~x23 & n6417 ) | ( n6412 & n6417 ) ;
  assign n6419 = ( n6412 & n6417 ) | ( n6412 & ~n6418 ) | ( n6417 & ~n6418 ) ;
  assign n6420 = ( x23 & n6418 ) | ( x23 & ~n6419 ) | ( n6418 & ~n6419 ) ;
  assign n6421 = ( n6409 & ~n6411 ) | ( n6409 & n6420 ) | ( ~n6411 & n6420 ) ;
  assign n6422 = ( ~n6306 & n6308 ) | ( ~n6306 & n6317 ) | ( n6308 & n6317 ) ;
  assign n6423 = ( n6306 & ~n6318 ) | ( n6306 & n6422 ) | ( ~n6318 & n6422 ) ;
  assign n6424 = n4290 & n4974 ;
  assign n6425 = n1852 & n5398 ;
  assign n6426 = n2023 | n4973 ;
  assign n6427 = n1926 & n4972 ;
  assign n6428 = ( ~n2023 & n6426 ) | ( ~n2023 & n6427 ) | ( n6426 & n6427 ) ;
  assign n6429 = ( ~n6424 & n6425 ) | ( ~n6424 & n6428 ) | ( n6425 & n6428 ) ;
  assign n6430 = ( ~x20 & n6424 ) | ( ~x20 & n6429 ) | ( n6424 & n6429 ) ;
  assign n6431 = ( n6424 & n6429 ) | ( n6424 & ~n6430 ) | ( n6429 & ~n6430 ) ;
  assign n6432 = ( x20 & n6430 ) | ( x20 & ~n6431 ) | ( n6430 & ~n6431 ) ;
  assign n6433 = ( n6421 & n6423 ) | ( n6421 & n6432 ) | ( n6423 & n6432 ) ;
  assign n6434 = ( ~n6318 & n6327 ) | ( ~n6318 & n6329 ) | ( n6327 & n6329 ) ;
  assign n6435 = ( n6318 & ~n6330 ) | ( n6318 & n6434 ) | ( ~n6330 & n6434 ) ;
  assign n6436 = ~n4302 & n4974 ;
  assign n6437 = ~n1750 & n5398 ;
  assign n6438 = n1926 & ~n4973 ;
  assign n6439 = n1852 & n4972 ;
  assign n6440 = ( n1926 & ~n6438 ) | ( n1926 & n6439 ) | ( ~n6438 & n6439 ) ;
  assign n6441 = ( ~n6436 & n6437 ) | ( ~n6436 & n6440 ) | ( n6437 & n6440 ) ;
  assign n6442 = ( ~x20 & n6436 ) | ( ~x20 & n6441 ) | ( n6436 & n6441 ) ;
  assign n6443 = ( n6436 & n6441 ) | ( n6436 & ~n6442 ) | ( n6441 & ~n6442 ) ;
  assign n6444 = ( x20 & n6442 ) | ( x20 & ~n6443 ) | ( n6442 & ~n6443 ) ;
  assign n6445 = ( n6433 & n6435 ) | ( n6433 & n6444 ) | ( n6435 & n6444 ) ;
  assign n6446 = ( n6330 & ~n6332 ) | ( n6330 & n6341 ) | ( ~n6332 & n6341 ) ;
  assign n6447 = ( n6332 & ~n6342 ) | ( n6332 & n6446 ) | ( ~n6342 & n6446 ) ;
  assign n6448 = ~n3955 & n5508 ;
  assign n6449 = ~n1338 & n5507 ;
  assign n6450 = n1458 & n5666 ;
  assign n6451 = n1576 & n5504 ;
  assign n6452 = n6450 | n6451 ;
  assign n6453 = ( ~n6448 & n6449 ) | ( ~n6448 & n6452 ) | ( n6449 & n6452 ) ;
  assign n6454 = ( ~x17 & n6448 ) | ( ~x17 & n6453 ) | ( n6448 & n6453 ) ;
  assign n6455 = ( n6448 & n6453 ) | ( n6448 & ~n6454 ) | ( n6453 & ~n6454 ) ;
  assign n6456 = ( x17 & n6454 ) | ( x17 & ~n6455 ) | ( n6454 & ~n6455 ) ;
  assign n6457 = ( n6445 & n6447 ) | ( n6445 & n6456 ) | ( n6447 & n6456 ) ;
  assign n6458 = ( n6342 & ~n6344 ) | ( n6342 & n6353 ) | ( ~n6344 & n6353 ) ;
  assign n6459 = ( n6344 & ~n6354 ) | ( n6344 & n6458 ) | ( ~n6354 & n6458 ) ;
  assign n6460 = ~n3665 & n5966 ;
  assign n6461 = ~n1290 & n5969 ;
  assign n6462 = ~n1246 & n5970 ;
  assign n6463 = ~n5963 & n5964 ;
  assign n6464 = ( ~n5960 & n5961 ) | ( ~n5960 & n6463 ) | ( n5961 & n6463 ) ;
  assign n6465 = ~n3658 & n6464 ;
  assign n6466 = n6462 | n6465 ;
  assign n6467 = ( ~n6460 & n6461 ) | ( ~n6460 & n6466 ) | ( n6461 & n6466 ) ;
  assign n6468 = ( ~x14 & n6460 ) | ( ~x14 & n6467 ) | ( n6460 & n6467 ) ;
  assign n6469 = ( n6460 & n6467 ) | ( n6460 & ~n6468 ) | ( n6467 & ~n6468 ) ;
  assign n6470 = ( x14 & n6468 ) | ( x14 & ~n6469 ) | ( n6468 & ~n6469 ) ;
  assign n6471 = ( n6457 & n6459 ) | ( n6457 & n6470 ) | ( n6459 & n6470 ) ;
  assign n6472 = n3692 & n6464 ;
  assign n6473 = ~n3658 & n5969 ;
  assign n6474 = ( n6464 & ~n6472 ) | ( n6464 & n6473 ) | ( ~n6472 & n6473 ) ;
  assign n6475 = ~n1290 & n5970 ;
  assign n6476 = n6474 | n6475 ;
  assign n6477 = ~n4182 & n5966 ;
  assign n6478 = ( x14 & n6476 ) | ( x14 & ~n6477 ) | ( n6476 & ~n6477 ) ;
  assign n6479 = ( ~x14 & n6476 ) | ( ~x14 & n6477 ) | ( n6476 & n6477 ) ;
  assign n6480 = ( ~n6476 & n6478 ) | ( ~n6476 & n6479 ) | ( n6478 & n6479 ) ;
  assign n6481 = ( ~n6354 & n6363 ) | ( ~n6354 & n6365 ) | ( n6363 & n6365 ) ;
  assign n6482 = ( n6354 & ~n6366 ) | ( n6354 & n6481 ) | ( ~n6366 & n6481 ) ;
  assign n6483 = ( n6471 & n6480 ) | ( n6471 & n6482 ) | ( n6480 & n6482 ) ;
  assign n6484 = n3800 & n5543 ;
  assign n6485 = ~n2910 & n3802 ;
  assign n6486 = n2965 & n3700 ;
  assign n6487 = n2843 & n3799 ;
  assign n6488 = ( n3700 & ~n6486 ) | ( n3700 & n6487 ) | ( ~n6486 & n6487 ) ;
  assign n6489 = ( ~n6484 & n6485 ) | ( ~n6484 & n6488 ) | ( n6485 & n6488 ) ;
  assign n6490 = ( ~x29 & n6484 ) | ( ~x29 & n6489 ) | ( n6484 & n6489 ) ;
  assign n6491 = ( n6484 & n6489 ) | ( n6484 & ~n6490 ) | ( n6489 & ~n6490 ) ;
  assign n6492 = ( x29 & n6490 ) | ( x29 & ~n6491 ) | ( n6490 & ~n6491 ) ;
  assign n6493 = ( ~n6258 & n6260 ) | ( ~n6258 & n6269 ) | ( n6260 & n6269 ) ;
  assign n6494 = ( n6258 & ~n6270 ) | ( n6258 & n6493 ) | ( ~n6270 & n6493 ) ;
  assign n6495 = n4202 & n5232 ;
  assign n6496 = ~n2810 & n4200 ;
  assign n6497 = n2635 & ~n4201 ;
  assign n6498 = ~n2725 & n4345 ;
  assign n6499 = ( n2635 & ~n6497 ) | ( n2635 & n6498 ) | ( ~n6497 & n6498 ) ;
  assign n6500 = ( ~n6495 & n6496 ) | ( ~n6495 & n6499 ) | ( n6496 & n6499 ) ;
  assign n6501 = ( ~x26 & n6495 ) | ( ~x26 & n6500 ) | ( n6495 & n6500 ) ;
  assign n6502 = ( n6495 & n6500 ) | ( n6495 & ~n6501 ) | ( n6500 & ~n6501 ) ;
  assign n6503 = ( x26 & n6501 ) | ( x26 & ~n6502 ) | ( n6501 & ~n6502 ) ;
  assign n6504 = ( n6492 & n6494 ) | ( n6492 & n6503 ) | ( n6494 & n6503 ) ;
  assign n6505 = ( ~n6385 & n6387 ) | ( ~n6385 & n6396 ) | ( n6387 & n6396 ) ;
  assign n6506 = ( ~n6396 & n6397 ) | ( ~n6396 & n6505 ) | ( n6397 & n6505 ) ;
  assign n6507 = n4713 & ~n4900 ;
  assign n6508 = n2396 & n4792 ;
  assign n6509 = ~n2298 & n4712 ;
  assign n6510 = ~n2491 & n4709 ;
  assign n6511 = n6509 | n6510 ;
  assign n6512 = ( ~n6507 & n6508 ) | ( ~n6507 & n6511 ) | ( n6508 & n6511 ) ;
  assign n6513 = ( ~x23 & n6507 ) | ( ~x23 & n6512 ) | ( n6507 & n6512 ) ;
  assign n6514 = ( n6507 & n6512 ) | ( n6507 & ~n6513 ) | ( n6512 & ~n6513 ) ;
  assign n6515 = ( x23 & n6513 ) | ( x23 & ~n6514 ) | ( n6513 & ~n6514 ) ;
  assign n6516 = ( n6504 & ~n6506 ) | ( n6504 & n6515 ) | ( ~n6506 & n6515 ) ;
  assign n6517 = n2298 | n4792 ;
  assign n6518 = n2270 & n4712 ;
  assign n6519 = ( ~n2298 & n6517 ) | ( ~n2298 & n6518 ) | ( n6517 & n6518 ) ;
  assign n6520 = ~n2396 & n4709 ;
  assign n6521 = ( n4709 & n6519 ) | ( n4709 & ~n6520 ) | ( n6519 & ~n6520 ) ;
  assign n6522 = ( n4713 & ~n4912 ) | ( n4713 & n6521 ) | ( ~n4912 & n6521 ) ;
  assign n6523 = n6521 & ~n6522 ;
  assign n6524 = ( ~x23 & n6522 ) | ( ~x23 & n6523 ) | ( n6522 & n6523 ) ;
  assign n6525 = ( n6522 & n6523 ) | ( n6522 & ~n6524 ) | ( n6523 & ~n6524 ) ;
  assign n6526 = ( x23 & n6524 ) | ( x23 & ~n6525 ) | ( n6524 & ~n6525 ) ;
  assign n6527 = ( ~n6397 & n6406 ) | ( ~n6397 & n6408 ) | ( n6406 & n6408 ) ;
  assign n6528 = ( n6397 & ~n6409 ) | ( n6397 & n6527 ) | ( ~n6409 & n6527 ) ;
  assign n6529 = ( n6516 & n6526 ) | ( n6516 & n6528 ) | ( n6526 & n6528 ) ;
  assign n6530 = ( ~n6409 & n6411 ) | ( ~n6409 & n6420 ) | ( n6411 & n6420 ) ;
  assign n6531 = ( ~n6420 & n6421 ) | ( ~n6420 & n6530 ) | ( n6421 & n6530 ) ;
  assign n6532 = ~n4457 & n4974 ;
  assign n6533 = n1926 & n5398 ;
  assign n6534 = n2089 & ~n4973 ;
  assign n6535 = ~n2023 & n4972 ;
  assign n6536 = ( n2089 & ~n6534 ) | ( n2089 & n6535 ) | ( ~n6534 & n6535 ) ;
  assign n6537 = ( ~n6532 & n6533 ) | ( ~n6532 & n6536 ) | ( n6533 & n6536 ) ;
  assign n6538 = ( ~x20 & n6532 ) | ( ~x20 & n6537 ) | ( n6532 & n6537 ) ;
  assign n6539 = ( n6532 & n6537 ) | ( n6532 & ~n6538 ) | ( n6537 & ~n6538 ) ;
  assign n6540 = ( x20 & n6538 ) | ( x20 & ~n6539 ) | ( n6538 & ~n6539 ) ;
  assign n6541 = ( n6529 & ~n6531 ) | ( n6529 & n6540 ) | ( ~n6531 & n6540 ) ;
  assign n6542 = ( ~n6421 & n6423 ) | ( ~n6421 & n6432 ) | ( n6423 & n6432 ) ;
  assign n6543 = ( n6421 & ~n6433 ) | ( n6421 & n6542 ) | ( ~n6433 & n6542 ) ;
  assign n6544 = n4326 & n5508 ;
  assign n6545 = n1576 & n5507 ;
  assign n6546 = n1750 | n5504 ;
  assign n6547 = ~n1669 & n5666 ;
  assign n6548 = ( ~n1750 & n6546 ) | ( ~n1750 & n6547 ) | ( n6546 & n6547 ) ;
  assign n6549 = ( ~n6544 & n6545 ) | ( ~n6544 & n6548 ) | ( n6545 & n6548 ) ;
  assign n6550 = ( ~x17 & n6544 ) | ( ~x17 & n6549 ) | ( n6544 & n6549 ) ;
  assign n6551 = ( n6544 & n6549 ) | ( n6544 & ~n6550 ) | ( n6549 & ~n6550 ) ;
  assign n6552 = ( x17 & n6550 ) | ( x17 & ~n6551 ) | ( n6550 & ~n6551 ) ;
  assign n6553 = ( n6541 & n6543 ) | ( n6541 & n6552 ) | ( n6543 & n6552 ) ;
  assign n6554 = ~n4159 & n5508 ;
  assign n6555 = n1458 & n5507 ;
  assign n6556 = ~n1669 & n5504 ;
  assign n6557 = n1576 & n5666 ;
  assign n6558 = n6556 | n6557 ;
  assign n6559 = ( ~n6554 & n6555 ) | ( ~n6554 & n6558 ) | ( n6555 & n6558 ) ;
  assign n6560 = ( ~x17 & n6554 ) | ( ~x17 & n6559 ) | ( n6554 & n6559 ) ;
  assign n6561 = ( n6554 & n6559 ) | ( n6554 & ~n6560 ) | ( n6559 & ~n6560 ) ;
  assign n6562 = ( x17 & n6560 ) | ( x17 & ~n6561 ) | ( n6560 & ~n6561 ) ;
  assign n6563 = ( ~n6433 & n6435 ) | ( ~n6433 & n6444 ) | ( n6435 & n6444 ) ;
  assign n6564 = ( n6433 & ~n6445 ) | ( n6433 & n6563 ) | ( ~n6445 & n6563 ) ;
  assign n6565 = ( n6553 & n6562 ) | ( n6553 & n6564 ) | ( n6562 & n6564 ) ;
  assign n6566 = ( n6445 & ~n6447 ) | ( n6445 & n6456 ) | ( ~n6447 & n6456 ) ;
  assign n6567 = ( n6447 & ~n6457 ) | ( n6447 & n6566 ) | ( ~n6457 & n6566 ) ;
  assign n6568 = n3621 & n5966 ;
  assign n6569 = ~n1290 & n6464 ;
  assign n6570 = n1267 & ~n5970 ;
  assign n6571 = ~n1246 & n5969 ;
  assign n6572 = ( n1267 & ~n6570 ) | ( n1267 & n6571 ) | ( ~n6570 & n6571 ) ;
  assign n6573 = ( ~n6568 & n6569 ) | ( ~n6568 & n6572 ) | ( n6569 & n6572 ) ;
  assign n6574 = ( ~x14 & n6568 ) | ( ~x14 & n6573 ) | ( n6568 & n6573 ) ;
  assign n6575 = ( n6568 & n6573 ) | ( n6568 & ~n6574 ) | ( n6573 & ~n6574 ) ;
  assign n6576 = ( x14 & n6574 ) | ( x14 & ~n6575 ) | ( n6574 & ~n6575 ) ;
  assign n6577 = ( n6565 & n6567 ) | ( n6565 & n6576 ) | ( n6567 & n6576 ) ;
  assign n6578 = x10 | x11 ;
  assign n6579 = x10 & x11 ;
  assign n6580 = n6578 & ~n6579 ;
  assign n6581 = x8 & x9 ;
  assign n6582 = x8 | x9 ;
  assign n6583 = ( n6580 & n6581 ) | ( n6580 & ~n6582 ) | ( n6581 & ~n6582 ) ;
  assign n6584 = n6580 & ~n6583 ;
  assign n6585 = x9 | x10 ;
  assign n6586 = x8 & ~x10 ;
  assign n6587 = ( ~n6582 & n6585 ) | ( ~n6582 & n6586 ) | ( n6585 & n6586 ) ;
  assign n6588 = n6583 & ~n6587 ;
  assign n6589 = ~n3692 & n6588 ;
  assign n6590 = ( n3691 & n3692 ) | ( n3691 & n6584 ) | ( n3692 & n6584 ) ;
  assign n6591 = ( n6584 & n6589 ) | ( n6584 & ~n6590 ) | ( n6589 & ~n6590 ) ;
  assign n6592 = x11 | n6591 ;
  assign n6593 = ( x11 & n6591 ) | ( x11 & ~n6592 ) | ( n6591 & ~n6592 ) ;
  assign n6594 = n6592 & ~n6593 ;
  assign n6595 = ( n6457 & ~n6459 ) | ( n6457 & n6470 ) | ( ~n6459 & n6470 ) ;
  assign n6596 = ( n6459 & ~n6471 ) | ( n6459 & n6595 ) | ( ~n6471 & n6595 ) ;
  assign n6597 = ( n6577 & n6594 ) | ( n6577 & n6596 ) | ( n6594 & n6596 ) ;
  assign n6598 = ( n58 & n96 ) | ( n58 & ~n3586 ) | ( n96 & ~n3586 ) ;
  assign n6599 = n3800 & n6061 ;
  assign n6600 = n3479 & n3802 ;
  assign n6601 = n3533 & n3700 ;
  assign n6602 = ~n3389 & n3799 ;
  assign n6603 = ( n3700 & ~n6601 ) | ( n3700 & n6602 ) | ( ~n6601 & n6602 ) ;
  assign n6604 = ( ~n6599 & n6600 ) | ( ~n6599 & n6603 ) | ( n6600 & n6603 ) ;
  assign n6605 = ( ~x29 & n6599 ) | ( ~x29 & n6604 ) | ( n6599 & n6604 ) ;
  assign n6606 = ( n6599 & n6604 ) | ( n6599 & ~n6605 ) | ( n6604 & ~n6605 ) ;
  assign n6607 = ( x29 & n6605 ) | ( x29 & ~n6606 ) | ( n6605 & ~n6606 ) ;
  assign n6608 = n3479 & n6009 ;
  assign n6609 = ( n3479 & n3800 ) | ( n3479 & n6009 ) | ( n3800 & n6009 ) ;
  assign n6610 = ~n3533 & n3802 ;
  assign n6611 = ( n3586 & n3694 ) | ( n3586 & n3699 ) | ( n3694 & n3699 ) ;
  assign n6612 = ( n3694 & n6610 ) | ( n3694 & ~n6611 ) | ( n6610 & ~n6611 ) ;
  assign n6613 = n3479 & ~n3799 ;
  assign n6614 = ( n3479 & n6612 ) | ( n3479 & ~n6613 ) | ( n6612 & ~n6613 ) ;
  assign n6615 = ( ~n6608 & n6609 ) | ( ~n6608 & n6614 ) | ( n6609 & n6614 ) ;
  assign n6616 = ~n3586 & n3697 ;
  assign n6617 = x29 & n6616 ;
  assign n6618 = n3533 & ~n3586 ;
  assign n6619 = ( n3800 & n6009 ) | ( n3800 & n6618 ) | ( n6009 & n6618 ) ;
  assign n6620 = ~n3533 & n3799 ;
  assign n6621 = n3586 | n3802 ;
  assign n6622 = ( ~n3586 & n6620 ) | ( ~n3586 & n6621 ) | ( n6620 & n6621 ) ;
  assign n6623 = n6619 | n6622 ;
  assign n6624 = ( x29 & n6617 ) | ( x29 & n6623 ) | ( n6617 & n6623 ) ;
  assign n6625 = n6615 | n6624 ;
  assign n6626 = x29 & ~n6625 ;
  assign n6627 = ( n6598 & n6607 ) | ( n6598 & n6626 ) | ( n6607 & n6626 ) ;
  assign n6628 = ( n1248 & n6009 ) | ( n1248 & n6618 ) | ( n6009 & n6618 ) ;
  assign n6629 = ( n1250 & ~n3586 ) | ( n1250 & n6628 ) | ( ~n3586 & n6628 ) ;
  assign n6630 = ( n606 & ~n3533 ) | ( n606 & n6628 ) | ( ~n3533 & n6628 ) ;
  assign n6631 = n6629 | n6630 ;
  assign n6632 = n3800 & ~n6104 ;
  assign n6633 = n3479 & n3700 ;
  assign n6634 = ~n3355 & n3799 ;
  assign n6635 = n3389 | n3802 ;
  assign n6636 = ( ~n3389 & n6634 ) | ( ~n3389 & n6635 ) | ( n6634 & n6635 ) ;
  assign n6637 = ( ~n6632 & n6633 ) | ( ~n6632 & n6636 ) | ( n6633 & n6636 ) ;
  assign n6638 = ( ~x29 & n6632 ) | ( ~x29 & n6637 ) | ( n6632 & n6637 ) ;
  assign n6639 = ( n6632 & n6637 ) | ( n6632 & ~n6638 ) | ( n6637 & ~n6638 ) ;
  assign n6640 = ( x29 & n6638 ) | ( x29 & ~n6639 ) | ( n6638 & ~n6639 ) ;
  assign n6641 = ( n6627 & n6631 ) | ( n6627 & n6640 ) | ( n6631 & n6640 ) ;
  assign n6642 = n3800 & ~n6154 ;
  assign n6643 = ~n3300 & n3799 ;
  assign n6644 = ~n3355 & n3802 ;
  assign n6645 = ( n3389 & n3694 ) | ( n3389 & n3699 ) | ( n3694 & n3699 ) ;
  assign n6646 = ( n3694 & n6644 ) | ( n3694 & ~n6645 ) | ( n6644 & ~n6645 ) ;
  assign n6647 = ( ~n6642 & n6643 ) | ( ~n6642 & n6646 ) | ( n6643 & n6646 ) ;
  assign n6648 = ( ~x29 & n6642 ) | ( ~x29 & n6647 ) | ( n6642 & n6647 ) ;
  assign n6649 = ( n6642 & n6647 ) | ( n6642 & ~n6648 ) | ( n6647 & ~n6648 ) ;
  assign n6650 = ( x29 & n6648 ) | ( x29 & ~n6649 ) | ( n6648 & ~n6649 ) ;
  assign n6651 = n6003 & n6011 ;
  assign n6652 = ( n6003 & n6012 ) | ( n6003 & ~n6651 ) | ( n6012 & ~n6651 ) ;
  assign n6653 = ( n6641 & n6650 ) | ( n6641 & ~n6652 ) | ( n6650 & ~n6652 ) ;
  assign n6654 = n3800 & n6200 ;
  assign n6655 = ~n3300 & n3802 ;
  assign n6656 = n3355 & n3700 ;
  assign n6657 = n3239 & n3799 ;
  assign n6658 = ( n3700 & ~n6656 ) | ( n3700 & n6657 ) | ( ~n6656 & n6657 ) ;
  assign n6659 = ( ~n6654 & n6655 ) | ( ~n6654 & n6658 ) | ( n6655 & n6658 ) ;
  assign n6660 = ( ~x29 & n6654 ) | ( ~x29 & n6659 ) | ( n6654 & n6659 ) ;
  assign n6661 = ( n6654 & n6659 ) | ( n6654 & ~n6660 ) | ( n6659 & ~n6660 ) ;
  assign n6662 = ( x29 & n6660 ) | ( x29 & ~n6661 ) | ( n6660 & ~n6661 ) ;
  assign n6663 = ( ~n6012 & n6054 ) | ( ~n6012 & n6063 ) | ( n6054 & n6063 ) ;
  assign n6664 = ( ~n6063 & n6064 ) | ( ~n6063 & n6663 ) | ( n6064 & n6663 ) ;
  assign n6665 = ( n6653 & n6662 ) | ( n6653 & ~n6664 ) | ( n6662 & ~n6664 ) ;
  assign n6666 = n3800 & ~n6243 ;
  assign n6667 = n3153 & n3799 ;
  assign n6668 = n3239 & n3802 ;
  assign n6669 = ( n3300 & n3694 ) | ( n3300 & n3699 ) | ( n3694 & n3699 ) ;
  assign n6670 = ( n3694 & n6668 ) | ( n3694 & ~n6669 ) | ( n6668 & ~n6669 ) ;
  assign n6671 = ( ~n6666 & n6667 ) | ( ~n6666 & n6670 ) | ( n6667 & n6670 ) ;
  assign n6672 = ( ~x29 & n6666 ) | ( ~x29 & n6671 ) | ( n6666 & n6671 ) ;
  assign n6673 = ( n6666 & n6671 ) | ( n6666 & ~n6672 ) | ( n6671 & ~n6672 ) ;
  assign n6674 = ( x29 & n6672 ) | ( x29 & ~n6673 ) | ( n6672 & ~n6673 ) ;
  assign n6675 = ( ~n6064 & n6097 ) | ( ~n6064 & n6106 ) | ( n6097 & n6106 ) ;
  assign n6676 = ( n6064 & ~n6107 ) | ( n6064 & n6675 ) | ( ~n6107 & n6675 ) ;
  assign n6677 = ( n6665 & n6674 ) | ( n6665 & n6676 ) | ( n6674 & n6676 ) ;
  assign n6678 = n3800 & n5710 ;
  assign n6679 = n3153 & n3802 ;
  assign n6680 = n3078 & n3799 ;
  assign n6681 = ( ~n3239 & n3694 ) | ( ~n3239 & n3699 ) | ( n3694 & n3699 ) ;
  assign n6682 = ( n3694 & n6680 ) | ( n3694 & ~n6681 ) | ( n6680 & ~n6681 ) ;
  assign n6683 = ( ~n6678 & n6679 ) | ( ~n6678 & n6682 ) | ( n6679 & n6682 ) ;
  assign n6684 = ( ~x29 & n6678 ) | ( ~x29 & n6683 ) | ( n6678 & n6683 ) ;
  assign n6685 = ( n6678 & n6683 ) | ( n6678 & ~n6684 ) | ( n6683 & ~n6684 ) ;
  assign n6686 = ( x29 & n6684 ) | ( x29 & ~n6685 ) | ( n6684 & ~n6685 ) ;
  assign n6687 = ( ~n6107 & n6147 ) | ( ~n6107 & n6156 ) | ( n6147 & n6156 ) ;
  assign n6688 = ( ~n6156 & n6157 ) | ( ~n6156 & n6687 ) | ( n6157 & n6687 ) ;
  assign n6689 = ( n6677 & n6686 ) | ( n6677 & ~n6688 ) | ( n6686 & ~n6688 ) ;
  assign n6690 = n3800 & ~n6267 ;
  assign n6691 = n3153 & n3700 ;
  assign n6692 = n3078 & ~n3802 ;
  assign n6693 = ~n3046 & n3799 ;
  assign n6694 = ( n3078 & ~n6692 ) | ( n3078 & n6693 ) | ( ~n6692 & n6693 ) ;
  assign n6695 = ( ~n6690 & n6691 ) | ( ~n6690 & n6694 ) | ( n6691 & n6694 ) ;
  assign n6696 = ( ~x29 & n6690 ) | ( ~x29 & n6695 ) | ( n6690 & n6695 ) ;
  assign n6697 = ( n6690 & n6695 ) | ( n6690 & ~n6696 ) | ( n6695 & ~n6696 ) ;
  assign n6698 = ( x29 & n6696 ) | ( x29 & ~n6697 ) | ( n6696 & ~n6697 ) ;
  assign n6699 = ( ~n6157 & n6193 ) | ( ~n6157 & n6202 ) | ( n6193 & n6202 ) ;
  assign n6700 = ( n6157 & ~n6203 ) | ( n6157 & n6699 ) | ( ~n6203 & n6699 ) ;
  assign n6701 = ( n6689 & n6698 ) | ( n6689 & n6700 ) | ( n6698 & n6700 ) ;
  assign n6702 = n3800 & n6279 ;
  assign n6703 = ~n2965 & n3799 ;
  assign n6704 = n3078 & n3700 ;
  assign n6705 = ~n3046 & n3802 ;
  assign n6706 = n6704 | n6705 ;
  assign n6707 = ( ~n6702 & n6703 ) | ( ~n6702 & n6706 ) | ( n6703 & n6706 ) ;
  assign n6708 = ( ~x29 & n6702 ) | ( ~x29 & n6707 ) | ( n6702 & n6707 ) ;
  assign n6709 = ( n6702 & n6707 ) | ( n6702 & ~n6708 ) | ( n6707 & ~n6708 ) ;
  assign n6710 = ( x29 & n6708 ) | ( x29 & ~n6709 ) | ( n6708 & ~n6709 ) ;
  assign n6711 = ( ~n6203 & n6236 ) | ( ~n6203 & n6245 ) | ( n6236 & n6245 ) ;
  assign n6712 = ( n6203 & ~n6246 ) | ( n6203 & n6711 ) | ( ~n6246 & n6711 ) ;
  assign n6713 = ( n6701 & n6710 ) | ( n6701 & n6712 ) | ( n6710 & n6712 ) ;
  assign n6714 = ( n6246 & ~n6248 ) | ( n6246 & n6257 ) | ( ~n6248 & n6257 ) ;
  assign n6715 = ( n6248 & ~n6258 ) | ( n6248 & n6714 ) | ( ~n6258 & n6714 ) ;
  assign n6716 = n4202 & ~n5586 ;
  assign n6717 = ~n2725 & n4201 ;
  assign n6718 = n2843 & n4200 ;
  assign n6719 = ~n2810 & n4345 ;
  assign n6720 = n6718 | n6719 ;
  assign n6721 = ( ~n6716 & n6717 ) | ( ~n6716 & n6720 ) | ( n6717 & n6720 ) ;
  assign n6722 = ( ~x26 & n6716 ) | ( ~x26 & n6721 ) | ( n6716 & n6721 ) ;
  assign n6723 = ( n6716 & n6721 ) | ( n6716 & ~n6722 ) | ( n6721 & ~n6722 ) ;
  assign n6724 = ( x26 & n6722 ) | ( x26 & ~n6723 ) | ( n6722 & ~n6723 ) ;
  assign n6725 = ( n6713 & n6715 ) | ( n6713 & n6724 ) | ( n6715 & n6724 ) ;
  assign n6726 = ( n6492 & ~n6494 ) | ( n6492 & n6503 ) | ( ~n6494 & n6503 ) ;
  assign n6727 = ( n6494 & ~n6504 ) | ( n6494 & n6726 ) | ( ~n6504 & n6726 ) ;
  assign n6728 = n4713 & ~n5084 ;
  assign n6729 = n2396 & n4712 ;
  assign n6730 = ~n2491 & n4792 ;
  assign n6731 = n2552 & n4709 ;
  assign n6732 = n6730 | n6731 ;
  assign n6733 = ( ~n6728 & n6729 ) | ( ~n6728 & n6732 ) | ( n6729 & n6732 ) ;
  assign n6734 = ( ~x23 & n6728 ) | ( ~x23 & n6733 ) | ( n6728 & n6733 ) ;
  assign n6735 = ( n6728 & n6733 ) | ( n6728 & ~n6734 ) | ( n6733 & ~n6734 ) ;
  assign n6736 = ( x23 & n6734 ) | ( x23 & ~n6735 ) | ( n6734 & ~n6735 ) ;
  assign n6737 = ( n6725 & n6727 ) | ( n6725 & n6736 ) | ( n6727 & n6736 ) ;
  assign n6738 = ( ~n6504 & n6506 ) | ( ~n6504 & n6515 ) | ( n6506 & n6515 ) ;
  assign n6739 = ( ~n6515 & n6516 ) | ( ~n6515 & n6738 ) | ( n6516 & n6738 ) ;
  assign n6740 = n4730 & n4974 ;
  assign n6741 = n2089 & n5398 ;
  assign n6742 = n2270 & ~n4973 ;
  assign n6743 = n2174 & n4972 ;
  assign n6744 = ( n2270 & ~n6742 ) | ( n2270 & n6743 ) | ( ~n6742 & n6743 ) ;
  assign n6745 = ( ~n6740 & n6741 ) | ( ~n6740 & n6744 ) | ( n6741 & n6744 ) ;
  assign n6746 = ( ~x20 & n6740 ) | ( ~x20 & n6745 ) | ( n6740 & n6745 ) ;
  assign n6747 = ( n6740 & n6745 ) | ( n6740 & ~n6746 ) | ( n6745 & ~n6746 ) ;
  assign n6748 = ( x20 & n6746 ) | ( x20 & ~n6747 ) | ( n6746 & ~n6747 ) ;
  assign n6749 = ( n6737 & ~n6739 ) | ( n6737 & n6748 ) | ( ~n6739 & n6748 ) ;
  assign n6750 = ( ~n6516 & n6526 ) | ( ~n6516 & n6528 ) | ( n6526 & n6528 ) ;
  assign n6751 = ( n6516 & ~n6529 ) | ( n6516 & n6750 ) | ( ~n6529 & n6750 ) ;
  assign n6752 = ~n4660 & n4974 ;
  assign n6753 = ~n2023 & n5398 ;
  assign n6754 = n2174 & ~n4973 ;
  assign n6755 = n2089 & n4972 ;
  assign n6756 = ( n2174 & ~n6754 ) | ( n2174 & n6755 ) | ( ~n6754 & n6755 ) ;
  assign n6757 = ( ~n6752 & n6753 ) | ( ~n6752 & n6756 ) | ( n6753 & n6756 ) ;
  assign n6758 = ( ~x20 & n6752 ) | ( ~x20 & n6757 ) | ( n6752 & n6757 ) ;
  assign n6759 = ( n6752 & n6757 ) | ( n6752 & ~n6758 ) | ( n6757 & ~n6758 ) ;
  assign n6760 = ( x20 & n6758 ) | ( x20 & ~n6759 ) | ( n6758 & ~n6759 ) ;
  assign n6761 = ( n6749 & n6751 ) | ( n6749 & n6760 ) | ( n6751 & n6760 ) ;
  assign n6762 = ( ~n6529 & n6531 ) | ( ~n6529 & n6540 ) | ( n6531 & n6540 ) ;
  assign n6763 = ( ~n6540 & n6541 ) | ( ~n6540 & n6762 ) | ( n6541 & n6762 ) ;
  assign n6764 = n4146 & n5508 ;
  assign n6765 = ~n1669 & n5507 ;
  assign n6766 = n1852 & ~n5504 ;
  assign n6767 = ~n1750 & n5666 ;
  assign n6768 = ( n1852 & ~n6766 ) | ( n1852 & n6767 ) | ( ~n6766 & n6767 ) ;
  assign n6769 = ( ~n6764 & n6765 ) | ( ~n6764 & n6768 ) | ( n6765 & n6768 ) ;
  assign n6770 = ( ~x17 & n6764 ) | ( ~x17 & n6769 ) | ( n6764 & n6769 ) ;
  assign n6771 = ( n6764 & n6769 ) | ( n6764 & ~n6770 ) | ( n6769 & ~n6770 ) ;
  assign n6772 = ( x17 & n6770 ) | ( x17 & ~n6771 ) | ( n6770 & ~n6771 ) ;
  assign n6773 = ( n6761 & ~n6763 ) | ( n6761 & n6772 ) | ( ~n6763 & n6772 ) ;
  assign n6774 = ( n6541 & ~n6543 ) | ( n6541 & n6552 ) | ( ~n6543 & n6552 ) ;
  assign n6775 = ( n6543 & ~n6553 ) | ( n6543 & n6774 ) | ( ~n6553 & n6774 ) ;
  assign n6776 = ~n3779 & n5966 ;
  assign n6777 = n1267 & n6464 ;
  assign n6778 = n1458 & ~n5970 ;
  assign n6779 = ~n1338 & n5969 ;
  assign n6780 = ( n1458 & ~n6778 ) | ( n1458 & n6779 ) | ( ~n6778 & n6779 ) ;
  assign n6781 = ( ~n6776 & n6777 ) | ( ~n6776 & n6780 ) | ( n6777 & n6780 ) ;
  assign n6782 = ( ~x14 & n6776 ) | ( ~x14 & n6781 ) | ( n6776 & n6781 ) ;
  assign n6783 = ( n6776 & n6781 ) | ( n6776 & ~n6782 ) | ( n6781 & ~n6782 ) ;
  assign n6784 = ( x14 & n6782 ) | ( x14 & ~n6783 ) | ( n6782 & ~n6783 ) ;
  assign n6785 = ( n6773 & n6775 ) | ( n6773 & n6784 ) | ( n6775 & n6784 ) ;
  assign n6786 = ( ~n6553 & n6562 ) | ( ~n6553 & n6564 ) | ( n6562 & n6564 ) ;
  assign n6787 = ( n6553 & ~n6565 ) | ( n6553 & n6786 ) | ( ~n6565 & n6786 ) ;
  assign n6788 = ~n3791 & n5966 ;
  assign n6789 = n1267 & n5969 ;
  assign n6790 = n1338 | n5970 ;
  assign n6791 = ~n1246 & n6464 ;
  assign n6792 = ( ~n1338 & n6790 ) | ( ~n1338 & n6791 ) | ( n6790 & n6791 ) ;
  assign n6793 = ( ~n6788 & n6789 ) | ( ~n6788 & n6792 ) | ( n6789 & n6792 ) ;
  assign n6794 = ( ~x14 & n6788 ) | ( ~x14 & n6793 ) | ( n6788 & n6793 ) ;
  assign n6795 = ( n6788 & n6793 ) | ( n6788 & ~n6794 ) | ( n6793 & ~n6794 ) ;
  assign n6796 = ( x14 & n6794 ) | ( x14 & ~n6795 ) | ( n6794 & ~n6795 ) ;
  assign n6797 = ( n6785 & n6787 ) | ( n6785 & n6796 ) | ( n6787 & n6796 ) ;
  assign n6798 = n3797 & n6584 ;
  assign n6799 = ~n3692 & n6587 ;
  assign n6800 = ~n3658 & n6588 ;
  assign n6801 = n6799 | n6800 ;
  assign n6802 = ( ~x11 & n6798 ) | ( ~x11 & n6801 ) | ( n6798 & n6801 ) ;
  assign n6803 = ( n6798 & n6801 ) | ( n6798 & ~n6802 ) | ( n6801 & ~n6802 ) ;
  assign n6804 = ( x11 & n6802 ) | ( x11 & ~n6803 ) | ( n6802 & ~n6803 ) ;
  assign n6805 = ( n6565 & ~n6567 ) | ( n6565 & n6576 ) | ( ~n6567 & n6576 ) ;
  assign n6806 = ( n6567 & ~n6577 ) | ( n6567 & n6805 ) | ( ~n6577 & n6805 ) ;
  assign n6807 = ( n6797 & n6804 ) | ( n6797 & n6806 ) | ( n6804 & n6806 ) ;
  assign n6808 = n4202 & n6061 ;
  assign n6809 = n3479 & n4345 ;
  assign n6810 = ~n3533 & n4200 ;
  assign n6811 = n3389 | n4201 ;
  assign n6812 = ( ~n3389 & n6810 ) | ( ~n3389 & n6811 ) | ( n6810 & n6811 ) ;
  assign n6813 = ( ~n6808 & n6809 ) | ( ~n6808 & n6812 ) | ( n6809 & n6812 ) ;
  assign n6814 = ( ~x26 & n6808 ) | ( ~x26 & n6813 ) | ( n6808 & n6813 ) ;
  assign n6815 = ( n6808 & n6813 ) | ( n6808 & ~n6814 ) | ( n6813 & ~n6814 ) ;
  assign n6816 = ( x26 & n6814 ) | ( x26 & ~n6815 ) | ( n6814 & ~n6815 ) ;
  assign n6817 = ( n3479 & n4202 ) | ( n3479 & n6009 ) | ( n4202 & n6009 ) ;
  assign n6818 = ~n3533 & n4345 ;
  assign n6819 = ~n3586 & n4200 ;
  assign n6820 = n6818 | n6819 ;
  assign n6821 = ~n3479 & n4201 ;
  assign n6822 = ( n4201 & n6820 ) | ( n4201 & ~n6821 ) | ( n6820 & ~n6821 ) ;
  assign n6823 = ( ~n6608 & n6817 ) | ( ~n6608 & n6822 ) | ( n6817 & n6822 ) ;
  assign n6824 = ~n3586 & n4195 ;
  assign n6825 = x26 & n6824 ;
  assign n6826 = ( n4202 & n6009 ) | ( n4202 & n6618 ) | ( n6009 & n6618 ) ;
  assign n6827 = ~n3533 & n4201 ;
  assign n6828 = ~n3586 & n4345 ;
  assign n6829 = n6827 | n6828 ;
  assign n6830 = n6826 | n6829 ;
  assign n6831 = ( x26 & n6825 ) | ( x26 & n6830 ) | ( n6825 & n6830 ) ;
  assign n6832 = n6823 | n6831 ;
  assign n6833 = x26 & ~n6832 ;
  assign n6834 = ( n6616 & n6816 ) | ( n6616 & n6833 ) | ( n6816 & n6833 ) ;
  assign n6835 = n4202 & ~n6104 ;
  assign n6836 = n3479 & n4200 ;
  assign n6837 = ~n3355 & n4201 ;
  assign n6838 = ~n3389 & n4345 ;
  assign n6839 = n6837 | n6838 ;
  assign n6840 = ( ~n6835 & n6836 ) | ( ~n6835 & n6839 ) | ( n6836 & n6839 ) ;
  assign n6841 = ( ~x26 & n6835 ) | ( ~x26 & n6840 ) | ( n6835 & n6840 ) ;
  assign n6842 = ( n6835 & n6840 ) | ( n6835 & ~n6841 ) | ( n6840 & ~n6841 ) ;
  assign n6843 = ( x26 & n6841 ) | ( x26 & ~n6842 ) | ( n6841 & ~n6842 ) ;
  assign n6844 = ( n6617 & n6619 ) | ( n6617 & n6622 ) | ( n6619 & n6622 ) ;
  assign n6845 = ~n6617 & n6623 ;
  assign n6846 = ( n6617 & ~n6844 ) | ( n6617 & n6845 ) | ( ~n6844 & n6845 ) ;
  assign n6847 = ( n6834 & n6843 ) | ( n6834 & n6846 ) | ( n6843 & n6846 ) ;
  assign n6848 = n4202 & ~n6154 ;
  assign n6849 = ~n3300 & n4201 ;
  assign n6850 = ~n3355 & n4345 ;
  assign n6851 = ~n3389 & n4200 ;
  assign n6852 = n6850 | n6851 ;
  assign n6853 = ( ~n6848 & n6849 ) | ( ~n6848 & n6852 ) | ( n6849 & n6852 ) ;
  assign n6854 = ( ~x26 & n6848 ) | ( ~x26 & n6853 ) | ( n6848 & n6853 ) ;
  assign n6855 = ( n6848 & n6853 ) | ( n6848 & ~n6854 ) | ( n6853 & ~n6854 ) ;
  assign n6856 = ( x26 & n6854 ) | ( x26 & ~n6855 ) | ( n6854 & ~n6855 ) ;
  assign n6857 = ( n6615 & n6624 ) | ( n6615 & ~n6625 ) | ( n6624 & ~n6625 ) ;
  assign n6858 = n6625 & ~n6857 ;
  assign n6859 = ( n6847 & n6856 ) | ( n6847 & n6858 ) | ( n6856 & n6858 ) ;
  assign n6860 = n4202 & n6200 ;
  assign n6861 = ~n3300 & n4345 ;
  assign n6862 = ~n3355 & n4200 ;
  assign n6863 = n3239 & ~n4201 ;
  assign n6864 = ( n3239 & n6862 ) | ( n3239 & ~n6863 ) | ( n6862 & ~n6863 ) ;
  assign n6865 = ( ~n6860 & n6861 ) | ( ~n6860 & n6864 ) | ( n6861 & n6864 ) ;
  assign n6866 = ( ~x26 & n6860 ) | ( ~x26 & n6865 ) | ( n6860 & n6865 ) ;
  assign n6867 = ( n6860 & n6865 ) | ( n6860 & ~n6866 ) | ( n6865 & ~n6866 ) ;
  assign n6868 = ( x26 & n6866 ) | ( x26 & ~n6867 ) | ( n6866 & ~n6867 ) ;
  assign n6869 = ( n6598 & n6607 ) | ( n6598 & ~n6626 ) | ( n6607 & ~n6626 ) ;
  assign n6870 = ( n6626 & ~n6627 ) | ( n6626 & n6869 ) | ( ~n6627 & n6869 ) ;
  assign n6871 = ( n6859 & n6868 ) | ( n6859 & n6870 ) | ( n6868 & n6870 ) ;
  assign n6872 = n4202 & ~n6243 ;
  assign n6873 = n3153 & n4201 ;
  assign n6874 = n3239 & n4345 ;
  assign n6875 = ~n3300 & n4200 ;
  assign n6876 = n6874 | n6875 ;
  assign n6877 = ( ~n6872 & n6873 ) | ( ~n6872 & n6876 ) | ( n6873 & n6876 ) ;
  assign n6878 = ( ~x26 & n6872 ) | ( ~x26 & n6877 ) | ( n6872 & n6877 ) ;
  assign n6879 = ( n6872 & n6877 ) | ( n6872 & ~n6878 ) | ( n6877 & ~n6878 ) ;
  assign n6880 = ( x26 & n6878 ) | ( x26 & ~n6879 ) | ( n6878 & ~n6879 ) ;
  assign n6881 = ( ~n6627 & n6631 ) | ( ~n6627 & n6640 ) | ( n6631 & n6640 ) ;
  assign n6882 = ( n6627 & ~n6641 ) | ( n6627 & n6881 ) | ( ~n6641 & n6881 ) ;
  assign n6883 = ( n6871 & n6880 ) | ( n6871 & n6882 ) | ( n6880 & n6882 ) ;
  assign n6884 = ( n6641 & ~n6650 ) | ( n6641 & n6652 ) | ( ~n6650 & n6652 ) ;
  assign n6885 = ( ~n6641 & n6653 ) | ( ~n6641 & n6884 ) | ( n6653 & n6884 ) ;
  assign n6886 = n4202 & n5710 ;
  assign n6887 = n3153 & n4345 ;
  assign n6888 = n3078 & n4201 ;
  assign n6889 = n3239 & n4200 ;
  assign n6890 = n6888 | n6889 ;
  assign n6891 = ( ~n6886 & n6887 ) | ( ~n6886 & n6890 ) | ( n6887 & n6890 ) ;
  assign n6892 = ( ~x26 & n6886 ) | ( ~x26 & n6891 ) | ( n6886 & n6891 ) ;
  assign n6893 = ( n6886 & n6891 ) | ( n6886 & ~n6892 ) | ( n6891 & ~n6892 ) ;
  assign n6894 = ( x26 & n6892 ) | ( x26 & ~n6893 ) | ( n6892 & ~n6893 ) ;
  assign n6895 = ( n6883 & ~n6885 ) | ( n6883 & n6894 ) | ( ~n6885 & n6894 ) ;
  assign n6896 = ( n6653 & ~n6662 ) | ( n6653 & n6664 ) | ( ~n6662 & n6664 ) ;
  assign n6897 = ( ~n6653 & n6665 ) | ( ~n6653 & n6896 ) | ( n6665 & n6896 ) ;
  assign n6898 = n4202 & ~n6267 ;
  assign n6899 = n3153 & n4200 ;
  assign n6900 = n3046 | n4201 ;
  assign n6901 = n3078 & n4345 ;
  assign n6902 = ( ~n3046 & n6900 ) | ( ~n3046 & n6901 ) | ( n6900 & n6901 ) ;
  assign n6903 = ( ~n6898 & n6899 ) | ( ~n6898 & n6902 ) | ( n6899 & n6902 ) ;
  assign n6904 = ( ~x26 & n6898 ) | ( ~x26 & n6903 ) | ( n6898 & n6903 ) ;
  assign n6905 = ( n6898 & n6903 ) | ( n6898 & ~n6904 ) | ( n6903 & ~n6904 ) ;
  assign n6906 = ( x26 & n6904 ) | ( x26 & ~n6905 ) | ( n6904 & ~n6905 ) ;
  assign n6907 = ( n6895 & ~n6897 ) | ( n6895 & n6906 ) | ( ~n6897 & n6906 ) ;
  assign n6908 = ( ~n6665 & n6674 ) | ( ~n6665 & n6676 ) | ( n6674 & n6676 ) ;
  assign n6909 = ( n6665 & ~n6677 ) | ( n6665 & n6908 ) | ( ~n6677 & n6908 ) ;
  assign n6910 = n4202 & n6279 ;
  assign n6911 = ~n2965 & n4201 ;
  assign n6912 = n3078 & n4200 ;
  assign n6913 = ~n3046 & n4345 ;
  assign n6914 = n6912 | n6913 ;
  assign n6915 = ( ~n6910 & n6911 ) | ( ~n6910 & n6914 ) | ( n6911 & n6914 ) ;
  assign n6916 = ( ~x26 & n6910 ) | ( ~x26 & n6915 ) | ( n6910 & n6915 ) ;
  assign n6917 = ( n6910 & n6915 ) | ( n6910 & ~n6916 ) | ( n6915 & ~n6916 ) ;
  assign n6918 = ( x26 & n6916 ) | ( x26 & ~n6917 ) | ( n6916 & ~n6917 ) ;
  assign n6919 = ( n6907 & n6909 ) | ( n6907 & n6918 ) | ( n6909 & n6918 ) ;
  assign n6920 = ( n6677 & ~n6686 ) | ( n6677 & n6688 ) | ( ~n6686 & n6688 ) ;
  assign n6921 = ( ~n6677 & n6689 ) | ( ~n6677 & n6920 ) | ( n6689 & n6920 ) ;
  assign n6922 = n4202 & ~n5768 ;
  assign n6923 = ~n2910 & n4201 ;
  assign n6924 = n3046 | n4200 ;
  assign n6925 = ~n2965 & n4345 ;
  assign n6926 = ( ~n3046 & n6924 ) | ( ~n3046 & n6925 ) | ( n6924 & n6925 ) ;
  assign n6927 = ( ~n6922 & n6923 ) | ( ~n6922 & n6926 ) | ( n6923 & n6926 ) ;
  assign n6928 = ( ~x26 & n6922 ) | ( ~x26 & n6927 ) | ( n6922 & n6927 ) ;
  assign n6929 = ( n6922 & n6927 ) | ( n6922 & ~n6928 ) | ( n6927 & ~n6928 ) ;
  assign n6930 = ( x26 & n6928 ) | ( x26 & ~n6929 ) | ( n6928 & ~n6929 ) ;
  assign n6931 = ( n6919 & ~n6921 ) | ( n6919 & n6930 ) | ( ~n6921 & n6930 ) ;
  assign n6932 = ( ~n6689 & n6698 ) | ( ~n6689 & n6700 ) | ( n6698 & n6700 ) ;
  assign n6933 = ( n6689 & ~n6701 ) | ( n6689 & n6932 ) | ( ~n6701 & n6932 ) ;
  assign n6934 = n4202 & n5543 ;
  assign n6935 = ~n2910 & n4345 ;
  assign n6936 = ~n2965 & n4200 ;
  assign n6937 = n2843 & ~n4201 ;
  assign n6938 = ( n2843 & n6936 ) | ( n2843 & ~n6937 ) | ( n6936 & ~n6937 ) ;
  assign n6939 = ( ~n6934 & n6935 ) | ( ~n6934 & n6938 ) | ( n6935 & n6938 ) ;
  assign n6940 = ( ~x26 & n6934 ) | ( ~x26 & n6939 ) | ( n6934 & n6939 ) ;
  assign n6941 = ( n6934 & n6939 ) | ( n6934 & ~n6940 ) | ( n6939 & ~n6940 ) ;
  assign n6942 = ( x26 & n6940 ) | ( x26 & ~n6941 ) | ( n6940 & ~n6941 ) ;
  assign n6943 = ( n6931 & n6933 ) | ( n6931 & n6942 ) | ( n6933 & n6942 ) ;
  assign n6944 = ( ~n6701 & n6710 ) | ( ~n6701 & n6712 ) | ( n6710 & n6712 ) ;
  assign n6945 = ( n6701 & ~n6713 ) | ( n6701 & n6944 ) | ( ~n6713 & n6944 ) ;
  assign n6946 = n4202 & n5791 ;
  assign n6947 = ~n2810 & n4201 ;
  assign n6948 = n2910 | n4200 ;
  assign n6949 = n2843 & n4345 ;
  assign n6950 = ( ~n2910 & n6948 ) | ( ~n2910 & n6949 ) | ( n6948 & n6949 ) ;
  assign n6951 = ( ~n6946 & n6947 ) | ( ~n6946 & n6950 ) | ( n6947 & n6950 ) ;
  assign n6952 = ( ~x26 & n6946 ) | ( ~x26 & n6951 ) | ( n6946 & n6951 ) ;
  assign n6953 = ( n6946 & n6951 ) | ( n6946 & ~n6952 ) | ( n6951 & ~n6952 ) ;
  assign n6954 = ( x26 & n6952 ) | ( x26 & ~n6953 ) | ( n6952 & ~n6953 ) ;
  assign n6955 = ( n6943 & n6945 ) | ( n6943 & n6954 ) | ( n6945 & n6954 ) ;
  assign n6956 = ( n6713 & ~n6715 ) | ( n6713 & n6724 ) | ( ~n6715 & n6724 ) ;
  assign n6957 = ( n6715 & ~n6725 ) | ( n6715 & n6956 ) | ( ~n6725 & n6956 ) ;
  assign n6958 = n4713 & ~n5270 ;
  assign n6959 = n2552 & n4792 ;
  assign n6960 = ~n2491 & n4712 ;
  assign n6961 = n2635 & n4709 ;
  assign n6962 = n6960 | n6961 ;
  assign n6963 = ( ~n6958 & n6959 ) | ( ~n6958 & n6962 ) | ( n6959 & n6962 ) ;
  assign n6964 = ( ~x23 & n6958 ) | ( ~x23 & n6963 ) | ( n6958 & n6963 ) ;
  assign n6965 = ( n6958 & n6963 ) | ( n6958 & ~n6964 ) | ( n6963 & ~n6964 ) ;
  assign n6966 = ( x23 & n6964 ) | ( x23 & ~n6965 ) | ( n6964 & ~n6965 ) ;
  assign n6967 = ( n6955 & n6957 ) | ( n6955 & n6966 ) | ( n6957 & n6966 ) ;
  assign n6968 = ( n6725 & ~n6727 ) | ( n6725 & n6736 ) | ( ~n6727 & n6736 ) ;
  assign n6969 = ( n6727 & ~n6737 ) | ( n6727 & n6968 ) | ( ~n6737 & n6968 ) ;
  assign n6970 = n4647 & n4974 ;
  assign n6971 = n2174 & n5398 ;
  assign n6972 = n2298 | n4973 ;
  assign n6973 = n2270 & n4972 ;
  assign n6974 = ( ~n2298 & n6972 ) | ( ~n2298 & n6973 ) | ( n6972 & n6973 ) ;
  assign n6975 = ( ~n6970 & n6971 ) | ( ~n6970 & n6974 ) | ( n6971 & n6974 ) ;
  assign n6976 = ( ~x20 & n6970 ) | ( ~x20 & n6975 ) | ( n6970 & n6975 ) ;
  assign n6977 = ( n6970 & n6975 ) | ( n6970 & ~n6976 ) | ( n6975 & ~n6976 ) ;
  assign n6978 = ( x20 & n6976 ) | ( x20 & ~n6977 ) | ( n6976 & ~n6977 ) ;
  assign n6979 = ( n6967 & n6969 ) | ( n6967 & n6978 ) | ( n6969 & n6978 ) ;
  assign n6980 = ( ~n6737 & n6739 ) | ( ~n6737 & n6748 ) | ( n6739 & n6748 ) ;
  assign n6981 = ( ~n6748 & n6749 ) | ( ~n6748 & n6980 ) | ( n6749 & n6980 ) ;
  assign n6982 = n4290 & n5508 ;
  assign n6983 = n1852 & n5507 ;
  assign n6984 = ~n2023 & n5504 ;
  assign n6985 = n1926 & n5666 ;
  assign n6986 = n6984 | n6985 ;
  assign n6987 = ( ~n6982 & n6983 ) | ( ~n6982 & n6986 ) | ( n6983 & n6986 ) ;
  assign n6988 = ( ~x17 & n6982 ) | ( ~x17 & n6987 ) | ( n6982 & n6987 ) ;
  assign n6989 = ( n6982 & n6987 ) | ( n6982 & ~n6988 ) | ( n6987 & ~n6988 ) ;
  assign n6990 = ( x17 & n6988 ) | ( x17 & ~n6989 ) | ( n6988 & ~n6989 ) ;
  assign n6991 = ( n6979 & ~n6981 ) | ( n6979 & n6990 ) | ( ~n6981 & n6990 ) ;
  assign n6992 = ~n4302 & n5508 ;
  assign n6993 = ~n1750 & n5507 ;
  assign n6994 = n1852 & n5666 ;
  assign n6995 = n1926 & n5504 ;
  assign n6996 = n6994 | n6995 ;
  assign n6997 = ( ~n6992 & n6993 ) | ( ~n6992 & n6996 ) | ( n6993 & n6996 ) ;
  assign n6998 = ( ~x17 & n6992 ) | ( ~x17 & n6997 ) | ( n6992 & n6997 ) ;
  assign n6999 = ( n6992 & n6997 ) | ( n6992 & ~n6998 ) | ( n6997 & ~n6998 ) ;
  assign n7000 = ( x17 & n6998 ) | ( x17 & ~n6999 ) | ( n6998 & ~n6999 ) ;
  assign n7001 = ( ~n6749 & n6751 ) | ( ~n6749 & n6760 ) | ( n6751 & n6760 ) ;
  assign n7002 = ( n6749 & ~n6761 ) | ( n6749 & n7001 ) | ( ~n6761 & n7001 ) ;
  assign n7003 = ( n6991 & n7000 ) | ( n6991 & n7002 ) | ( n7000 & n7002 ) ;
  assign n7004 = ( ~n6761 & n6763 ) | ( ~n6761 & n6772 ) | ( n6763 & n6772 ) ;
  assign n7005 = ( ~n6772 & n6773 ) | ( ~n6772 & n7004 ) | ( n6773 & n7004 ) ;
  assign n7006 = ~n3955 & n5966 ;
  assign n7007 = ~n1338 & n6464 ;
  assign n7008 = n1458 & n5969 ;
  assign n7009 = n1576 & n5970 ;
  assign n7010 = n7008 | n7009 ;
  assign n7011 = ( ~n7006 & n7007 ) | ( ~n7006 & n7010 ) | ( n7007 & n7010 ) ;
  assign n7012 = ( ~x14 & n7006 ) | ( ~x14 & n7011 ) | ( n7006 & n7011 ) ;
  assign n7013 = ( n7006 & n7011 ) | ( n7006 & ~n7012 ) | ( n7011 & ~n7012 ) ;
  assign n7014 = ( x14 & n7012 ) | ( x14 & ~n7013 ) | ( n7012 & ~n7013 ) ;
  assign n7015 = ( n7003 & ~n7005 ) | ( n7003 & n7014 ) | ( ~n7005 & n7014 ) ;
  assign n7016 = ( ~n6773 & n6775 ) | ( ~n6773 & n6784 ) | ( n6775 & n6784 ) ;
  assign n7017 = ( n6773 & ~n6785 ) | ( n6773 & n7016 ) | ( ~n6785 & n7016 ) ;
  assign n7018 = ~n3665 & n6584 ;
  assign n7019 = ~n1290 & n6587 ;
  assign n7020 = ~n1246 & n6588 ;
  assign n7021 = ~n6581 & n6582 ;
  assign n7022 = ( ~n6578 & n6579 ) | ( ~n6578 & n7021 ) | ( n6579 & n7021 ) ;
  assign n7023 = ~n3658 & n7022 ;
  assign n7024 = n7020 | n7023 ;
  assign n7025 = ( ~n7018 & n7019 ) | ( ~n7018 & n7024 ) | ( n7019 & n7024 ) ;
  assign n7026 = ( ~x11 & n7018 ) | ( ~x11 & n7025 ) | ( n7018 & n7025 ) ;
  assign n7027 = ( n7018 & n7025 ) | ( n7018 & ~n7026 ) | ( n7025 & ~n7026 ) ;
  assign n7028 = ( x11 & n7026 ) | ( x11 & ~n7027 ) | ( n7026 & ~n7027 ) ;
  assign n7029 = ( n7015 & n7017 ) | ( n7015 & n7028 ) | ( n7017 & n7028 ) ;
  assign n7030 = n3692 & n7022 ;
  assign n7031 = ~n3658 & n6587 ;
  assign n7032 = ( n7022 & ~n7030 ) | ( n7022 & n7031 ) | ( ~n7030 & n7031 ) ;
  assign n7033 = ~n1290 & n6588 ;
  assign n7034 = n7032 | n7033 ;
  assign n7035 = ~n4182 & n6584 ;
  assign n7036 = ( x11 & n7034 ) | ( x11 & ~n7035 ) | ( n7034 & ~n7035 ) ;
  assign n7037 = ( ~x11 & n7034 ) | ( ~x11 & n7035 ) | ( n7034 & n7035 ) ;
  assign n7038 = ( ~n7034 & n7036 ) | ( ~n7034 & n7037 ) | ( n7036 & n7037 ) ;
  assign n7039 = ( ~n6785 & n6787 ) | ( ~n6785 & n6796 ) | ( n6787 & n6796 ) ;
  assign n7040 = ( n6785 & ~n6797 ) | ( n6785 & n7039 ) | ( ~n6797 & n7039 ) ;
  assign n7041 = ( n7029 & n7038 ) | ( n7029 & n7040 ) | ( n7038 & n7040 ) ;
  assign n7042 = n4713 & n6061 ;
  assign n7043 = n3479 & n4792 ;
  assign n7044 = n3533 | n4709 ;
  assign n7045 = ~n3389 & n4712 ;
  assign n7046 = ( ~n3533 & n7044 ) | ( ~n3533 & n7045 ) | ( n7044 & n7045 ) ;
  assign n7047 = ( ~n7042 & n7043 ) | ( ~n7042 & n7046 ) | ( n7043 & n7046 ) ;
  assign n7048 = ( ~x23 & n7042 ) | ( ~x23 & n7047 ) | ( n7042 & n7047 ) ;
  assign n7049 = ( n7042 & n7047 ) | ( n7042 & ~n7048 ) | ( n7047 & ~n7048 ) ;
  assign n7050 = ( x23 & n7048 ) | ( x23 & ~n7049 ) | ( n7048 & ~n7049 ) ;
  assign n7051 = ( n3479 & n4713 ) | ( n3479 & n6009 ) | ( n4713 & n6009 ) ;
  assign n7052 = ~n3533 & n4792 ;
  assign n7053 = ~n3586 & n4709 ;
  assign n7054 = n7052 | n7053 ;
  assign n7055 = ~n3479 & n4712 ;
  assign n7056 = ( n4712 & n7054 ) | ( n4712 & ~n7055 ) | ( n7054 & ~n7055 ) ;
  assign n7057 = ( ~n6608 & n7051 ) | ( ~n6608 & n7056 ) | ( n7051 & n7056 ) ;
  assign n7058 = ~n3586 & n4711 ;
  assign n7059 = x23 & n7058 ;
  assign n7060 = ( n4713 & n6009 ) | ( n4713 & n6618 ) | ( n6009 & n6618 ) ;
  assign n7061 = ~n3533 & n4712 ;
  assign n7062 = n3586 | n4792 ;
  assign n7063 = ( ~n3586 & n7061 ) | ( ~n3586 & n7062 ) | ( n7061 & n7062 ) ;
  assign n7064 = n7060 | n7063 ;
  assign n7065 = ( x23 & n7059 ) | ( x23 & n7064 ) | ( n7059 & n7064 ) ;
  assign n7066 = n7057 | n7065 ;
  assign n7067 = x23 & ~n7066 ;
  assign n7068 = ( n6824 & n7050 ) | ( n6824 & n7067 ) | ( n7050 & n7067 ) ;
  assign n7069 = ~n3355 & n4712 ;
  assign n7070 = n3389 | n4792 ;
  assign n7071 = ( ~n3389 & n7069 ) | ( ~n3389 & n7070 ) | ( n7069 & n7070 ) ;
  assign n7072 = ~n3479 & n4709 ;
  assign n7073 = ( n4709 & n7071 ) | ( n4709 & ~n7072 ) | ( n7071 & ~n7072 ) ;
  assign n7074 = ( n4713 & ~n6104 ) | ( n4713 & n7073 ) | ( ~n6104 & n7073 ) ;
  assign n7075 = n7073 & ~n7074 ;
  assign n7076 = ( ~x23 & n7074 ) | ( ~x23 & n7075 ) | ( n7074 & n7075 ) ;
  assign n7077 = ( n7074 & n7075 ) | ( n7074 & ~n7076 ) | ( n7075 & ~n7076 ) ;
  assign n7078 = ( x23 & n7076 ) | ( x23 & ~n7077 ) | ( n7076 & ~n7077 ) ;
  assign n7079 = ( n6825 & n6826 ) | ( n6825 & n6829 ) | ( n6826 & n6829 ) ;
  assign n7080 = ~n6825 & n6830 ;
  assign n7081 = ( n6825 & ~n7079 ) | ( n6825 & n7080 ) | ( ~n7079 & n7080 ) ;
  assign n7082 = ( n7068 & n7078 ) | ( n7068 & n7081 ) | ( n7078 & n7081 ) ;
  assign n7083 = n4713 & ~n6154 ;
  assign n7084 = ~n3300 & n4712 ;
  assign n7085 = ~n3355 & n4792 ;
  assign n7086 = ~n3389 & n4709 ;
  assign n7087 = n7085 | n7086 ;
  assign n7088 = ( ~n7083 & n7084 ) | ( ~n7083 & n7087 ) | ( n7084 & n7087 ) ;
  assign n7089 = ( ~x23 & n7083 ) | ( ~x23 & n7088 ) | ( n7083 & n7088 ) ;
  assign n7090 = ( n7083 & n7088 ) | ( n7083 & ~n7089 ) | ( n7088 & ~n7089 ) ;
  assign n7091 = ( x23 & n7089 ) | ( x23 & ~n7090 ) | ( n7089 & ~n7090 ) ;
  assign n7092 = ( n6823 & n6831 ) | ( n6823 & ~n6832 ) | ( n6831 & ~n6832 ) ;
  assign n7093 = n6832 & ~n7092 ;
  assign n7094 = ( n7082 & n7091 ) | ( n7082 & n7093 ) | ( n7091 & n7093 ) ;
  assign n7095 = n4713 & n6200 ;
  assign n7096 = ~n3300 & n4792 ;
  assign n7097 = n3355 | n4709 ;
  assign n7098 = n3239 & n4712 ;
  assign n7099 = ( ~n3355 & n7097 ) | ( ~n3355 & n7098 ) | ( n7097 & n7098 ) ;
  assign n7100 = ( ~n7095 & n7096 ) | ( ~n7095 & n7099 ) | ( n7096 & n7099 ) ;
  assign n7101 = ( ~x23 & n7095 ) | ( ~x23 & n7100 ) | ( n7095 & n7100 ) ;
  assign n7102 = ( n7095 & n7100 ) | ( n7095 & ~n7101 ) | ( n7100 & ~n7101 ) ;
  assign n7103 = ( x23 & n7101 ) | ( x23 & ~n7102 ) | ( n7101 & ~n7102 ) ;
  assign n7104 = ( n6616 & n6816 ) | ( n6616 & ~n6833 ) | ( n6816 & ~n6833 ) ;
  assign n7105 = ( n6833 & ~n6834 ) | ( n6833 & n7104 ) | ( ~n6834 & n7104 ) ;
  assign n7106 = ( n7094 & n7103 ) | ( n7094 & n7105 ) | ( n7103 & n7105 ) ;
  assign n7107 = n4713 & ~n6243 ;
  assign n7108 = n3153 & n4712 ;
  assign n7109 = n3239 & n4792 ;
  assign n7110 = ~n3300 & n4709 ;
  assign n7111 = n7109 | n7110 ;
  assign n7112 = ( ~n7107 & n7108 ) | ( ~n7107 & n7111 ) | ( n7108 & n7111 ) ;
  assign n7113 = ( ~x23 & n7107 ) | ( ~x23 & n7112 ) | ( n7107 & n7112 ) ;
  assign n7114 = ( n7107 & n7112 ) | ( n7107 & ~n7113 ) | ( n7112 & ~n7113 ) ;
  assign n7115 = ( x23 & n7113 ) | ( x23 & ~n7114 ) | ( n7113 & ~n7114 ) ;
  assign n7116 = ( ~n6834 & n6843 ) | ( ~n6834 & n6846 ) | ( n6843 & n6846 ) ;
  assign n7117 = ( n6834 & ~n6847 ) | ( n6834 & n7116 ) | ( ~n6847 & n7116 ) ;
  assign n7118 = ( n7106 & n7115 ) | ( n7106 & n7117 ) | ( n7115 & n7117 ) ;
  assign n7119 = ( ~n6847 & n6856 ) | ( ~n6847 & n6858 ) | ( n6856 & n6858 ) ;
  assign n7120 = ( n6847 & ~n6859 ) | ( n6847 & n7119 ) | ( ~n6859 & n7119 ) ;
  assign n7121 = n4713 & n5710 ;
  assign n7122 = n3153 & n4792 ;
  assign n7123 = n3078 & n4712 ;
  assign n7124 = n3239 & n4709 ;
  assign n7125 = n7123 | n7124 ;
  assign n7126 = ( ~n7121 & n7122 ) | ( ~n7121 & n7125 ) | ( n7122 & n7125 ) ;
  assign n7127 = ( ~x23 & n7121 ) | ( ~x23 & n7126 ) | ( n7121 & n7126 ) ;
  assign n7128 = ( n7121 & n7126 ) | ( n7121 & ~n7127 ) | ( n7126 & ~n7127 ) ;
  assign n7129 = ( x23 & n7127 ) | ( x23 & ~n7128 ) | ( n7127 & ~n7128 ) ;
  assign n7130 = ( n7118 & n7120 ) | ( n7118 & n7129 ) | ( n7120 & n7129 ) ;
  assign n7131 = ( ~n6859 & n6868 ) | ( ~n6859 & n6870 ) | ( n6868 & n6870 ) ;
  assign n7132 = ( n6859 & ~n6871 ) | ( n6859 & n7131 ) | ( ~n6871 & n7131 ) ;
  assign n7133 = n3078 & ~n4792 ;
  assign n7134 = ~n3046 & n4712 ;
  assign n7135 = ( n3078 & ~n7133 ) | ( n3078 & n7134 ) | ( ~n7133 & n7134 ) ;
  assign n7136 = ~n3153 & n4709 ;
  assign n7137 = ( n4709 & n7135 ) | ( n4709 & ~n7136 ) | ( n7135 & ~n7136 ) ;
  assign n7138 = ( n4713 & ~n6267 ) | ( n4713 & n7137 ) | ( ~n6267 & n7137 ) ;
  assign n7139 = n7137 & ~n7138 ;
  assign n7140 = ( ~x23 & n7138 ) | ( ~x23 & n7139 ) | ( n7138 & n7139 ) ;
  assign n7141 = ( n7138 & n7139 ) | ( n7138 & ~n7140 ) | ( n7139 & ~n7140 ) ;
  assign n7142 = ( x23 & n7140 ) | ( x23 & ~n7141 ) | ( n7140 & ~n7141 ) ;
  assign n7143 = ( n7130 & n7132 ) | ( n7130 & n7142 ) | ( n7132 & n7142 ) ;
  assign n7144 = n4713 & n6279 ;
  assign n7145 = ~n2965 & n4712 ;
  assign n7146 = n3078 & n4709 ;
  assign n7147 = ~n3046 & n4792 ;
  assign n7148 = n7146 | n7147 ;
  assign n7149 = ( ~n7144 & n7145 ) | ( ~n7144 & n7148 ) | ( n7145 & n7148 ) ;
  assign n7150 = ( ~x23 & n7144 ) | ( ~x23 & n7149 ) | ( n7144 & n7149 ) ;
  assign n7151 = ( n7144 & n7149 ) | ( n7144 & ~n7150 ) | ( n7149 & ~n7150 ) ;
  assign n7152 = ( x23 & n7150 ) | ( x23 & ~n7151 ) | ( n7150 & ~n7151 ) ;
  assign n7153 = ( ~n6871 & n6880 ) | ( ~n6871 & n6882 ) | ( n6880 & n6882 ) ;
  assign n7154 = ( n6871 & ~n6883 ) | ( n6871 & n7153 ) | ( ~n6883 & n7153 ) ;
  assign n7155 = ( n7143 & n7152 ) | ( n7143 & n7154 ) | ( n7152 & n7154 ) ;
  assign n7156 = n4713 & ~n5768 ;
  assign n7157 = ~n2910 & n4712 ;
  assign n7158 = n3046 | n4709 ;
  assign n7159 = ~n2965 & n4792 ;
  assign n7160 = ( ~n3046 & n7158 ) | ( ~n3046 & n7159 ) | ( n7158 & n7159 ) ;
  assign n7161 = ( ~n7156 & n7157 ) | ( ~n7156 & n7160 ) | ( n7157 & n7160 ) ;
  assign n7162 = ( ~x23 & n7156 ) | ( ~x23 & n7161 ) | ( n7156 & n7161 ) ;
  assign n7163 = ( n7156 & n7161 ) | ( n7156 & ~n7162 ) | ( n7161 & ~n7162 ) ;
  assign n7164 = ( x23 & n7162 ) | ( x23 & ~n7163 ) | ( n7162 & ~n7163 ) ;
  assign n7165 = ( ~n6883 & n6885 ) | ( ~n6883 & n6894 ) | ( n6885 & n6894 ) ;
  assign n7166 = ( ~n6894 & n6895 ) | ( ~n6894 & n7165 ) | ( n6895 & n7165 ) ;
  assign n7167 = ( n7155 & n7164 ) | ( n7155 & ~n7166 ) | ( n7164 & ~n7166 ) ;
  assign n7168 = n4713 & n5543 ;
  assign n7169 = ~n2910 & n4792 ;
  assign n7170 = n2965 | n4709 ;
  assign n7171 = n2843 & n4712 ;
  assign n7172 = ( ~n2965 & n7170 ) | ( ~n2965 & n7171 ) | ( n7170 & n7171 ) ;
  assign n7173 = ( ~n7168 & n7169 ) | ( ~n7168 & n7172 ) | ( n7169 & n7172 ) ;
  assign n7174 = ( ~x23 & n7168 ) | ( ~x23 & n7173 ) | ( n7168 & n7173 ) ;
  assign n7175 = ( n7168 & n7173 ) | ( n7168 & ~n7174 ) | ( n7173 & ~n7174 ) ;
  assign n7176 = ( x23 & n7174 ) | ( x23 & ~n7175 ) | ( n7174 & ~n7175 ) ;
  assign n7177 = ( ~n6895 & n6897 ) | ( ~n6895 & n6906 ) | ( n6897 & n6906 ) ;
  assign n7178 = ( ~n6906 & n6907 ) | ( ~n6906 & n7177 ) | ( n6907 & n7177 ) ;
  assign n7179 = ( n7167 & n7176 ) | ( n7167 & ~n7178 ) | ( n7176 & ~n7178 ) ;
  assign n7180 = n4713 & n5791 ;
  assign n7181 = ~n2810 & n4712 ;
  assign n7182 = n2910 | n4709 ;
  assign n7183 = n2843 & n4792 ;
  assign n7184 = ( ~n2910 & n7182 ) | ( ~n2910 & n7183 ) | ( n7182 & n7183 ) ;
  assign n7185 = ( ~n7180 & n7181 ) | ( ~n7180 & n7184 ) | ( n7181 & n7184 ) ;
  assign n7186 = ( ~x23 & n7180 ) | ( ~x23 & n7185 ) | ( n7180 & n7185 ) ;
  assign n7187 = ( n7180 & n7185 ) | ( n7180 & ~n7186 ) | ( n7185 & ~n7186 ) ;
  assign n7188 = ( x23 & n7186 ) | ( x23 & ~n7187 ) | ( n7186 & ~n7187 ) ;
  assign n7189 = ( ~n6907 & n6909 ) | ( ~n6907 & n6918 ) | ( n6909 & n6918 ) ;
  assign n7190 = ( n6907 & ~n6919 ) | ( n6907 & n7189 ) | ( ~n6919 & n7189 ) ;
  assign n7191 = ( n7179 & n7188 ) | ( n7179 & n7190 ) | ( n7188 & n7190 ) ;
  assign n7192 = n4713 & ~n5586 ;
  assign n7193 = ~n2725 & n4712 ;
  assign n7194 = n2843 & n4709 ;
  assign n7195 = ~n2810 & n4792 ;
  assign n7196 = n7194 | n7195 ;
  assign n7197 = ( ~n7192 & n7193 ) | ( ~n7192 & n7196 ) | ( n7193 & n7196 ) ;
  assign n7198 = ( ~x23 & n7192 ) | ( ~x23 & n7197 ) | ( n7192 & n7197 ) ;
  assign n7199 = ( n7192 & n7197 ) | ( n7192 & ~n7198 ) | ( n7197 & ~n7198 ) ;
  assign n7200 = ( x23 & n7198 ) | ( x23 & ~n7199 ) | ( n7198 & ~n7199 ) ;
  assign n7201 = ( ~n6919 & n6921 ) | ( ~n6919 & n6930 ) | ( n6921 & n6930 ) ;
  assign n7202 = ( ~n6930 & n6931 ) | ( ~n6930 & n7201 ) | ( n6931 & n7201 ) ;
  assign n7203 = ( n7191 & n7200 ) | ( n7191 & ~n7202 ) | ( n7200 & ~n7202 ) ;
  assign n7204 = n2725 | n4792 ;
  assign n7205 = n2635 & n4712 ;
  assign n7206 = ( ~n2725 & n7204 ) | ( ~n2725 & n7205 ) | ( n7204 & n7205 ) ;
  assign n7207 = n2810 & n4709 ;
  assign n7208 = ( n4709 & n7206 ) | ( n4709 & ~n7207 ) | ( n7206 & ~n7207 ) ;
  assign n7209 = ( n4711 & n4712 ) | ( n4711 & n5232 ) | ( n4712 & n5232 ) ;
  assign n7210 = ( ~n4712 & n7208 ) | ( ~n4712 & n7209 ) | ( n7208 & n7209 ) ;
  assign n7211 = x23 | n7210 ;
  assign n7212 = ( x23 & n7210 ) | ( x23 & ~n7211 ) | ( n7210 & ~n7211 ) ;
  assign n7213 = n7211 & ~n7212 ;
  assign n7214 = ( ~n6931 & n6933 ) | ( ~n6931 & n6942 ) | ( n6933 & n6942 ) ;
  assign n7215 = ( n6931 & ~n6943 ) | ( n6931 & n7214 ) | ( ~n6943 & n7214 ) ;
  assign n7216 = ( n7203 & n7213 ) | ( n7203 & n7215 ) | ( n7213 & n7215 ) ;
  assign n7217 = n4713 & ~n5425 ;
  assign n7218 = n2552 & n4712 ;
  assign n7219 = ~n2725 & n4709 ;
  assign n7220 = n2635 & n4792 ;
  assign n7221 = n7219 | n7220 ;
  assign n7222 = ( ~n7217 & n7218 ) | ( ~n7217 & n7221 ) | ( n7218 & n7221 ) ;
  assign n7223 = ( ~x23 & n7217 ) | ( ~x23 & n7222 ) | ( n7217 & n7222 ) ;
  assign n7224 = ( n7217 & n7222 ) | ( n7217 & ~n7223 ) | ( n7222 & ~n7223 ) ;
  assign n7225 = ( x23 & n7223 ) | ( x23 & ~n7224 ) | ( n7223 & ~n7224 ) ;
  assign n7226 = ( ~n6943 & n6945 ) | ( ~n6943 & n6954 ) | ( n6945 & n6954 ) ;
  assign n7227 = ( n6943 & ~n6955 ) | ( n6943 & n7226 ) | ( ~n6955 & n7226 ) ;
  assign n7228 = ( n7216 & n7225 ) | ( n7216 & n7227 ) | ( n7225 & n7227 ) ;
  assign n7229 = ( n6955 & ~n6957 ) | ( n6955 & n6966 ) | ( ~n6957 & n6966 ) ;
  assign n7230 = ( n6957 & ~n6967 ) | ( n6957 & n7229 ) | ( ~n6967 & n7229 ) ;
  assign n7231 = n2298 | n4972 ;
  assign n7232 = n2270 & n5398 ;
  assign n7233 = ( ~n2298 & n7231 ) | ( ~n2298 & n7232 ) | ( n7231 & n7232 ) ;
  assign n7234 = n2396 & ~n4973 ;
  assign n7235 = ( n2396 & n7233 ) | ( n2396 & ~n7234 ) | ( n7233 & ~n7234 ) ;
  assign n7236 = ( ~n4912 & n4974 ) | ( ~n4912 & n7235 ) | ( n4974 & n7235 ) ;
  assign n7237 = n7235 & ~n7236 ;
  assign n7238 = ( ~x20 & n7236 ) | ( ~x20 & n7237 ) | ( n7236 & n7237 ) ;
  assign n7239 = ( n7236 & n7237 ) | ( n7236 & ~n7238 ) | ( n7237 & ~n7238 ) ;
  assign n7240 = ( x20 & n7238 ) | ( x20 & ~n7239 ) | ( n7238 & ~n7239 ) ;
  assign n7241 = ( n7228 & n7230 ) | ( n7228 & n7240 ) | ( n7230 & n7240 ) ;
  assign n7242 = ( n6967 & ~n6969 ) | ( n6967 & n6978 ) | ( ~n6969 & n6978 ) ;
  assign n7243 = ( n6969 & ~n6979 ) | ( n6969 & n7242 ) | ( ~n6979 & n7242 ) ;
  assign n7244 = ~n4457 & n5508 ;
  assign n7245 = n1926 & n5507 ;
  assign n7246 = ~n2023 & n5666 ;
  assign n7247 = n2089 & n5504 ;
  assign n7248 = n7246 | n7247 ;
  assign n7249 = ( ~n7244 & n7245 ) | ( ~n7244 & n7248 ) | ( n7245 & n7248 ) ;
  assign n7250 = ( ~x17 & n7244 ) | ( ~x17 & n7249 ) | ( n7244 & n7249 ) ;
  assign n7251 = ( n7244 & n7249 ) | ( n7244 & ~n7250 ) | ( n7249 & ~n7250 ) ;
  assign n7252 = ( x17 & n7250 ) | ( x17 & ~n7251 ) | ( n7250 & ~n7251 ) ;
  assign n7253 = ( n7241 & n7243 ) | ( n7241 & n7252 ) | ( n7243 & n7252 ) ;
  assign n7254 = ( ~n6979 & n6981 ) | ( ~n6979 & n6990 ) | ( n6981 & n6990 ) ;
  assign n7255 = ( ~n6990 & n6991 ) | ( ~n6990 & n7254 ) | ( n6991 & n7254 ) ;
  assign n7256 = n4326 & n5966 ;
  assign n7257 = n1576 & n6464 ;
  assign n7258 = n1750 | n5970 ;
  assign n7259 = ~n1669 & n5969 ;
  assign n7260 = ( ~n1750 & n7258 ) | ( ~n1750 & n7259 ) | ( n7258 & n7259 ) ;
  assign n7261 = ( ~n7256 & n7257 ) | ( ~n7256 & n7260 ) | ( n7257 & n7260 ) ;
  assign n7262 = ( ~x14 & n7256 ) | ( ~x14 & n7261 ) | ( n7256 & n7261 ) ;
  assign n7263 = ( n7256 & n7261 ) | ( n7256 & ~n7262 ) | ( n7261 & ~n7262 ) ;
  assign n7264 = ( x14 & n7262 ) | ( x14 & ~n7263 ) | ( n7262 & ~n7263 ) ;
  assign n7265 = ( n7253 & ~n7255 ) | ( n7253 & n7264 ) | ( ~n7255 & n7264 ) ;
  assign n7266 = ( ~n6991 & n7000 ) | ( ~n6991 & n7002 ) | ( n7000 & n7002 ) ;
  assign n7267 = ( n6991 & ~n7003 ) | ( n6991 & n7266 ) | ( ~n7003 & n7266 ) ;
  assign n7268 = ~n4159 & n5966 ;
  assign n7269 = n1458 & n6464 ;
  assign n7270 = n1669 | n5970 ;
  assign n7271 = n1576 & n5969 ;
  assign n7272 = ( ~n1669 & n7270 ) | ( ~n1669 & n7271 ) | ( n7270 & n7271 ) ;
  assign n7273 = ( ~n7268 & n7269 ) | ( ~n7268 & n7272 ) | ( n7269 & n7272 ) ;
  assign n7274 = ( ~x14 & n7268 ) | ( ~x14 & n7273 ) | ( n7268 & n7273 ) ;
  assign n7275 = ( n7268 & n7273 ) | ( n7268 & ~n7274 ) | ( n7273 & ~n7274 ) ;
  assign n7276 = ( x14 & n7274 ) | ( x14 & ~n7275 ) | ( n7274 & ~n7275 ) ;
  assign n7277 = ( n7265 & n7267 ) | ( n7265 & n7276 ) | ( n7267 & n7276 ) ;
  assign n7278 = ( ~n7003 & n7005 ) | ( ~n7003 & n7014 ) | ( n7005 & n7014 ) ;
  assign n7279 = ( ~n7014 & n7015 ) | ( ~n7014 & n7278 ) | ( n7015 & n7278 ) ;
  assign n7280 = n3621 & n6584 ;
  assign n7281 = ~n1290 & n7022 ;
  assign n7282 = n1267 & ~n6588 ;
  assign n7283 = ~n1246 & n6587 ;
  assign n7284 = ( n1267 & ~n7282 ) | ( n1267 & n7283 ) | ( ~n7282 & n7283 ) ;
  assign n7285 = ( ~n7280 & n7281 ) | ( ~n7280 & n7284 ) | ( n7281 & n7284 ) ;
  assign n7286 = ( ~x11 & n7280 ) | ( ~x11 & n7285 ) | ( n7280 & n7285 ) ;
  assign n7287 = ( n7280 & n7285 ) | ( n7280 & ~n7286 ) | ( n7285 & ~n7286 ) ;
  assign n7288 = ( x11 & n7286 ) | ( x11 & ~n7287 ) | ( n7286 & ~n7287 ) ;
  assign n7289 = ( n7277 & ~n7279 ) | ( n7277 & n7288 ) | ( ~n7279 & n7288 ) ;
  assign n7290 = x7 | x8 ;
  assign n7291 = x7 & x8 ;
  assign n7292 = n7290 & ~n7291 ;
  assign n7293 = x5 & x6 ;
  assign n7294 = x5 | x6 ;
  assign n7295 = ( n7292 & n7293 ) | ( n7292 & ~n7294 ) | ( n7293 & ~n7294 ) ;
  assign n7296 = n7292 & ~n7295 ;
  assign n7297 = x6 | x7 ;
  assign n7298 = x5 & ~x7 ;
  assign n7299 = ( ~n7294 & n7297 ) | ( ~n7294 & n7298 ) | ( n7297 & n7298 ) ;
  assign n7300 = n7295 & ~n7299 ;
  assign n7301 = ~n3692 & n7300 ;
  assign n7302 = ( n3691 & n3692 ) | ( n3691 & n7296 ) | ( n3692 & n7296 ) ;
  assign n7303 = ( n7296 & n7301 ) | ( n7296 & ~n7302 ) | ( n7301 & ~n7302 ) ;
  assign n7304 = x8 | n7303 ;
  assign n7305 = ( x8 & n7303 ) | ( x8 & ~n7304 ) | ( n7303 & ~n7304 ) ;
  assign n7306 = n7304 & ~n7305 ;
  assign n7307 = ( n7015 & ~n7017 ) | ( n7015 & n7028 ) | ( ~n7017 & n7028 ) ;
  assign n7308 = ( n7017 & ~n7029 ) | ( n7017 & n7307 ) | ( ~n7029 & n7307 ) ;
  assign n7309 = ( n7289 & n7306 ) | ( n7289 & n7308 ) | ( n7306 & n7308 ) ;
  assign n7310 = n4974 & n6061 ;
  assign n7311 = n3479 & n4972 ;
  assign n7312 = n3533 | n4973 ;
  assign n7313 = ~n3389 & n5398 ;
  assign n7314 = ( ~n3533 & n7312 ) | ( ~n3533 & n7313 ) | ( n7312 & n7313 ) ;
  assign n7315 = ( ~n7310 & n7311 ) | ( ~n7310 & n7314 ) | ( n7311 & n7314 ) ;
  assign n7316 = ( ~x20 & n7310 ) | ( ~x20 & n7315 ) | ( n7310 & n7315 ) ;
  assign n7317 = ( n7310 & n7315 ) | ( n7310 & ~n7316 ) | ( n7315 & ~n7316 ) ;
  assign n7318 = ( x20 & n7316 ) | ( x20 & ~n7317 ) | ( n7316 & ~n7317 ) ;
  assign n7319 = ( n3479 & n4974 ) | ( n3479 & n6009 ) | ( n4974 & n6009 ) ;
  assign n7320 = ~n3533 & n4972 ;
  assign n7321 = ~n3586 & n4973 ;
  assign n7322 = n7320 | n7321 ;
  assign n7323 = ~n3479 & n5398 ;
  assign n7324 = ( n5398 & n7322 ) | ( n5398 & ~n7323 ) | ( n7322 & ~n7323 ) ;
  assign n7325 = ( ~n6608 & n7319 ) | ( ~n6608 & n7324 ) | ( n7319 & n7324 ) ;
  assign n7326 = ~n3586 & n5397 ;
  assign n7327 = x20 & n7326 ;
  assign n7328 = ( n4974 & n6009 ) | ( n4974 & n6618 ) | ( n6009 & n6618 ) ;
  assign n7329 = ~n3533 & n5398 ;
  assign n7330 = n3586 | n4972 ;
  assign n7331 = ( ~n3586 & n7329 ) | ( ~n3586 & n7330 ) | ( n7329 & n7330 ) ;
  assign n7332 = n7328 | n7331 ;
  assign n7333 = ( x20 & n7327 ) | ( x20 & n7332 ) | ( n7327 & n7332 ) ;
  assign n7334 = n7325 | n7333 ;
  assign n7335 = x20 & ~n7334 ;
  assign n7336 = ( n7058 & n7318 ) | ( n7058 & n7335 ) | ( n7318 & n7335 ) ;
  assign n7337 = n3389 | n4972 ;
  assign n7338 = ~n3355 & n5398 ;
  assign n7339 = ( ~n3389 & n7337 ) | ( ~n3389 & n7338 ) | ( n7337 & n7338 ) ;
  assign n7340 = n3479 & ~n4973 ;
  assign n7341 = ( n3479 & n7339 ) | ( n3479 & ~n7340 ) | ( n7339 & ~n7340 ) ;
  assign n7342 = ( n4974 & ~n6104 ) | ( n4974 & n7341 ) | ( ~n6104 & n7341 ) ;
  assign n7343 = n7341 & ~n7342 ;
  assign n7344 = ( ~x20 & n7342 ) | ( ~x20 & n7343 ) | ( n7342 & n7343 ) ;
  assign n7345 = ( n7342 & n7343 ) | ( n7342 & ~n7344 ) | ( n7343 & ~n7344 ) ;
  assign n7346 = ( x20 & n7344 ) | ( x20 & ~n7345 ) | ( n7344 & ~n7345 ) ;
  assign n7347 = ( n7059 & n7060 ) | ( n7059 & n7063 ) | ( n7060 & n7063 ) ;
  assign n7348 = ~n7059 & n7064 ;
  assign n7349 = ( n7059 & ~n7347 ) | ( n7059 & n7348 ) | ( ~n7347 & n7348 ) ;
  assign n7350 = ( n7336 & n7346 ) | ( n7336 & n7349 ) | ( n7346 & n7349 ) ;
  assign n7351 = n4974 & ~n6154 ;
  assign n7352 = ~n3300 & n5398 ;
  assign n7353 = n3389 | n4973 ;
  assign n7354 = ~n3355 & n4972 ;
  assign n7355 = ( ~n3389 & n7353 ) | ( ~n3389 & n7354 ) | ( n7353 & n7354 ) ;
  assign n7356 = ( ~n7351 & n7352 ) | ( ~n7351 & n7355 ) | ( n7352 & n7355 ) ;
  assign n7357 = ( ~x20 & n7351 ) | ( ~x20 & n7356 ) | ( n7351 & n7356 ) ;
  assign n7358 = ( n7351 & n7356 ) | ( n7351 & ~n7357 ) | ( n7356 & ~n7357 ) ;
  assign n7359 = ( x20 & n7357 ) | ( x20 & ~n7358 ) | ( n7357 & ~n7358 ) ;
  assign n7360 = ( n7057 & n7065 ) | ( n7057 & ~n7066 ) | ( n7065 & ~n7066 ) ;
  assign n7361 = n7066 & ~n7360 ;
  assign n7362 = ( n7350 & n7359 ) | ( n7350 & n7361 ) | ( n7359 & n7361 ) ;
  assign n7363 = n4974 & n6200 ;
  assign n7364 = ~n3300 & n4972 ;
  assign n7365 = n3355 | n4973 ;
  assign n7366 = n3239 & n5398 ;
  assign n7367 = ( ~n3355 & n7365 ) | ( ~n3355 & n7366 ) | ( n7365 & n7366 ) ;
  assign n7368 = ( ~n7363 & n7364 ) | ( ~n7363 & n7367 ) | ( n7364 & n7367 ) ;
  assign n7369 = ( ~x20 & n7363 ) | ( ~x20 & n7368 ) | ( n7363 & n7368 ) ;
  assign n7370 = ( n7363 & n7368 ) | ( n7363 & ~n7369 ) | ( n7368 & ~n7369 ) ;
  assign n7371 = ( x20 & n7369 ) | ( x20 & ~n7370 ) | ( n7369 & ~n7370 ) ;
  assign n7372 = ( n6824 & n7050 ) | ( n6824 & ~n7067 ) | ( n7050 & ~n7067 ) ;
  assign n7373 = ( n7067 & ~n7068 ) | ( n7067 & n7372 ) | ( ~n7068 & n7372 ) ;
  assign n7374 = ( n7362 & n7371 ) | ( n7362 & n7373 ) | ( n7371 & n7373 ) ;
  assign n7375 = n4974 & ~n6243 ;
  assign n7376 = n3153 & n5398 ;
  assign n7377 = n3300 | n4973 ;
  assign n7378 = n3239 & n4972 ;
  assign n7379 = ( ~n3300 & n7377 ) | ( ~n3300 & n7378 ) | ( n7377 & n7378 ) ;
  assign n7380 = ( ~n7375 & n7376 ) | ( ~n7375 & n7379 ) | ( n7376 & n7379 ) ;
  assign n7381 = ( ~x20 & n7375 ) | ( ~x20 & n7380 ) | ( n7375 & n7380 ) ;
  assign n7382 = ( n7375 & n7380 ) | ( n7375 & ~n7381 ) | ( n7380 & ~n7381 ) ;
  assign n7383 = ( x20 & n7381 ) | ( x20 & ~n7382 ) | ( n7381 & ~n7382 ) ;
  assign n7384 = ( ~n7068 & n7078 ) | ( ~n7068 & n7081 ) | ( n7078 & n7081 ) ;
  assign n7385 = ( n7068 & ~n7082 ) | ( n7068 & n7384 ) | ( ~n7082 & n7384 ) ;
  assign n7386 = ( n7374 & n7383 ) | ( n7374 & n7385 ) | ( n7383 & n7385 ) ;
  assign n7387 = ( ~n7082 & n7091 ) | ( ~n7082 & n7093 ) | ( n7091 & n7093 ) ;
  assign n7388 = ( n7082 & ~n7094 ) | ( n7082 & n7387 ) | ( ~n7094 & n7387 ) ;
  assign n7389 = n4974 & n5710 ;
  assign n7390 = n3153 & n4972 ;
  assign n7391 = n3239 & ~n4973 ;
  assign n7392 = n3078 & n5398 ;
  assign n7393 = ( n3239 & ~n7391 ) | ( n3239 & n7392 ) | ( ~n7391 & n7392 ) ;
  assign n7394 = ( ~n7389 & n7390 ) | ( ~n7389 & n7393 ) | ( n7390 & n7393 ) ;
  assign n7395 = ( ~x20 & n7389 ) | ( ~x20 & n7394 ) | ( n7389 & n7394 ) ;
  assign n7396 = ( n7389 & n7394 ) | ( n7389 & ~n7395 ) | ( n7394 & ~n7395 ) ;
  assign n7397 = ( x20 & n7395 ) | ( x20 & ~n7396 ) | ( n7395 & ~n7396 ) ;
  assign n7398 = ( n7386 & n7388 ) | ( n7386 & n7397 ) | ( n7388 & n7397 ) ;
  assign n7399 = ( ~n7094 & n7103 ) | ( ~n7094 & n7105 ) | ( n7103 & n7105 ) ;
  assign n7400 = ( n7094 & ~n7106 ) | ( n7094 & n7399 ) | ( ~n7106 & n7399 ) ;
  assign n7401 = n3078 & ~n4972 ;
  assign n7402 = ~n3046 & n5398 ;
  assign n7403 = ( n3078 & ~n7401 ) | ( n3078 & n7402 ) | ( ~n7401 & n7402 ) ;
  assign n7404 = n3153 & ~n4973 ;
  assign n7405 = ( n3153 & n7403 ) | ( n3153 & ~n7404 ) | ( n7403 & ~n7404 ) ;
  assign n7406 = ( n4974 & ~n6267 ) | ( n4974 & n7405 ) | ( ~n6267 & n7405 ) ;
  assign n7407 = n7405 & ~n7406 ;
  assign n7408 = ( ~x20 & n7406 ) | ( ~x20 & n7407 ) | ( n7406 & n7407 ) ;
  assign n7409 = ( n7406 & n7407 ) | ( n7406 & ~n7408 ) | ( n7407 & ~n7408 ) ;
  assign n7410 = ( x20 & n7408 ) | ( x20 & ~n7409 ) | ( n7408 & ~n7409 ) ;
  assign n7411 = ( n7398 & n7400 ) | ( n7398 & n7410 ) | ( n7400 & n7410 ) ;
  assign n7412 = ( ~n7106 & n7115 ) | ( ~n7106 & n7117 ) | ( n7115 & n7117 ) ;
  assign n7413 = ( n7106 & ~n7118 ) | ( n7106 & n7412 ) | ( ~n7118 & n7412 ) ;
  assign n7414 = n4974 & n6279 ;
  assign n7415 = ~n2965 & n5398 ;
  assign n7416 = n3078 & ~n4973 ;
  assign n7417 = ~n3046 & n4972 ;
  assign n7418 = ( n3078 & ~n7416 ) | ( n3078 & n7417 ) | ( ~n7416 & n7417 ) ;
  assign n7419 = ( ~n7414 & n7415 ) | ( ~n7414 & n7418 ) | ( n7415 & n7418 ) ;
  assign n7420 = ( ~x20 & n7414 ) | ( ~x20 & n7419 ) | ( n7414 & n7419 ) ;
  assign n7421 = ( n7414 & n7419 ) | ( n7414 & ~n7420 ) | ( n7419 & ~n7420 ) ;
  assign n7422 = ( x20 & n7420 ) | ( x20 & ~n7421 ) | ( n7420 & ~n7421 ) ;
  assign n7423 = ( n7411 & n7413 ) | ( n7411 & n7422 ) | ( n7413 & n7422 ) ;
  assign n7424 = n4974 & ~n5768 ;
  assign n7425 = ~n2910 & n5398 ;
  assign n7426 = n3046 | n4973 ;
  assign n7427 = ~n2965 & n4972 ;
  assign n7428 = ( ~n3046 & n7426 ) | ( ~n3046 & n7427 ) | ( n7426 & n7427 ) ;
  assign n7429 = ( ~n7424 & n7425 ) | ( ~n7424 & n7428 ) | ( n7425 & n7428 ) ;
  assign n7430 = ( ~x20 & n7424 ) | ( ~x20 & n7429 ) | ( n7424 & n7429 ) ;
  assign n7431 = ( n7424 & n7429 ) | ( n7424 & ~n7430 ) | ( n7429 & ~n7430 ) ;
  assign n7432 = ( x20 & n7430 ) | ( x20 & ~n7431 ) | ( n7430 & ~n7431 ) ;
  assign n7433 = ( ~n7118 & n7120 ) | ( ~n7118 & n7129 ) | ( n7120 & n7129 ) ;
  assign n7434 = ( n7118 & ~n7130 ) | ( n7118 & n7433 ) | ( ~n7130 & n7433 ) ;
  assign n7435 = ( n7423 & n7432 ) | ( n7423 & n7434 ) | ( n7432 & n7434 ) ;
  assign n7436 = n4974 & n5543 ;
  assign n7437 = ~n2910 & n4972 ;
  assign n7438 = n2965 | n4973 ;
  assign n7439 = n2843 & n5398 ;
  assign n7440 = ( ~n2965 & n7438 ) | ( ~n2965 & n7439 ) | ( n7438 & n7439 ) ;
  assign n7441 = ( ~n7436 & n7437 ) | ( ~n7436 & n7440 ) | ( n7437 & n7440 ) ;
  assign n7442 = ( ~x20 & n7436 ) | ( ~x20 & n7441 ) | ( n7436 & n7441 ) ;
  assign n7443 = ( n7436 & n7441 ) | ( n7436 & ~n7442 ) | ( n7441 & ~n7442 ) ;
  assign n7444 = ( x20 & n7442 ) | ( x20 & ~n7443 ) | ( n7442 & ~n7443 ) ;
  assign n7445 = ( ~n7130 & n7132 ) | ( ~n7130 & n7142 ) | ( n7132 & n7142 ) ;
  assign n7446 = ( n7130 & ~n7143 ) | ( n7130 & n7445 ) | ( ~n7143 & n7445 ) ;
  assign n7447 = ( n7435 & n7444 ) | ( n7435 & n7446 ) | ( n7444 & n7446 ) ;
  assign n7448 = ( ~n7143 & n7152 ) | ( ~n7143 & n7154 ) | ( n7152 & n7154 ) ;
  assign n7449 = ( n7143 & ~n7155 ) | ( n7143 & n7448 ) | ( ~n7155 & n7448 ) ;
  assign n7450 = n4974 & n5791 ;
  assign n7451 = ~n2810 & n5398 ;
  assign n7452 = n2910 | n4973 ;
  assign n7453 = n2843 & n4972 ;
  assign n7454 = ( ~n2910 & n7452 ) | ( ~n2910 & n7453 ) | ( n7452 & n7453 ) ;
  assign n7455 = ( ~n7450 & n7451 ) | ( ~n7450 & n7454 ) | ( n7451 & n7454 ) ;
  assign n7456 = ( ~x20 & n7450 ) | ( ~x20 & n7455 ) | ( n7450 & n7455 ) ;
  assign n7457 = ( n7450 & n7455 ) | ( n7450 & ~n7456 ) | ( n7455 & ~n7456 ) ;
  assign n7458 = ( x20 & n7456 ) | ( x20 & ~n7457 ) | ( n7456 & ~n7457 ) ;
  assign n7459 = ( n7447 & n7449 ) | ( n7447 & n7458 ) | ( n7449 & n7458 ) ;
  assign n7460 = ( n7155 & ~n7164 ) | ( n7155 & n7166 ) | ( ~n7164 & n7166 ) ;
  assign n7461 = ( ~n7155 & n7167 ) | ( ~n7155 & n7460 ) | ( n7167 & n7460 ) ;
  assign n7462 = n4974 & ~n5586 ;
  assign n7463 = ~n2725 & n5398 ;
  assign n7464 = n2843 & ~n4973 ;
  assign n7465 = ~n2810 & n4972 ;
  assign n7466 = ( n2843 & ~n7464 ) | ( n2843 & n7465 ) | ( ~n7464 & n7465 ) ;
  assign n7467 = ( ~n7462 & n7463 ) | ( ~n7462 & n7466 ) | ( n7463 & n7466 ) ;
  assign n7468 = ( ~x20 & n7462 ) | ( ~x20 & n7467 ) | ( n7462 & n7467 ) ;
  assign n7469 = ( n7462 & n7467 ) | ( n7462 & ~n7468 ) | ( n7467 & ~n7468 ) ;
  assign n7470 = ( x20 & n7468 ) | ( x20 & ~n7469 ) | ( n7468 & ~n7469 ) ;
  assign n7471 = ( n7459 & ~n7461 ) | ( n7459 & n7470 ) | ( ~n7461 & n7470 ) ;
  assign n7472 = ( n7167 & ~n7176 ) | ( n7167 & n7178 ) | ( ~n7176 & n7178 ) ;
  assign n7473 = ( ~n7167 & n7179 ) | ( ~n7167 & n7472 ) | ( n7179 & n7472 ) ;
  assign n7474 = n2725 | n4972 ;
  assign n7475 = n2635 & n5398 ;
  assign n7476 = ( ~n2725 & n7474 ) | ( ~n2725 & n7475 ) | ( n7474 & n7475 ) ;
  assign n7477 = n2810 | n4973 ;
  assign n7478 = ( ~n2810 & n7476 ) | ( ~n2810 & n7477 ) | ( n7476 & n7477 ) ;
  assign n7479 = ( n4966 & n4969 ) | ( n4966 & n5232 ) | ( n4969 & n5232 ) ;
  assign n7480 = ( ~n4969 & n7478 ) | ( ~n4969 & n7479 ) | ( n7478 & n7479 ) ;
  assign n7481 = x20 | n7480 ;
  assign n7482 = ( x20 & n7480 ) | ( x20 & ~n7481 ) | ( n7480 & ~n7481 ) ;
  assign n7483 = n7481 & ~n7482 ;
  assign n7484 = ( n7471 & ~n7473 ) | ( n7471 & n7483 ) | ( ~n7473 & n7483 ) ;
  assign n7485 = ( ~n7179 & n7188 ) | ( ~n7179 & n7190 ) | ( n7188 & n7190 ) ;
  assign n7486 = ( n7179 & ~n7191 ) | ( n7179 & n7485 ) | ( ~n7191 & n7485 ) ;
  assign n7487 = n4974 & ~n5425 ;
  assign n7488 = n2552 & n5398 ;
  assign n7489 = n2725 | n4973 ;
  assign n7490 = n2635 & n4972 ;
  assign n7491 = ( ~n2725 & n7489 ) | ( ~n2725 & n7490 ) | ( n7489 & n7490 ) ;
  assign n7492 = ( ~n7487 & n7488 ) | ( ~n7487 & n7491 ) | ( n7488 & n7491 ) ;
  assign n7493 = ( ~x20 & n7487 ) | ( ~x20 & n7492 ) | ( n7487 & n7492 ) ;
  assign n7494 = ( n7487 & n7492 ) | ( n7487 & ~n7493 ) | ( n7492 & ~n7493 ) ;
  assign n7495 = ( x20 & n7493 ) | ( x20 & ~n7494 ) | ( n7493 & ~n7494 ) ;
  assign n7496 = ( n7484 & n7486 ) | ( n7484 & n7495 ) | ( n7486 & n7495 ) ;
  assign n7497 = ( n7191 & ~n7200 ) | ( n7191 & n7202 ) | ( ~n7200 & n7202 ) ;
  assign n7498 = ( ~n7191 & n7203 ) | ( ~n7191 & n7497 ) | ( n7203 & n7497 ) ;
  assign n7499 = n4974 & ~n5270 ;
  assign n7500 = n2552 & n4972 ;
  assign n7501 = n2635 & ~n4973 ;
  assign n7502 = ~n2491 & n5398 ;
  assign n7503 = ( n2635 & ~n7501 ) | ( n2635 & n7502 ) | ( ~n7501 & n7502 ) ;
  assign n7504 = ( ~n7499 & n7500 ) | ( ~n7499 & n7503 ) | ( n7500 & n7503 ) ;
  assign n7505 = ( ~x20 & n7499 ) | ( ~x20 & n7504 ) | ( n7499 & n7504 ) ;
  assign n7506 = ( n7499 & n7504 ) | ( n7499 & ~n7505 ) | ( n7504 & ~n7505 ) ;
  assign n7507 = ( x20 & n7505 ) | ( x20 & ~n7506 ) | ( n7505 & ~n7506 ) ;
  assign n7508 = ( n7496 & ~n7498 ) | ( n7496 & n7507 ) | ( ~n7498 & n7507 ) ;
  assign n7509 = ( ~n7203 & n7213 ) | ( ~n7203 & n7215 ) | ( n7213 & n7215 ) ;
  assign n7510 = ( n7203 & ~n7216 ) | ( n7203 & n7509 ) | ( ~n7216 & n7509 ) ;
  assign n7511 = n4974 & ~n5084 ;
  assign n7512 = n2396 & n5398 ;
  assign n7513 = n2552 & ~n4973 ;
  assign n7514 = ~n2491 & n4972 ;
  assign n7515 = ( n2552 & ~n7513 ) | ( n2552 & n7514 ) | ( ~n7513 & n7514 ) ;
  assign n7516 = ( ~n7511 & n7512 ) | ( ~n7511 & n7515 ) | ( n7512 & n7515 ) ;
  assign n7517 = ( ~x20 & n7511 ) | ( ~x20 & n7516 ) | ( n7511 & n7516 ) ;
  assign n7518 = ( n7511 & n7516 ) | ( n7511 & ~n7517 ) | ( n7516 & ~n7517 ) ;
  assign n7519 = ( x20 & n7517 ) | ( x20 & ~n7518 ) | ( n7517 & ~n7518 ) ;
  assign n7520 = ( n7508 & n7510 ) | ( n7508 & n7519 ) | ( n7510 & n7519 ) ;
  assign n7521 = ( ~n7216 & n7225 ) | ( ~n7216 & n7227 ) | ( n7225 & n7227 ) ;
  assign n7522 = ( n7216 & ~n7228 ) | ( n7216 & n7521 ) | ( ~n7228 & n7521 ) ;
  assign n7523 = ~n4900 & n4974 ;
  assign n7524 = n2396 & n4972 ;
  assign n7525 = ~n2298 & n5398 ;
  assign n7526 = ~n2491 & n4973 ;
  assign n7527 = n7525 | n7526 ;
  assign n7528 = ( ~n7523 & n7524 ) | ( ~n7523 & n7527 ) | ( n7524 & n7527 ) ;
  assign n7529 = ( ~x20 & n7523 ) | ( ~x20 & n7528 ) | ( n7523 & n7528 ) ;
  assign n7530 = ( n7523 & n7528 ) | ( n7523 & ~n7529 ) | ( n7528 & ~n7529 ) ;
  assign n7531 = ( x20 & n7529 ) | ( x20 & ~n7530 ) | ( n7529 & ~n7530 ) ;
  assign n7532 = ( n7520 & n7522 ) | ( n7520 & n7531 ) | ( n7522 & n7531 ) ;
  assign n7533 = ( n7228 & ~n7230 ) | ( n7228 & n7240 ) | ( ~n7230 & n7240 ) ;
  assign n7534 = ( n7230 & ~n7241 ) | ( n7230 & n7533 ) | ( ~n7241 & n7533 ) ;
  assign n7535 = ~n4660 & n5508 ;
  assign n7536 = ~n2023 & n5507 ;
  assign n7537 = n2174 & n5504 ;
  assign n7538 = n2089 & n5666 ;
  assign n7539 = n7537 | n7538 ;
  assign n7540 = ( ~n7535 & n7536 ) | ( ~n7535 & n7539 ) | ( n7536 & n7539 ) ;
  assign n7541 = ( ~x17 & n7535 ) | ( ~x17 & n7540 ) | ( n7535 & n7540 ) ;
  assign n7542 = ( n7535 & n7540 ) | ( n7535 & ~n7541 ) | ( n7540 & ~n7541 ) ;
  assign n7543 = ( x17 & n7541 ) | ( x17 & ~n7542 ) | ( n7541 & ~n7542 ) ;
  assign n7544 = ( n7532 & n7534 ) | ( n7532 & n7543 ) | ( n7534 & n7543 ) ;
  assign n7545 = ( n7241 & ~n7243 ) | ( n7241 & n7252 ) | ( ~n7243 & n7252 ) ;
  assign n7546 = ( n7243 & ~n7253 ) | ( n7243 & n7545 ) | ( ~n7253 & n7545 ) ;
  assign n7547 = n4146 & n5966 ;
  assign n7548 = ~n1669 & n6464 ;
  assign n7549 = n1852 & ~n5970 ;
  assign n7550 = ~n1750 & n5969 ;
  assign n7551 = ( n1852 & ~n7549 ) | ( n1852 & n7550 ) | ( ~n7549 & n7550 ) ;
  assign n7552 = ( ~n7547 & n7548 ) | ( ~n7547 & n7551 ) | ( n7548 & n7551 ) ;
  assign n7553 = ( ~x14 & n7547 ) | ( ~x14 & n7552 ) | ( n7547 & n7552 ) ;
  assign n7554 = ( n7547 & n7552 ) | ( n7547 & ~n7553 ) | ( n7552 & ~n7553 ) ;
  assign n7555 = ( x14 & n7553 ) | ( x14 & ~n7554 ) | ( n7553 & ~n7554 ) ;
  assign n7556 = ( n7544 & n7546 ) | ( n7544 & n7555 ) | ( n7546 & n7555 ) ;
  assign n7557 = ( ~n7253 & n7255 ) | ( ~n7253 & n7264 ) | ( n7255 & n7264 ) ;
  assign n7558 = ( ~n7264 & n7265 ) | ( ~n7264 & n7557 ) | ( n7265 & n7557 ) ;
  assign n7559 = ~n3779 & n6584 ;
  assign n7560 = n1267 & n7022 ;
  assign n7561 = n1458 & ~n6588 ;
  assign n7562 = ~n1338 & n6587 ;
  assign n7563 = ( n1458 & ~n7561 ) | ( n1458 & n7562 ) | ( ~n7561 & n7562 ) ;
  assign n7564 = ( ~n7559 & n7560 ) | ( ~n7559 & n7563 ) | ( n7560 & n7563 ) ;
  assign n7565 = ( ~x11 & n7559 ) | ( ~x11 & n7564 ) | ( n7559 & n7564 ) ;
  assign n7566 = ( n7559 & n7564 ) | ( n7559 & ~n7565 ) | ( n7564 & ~n7565 ) ;
  assign n7567 = ( x11 & n7565 ) | ( x11 & ~n7566 ) | ( n7565 & ~n7566 ) ;
  assign n7568 = ( n7556 & ~n7558 ) | ( n7556 & n7567 ) | ( ~n7558 & n7567 ) ;
  assign n7569 = ~n3791 & n6584 ;
  assign n7570 = n1267 & n6587 ;
  assign n7571 = n1338 | n6588 ;
  assign n7572 = ~n1246 & n7022 ;
  assign n7573 = ( ~n1338 & n7571 ) | ( ~n1338 & n7572 ) | ( n7571 & n7572 ) ;
  assign n7574 = ( ~n7569 & n7570 ) | ( ~n7569 & n7573 ) | ( n7570 & n7573 ) ;
  assign n7575 = ( ~x11 & n7569 ) | ( ~x11 & n7574 ) | ( n7569 & n7574 ) ;
  assign n7576 = ( n7569 & n7574 ) | ( n7569 & ~n7575 ) | ( n7574 & ~n7575 ) ;
  assign n7577 = ( x11 & n7575 ) | ( x11 & ~n7576 ) | ( n7575 & ~n7576 ) ;
  assign n7578 = ( ~n7265 & n7267 ) | ( ~n7265 & n7276 ) | ( n7267 & n7276 ) ;
  assign n7579 = ( n7265 & ~n7277 ) | ( n7265 & n7578 ) | ( ~n7277 & n7578 ) ;
  assign n7580 = ( n7568 & n7577 ) | ( n7568 & n7579 ) | ( n7577 & n7579 ) ;
  assign n7581 = n3797 & n7296 ;
  assign n7582 = ~n3692 & n7299 ;
  assign n7583 = ~n3658 & n7300 ;
  assign n7584 = n7582 | n7583 ;
  assign n7585 = ( ~x8 & n7581 ) | ( ~x8 & n7584 ) | ( n7581 & n7584 ) ;
  assign n7586 = ( n7581 & n7584 ) | ( n7581 & ~n7585 ) | ( n7584 & ~n7585 ) ;
  assign n7587 = ( x8 & n7585 ) | ( x8 & ~n7586 ) | ( n7585 & ~n7586 ) ;
  assign n7588 = ( ~n7277 & n7279 ) | ( ~n7277 & n7288 ) | ( n7279 & n7288 ) ;
  assign n7589 = ( ~n7288 & n7289 ) | ( ~n7288 & n7588 ) | ( n7289 & n7588 ) ;
  assign n7590 = ( n7580 & n7587 ) | ( n7580 & ~n7589 ) | ( n7587 & ~n7589 ) ;
  assign n7591 = n5508 & n6061 ;
  assign n7592 = n3479 & n5666 ;
  assign n7593 = n3533 | n5504 ;
  assign n7594 = ~n3389 & n5507 ;
  assign n7595 = ( ~n3533 & n7593 ) | ( ~n3533 & n7594 ) | ( n7593 & n7594 ) ;
  assign n7596 = ( ~n7591 & n7592 ) | ( ~n7591 & n7595 ) | ( n7592 & n7595 ) ;
  assign n7597 = ( ~x17 & n7591 ) | ( ~x17 & n7596 ) | ( n7591 & n7596 ) ;
  assign n7598 = ( n7591 & n7596 ) | ( n7591 & ~n7597 ) | ( n7596 & ~n7597 ) ;
  assign n7599 = ( x17 & n7597 ) | ( x17 & ~n7598 ) | ( n7597 & ~n7598 ) ;
  assign n7600 = ( n3479 & n5508 ) | ( n3479 & n6009 ) | ( n5508 & n6009 ) ;
  assign n7601 = ~n3533 & n5666 ;
  assign n7602 = ~n3586 & n5504 ;
  assign n7603 = n7601 | n7602 ;
  assign n7604 = ~n3479 & n5507 ;
  assign n7605 = ( n5507 & n7603 ) | ( n5507 & ~n7604 ) | ( n7603 & ~n7604 ) ;
  assign n7606 = ( ~n6608 & n7600 ) | ( ~n6608 & n7605 ) | ( n7600 & n7605 ) ;
  assign n7607 = ~n3586 & n5506 ;
  assign n7608 = x17 & n7607 ;
  assign n7609 = ( n5508 & n6009 ) | ( n5508 & n6618 ) | ( n6009 & n6618 ) ;
  assign n7610 = ~n3533 & n5507 ;
  assign n7611 = n3586 | n5666 ;
  assign n7612 = ( ~n3586 & n7610 ) | ( ~n3586 & n7611 ) | ( n7610 & n7611 ) ;
  assign n7613 = n7609 | n7612 ;
  assign n7614 = ( x17 & n7608 ) | ( x17 & n7613 ) | ( n7608 & n7613 ) ;
  assign n7615 = n7606 | n7614 ;
  assign n7616 = x17 & ~n7615 ;
  assign n7617 = ( n7326 & n7599 ) | ( n7326 & n7616 ) | ( n7599 & n7616 ) ;
  assign n7618 = ~n3355 & n5507 ;
  assign n7619 = n3389 | n5666 ;
  assign n7620 = ( ~n3389 & n7618 ) | ( ~n3389 & n7619 ) | ( n7618 & n7619 ) ;
  assign n7621 = ~n3479 & n5504 ;
  assign n7622 = ( n5504 & n7620 ) | ( n5504 & ~n7621 ) | ( n7620 & ~n7621 ) ;
  assign n7623 = ( n5508 & ~n6104 ) | ( n5508 & n7622 ) | ( ~n6104 & n7622 ) ;
  assign n7624 = n7622 & ~n7623 ;
  assign n7625 = ( ~x17 & n7623 ) | ( ~x17 & n7624 ) | ( n7623 & n7624 ) ;
  assign n7626 = ( n7623 & n7624 ) | ( n7623 & ~n7625 ) | ( n7624 & ~n7625 ) ;
  assign n7627 = ( x17 & n7625 ) | ( x17 & ~n7626 ) | ( n7625 & ~n7626 ) ;
  assign n7628 = ( n7327 & n7328 ) | ( n7327 & n7331 ) | ( n7328 & n7331 ) ;
  assign n7629 = ~n7327 & n7332 ;
  assign n7630 = ( n7327 & ~n7628 ) | ( n7327 & n7629 ) | ( ~n7628 & n7629 ) ;
  assign n7631 = ( n7617 & n7627 ) | ( n7617 & n7630 ) | ( n7627 & n7630 ) ;
  assign n7632 = n5508 & ~n6154 ;
  assign n7633 = ~n3300 & n5507 ;
  assign n7634 = ~n3355 & n5666 ;
  assign n7635 = ~n3389 & n5504 ;
  assign n7636 = n7634 | n7635 ;
  assign n7637 = ( ~n7632 & n7633 ) | ( ~n7632 & n7636 ) | ( n7633 & n7636 ) ;
  assign n7638 = ( ~x17 & n7632 ) | ( ~x17 & n7637 ) | ( n7632 & n7637 ) ;
  assign n7639 = ( n7632 & n7637 ) | ( n7632 & ~n7638 ) | ( n7637 & ~n7638 ) ;
  assign n7640 = ( x17 & n7638 ) | ( x17 & ~n7639 ) | ( n7638 & ~n7639 ) ;
  assign n7641 = ( n7325 & n7333 ) | ( n7325 & ~n7334 ) | ( n7333 & ~n7334 ) ;
  assign n7642 = n7334 & ~n7641 ;
  assign n7643 = ( n7631 & n7640 ) | ( n7631 & n7642 ) | ( n7640 & n7642 ) ;
  assign n7644 = n5508 & n6200 ;
  assign n7645 = ~n3300 & n5666 ;
  assign n7646 = n3355 | n5504 ;
  assign n7647 = n3239 & n5507 ;
  assign n7648 = ( ~n3355 & n7646 ) | ( ~n3355 & n7647 ) | ( n7646 & n7647 ) ;
  assign n7649 = ( ~n7644 & n7645 ) | ( ~n7644 & n7648 ) | ( n7645 & n7648 ) ;
  assign n7650 = ( ~x17 & n7644 ) | ( ~x17 & n7649 ) | ( n7644 & n7649 ) ;
  assign n7651 = ( n7644 & n7649 ) | ( n7644 & ~n7650 ) | ( n7649 & ~n7650 ) ;
  assign n7652 = ( x17 & n7650 ) | ( x17 & ~n7651 ) | ( n7650 & ~n7651 ) ;
  assign n7653 = ( n7058 & n7318 ) | ( n7058 & ~n7335 ) | ( n7318 & ~n7335 ) ;
  assign n7654 = ( n7335 & ~n7336 ) | ( n7335 & n7653 ) | ( ~n7336 & n7653 ) ;
  assign n7655 = ( n7643 & n7652 ) | ( n7643 & n7654 ) | ( n7652 & n7654 ) ;
  assign n7656 = n5508 & ~n6243 ;
  assign n7657 = n3153 & n5507 ;
  assign n7658 = n3239 & n5666 ;
  assign n7659 = ~n3300 & n5504 ;
  assign n7660 = n7658 | n7659 ;
  assign n7661 = ( ~n7656 & n7657 ) | ( ~n7656 & n7660 ) | ( n7657 & n7660 ) ;
  assign n7662 = ( ~x17 & n7656 ) | ( ~x17 & n7661 ) | ( n7656 & n7661 ) ;
  assign n7663 = ( n7656 & n7661 ) | ( n7656 & ~n7662 ) | ( n7661 & ~n7662 ) ;
  assign n7664 = ( x17 & n7662 ) | ( x17 & ~n7663 ) | ( n7662 & ~n7663 ) ;
  assign n7665 = ( ~n7336 & n7346 ) | ( ~n7336 & n7349 ) | ( n7346 & n7349 ) ;
  assign n7666 = ( n7336 & ~n7350 ) | ( n7336 & n7665 ) | ( ~n7350 & n7665 ) ;
  assign n7667 = ( n7655 & n7664 ) | ( n7655 & n7666 ) | ( n7664 & n7666 ) ;
  assign n7668 = ( ~n7350 & n7359 ) | ( ~n7350 & n7361 ) | ( n7359 & n7361 ) ;
  assign n7669 = ( n7350 & ~n7362 ) | ( n7350 & n7668 ) | ( ~n7362 & n7668 ) ;
  assign n7670 = n5508 & n5710 ;
  assign n7671 = n3153 & n5666 ;
  assign n7672 = n3078 & n5507 ;
  assign n7673 = n3239 & n5504 ;
  assign n7674 = n7672 | n7673 ;
  assign n7675 = ( ~n7670 & n7671 ) | ( ~n7670 & n7674 ) | ( n7671 & n7674 ) ;
  assign n7676 = ( ~x17 & n7670 ) | ( ~x17 & n7675 ) | ( n7670 & n7675 ) ;
  assign n7677 = ( n7670 & n7675 ) | ( n7670 & ~n7676 ) | ( n7675 & ~n7676 ) ;
  assign n7678 = ( x17 & n7676 ) | ( x17 & ~n7677 ) | ( n7676 & ~n7677 ) ;
  assign n7679 = ( n7667 & n7669 ) | ( n7667 & n7678 ) | ( n7669 & n7678 ) ;
  assign n7680 = ( ~n7362 & n7371 ) | ( ~n7362 & n7373 ) | ( n7371 & n7373 ) ;
  assign n7681 = ( n7362 & ~n7374 ) | ( n7362 & n7680 ) | ( ~n7374 & n7680 ) ;
  assign n7682 = n3078 & ~n5666 ;
  assign n7683 = ~n3046 & n5507 ;
  assign n7684 = ( n3078 & ~n7682 ) | ( n3078 & n7683 ) | ( ~n7682 & n7683 ) ;
  assign n7685 = ~n3153 & n5504 ;
  assign n7686 = ( n5504 & n7684 ) | ( n5504 & ~n7685 ) | ( n7684 & ~n7685 ) ;
  assign n7687 = ( n5508 & ~n6267 ) | ( n5508 & n7686 ) | ( ~n6267 & n7686 ) ;
  assign n7688 = n7686 & ~n7687 ;
  assign n7689 = ( ~x17 & n7687 ) | ( ~x17 & n7688 ) | ( n7687 & n7688 ) ;
  assign n7690 = ( n7687 & n7688 ) | ( n7687 & ~n7689 ) | ( n7688 & ~n7689 ) ;
  assign n7691 = ( x17 & n7689 ) | ( x17 & ~n7690 ) | ( n7689 & ~n7690 ) ;
  assign n7692 = ( n7679 & n7681 ) | ( n7679 & n7691 ) | ( n7681 & n7691 ) ;
  assign n7693 = ( ~n7374 & n7383 ) | ( ~n7374 & n7385 ) | ( n7383 & n7385 ) ;
  assign n7694 = ( n7374 & ~n7386 ) | ( n7374 & n7693 ) | ( ~n7386 & n7693 ) ;
  assign n7695 = n5508 & n6279 ;
  assign n7696 = ~n2965 & n5507 ;
  assign n7697 = n3078 & n5504 ;
  assign n7698 = ~n3046 & n5666 ;
  assign n7699 = n7697 | n7698 ;
  assign n7700 = ( ~n7695 & n7696 ) | ( ~n7695 & n7699 ) | ( n7696 & n7699 ) ;
  assign n7701 = ( ~x17 & n7695 ) | ( ~x17 & n7700 ) | ( n7695 & n7700 ) ;
  assign n7702 = ( n7695 & n7700 ) | ( n7695 & ~n7701 ) | ( n7700 & ~n7701 ) ;
  assign n7703 = ( x17 & n7701 ) | ( x17 & ~n7702 ) | ( n7701 & ~n7702 ) ;
  assign n7704 = ( n7692 & n7694 ) | ( n7692 & n7703 ) | ( n7694 & n7703 ) ;
  assign n7705 = n5508 & ~n5768 ;
  assign n7706 = ~n2910 & n5507 ;
  assign n7707 = n3046 | n5504 ;
  assign n7708 = ~n2965 & n5666 ;
  assign n7709 = ( ~n3046 & n7707 ) | ( ~n3046 & n7708 ) | ( n7707 & n7708 ) ;
  assign n7710 = ( ~n7705 & n7706 ) | ( ~n7705 & n7709 ) | ( n7706 & n7709 ) ;
  assign n7711 = ( ~x17 & n7705 ) | ( ~x17 & n7710 ) | ( n7705 & n7710 ) ;
  assign n7712 = ( n7705 & n7710 ) | ( n7705 & ~n7711 ) | ( n7710 & ~n7711 ) ;
  assign n7713 = ( x17 & n7711 ) | ( x17 & ~n7712 ) | ( n7711 & ~n7712 ) ;
  assign n7714 = ( ~n7386 & n7388 ) | ( ~n7386 & n7397 ) | ( n7388 & n7397 ) ;
  assign n7715 = ( n7386 & ~n7398 ) | ( n7386 & n7714 ) | ( ~n7398 & n7714 ) ;
  assign n7716 = ( n7704 & n7713 ) | ( n7704 & n7715 ) | ( n7713 & n7715 ) ;
  assign n7717 = n5508 & n5543 ;
  assign n7718 = ~n2910 & n5666 ;
  assign n7719 = n2965 | n5504 ;
  assign n7720 = n2843 & n5507 ;
  assign n7721 = ( ~n2965 & n7719 ) | ( ~n2965 & n7720 ) | ( n7719 & n7720 ) ;
  assign n7722 = ( ~n7717 & n7718 ) | ( ~n7717 & n7721 ) | ( n7718 & n7721 ) ;
  assign n7723 = ( ~x17 & n7717 ) | ( ~x17 & n7722 ) | ( n7717 & n7722 ) ;
  assign n7724 = ( n7717 & n7722 ) | ( n7717 & ~n7723 ) | ( n7722 & ~n7723 ) ;
  assign n7725 = ( x17 & n7723 ) | ( x17 & ~n7724 ) | ( n7723 & ~n7724 ) ;
  assign n7726 = ( ~n7398 & n7400 ) | ( ~n7398 & n7410 ) | ( n7400 & n7410 ) ;
  assign n7727 = ( n7398 & ~n7411 ) | ( n7398 & n7726 ) | ( ~n7411 & n7726 ) ;
  assign n7728 = ( n7716 & n7725 ) | ( n7716 & n7727 ) | ( n7725 & n7727 ) ;
  assign n7729 = n5508 & n5791 ;
  assign n7730 = ~n2810 & n5507 ;
  assign n7731 = n2910 | n5504 ;
  assign n7732 = n2843 & n5666 ;
  assign n7733 = ( ~n2910 & n7731 ) | ( ~n2910 & n7732 ) | ( n7731 & n7732 ) ;
  assign n7734 = ( ~n7729 & n7730 ) | ( ~n7729 & n7733 ) | ( n7730 & n7733 ) ;
  assign n7735 = ( ~x17 & n7729 ) | ( ~x17 & n7734 ) | ( n7729 & n7734 ) ;
  assign n7736 = ( n7729 & n7734 ) | ( n7729 & ~n7735 ) | ( n7734 & ~n7735 ) ;
  assign n7737 = ( x17 & n7735 ) | ( x17 & ~n7736 ) | ( n7735 & ~n7736 ) ;
  assign n7738 = ( ~n7411 & n7413 ) | ( ~n7411 & n7422 ) | ( n7413 & n7422 ) ;
  assign n7739 = ( n7411 & ~n7423 ) | ( n7411 & n7738 ) | ( ~n7423 & n7738 ) ;
  assign n7740 = ( n7728 & n7737 ) | ( n7728 & n7739 ) | ( n7737 & n7739 ) ;
  assign n7741 = ( ~n7423 & n7432 ) | ( ~n7423 & n7434 ) | ( n7432 & n7434 ) ;
  assign n7742 = ( n7423 & ~n7435 ) | ( n7423 & n7741 ) | ( ~n7435 & n7741 ) ;
  assign n7743 = n5508 & ~n5586 ;
  assign n7744 = ~n2725 & n5507 ;
  assign n7745 = n2843 & n5504 ;
  assign n7746 = ~n2810 & n5666 ;
  assign n7747 = n7745 | n7746 ;
  assign n7748 = ( ~n7743 & n7744 ) | ( ~n7743 & n7747 ) | ( n7744 & n7747 ) ;
  assign n7749 = ( ~x17 & n7743 ) | ( ~x17 & n7748 ) | ( n7743 & n7748 ) ;
  assign n7750 = ( n7743 & n7748 ) | ( n7743 & ~n7749 ) | ( n7748 & ~n7749 ) ;
  assign n7751 = ( x17 & n7749 ) | ( x17 & ~n7750 ) | ( n7749 & ~n7750 ) ;
  assign n7752 = ( n7740 & n7742 ) | ( n7740 & n7751 ) | ( n7742 & n7751 ) ;
  assign n7753 = ( ~n7435 & n7444 ) | ( ~n7435 & n7446 ) | ( n7444 & n7446 ) ;
  assign n7754 = ( n7435 & ~n7447 ) | ( n7435 & n7753 ) | ( ~n7447 & n7753 ) ;
  assign n7755 = n2725 | n5666 ;
  assign n7756 = n2635 & n5507 ;
  assign n7757 = ( ~n2725 & n7755 ) | ( ~n2725 & n7756 ) | ( n7755 & n7756 ) ;
  assign n7758 = ~n2810 & n5504 ;
  assign n7759 = n7757 | n7758 ;
  assign n7760 = n5232 & n5508 ;
  assign n7761 = ( x17 & n7759 ) | ( x17 & ~n7760 ) | ( n7759 & ~n7760 ) ;
  assign n7762 = ( ~x17 & n7759 ) | ( ~x17 & n7760 ) | ( n7759 & n7760 ) ;
  assign n7763 = ( ~n7759 & n7761 ) | ( ~n7759 & n7762 ) | ( n7761 & n7762 ) ;
  assign n7764 = ( n7752 & n7754 ) | ( n7752 & n7763 ) | ( n7754 & n7763 ) ;
  assign n7765 = ~n5425 & n5508 ;
  assign n7766 = n2552 & n5507 ;
  assign n7767 = ~n2725 & n5504 ;
  assign n7768 = n2635 & n5666 ;
  assign n7769 = n7767 | n7768 ;
  assign n7770 = ( ~n7765 & n7766 ) | ( ~n7765 & n7769 ) | ( n7766 & n7769 ) ;
  assign n7771 = ( ~x17 & n7765 ) | ( ~x17 & n7770 ) | ( n7765 & n7770 ) ;
  assign n7772 = ( n7765 & n7770 ) | ( n7765 & ~n7771 ) | ( n7770 & ~n7771 ) ;
  assign n7773 = ( x17 & n7771 ) | ( x17 & ~n7772 ) | ( n7771 & ~n7772 ) ;
  assign n7774 = ( ~n7447 & n7449 ) | ( ~n7447 & n7458 ) | ( n7449 & n7458 ) ;
  assign n7775 = ( n7447 & ~n7459 ) | ( n7447 & n7774 ) | ( ~n7459 & n7774 ) ;
  assign n7776 = ( n7764 & n7773 ) | ( n7764 & n7775 ) | ( n7773 & n7775 ) ;
  assign n7777 = ~n5270 & n5508 ;
  assign n7778 = n2552 & n5666 ;
  assign n7779 = ~n2491 & n5507 ;
  assign n7780 = n2635 & n5504 ;
  assign n7781 = n7779 | n7780 ;
  assign n7782 = ( ~n7777 & n7778 ) | ( ~n7777 & n7781 ) | ( n7778 & n7781 ) ;
  assign n7783 = ( ~x17 & n7777 ) | ( ~x17 & n7782 ) | ( n7777 & n7782 ) ;
  assign n7784 = ( n7777 & n7782 ) | ( n7777 & ~n7783 ) | ( n7782 & ~n7783 ) ;
  assign n7785 = ( x17 & n7783 ) | ( x17 & ~n7784 ) | ( n7783 & ~n7784 ) ;
  assign n7786 = ( ~n7459 & n7461 ) | ( ~n7459 & n7470 ) | ( n7461 & n7470 ) ;
  assign n7787 = ( ~n7470 & n7471 ) | ( ~n7470 & n7786 ) | ( n7471 & n7786 ) ;
  assign n7788 = ( n7776 & n7785 ) | ( n7776 & ~n7787 ) | ( n7785 & ~n7787 ) ;
  assign n7789 = ~n5084 & n5508 ;
  assign n7790 = n2396 & n5507 ;
  assign n7791 = ~n2491 & n5666 ;
  assign n7792 = n2552 & n5504 ;
  assign n7793 = n7791 | n7792 ;
  assign n7794 = ( ~n7789 & n7790 ) | ( ~n7789 & n7793 ) | ( n7790 & n7793 ) ;
  assign n7795 = ( ~x17 & n7789 ) | ( ~x17 & n7794 ) | ( n7789 & n7794 ) ;
  assign n7796 = ( n7789 & n7794 ) | ( n7789 & ~n7795 ) | ( n7794 & ~n7795 ) ;
  assign n7797 = ( x17 & n7795 ) | ( x17 & ~n7796 ) | ( n7795 & ~n7796 ) ;
  assign n7798 = ( ~n7471 & n7473 ) | ( ~n7471 & n7483 ) | ( n7473 & n7483 ) ;
  assign n7799 = ( ~n7483 & n7484 ) | ( ~n7483 & n7798 ) | ( n7484 & n7798 ) ;
  assign n7800 = ( n7788 & n7797 ) | ( n7788 & ~n7799 ) | ( n7797 & ~n7799 ) ;
  assign n7801 = ~n4900 & n5508 ;
  assign n7802 = n2396 & n5666 ;
  assign n7803 = ~n2298 & n5507 ;
  assign n7804 = ~n2491 & n5504 ;
  assign n7805 = n7803 | n7804 ;
  assign n7806 = ( ~n7801 & n7802 ) | ( ~n7801 & n7805 ) | ( n7802 & n7805 ) ;
  assign n7807 = ( ~x17 & n7801 ) | ( ~x17 & n7806 ) | ( n7801 & n7806 ) ;
  assign n7808 = ( n7801 & n7806 ) | ( n7801 & ~n7807 ) | ( n7806 & ~n7807 ) ;
  assign n7809 = ( x17 & n7807 ) | ( x17 & ~n7808 ) | ( n7807 & ~n7808 ) ;
  assign n7810 = ( ~n7484 & n7486 ) | ( ~n7484 & n7495 ) | ( n7486 & n7495 ) ;
  assign n7811 = ( n7484 & ~n7496 ) | ( n7484 & n7810 ) | ( ~n7496 & n7810 ) ;
  assign n7812 = ( n7800 & n7809 ) | ( n7800 & n7811 ) | ( n7809 & n7811 ) ;
  assign n7813 = n2298 | n5666 ;
  assign n7814 = n2270 & n5507 ;
  assign n7815 = ( ~n2298 & n7813 ) | ( ~n2298 & n7814 ) | ( n7813 & n7814 ) ;
  assign n7816 = n2396 & n5504 ;
  assign n7817 = n7815 | n7816 ;
  assign n7818 = ~n4912 & n5508 ;
  assign n7819 = ( x17 & n7817 ) | ( x17 & ~n7818 ) | ( n7817 & ~n7818 ) ;
  assign n7820 = ( ~x17 & n7817 ) | ( ~x17 & n7818 ) | ( n7817 & n7818 ) ;
  assign n7821 = ( ~n7817 & n7819 ) | ( ~n7817 & n7820 ) | ( n7819 & n7820 ) ;
  assign n7822 = ( ~n7496 & n7498 ) | ( ~n7496 & n7507 ) | ( n7498 & n7507 ) ;
  assign n7823 = ( ~n7507 & n7508 ) | ( ~n7507 & n7822 ) | ( n7508 & n7822 ) ;
  assign n7824 = ( n7812 & n7821 ) | ( n7812 & ~n7823 ) | ( n7821 & ~n7823 ) ;
  assign n7825 = n4647 & n5508 ;
  assign n7826 = n2174 & n5507 ;
  assign n7827 = n2298 | n5504 ;
  assign n7828 = n2270 & n5666 ;
  assign n7829 = ( ~n2298 & n7827 ) | ( ~n2298 & n7828 ) | ( n7827 & n7828 ) ;
  assign n7830 = ( ~n7825 & n7826 ) | ( ~n7825 & n7829 ) | ( n7826 & n7829 ) ;
  assign n7831 = ( ~x17 & n7825 ) | ( ~x17 & n7830 ) | ( n7825 & n7830 ) ;
  assign n7832 = ( n7825 & n7830 ) | ( n7825 & ~n7831 ) | ( n7830 & ~n7831 ) ;
  assign n7833 = ( x17 & n7831 ) | ( x17 & ~n7832 ) | ( n7831 & ~n7832 ) ;
  assign n7834 = ( ~n7508 & n7510 ) | ( ~n7508 & n7519 ) | ( n7510 & n7519 ) ;
  assign n7835 = ( n7508 & ~n7520 ) | ( n7508 & n7834 ) | ( ~n7520 & n7834 ) ;
  assign n7836 = ( n7824 & n7833 ) | ( n7824 & n7835 ) | ( n7833 & n7835 ) ;
  assign n7837 = n4730 & n5508 ;
  assign n7838 = n2089 & n5507 ;
  assign n7839 = n2270 & n5504 ;
  assign n7840 = n2174 & n5666 ;
  assign n7841 = n7839 | n7840 ;
  assign n7842 = ( ~n7837 & n7838 ) | ( ~n7837 & n7841 ) | ( n7838 & n7841 ) ;
  assign n7843 = ( ~x17 & n7837 ) | ( ~x17 & n7842 ) | ( n7837 & n7842 ) ;
  assign n7844 = ( n7837 & n7842 ) | ( n7837 & ~n7843 ) | ( n7842 & ~n7843 ) ;
  assign n7845 = ( x17 & n7843 ) | ( x17 & ~n7844 ) | ( n7843 & ~n7844 ) ;
  assign n7846 = ( ~n7520 & n7522 ) | ( ~n7520 & n7531 ) | ( n7522 & n7531 ) ;
  assign n7847 = ( n7520 & ~n7532 ) | ( n7520 & n7846 ) | ( ~n7532 & n7846 ) ;
  assign n7848 = ( n7836 & n7845 ) | ( n7836 & n7847 ) | ( n7845 & n7847 ) ;
  assign n7849 = ( n7532 & ~n7534 ) | ( n7532 & n7543 ) | ( ~n7534 & n7543 ) ;
  assign n7850 = ( n7534 & ~n7544 ) | ( n7534 & n7849 ) | ( ~n7544 & n7849 ) ;
  assign n7851 = ~n4302 & n5966 ;
  assign n7852 = ~n1750 & n6464 ;
  assign n7853 = n1926 & ~n5970 ;
  assign n7854 = n1852 & n5969 ;
  assign n7855 = ( n1926 & ~n7853 ) | ( n1926 & n7854 ) | ( ~n7853 & n7854 ) ;
  assign n7856 = ( ~n7851 & n7852 ) | ( ~n7851 & n7855 ) | ( n7852 & n7855 ) ;
  assign n7857 = ( ~x14 & n7851 ) | ( ~x14 & n7856 ) | ( n7851 & n7856 ) ;
  assign n7858 = ( n7851 & n7856 ) | ( n7851 & ~n7857 ) | ( n7856 & ~n7857 ) ;
  assign n7859 = ( x14 & n7857 ) | ( x14 & ~n7858 ) | ( n7857 & ~n7858 ) ;
  assign n7860 = ( n7848 & n7850 ) | ( n7848 & n7859 ) | ( n7850 & n7859 ) ;
  assign n7861 = ( n7544 & ~n7546 ) | ( n7544 & n7555 ) | ( ~n7546 & n7555 ) ;
  assign n7862 = ( n7546 & ~n7556 ) | ( n7546 & n7861 ) | ( ~n7556 & n7861 ) ;
  assign n7863 = ~n3955 & n6584 ;
  assign n7864 = ~n1338 & n7022 ;
  assign n7865 = n1458 & n6587 ;
  assign n7866 = n1576 & n6588 ;
  assign n7867 = n7865 | n7866 ;
  assign n7868 = ( ~n7863 & n7864 ) | ( ~n7863 & n7867 ) | ( n7864 & n7867 ) ;
  assign n7869 = ( ~x11 & n7863 ) | ( ~x11 & n7868 ) | ( n7863 & n7868 ) ;
  assign n7870 = ( n7863 & n7868 ) | ( n7863 & ~n7869 ) | ( n7868 & ~n7869 ) ;
  assign n7871 = ( x11 & n7869 ) | ( x11 & ~n7870 ) | ( n7869 & ~n7870 ) ;
  assign n7872 = ( n7860 & n7862 ) | ( n7860 & n7871 ) | ( n7862 & n7871 ) ;
  assign n7873 = ( ~n7556 & n7558 ) | ( ~n7556 & n7567 ) | ( n7558 & n7567 ) ;
  assign n7874 = ( ~n7567 & n7568 ) | ( ~n7567 & n7873 ) | ( n7568 & n7873 ) ;
  assign n7875 = ~n3665 & n7296 ;
  assign n7876 = ~n1290 & n7299 ;
  assign n7877 = ~n1246 & n7300 ;
  assign n7878 = ~n7293 & n7294 ;
  assign n7879 = ( ~n7290 & n7291 ) | ( ~n7290 & n7878 ) | ( n7291 & n7878 ) ;
  assign n7880 = ~n3658 & n7879 ;
  assign n7881 = n7877 | n7880 ;
  assign n7882 = ( ~n7875 & n7876 ) | ( ~n7875 & n7881 ) | ( n7876 & n7881 ) ;
  assign n7883 = ( ~x8 & n7875 ) | ( ~x8 & n7882 ) | ( n7875 & n7882 ) ;
  assign n7884 = ( n7875 & n7882 ) | ( n7875 & ~n7883 ) | ( n7882 & ~n7883 ) ;
  assign n7885 = ( x8 & n7883 ) | ( x8 & ~n7884 ) | ( n7883 & ~n7884 ) ;
  assign n7886 = ( n7872 & ~n7874 ) | ( n7872 & n7885 ) | ( ~n7874 & n7885 ) ;
  assign n7887 = n3692 & n7879 ;
  assign n7888 = ~n3658 & n7299 ;
  assign n7889 = ( n7879 & ~n7887 ) | ( n7879 & n7888 ) | ( ~n7887 & n7888 ) ;
  assign n7890 = ~n1290 & n7300 ;
  assign n7891 = n7889 | n7890 ;
  assign n7892 = ~n4182 & n7296 ;
  assign n7893 = ( x8 & n7891 ) | ( x8 & ~n7892 ) | ( n7891 & ~n7892 ) ;
  assign n7894 = ( ~x8 & n7891 ) | ( ~x8 & n7892 ) | ( n7891 & n7892 ) ;
  assign n7895 = ( ~n7891 & n7893 ) | ( ~n7891 & n7894 ) | ( n7893 & n7894 ) ;
  assign n7896 = ( n7568 & ~n7577 ) | ( n7568 & n7579 ) | ( ~n7577 & n7579 ) ;
  assign n7897 = ( n7577 & ~n7580 ) | ( n7577 & n7896 ) | ( ~n7580 & n7896 ) ;
  assign n7898 = ( n7886 & n7895 ) | ( n7886 & n7897 ) | ( n7895 & n7897 ) ;
  assign n7899 = n5966 & n6061 ;
  assign n7900 = n3479 & n5969 ;
  assign n7901 = n3533 | n5970 ;
  assign n7902 = ~n3389 & n6464 ;
  assign n7903 = ( ~n3533 & n7901 ) | ( ~n3533 & n7902 ) | ( n7901 & n7902 ) ;
  assign n7904 = ( ~n7899 & n7900 ) | ( ~n7899 & n7903 ) | ( n7900 & n7903 ) ;
  assign n7905 = ( ~x14 & n7899 ) | ( ~x14 & n7904 ) | ( n7899 & n7904 ) ;
  assign n7906 = ( n7899 & n7904 ) | ( n7899 & ~n7905 ) | ( n7904 & ~n7905 ) ;
  assign n7907 = ( x14 & n7905 ) | ( x14 & ~n7906 ) | ( n7905 & ~n7906 ) ;
  assign n7908 = ( n3479 & n5966 ) | ( n3479 & n6009 ) | ( n5966 & n6009 ) ;
  assign n7909 = ~n3533 & n5969 ;
  assign n7910 = ~n3586 & n5970 ;
  assign n7911 = n7909 | n7910 ;
  assign n7912 = ~n3479 & n6464 ;
  assign n7913 = ( n6464 & n7911 ) | ( n6464 & ~n7912 ) | ( n7911 & ~n7912 ) ;
  assign n7914 = ( ~n6608 & n7908 ) | ( ~n6608 & n7913 ) | ( n7908 & n7913 ) ;
  assign n7915 = ~n3586 & n6463 ;
  assign n7916 = x14 & n7915 ;
  assign n7917 = ( n5966 & n6009 ) | ( n5966 & n6618 ) | ( n6009 & n6618 ) ;
  assign n7918 = ~n3533 & n6464 ;
  assign n7919 = n3586 | n5969 ;
  assign n7920 = ( ~n3586 & n7918 ) | ( ~n3586 & n7919 ) | ( n7918 & n7919 ) ;
  assign n7921 = n7917 | n7920 ;
  assign n7922 = ( x14 & n7916 ) | ( x14 & n7921 ) | ( n7916 & n7921 ) ;
  assign n7923 = n7914 | n7922 ;
  assign n7924 = x14 & ~n7923 ;
  assign n7925 = ( n7607 & n7907 ) | ( n7607 & n7924 ) | ( n7907 & n7924 ) ;
  assign n7926 = n3389 | n5969 ;
  assign n7927 = ~n3355 & n6464 ;
  assign n7928 = ( ~n3389 & n7926 ) | ( ~n3389 & n7927 ) | ( n7926 & n7927 ) ;
  assign n7929 = n3479 & ~n5970 ;
  assign n7930 = ( n3479 & n7928 ) | ( n3479 & ~n7929 ) | ( n7928 & ~n7929 ) ;
  assign n7931 = ( n5966 & ~n6104 ) | ( n5966 & n7930 ) | ( ~n6104 & n7930 ) ;
  assign n7932 = n7930 & ~n7931 ;
  assign n7933 = ( ~x14 & n7931 ) | ( ~x14 & n7932 ) | ( n7931 & n7932 ) ;
  assign n7934 = ( n7931 & n7932 ) | ( n7931 & ~n7933 ) | ( n7932 & ~n7933 ) ;
  assign n7935 = ( x14 & n7933 ) | ( x14 & ~n7934 ) | ( n7933 & ~n7934 ) ;
  assign n7936 = ( n7608 & n7609 ) | ( n7608 & n7612 ) | ( n7609 & n7612 ) ;
  assign n7937 = ~n7608 & n7613 ;
  assign n7938 = ( n7608 & ~n7936 ) | ( n7608 & n7937 ) | ( ~n7936 & n7937 ) ;
  assign n7939 = ( n7925 & n7935 ) | ( n7925 & n7938 ) | ( n7935 & n7938 ) ;
  assign n7940 = n5966 & ~n6154 ;
  assign n7941 = ~n3300 & n6464 ;
  assign n7942 = n3389 | n5970 ;
  assign n7943 = ~n3355 & n5969 ;
  assign n7944 = ( ~n3389 & n7942 ) | ( ~n3389 & n7943 ) | ( n7942 & n7943 ) ;
  assign n7945 = ( ~n7940 & n7941 ) | ( ~n7940 & n7944 ) | ( n7941 & n7944 ) ;
  assign n7946 = ( ~x14 & n7940 ) | ( ~x14 & n7945 ) | ( n7940 & n7945 ) ;
  assign n7947 = ( n7940 & n7945 ) | ( n7940 & ~n7946 ) | ( n7945 & ~n7946 ) ;
  assign n7948 = ( x14 & n7946 ) | ( x14 & ~n7947 ) | ( n7946 & ~n7947 ) ;
  assign n7949 = ( n7606 & n7614 ) | ( n7606 & ~n7615 ) | ( n7614 & ~n7615 ) ;
  assign n7950 = n7615 & ~n7949 ;
  assign n7951 = ( n7939 & n7948 ) | ( n7939 & n7950 ) | ( n7948 & n7950 ) ;
  assign n7952 = n5966 & n6200 ;
  assign n7953 = ~n3300 & n5969 ;
  assign n7954 = n3355 | n5970 ;
  assign n7955 = n3239 & n6464 ;
  assign n7956 = ( ~n3355 & n7954 ) | ( ~n3355 & n7955 ) | ( n7954 & n7955 ) ;
  assign n7957 = ( ~n7952 & n7953 ) | ( ~n7952 & n7956 ) | ( n7953 & n7956 ) ;
  assign n7958 = ( ~x14 & n7952 ) | ( ~x14 & n7957 ) | ( n7952 & n7957 ) ;
  assign n7959 = ( n7952 & n7957 ) | ( n7952 & ~n7958 ) | ( n7957 & ~n7958 ) ;
  assign n7960 = ( x14 & n7958 ) | ( x14 & ~n7959 ) | ( n7958 & ~n7959 ) ;
  assign n7961 = ( n7326 & n7599 ) | ( n7326 & ~n7616 ) | ( n7599 & ~n7616 ) ;
  assign n7962 = ( n7616 & ~n7617 ) | ( n7616 & n7961 ) | ( ~n7617 & n7961 ) ;
  assign n7963 = ( n7951 & n7960 ) | ( n7951 & n7962 ) | ( n7960 & n7962 ) ;
  assign n7964 = n5966 & ~n6243 ;
  assign n7965 = n3153 & n6464 ;
  assign n7966 = n3300 | n5970 ;
  assign n7967 = n3239 & n5969 ;
  assign n7968 = ( ~n3300 & n7966 ) | ( ~n3300 & n7967 ) | ( n7966 & n7967 ) ;
  assign n7969 = ( ~n7964 & n7965 ) | ( ~n7964 & n7968 ) | ( n7965 & n7968 ) ;
  assign n7970 = ( ~x14 & n7964 ) | ( ~x14 & n7969 ) | ( n7964 & n7969 ) ;
  assign n7971 = ( n7964 & n7969 ) | ( n7964 & ~n7970 ) | ( n7969 & ~n7970 ) ;
  assign n7972 = ( x14 & n7970 ) | ( x14 & ~n7971 ) | ( n7970 & ~n7971 ) ;
  assign n7973 = ( ~n7617 & n7627 ) | ( ~n7617 & n7630 ) | ( n7627 & n7630 ) ;
  assign n7974 = ( n7617 & ~n7631 ) | ( n7617 & n7973 ) | ( ~n7631 & n7973 ) ;
  assign n7975 = ( n7963 & n7972 ) | ( n7963 & n7974 ) | ( n7972 & n7974 ) ;
  assign n7976 = ( ~n7631 & n7640 ) | ( ~n7631 & n7642 ) | ( n7640 & n7642 ) ;
  assign n7977 = ( n7631 & ~n7643 ) | ( n7631 & n7976 ) | ( ~n7643 & n7976 ) ;
  assign n7978 = n5710 & n5966 ;
  assign n7979 = n3153 & n5969 ;
  assign n7980 = n3239 & ~n5970 ;
  assign n7981 = n3078 & n6464 ;
  assign n7982 = ( n3239 & ~n7980 ) | ( n3239 & n7981 ) | ( ~n7980 & n7981 ) ;
  assign n7983 = ( ~n7978 & n7979 ) | ( ~n7978 & n7982 ) | ( n7979 & n7982 ) ;
  assign n7984 = ( ~x14 & n7978 ) | ( ~x14 & n7983 ) | ( n7978 & n7983 ) ;
  assign n7985 = ( n7978 & n7983 ) | ( n7978 & ~n7984 ) | ( n7983 & ~n7984 ) ;
  assign n7986 = ( x14 & n7984 ) | ( x14 & ~n7985 ) | ( n7984 & ~n7985 ) ;
  assign n7987 = ( n7975 & n7977 ) | ( n7975 & n7986 ) | ( n7977 & n7986 ) ;
  assign n7988 = ( ~n7643 & n7652 ) | ( ~n7643 & n7654 ) | ( n7652 & n7654 ) ;
  assign n7989 = ( n7643 & ~n7655 ) | ( n7643 & n7988 ) | ( ~n7655 & n7988 ) ;
  assign n7990 = n3078 & ~n5969 ;
  assign n7991 = ~n3046 & n6464 ;
  assign n7992 = ( n3078 & ~n7990 ) | ( n3078 & n7991 ) | ( ~n7990 & n7991 ) ;
  assign n7993 = n3153 & ~n5970 ;
  assign n7994 = ( n3153 & n7992 ) | ( n3153 & ~n7993 ) | ( n7992 & ~n7993 ) ;
  assign n7995 = ( n5966 & ~n6267 ) | ( n5966 & n7994 ) | ( ~n6267 & n7994 ) ;
  assign n7996 = n7994 & ~n7995 ;
  assign n7997 = ( ~x14 & n7995 ) | ( ~x14 & n7996 ) | ( n7995 & n7996 ) ;
  assign n7998 = ( n7995 & n7996 ) | ( n7995 & ~n7997 ) | ( n7996 & ~n7997 ) ;
  assign n7999 = ( x14 & n7997 ) | ( x14 & ~n7998 ) | ( n7997 & ~n7998 ) ;
  assign n8000 = ( n7987 & n7989 ) | ( n7987 & n7999 ) | ( n7989 & n7999 ) ;
  assign n8001 = ( ~n7655 & n7664 ) | ( ~n7655 & n7666 ) | ( n7664 & n7666 ) ;
  assign n8002 = ( n7655 & ~n7667 ) | ( n7655 & n8001 ) | ( ~n7667 & n8001 ) ;
  assign n8003 = n5966 & n6279 ;
  assign n8004 = ~n2965 & n6464 ;
  assign n8005 = n3078 & ~n5970 ;
  assign n8006 = ~n3046 & n5969 ;
  assign n8007 = ( n3078 & ~n8005 ) | ( n3078 & n8006 ) | ( ~n8005 & n8006 ) ;
  assign n8008 = ( ~n8003 & n8004 ) | ( ~n8003 & n8007 ) | ( n8004 & n8007 ) ;
  assign n8009 = ( ~x14 & n8003 ) | ( ~x14 & n8008 ) | ( n8003 & n8008 ) ;
  assign n8010 = ( n8003 & n8008 ) | ( n8003 & ~n8009 ) | ( n8008 & ~n8009 ) ;
  assign n8011 = ( x14 & n8009 ) | ( x14 & ~n8010 ) | ( n8009 & ~n8010 ) ;
  assign n8012 = ( n8000 & n8002 ) | ( n8000 & n8011 ) | ( n8002 & n8011 ) ;
  assign n8013 = ~n5768 & n5966 ;
  assign n8014 = ~n2910 & n6464 ;
  assign n8015 = n3046 | n5970 ;
  assign n8016 = ~n2965 & n5969 ;
  assign n8017 = ( ~n3046 & n8015 ) | ( ~n3046 & n8016 ) | ( n8015 & n8016 ) ;
  assign n8018 = ( ~n8013 & n8014 ) | ( ~n8013 & n8017 ) | ( n8014 & n8017 ) ;
  assign n8019 = ( ~x14 & n8013 ) | ( ~x14 & n8018 ) | ( n8013 & n8018 ) ;
  assign n8020 = ( n8013 & n8018 ) | ( n8013 & ~n8019 ) | ( n8018 & ~n8019 ) ;
  assign n8021 = ( x14 & n8019 ) | ( x14 & ~n8020 ) | ( n8019 & ~n8020 ) ;
  assign n8022 = ( ~n7667 & n7669 ) | ( ~n7667 & n7678 ) | ( n7669 & n7678 ) ;
  assign n8023 = ( n7667 & ~n7679 ) | ( n7667 & n8022 ) | ( ~n7679 & n8022 ) ;
  assign n8024 = ( n8012 & n8021 ) | ( n8012 & n8023 ) | ( n8021 & n8023 ) ;
  assign n8025 = n5543 & n5966 ;
  assign n8026 = ~n2910 & n5969 ;
  assign n8027 = n2965 | n5970 ;
  assign n8028 = n2843 & n6464 ;
  assign n8029 = ( ~n2965 & n8027 ) | ( ~n2965 & n8028 ) | ( n8027 & n8028 ) ;
  assign n8030 = ( ~n8025 & n8026 ) | ( ~n8025 & n8029 ) | ( n8026 & n8029 ) ;
  assign n8031 = ( ~x14 & n8025 ) | ( ~x14 & n8030 ) | ( n8025 & n8030 ) ;
  assign n8032 = ( n8025 & n8030 ) | ( n8025 & ~n8031 ) | ( n8030 & ~n8031 ) ;
  assign n8033 = ( x14 & n8031 ) | ( x14 & ~n8032 ) | ( n8031 & ~n8032 ) ;
  assign n8034 = ( ~n7679 & n7681 ) | ( ~n7679 & n7691 ) | ( n7681 & n7691 ) ;
  assign n8035 = ( n7679 & ~n7692 ) | ( n7679 & n8034 ) | ( ~n7692 & n8034 ) ;
  assign n8036 = ( n8024 & n8033 ) | ( n8024 & n8035 ) | ( n8033 & n8035 ) ;
  assign n8037 = n5791 & n5966 ;
  assign n8038 = ~n2810 & n6464 ;
  assign n8039 = n2910 | n5970 ;
  assign n8040 = n2843 & n5969 ;
  assign n8041 = ( ~n2910 & n8039 ) | ( ~n2910 & n8040 ) | ( n8039 & n8040 ) ;
  assign n8042 = ( ~n8037 & n8038 ) | ( ~n8037 & n8041 ) | ( n8038 & n8041 ) ;
  assign n8043 = ( ~x14 & n8037 ) | ( ~x14 & n8042 ) | ( n8037 & n8042 ) ;
  assign n8044 = ( n8037 & n8042 ) | ( n8037 & ~n8043 ) | ( n8042 & ~n8043 ) ;
  assign n8045 = ( x14 & n8043 ) | ( x14 & ~n8044 ) | ( n8043 & ~n8044 ) ;
  assign n8046 = ( ~n7692 & n7694 ) | ( ~n7692 & n7703 ) | ( n7694 & n7703 ) ;
  assign n8047 = ( n7692 & ~n7704 ) | ( n7692 & n8046 ) | ( ~n7704 & n8046 ) ;
  assign n8048 = ( n8036 & n8045 ) | ( n8036 & n8047 ) | ( n8045 & n8047 ) ;
  assign n8049 = ( ~n7704 & n7713 ) | ( ~n7704 & n7715 ) | ( n7713 & n7715 ) ;
  assign n8050 = ( n7704 & ~n7716 ) | ( n7704 & n8049 ) | ( ~n7716 & n8049 ) ;
  assign n8051 = ~n5586 & n5966 ;
  assign n8052 = ~n2725 & n6464 ;
  assign n8053 = n2843 & ~n5970 ;
  assign n8054 = ~n2810 & n5969 ;
  assign n8055 = ( n2843 & ~n8053 ) | ( n2843 & n8054 ) | ( ~n8053 & n8054 ) ;
  assign n8056 = ( ~n8051 & n8052 ) | ( ~n8051 & n8055 ) | ( n8052 & n8055 ) ;
  assign n8057 = ( ~x14 & n8051 ) | ( ~x14 & n8056 ) | ( n8051 & n8056 ) ;
  assign n8058 = ( n8051 & n8056 ) | ( n8051 & ~n8057 ) | ( n8056 & ~n8057 ) ;
  assign n8059 = ( x14 & n8057 ) | ( x14 & ~n8058 ) | ( n8057 & ~n8058 ) ;
  assign n8060 = ( n8048 & n8050 ) | ( n8048 & n8059 ) | ( n8050 & n8059 ) ;
  assign n8061 = ( ~n7716 & n7725 ) | ( ~n7716 & n7727 ) | ( n7725 & n7727 ) ;
  assign n8062 = ( n7716 & ~n7728 ) | ( n7716 & n8061 ) | ( ~n7728 & n8061 ) ;
  assign n8063 = n2725 | n5969 ;
  assign n8064 = n2635 & n6464 ;
  assign n8065 = ( ~n2725 & n8063 ) | ( ~n2725 & n8064 ) | ( n8063 & n8064 ) ;
  assign n8066 = ~n2810 & n5970 ;
  assign n8067 = n8065 | n8066 ;
  assign n8068 = n5232 & n5966 ;
  assign n8069 = ( x14 & n8067 ) | ( x14 & ~n8068 ) | ( n8067 & ~n8068 ) ;
  assign n8070 = ( ~x14 & n8067 ) | ( ~x14 & n8068 ) | ( n8067 & n8068 ) ;
  assign n8071 = ( ~n8067 & n8069 ) | ( ~n8067 & n8070 ) | ( n8069 & n8070 ) ;
  assign n8072 = ( n8060 & n8062 ) | ( n8060 & n8071 ) | ( n8062 & n8071 ) ;
  assign n8073 = ( ~n7728 & n7737 ) | ( ~n7728 & n7739 ) | ( n7737 & n7739 ) ;
  assign n8074 = ( n7728 & ~n7740 ) | ( n7728 & n8073 ) | ( ~n7740 & n8073 ) ;
  assign n8075 = ~n5425 & n5966 ;
  assign n8076 = n2552 & n6464 ;
  assign n8077 = n2725 | n5970 ;
  assign n8078 = n2635 & n5969 ;
  assign n8079 = ( ~n2725 & n8077 ) | ( ~n2725 & n8078 ) | ( n8077 & n8078 ) ;
  assign n8080 = ( ~n8075 & n8076 ) | ( ~n8075 & n8079 ) | ( n8076 & n8079 ) ;
  assign n8081 = ( ~x14 & n8075 ) | ( ~x14 & n8080 ) | ( n8075 & n8080 ) ;
  assign n8082 = ( n8075 & n8080 ) | ( n8075 & ~n8081 ) | ( n8080 & ~n8081 ) ;
  assign n8083 = ( x14 & n8081 ) | ( x14 & ~n8082 ) | ( n8081 & ~n8082 ) ;
  assign n8084 = ( n8072 & n8074 ) | ( n8072 & n8083 ) | ( n8074 & n8083 ) ;
  assign n8085 = ~n5270 & n5966 ;
  assign n8086 = n2552 & n5969 ;
  assign n8087 = n2635 & ~n5970 ;
  assign n8088 = ~n2491 & n6464 ;
  assign n8089 = ( n2635 & ~n8087 ) | ( n2635 & n8088 ) | ( ~n8087 & n8088 ) ;
  assign n8090 = ( ~n8085 & n8086 ) | ( ~n8085 & n8089 ) | ( n8086 & n8089 ) ;
  assign n8091 = ( ~x14 & n8085 ) | ( ~x14 & n8090 ) | ( n8085 & n8090 ) ;
  assign n8092 = ( n8085 & n8090 ) | ( n8085 & ~n8091 ) | ( n8090 & ~n8091 ) ;
  assign n8093 = ( x14 & n8091 ) | ( x14 & ~n8092 ) | ( n8091 & ~n8092 ) ;
  assign n8094 = ( ~n7740 & n7742 ) | ( ~n7740 & n7751 ) | ( n7742 & n7751 ) ;
  assign n8095 = ( n7740 & ~n7752 ) | ( n7740 & n8094 ) | ( ~n7752 & n8094 ) ;
  assign n8096 = ( n8084 & n8093 ) | ( n8084 & n8095 ) | ( n8093 & n8095 ) ;
  assign n8097 = ~n5084 & n5966 ;
  assign n8098 = n2396 & n6464 ;
  assign n8099 = n2552 & ~n5970 ;
  assign n8100 = ~n2491 & n5969 ;
  assign n8101 = ( n2552 & ~n8099 ) | ( n2552 & n8100 ) | ( ~n8099 & n8100 ) ;
  assign n8102 = ( ~n8097 & n8098 ) | ( ~n8097 & n8101 ) | ( n8098 & n8101 ) ;
  assign n8103 = ( ~x14 & n8097 ) | ( ~x14 & n8102 ) | ( n8097 & n8102 ) ;
  assign n8104 = ( n8097 & n8102 ) | ( n8097 & ~n8103 ) | ( n8102 & ~n8103 ) ;
  assign n8105 = ( x14 & n8103 ) | ( x14 & ~n8104 ) | ( n8103 & ~n8104 ) ;
  assign n8106 = ( ~n7752 & n7754 ) | ( ~n7752 & n7763 ) | ( n7754 & n7763 ) ;
  assign n8107 = ( n7752 & ~n7764 ) | ( n7752 & n8106 ) | ( ~n7764 & n8106 ) ;
  assign n8108 = ( n8096 & n8105 ) | ( n8096 & n8107 ) | ( n8105 & n8107 ) ;
  assign n8109 = ( ~n7764 & n7773 ) | ( ~n7764 & n7775 ) | ( n7773 & n7775 ) ;
  assign n8110 = ( n7764 & ~n7776 ) | ( n7764 & n8109 ) | ( ~n7776 & n8109 ) ;
  assign n8111 = ~n4900 & n5966 ;
  assign n8112 = n2396 & n5969 ;
  assign n8113 = ~n2298 & n6464 ;
  assign n8114 = ~n2491 & n5970 ;
  assign n8115 = n8113 | n8114 ;
  assign n8116 = ( ~n8111 & n8112 ) | ( ~n8111 & n8115 ) | ( n8112 & n8115 ) ;
  assign n8117 = ( ~x14 & n8111 ) | ( ~x14 & n8116 ) | ( n8111 & n8116 ) ;
  assign n8118 = ( n8111 & n8116 ) | ( n8111 & ~n8117 ) | ( n8116 & ~n8117 ) ;
  assign n8119 = ( x14 & n8117 ) | ( x14 & ~n8118 ) | ( n8117 & ~n8118 ) ;
  assign n8120 = ( n8108 & n8110 ) | ( n8108 & n8119 ) | ( n8110 & n8119 ) ;
  assign n8121 = ( n7776 & ~n7785 ) | ( n7776 & n7787 ) | ( ~n7785 & n7787 ) ;
  assign n8122 = ( ~n7776 & n7788 ) | ( ~n7776 & n8121 ) | ( n7788 & n8121 ) ;
  assign n8123 = n2298 | n5969 ;
  assign n8124 = n2270 & n6464 ;
  assign n8125 = ( ~n2298 & n8123 ) | ( ~n2298 & n8124 ) | ( n8123 & n8124 ) ;
  assign n8126 = n2396 & n5970 ;
  assign n8127 = n8125 | n8126 ;
  assign n8128 = ~n4912 & n5966 ;
  assign n8129 = ( x14 & n8127 ) | ( x14 & ~n8128 ) | ( n8127 & ~n8128 ) ;
  assign n8130 = ( ~x14 & n8127 ) | ( ~x14 & n8128 ) | ( n8127 & n8128 ) ;
  assign n8131 = ( ~n8127 & n8129 ) | ( ~n8127 & n8130 ) | ( n8129 & n8130 ) ;
  assign n8132 = ( n8120 & ~n8122 ) | ( n8120 & n8131 ) | ( ~n8122 & n8131 ) ;
  assign n8133 = ( n7788 & ~n7797 ) | ( n7788 & n7799 ) | ( ~n7797 & n7799 ) ;
  assign n8134 = ( ~n7788 & n7800 ) | ( ~n7788 & n8133 ) | ( n7800 & n8133 ) ;
  assign n8135 = n4647 & n5966 ;
  assign n8136 = n2174 & n6464 ;
  assign n8137 = n2298 | n5970 ;
  assign n8138 = n2270 & n5969 ;
  assign n8139 = ( ~n2298 & n8137 ) | ( ~n2298 & n8138 ) | ( n8137 & n8138 ) ;
  assign n8140 = ( ~n8135 & n8136 ) | ( ~n8135 & n8139 ) | ( n8136 & n8139 ) ;
  assign n8141 = ( ~x14 & n8135 ) | ( ~x14 & n8140 ) | ( n8135 & n8140 ) ;
  assign n8142 = ( n8135 & n8140 ) | ( n8135 & ~n8141 ) | ( n8140 & ~n8141 ) ;
  assign n8143 = ( x14 & n8141 ) | ( x14 & ~n8142 ) | ( n8141 & ~n8142 ) ;
  assign n8144 = ( n8132 & ~n8134 ) | ( n8132 & n8143 ) | ( ~n8134 & n8143 ) ;
  assign n8145 = ( ~n7800 & n7809 ) | ( ~n7800 & n7811 ) | ( n7809 & n7811 ) ;
  assign n8146 = ( n7800 & ~n7812 ) | ( n7800 & n8145 ) | ( ~n7812 & n8145 ) ;
  assign n8147 = n4730 & n5966 ;
  assign n8148 = n2089 & n6464 ;
  assign n8149 = n2270 & ~n5970 ;
  assign n8150 = n2174 & n5969 ;
  assign n8151 = ( n2270 & ~n8149 ) | ( n2270 & n8150 ) | ( ~n8149 & n8150 ) ;
  assign n8152 = ( ~n8147 & n8148 ) | ( ~n8147 & n8151 ) | ( n8148 & n8151 ) ;
  assign n8153 = ( ~x14 & n8147 ) | ( ~x14 & n8152 ) | ( n8147 & n8152 ) ;
  assign n8154 = ( n8147 & n8152 ) | ( n8147 & ~n8153 ) | ( n8152 & ~n8153 ) ;
  assign n8155 = ( x14 & n8153 ) | ( x14 & ~n8154 ) | ( n8153 & ~n8154 ) ;
  assign n8156 = ( n8144 & n8146 ) | ( n8144 & n8155 ) | ( n8146 & n8155 ) ;
  assign n8157 = ( n7812 & ~n7821 ) | ( n7812 & n7823 ) | ( ~n7821 & n7823 ) ;
  assign n8158 = ( ~n7812 & n7824 ) | ( ~n7812 & n8157 ) | ( n7824 & n8157 ) ;
  assign n8159 = ~n4660 & n5966 ;
  assign n8160 = ~n2023 & n6464 ;
  assign n8161 = n2174 & ~n5970 ;
  assign n8162 = n2089 & n5969 ;
  assign n8163 = ( n2174 & ~n8161 ) | ( n2174 & n8162 ) | ( ~n8161 & n8162 ) ;
  assign n8164 = ( ~n8159 & n8160 ) | ( ~n8159 & n8163 ) | ( n8160 & n8163 ) ;
  assign n8165 = ( ~x14 & n8159 ) | ( ~x14 & n8164 ) | ( n8159 & n8164 ) ;
  assign n8166 = ( n8159 & n8164 ) | ( n8159 & ~n8165 ) | ( n8164 & ~n8165 ) ;
  assign n8167 = ( x14 & n8165 ) | ( x14 & ~n8166 ) | ( n8165 & ~n8166 ) ;
  assign n8168 = ( n8156 & ~n8158 ) | ( n8156 & n8167 ) | ( ~n8158 & n8167 ) ;
  assign n8169 = ( ~n7824 & n7833 ) | ( ~n7824 & n7835 ) | ( n7833 & n7835 ) ;
  assign n8170 = ( n7824 & ~n7836 ) | ( n7824 & n8169 ) | ( ~n7836 & n8169 ) ;
  assign n8171 = ~n4457 & n5966 ;
  assign n8172 = n1926 & n6464 ;
  assign n8173 = n2089 & ~n5970 ;
  assign n8174 = ~n2023 & n5969 ;
  assign n8175 = ( n2089 & ~n8173 ) | ( n2089 & n8174 ) | ( ~n8173 & n8174 ) ;
  assign n8176 = ( ~n8171 & n8172 ) | ( ~n8171 & n8175 ) | ( n8172 & n8175 ) ;
  assign n8177 = ( ~x14 & n8171 ) | ( ~x14 & n8176 ) | ( n8171 & n8176 ) ;
  assign n8178 = ( n8171 & n8176 ) | ( n8171 & ~n8177 ) | ( n8176 & ~n8177 ) ;
  assign n8179 = ( x14 & n8177 ) | ( x14 & ~n8178 ) | ( n8177 & ~n8178 ) ;
  assign n8180 = ( n8168 & n8170 ) | ( n8168 & n8179 ) | ( n8170 & n8179 ) ;
  assign n8181 = ( ~n7836 & n7845 ) | ( ~n7836 & n7847 ) | ( n7845 & n7847 ) ;
  assign n8182 = ( n7836 & ~n7848 ) | ( n7836 & n8181 ) | ( ~n7848 & n8181 ) ;
  assign n8183 = n4290 & n5966 ;
  assign n8184 = n1852 & n6464 ;
  assign n8185 = n2023 | n5970 ;
  assign n8186 = n1926 & n5969 ;
  assign n8187 = ( ~n2023 & n8185 ) | ( ~n2023 & n8186 ) | ( n8185 & n8186 ) ;
  assign n8188 = ( ~n8183 & n8184 ) | ( ~n8183 & n8187 ) | ( n8184 & n8187 ) ;
  assign n8189 = ( ~x14 & n8183 ) | ( ~x14 & n8188 ) | ( n8183 & n8188 ) ;
  assign n8190 = ( n8183 & n8188 ) | ( n8183 & ~n8189 ) | ( n8188 & ~n8189 ) ;
  assign n8191 = ( x14 & n8189 ) | ( x14 & ~n8190 ) | ( n8189 & ~n8190 ) ;
  assign n8192 = ( n8180 & n8182 ) | ( n8180 & n8191 ) | ( n8182 & n8191 ) ;
  assign n8193 = ( n7848 & ~n7850 ) | ( n7848 & n7859 ) | ( ~n7850 & n7859 ) ;
  assign n8194 = ( n7850 & ~n7860 ) | ( n7850 & n8193 ) | ( ~n7860 & n8193 ) ;
  assign n8195 = ~n4159 & n6584 ;
  assign n8196 = n1458 & n7022 ;
  assign n8197 = n1669 | n6588 ;
  assign n8198 = n1576 & n6587 ;
  assign n8199 = ( ~n1669 & n8197 ) | ( ~n1669 & n8198 ) | ( n8197 & n8198 ) ;
  assign n8200 = ( ~n8195 & n8196 ) | ( ~n8195 & n8199 ) | ( n8196 & n8199 ) ;
  assign n8201 = ( ~x11 & n8195 ) | ( ~x11 & n8200 ) | ( n8195 & n8200 ) ;
  assign n8202 = ( n8195 & n8200 ) | ( n8195 & ~n8201 ) | ( n8200 & ~n8201 ) ;
  assign n8203 = ( x11 & n8201 ) | ( x11 & ~n8202 ) | ( n8201 & ~n8202 ) ;
  assign n8204 = ( n8192 & n8194 ) | ( n8192 & n8203 ) | ( n8194 & n8203 ) ;
  assign n8205 = ( n7860 & ~n7862 ) | ( n7860 & n7871 ) | ( ~n7862 & n7871 ) ;
  assign n8206 = ( n7862 & ~n7872 ) | ( n7862 & n8205 ) | ( ~n7872 & n8205 ) ;
  assign n8207 = n3621 & n7296 ;
  assign n8208 = ~n1290 & n7879 ;
  assign n8209 = n1267 & ~n7300 ;
  assign n8210 = ~n1246 & n7299 ;
  assign n8211 = ( n1267 & ~n8209 ) | ( n1267 & n8210 ) | ( ~n8209 & n8210 ) ;
  assign n8212 = ( ~n8207 & n8208 ) | ( ~n8207 & n8211 ) | ( n8208 & n8211 ) ;
  assign n8213 = ( ~x8 & n8207 ) | ( ~x8 & n8212 ) | ( n8207 & n8212 ) ;
  assign n8214 = ( n8207 & n8212 ) | ( n8207 & ~n8213 ) | ( n8212 & ~n8213 ) ;
  assign n8215 = ( x8 & n8213 ) | ( x8 & ~n8214 ) | ( n8213 & ~n8214 ) ;
  assign n8216 = ( n8204 & n8206 ) | ( n8204 & n8215 ) | ( n8206 & n8215 ) ;
  assign n8217 = x2 | x3 ;
  assign n8218 = x2 & x3 ;
  assign n8219 = x4 | x5 ;
  assign n8220 = x4 & x5 ;
  assign n8221 = n8219 & ~n8220 ;
  assign n8222 = ( ~n8217 & n8218 ) | ( ~n8217 & n8221 ) | ( n8218 & n8221 ) ;
  assign n8223 = x3 | x4 ;
  assign n8224 = x2 & ~x4 ;
  assign n8225 = ( ~n8217 & n8223 ) | ( ~n8217 & n8224 ) | ( n8223 & n8224 ) ;
  assign n8226 = n8222 & ~n8225 ;
  assign n8227 = ~n3692 & n8226 ;
  assign n8228 = n8217 & ~n8218 ;
  assign n8229 = ( ~n8219 & n8220 ) | ( ~n8219 & n8228 ) | ( n8220 & n8228 ) ;
  assign n8230 = n8228 & ~n8229 ;
  assign n8231 = ~n3691 & n8230 ;
  assign n8232 = ( ~n3692 & n8227 ) | ( ~n3692 & n8231 ) | ( n8227 & n8231 ) ;
  assign n8233 = x5 | n8232 ;
  assign n8234 = ( x5 & n8232 ) | ( x5 & ~n8233 ) | ( n8232 & ~n8233 ) ;
  assign n8235 = n8233 & ~n8234 ;
  assign n8236 = ( ~n7872 & n7874 ) | ( ~n7872 & n7885 ) | ( n7874 & n7885 ) ;
  assign n8237 = ( ~n7885 & n7886 ) | ( ~n7885 & n8236 ) | ( n7886 & n8236 ) ;
  assign n8238 = ( n8216 & n8235 ) | ( n8216 & ~n8237 ) | ( n8235 & ~n8237 ) ;
  assign n8239 = n6061 & n6584 ;
  assign n8240 = n3479 & n6587 ;
  assign n8241 = n3533 | n6588 ;
  assign n8242 = ~n3389 & n7022 ;
  assign n8243 = ( ~n3533 & n8241 ) | ( ~n3533 & n8242 ) | ( n8241 & n8242 ) ;
  assign n8244 = ( ~n8239 & n8240 ) | ( ~n8239 & n8243 ) | ( n8240 & n8243 ) ;
  assign n8245 = ( ~x11 & n8239 ) | ( ~x11 & n8244 ) | ( n8239 & n8244 ) ;
  assign n8246 = ( n8239 & n8244 ) | ( n8239 & ~n8245 ) | ( n8244 & ~n8245 ) ;
  assign n8247 = ( x11 & n8245 ) | ( x11 & ~n8246 ) | ( n8245 & ~n8246 ) ;
  assign n8248 = ( n3479 & n6009 ) | ( n3479 & n6584 ) | ( n6009 & n6584 ) ;
  assign n8249 = ~n3533 & n6587 ;
  assign n8250 = ~n3586 & n6588 ;
  assign n8251 = n8249 | n8250 ;
  assign n8252 = ~n3479 & n7022 ;
  assign n8253 = ( n7022 & n8251 ) | ( n7022 & ~n8252 ) | ( n8251 & ~n8252 ) ;
  assign n8254 = ( ~n6608 & n8248 ) | ( ~n6608 & n8253 ) | ( n8248 & n8253 ) ;
  assign n8255 = ~n3586 & n7021 ;
  assign n8256 = x11 & n8255 ;
  assign n8257 = ( n6009 & n6584 ) | ( n6009 & n6618 ) | ( n6584 & n6618 ) ;
  assign n8258 = ~n3533 & n7022 ;
  assign n8259 = n3586 | n6587 ;
  assign n8260 = ( ~n3586 & n8258 ) | ( ~n3586 & n8259 ) | ( n8258 & n8259 ) ;
  assign n8261 = n8257 | n8260 ;
  assign n8262 = ( x11 & n8256 ) | ( x11 & n8261 ) | ( n8256 & n8261 ) ;
  assign n8263 = n8254 | n8262 ;
  assign n8264 = x11 & ~n8263 ;
  assign n8265 = ( n7915 & n8247 ) | ( n7915 & n8264 ) | ( n8247 & n8264 ) ;
  assign n8266 = n3389 | n6587 ;
  assign n8267 = ~n3355 & n7022 ;
  assign n8268 = ( ~n3389 & n8266 ) | ( ~n3389 & n8267 ) | ( n8266 & n8267 ) ;
  assign n8269 = n3479 & n6588 ;
  assign n8270 = n8268 | n8269 ;
  assign n8271 = ~n6104 & n6584 ;
  assign n8272 = ( x11 & n8270 ) | ( x11 & ~n8271 ) | ( n8270 & ~n8271 ) ;
  assign n8273 = ( ~x11 & n8270 ) | ( ~x11 & n8271 ) | ( n8270 & n8271 ) ;
  assign n8274 = ( ~n8270 & n8272 ) | ( ~n8270 & n8273 ) | ( n8272 & n8273 ) ;
  assign n8275 = ( n7916 & n7917 ) | ( n7916 & n7920 ) | ( n7917 & n7920 ) ;
  assign n8276 = ~n7916 & n7921 ;
  assign n8277 = ( n7916 & ~n8275 ) | ( n7916 & n8276 ) | ( ~n8275 & n8276 ) ;
  assign n8278 = ( n8265 & n8274 ) | ( n8265 & n8277 ) | ( n8274 & n8277 ) ;
  assign n8279 = ~n6154 & n6584 ;
  assign n8280 = ~n3300 & n7022 ;
  assign n8281 = n3389 | n6588 ;
  assign n8282 = ~n3355 & n6587 ;
  assign n8283 = ( ~n3389 & n8281 ) | ( ~n3389 & n8282 ) | ( n8281 & n8282 ) ;
  assign n8284 = ( ~n8279 & n8280 ) | ( ~n8279 & n8283 ) | ( n8280 & n8283 ) ;
  assign n8285 = ( ~x11 & n8279 ) | ( ~x11 & n8284 ) | ( n8279 & n8284 ) ;
  assign n8286 = ( n8279 & n8284 ) | ( n8279 & ~n8285 ) | ( n8284 & ~n8285 ) ;
  assign n8287 = ( x11 & n8285 ) | ( x11 & ~n8286 ) | ( n8285 & ~n8286 ) ;
  assign n8288 = ( n7914 & n7922 ) | ( n7914 & ~n7923 ) | ( n7922 & ~n7923 ) ;
  assign n8289 = n7923 & ~n8288 ;
  assign n8290 = ( n8278 & n8287 ) | ( n8278 & n8289 ) | ( n8287 & n8289 ) ;
  assign n8291 = n6200 & n6584 ;
  assign n8292 = ~n3300 & n6587 ;
  assign n8293 = n3355 | n6588 ;
  assign n8294 = n3239 & n7022 ;
  assign n8295 = ( ~n3355 & n8293 ) | ( ~n3355 & n8294 ) | ( n8293 & n8294 ) ;
  assign n8296 = ( ~n8291 & n8292 ) | ( ~n8291 & n8295 ) | ( n8292 & n8295 ) ;
  assign n8297 = ( ~x11 & n8291 ) | ( ~x11 & n8296 ) | ( n8291 & n8296 ) ;
  assign n8298 = ( n8291 & n8296 ) | ( n8291 & ~n8297 ) | ( n8296 & ~n8297 ) ;
  assign n8299 = ( x11 & n8297 ) | ( x11 & ~n8298 ) | ( n8297 & ~n8298 ) ;
  assign n8300 = ( n7607 & n7907 ) | ( n7607 & ~n7924 ) | ( n7907 & ~n7924 ) ;
  assign n8301 = ( n7924 & ~n7925 ) | ( n7924 & n8300 ) | ( ~n7925 & n8300 ) ;
  assign n8302 = ( n8290 & n8299 ) | ( n8290 & n8301 ) | ( n8299 & n8301 ) ;
  assign n8303 = ~n6243 & n6584 ;
  assign n8304 = n3153 & n7022 ;
  assign n8305 = n3300 | n6588 ;
  assign n8306 = n3239 & n6587 ;
  assign n8307 = ( ~n3300 & n8305 ) | ( ~n3300 & n8306 ) | ( n8305 & n8306 ) ;
  assign n8308 = ( ~n8303 & n8304 ) | ( ~n8303 & n8307 ) | ( n8304 & n8307 ) ;
  assign n8309 = ( ~x11 & n8303 ) | ( ~x11 & n8308 ) | ( n8303 & n8308 ) ;
  assign n8310 = ( n8303 & n8308 ) | ( n8303 & ~n8309 ) | ( n8308 & ~n8309 ) ;
  assign n8311 = ( x11 & n8309 ) | ( x11 & ~n8310 ) | ( n8309 & ~n8310 ) ;
  assign n8312 = ( ~n7925 & n7935 ) | ( ~n7925 & n7938 ) | ( n7935 & n7938 ) ;
  assign n8313 = ( n7925 & ~n7939 ) | ( n7925 & n8312 ) | ( ~n7939 & n8312 ) ;
  assign n8314 = ( n8302 & n8311 ) | ( n8302 & n8313 ) | ( n8311 & n8313 ) ;
  assign n8315 = ( ~n7939 & n7948 ) | ( ~n7939 & n7950 ) | ( n7948 & n7950 ) ;
  assign n8316 = ( n7939 & ~n7951 ) | ( n7939 & n8315 ) | ( ~n7951 & n8315 ) ;
  assign n8317 = n5710 & n6584 ;
  assign n8318 = n3153 & n6587 ;
  assign n8319 = n3239 & ~n6588 ;
  assign n8320 = n3078 & n7022 ;
  assign n8321 = ( n3239 & ~n8319 ) | ( n3239 & n8320 ) | ( ~n8319 & n8320 ) ;
  assign n8322 = ( ~n8317 & n8318 ) | ( ~n8317 & n8321 ) | ( n8318 & n8321 ) ;
  assign n8323 = ( ~x11 & n8317 ) | ( ~x11 & n8322 ) | ( n8317 & n8322 ) ;
  assign n8324 = ( n8317 & n8322 ) | ( n8317 & ~n8323 ) | ( n8322 & ~n8323 ) ;
  assign n8325 = ( x11 & n8323 ) | ( x11 & ~n8324 ) | ( n8323 & ~n8324 ) ;
  assign n8326 = ( n8314 & n8316 ) | ( n8314 & n8325 ) | ( n8316 & n8325 ) ;
  assign n8327 = ( ~n7951 & n7960 ) | ( ~n7951 & n7962 ) | ( n7960 & n7962 ) ;
  assign n8328 = ( n7951 & ~n7963 ) | ( n7951 & n8327 ) | ( ~n7963 & n8327 ) ;
  assign n8329 = n3078 & ~n6587 ;
  assign n8330 = ~n3046 & n7022 ;
  assign n8331 = ( n3078 & ~n8329 ) | ( n3078 & n8330 ) | ( ~n8329 & n8330 ) ;
  assign n8332 = n3153 & n6588 ;
  assign n8333 = n8331 | n8332 ;
  assign n8334 = ~n6267 & n6584 ;
  assign n8335 = ( x11 & n8333 ) | ( x11 & ~n8334 ) | ( n8333 & ~n8334 ) ;
  assign n8336 = ( ~x11 & n8333 ) | ( ~x11 & n8334 ) | ( n8333 & n8334 ) ;
  assign n8337 = ( ~n8333 & n8335 ) | ( ~n8333 & n8336 ) | ( n8335 & n8336 ) ;
  assign n8338 = ( n8326 & n8328 ) | ( n8326 & n8337 ) | ( n8328 & n8337 ) ;
  assign n8339 = ( ~n7963 & n7972 ) | ( ~n7963 & n7974 ) | ( n7972 & n7974 ) ;
  assign n8340 = ( n7963 & ~n7975 ) | ( n7963 & n8339 ) | ( ~n7975 & n8339 ) ;
  assign n8341 = n6279 & n6584 ;
  assign n8342 = ~n2965 & n7022 ;
  assign n8343 = n3078 & ~n6588 ;
  assign n8344 = ~n3046 & n6587 ;
  assign n8345 = ( n3078 & ~n8343 ) | ( n3078 & n8344 ) | ( ~n8343 & n8344 ) ;
  assign n8346 = ( ~n8341 & n8342 ) | ( ~n8341 & n8345 ) | ( n8342 & n8345 ) ;
  assign n8347 = ( ~x11 & n8341 ) | ( ~x11 & n8346 ) | ( n8341 & n8346 ) ;
  assign n8348 = ( n8341 & n8346 ) | ( n8341 & ~n8347 ) | ( n8346 & ~n8347 ) ;
  assign n8349 = ( x11 & n8347 ) | ( x11 & ~n8348 ) | ( n8347 & ~n8348 ) ;
  assign n8350 = ( n8338 & n8340 ) | ( n8338 & n8349 ) | ( n8340 & n8349 ) ;
  assign n8351 = ~n5768 & n6584 ;
  assign n8352 = ~n2910 & n7022 ;
  assign n8353 = n3046 | n6588 ;
  assign n8354 = ~n2965 & n6587 ;
  assign n8355 = ( ~n3046 & n8353 ) | ( ~n3046 & n8354 ) | ( n8353 & n8354 ) ;
  assign n8356 = ( ~n8351 & n8352 ) | ( ~n8351 & n8355 ) | ( n8352 & n8355 ) ;
  assign n8357 = ( ~x11 & n8351 ) | ( ~x11 & n8356 ) | ( n8351 & n8356 ) ;
  assign n8358 = ( n8351 & n8356 ) | ( n8351 & ~n8357 ) | ( n8356 & ~n8357 ) ;
  assign n8359 = ( x11 & n8357 ) | ( x11 & ~n8358 ) | ( n8357 & ~n8358 ) ;
  assign n8360 = ( ~n7975 & n7977 ) | ( ~n7975 & n7986 ) | ( n7977 & n7986 ) ;
  assign n8361 = ( n7975 & ~n7987 ) | ( n7975 & n8360 ) | ( ~n7987 & n8360 ) ;
  assign n8362 = ( n8350 & n8359 ) | ( n8350 & n8361 ) | ( n8359 & n8361 ) ;
  assign n8363 = n5543 & n6584 ;
  assign n8364 = ~n2910 & n6587 ;
  assign n8365 = n2965 | n6588 ;
  assign n8366 = n2843 & n7022 ;
  assign n8367 = ( ~n2965 & n8365 ) | ( ~n2965 & n8366 ) | ( n8365 & n8366 ) ;
  assign n8368 = ( ~n8363 & n8364 ) | ( ~n8363 & n8367 ) | ( n8364 & n8367 ) ;
  assign n8369 = ( ~x11 & n8363 ) | ( ~x11 & n8368 ) | ( n8363 & n8368 ) ;
  assign n8370 = ( n8363 & n8368 ) | ( n8363 & ~n8369 ) | ( n8368 & ~n8369 ) ;
  assign n8371 = ( x11 & n8369 ) | ( x11 & ~n8370 ) | ( n8369 & ~n8370 ) ;
  assign n8372 = ( ~n7987 & n7989 ) | ( ~n7987 & n7999 ) | ( n7989 & n7999 ) ;
  assign n8373 = ( n7987 & ~n8000 ) | ( n7987 & n8372 ) | ( ~n8000 & n8372 ) ;
  assign n8374 = ( n8362 & n8371 ) | ( n8362 & n8373 ) | ( n8371 & n8373 ) ;
  assign n8375 = n5791 & n6584 ;
  assign n8376 = ~n2810 & n7022 ;
  assign n8377 = n2910 | n6588 ;
  assign n8378 = n2843 & n6587 ;
  assign n8379 = ( ~n2910 & n8377 ) | ( ~n2910 & n8378 ) | ( n8377 & n8378 ) ;
  assign n8380 = ( ~n8375 & n8376 ) | ( ~n8375 & n8379 ) | ( n8376 & n8379 ) ;
  assign n8381 = ( ~x11 & n8375 ) | ( ~x11 & n8380 ) | ( n8375 & n8380 ) ;
  assign n8382 = ( n8375 & n8380 ) | ( n8375 & ~n8381 ) | ( n8380 & ~n8381 ) ;
  assign n8383 = ( x11 & n8381 ) | ( x11 & ~n8382 ) | ( n8381 & ~n8382 ) ;
  assign n8384 = ( ~n8000 & n8002 ) | ( ~n8000 & n8011 ) | ( n8002 & n8011 ) ;
  assign n8385 = ( n8000 & ~n8012 ) | ( n8000 & n8384 ) | ( ~n8012 & n8384 ) ;
  assign n8386 = ( n8374 & n8383 ) | ( n8374 & n8385 ) | ( n8383 & n8385 ) ;
  assign n8387 = ( ~n8012 & n8021 ) | ( ~n8012 & n8023 ) | ( n8021 & n8023 ) ;
  assign n8388 = ( n8012 & ~n8024 ) | ( n8012 & n8387 ) | ( ~n8024 & n8387 ) ;
  assign n8389 = ~n5586 & n6584 ;
  assign n8390 = ~n2725 & n7022 ;
  assign n8391 = n2843 & ~n6588 ;
  assign n8392 = ~n2810 & n6587 ;
  assign n8393 = ( n2843 & ~n8391 ) | ( n2843 & n8392 ) | ( ~n8391 & n8392 ) ;
  assign n8394 = ( ~n8389 & n8390 ) | ( ~n8389 & n8393 ) | ( n8390 & n8393 ) ;
  assign n8395 = ( ~x11 & n8389 ) | ( ~x11 & n8394 ) | ( n8389 & n8394 ) ;
  assign n8396 = ( n8389 & n8394 ) | ( n8389 & ~n8395 ) | ( n8394 & ~n8395 ) ;
  assign n8397 = ( x11 & n8395 ) | ( x11 & ~n8396 ) | ( n8395 & ~n8396 ) ;
  assign n8398 = ( n8386 & n8388 ) | ( n8386 & n8397 ) | ( n8388 & n8397 ) ;
  assign n8399 = ( ~n8024 & n8033 ) | ( ~n8024 & n8035 ) | ( n8033 & n8035 ) ;
  assign n8400 = ( n8024 & ~n8036 ) | ( n8024 & n8399 ) | ( ~n8036 & n8399 ) ;
  assign n8401 = n2725 | n6587 ;
  assign n8402 = n2635 & n7022 ;
  assign n8403 = ( ~n2725 & n8401 ) | ( ~n2725 & n8402 ) | ( n8401 & n8402 ) ;
  assign n8404 = ~n2810 & n6588 ;
  assign n8405 = n8403 | n8404 ;
  assign n8406 = n5232 & n6584 ;
  assign n8407 = ( x11 & n8405 ) | ( x11 & ~n8406 ) | ( n8405 & ~n8406 ) ;
  assign n8408 = ( ~x11 & n8405 ) | ( ~x11 & n8406 ) | ( n8405 & n8406 ) ;
  assign n8409 = ( ~n8405 & n8407 ) | ( ~n8405 & n8408 ) | ( n8407 & n8408 ) ;
  assign n8410 = ( n8398 & n8400 ) | ( n8398 & n8409 ) | ( n8400 & n8409 ) ;
  assign n8411 = ( ~n8036 & n8045 ) | ( ~n8036 & n8047 ) | ( n8045 & n8047 ) ;
  assign n8412 = ( n8036 & ~n8048 ) | ( n8036 & n8411 ) | ( ~n8048 & n8411 ) ;
  assign n8413 = ~n5425 & n6584 ;
  assign n8414 = n2552 & n7022 ;
  assign n8415 = n2725 | n6588 ;
  assign n8416 = n2635 & n6587 ;
  assign n8417 = ( ~n2725 & n8415 ) | ( ~n2725 & n8416 ) | ( n8415 & n8416 ) ;
  assign n8418 = ( ~n8413 & n8414 ) | ( ~n8413 & n8417 ) | ( n8414 & n8417 ) ;
  assign n8419 = ( ~x11 & n8413 ) | ( ~x11 & n8418 ) | ( n8413 & n8418 ) ;
  assign n8420 = ( n8413 & n8418 ) | ( n8413 & ~n8419 ) | ( n8418 & ~n8419 ) ;
  assign n8421 = ( x11 & n8419 ) | ( x11 & ~n8420 ) | ( n8419 & ~n8420 ) ;
  assign n8422 = ( n8410 & n8412 ) | ( n8410 & n8421 ) | ( n8412 & n8421 ) ;
  assign n8423 = ~n5270 & n6584 ;
  assign n8424 = n2552 & n6587 ;
  assign n8425 = n2635 & ~n6588 ;
  assign n8426 = ~n2491 & n7022 ;
  assign n8427 = ( n2635 & ~n8425 ) | ( n2635 & n8426 ) | ( ~n8425 & n8426 ) ;
  assign n8428 = ( ~n8423 & n8424 ) | ( ~n8423 & n8427 ) | ( n8424 & n8427 ) ;
  assign n8429 = ( ~x11 & n8423 ) | ( ~x11 & n8428 ) | ( n8423 & n8428 ) ;
  assign n8430 = ( n8423 & n8428 ) | ( n8423 & ~n8429 ) | ( n8428 & ~n8429 ) ;
  assign n8431 = ( x11 & n8429 ) | ( x11 & ~n8430 ) | ( n8429 & ~n8430 ) ;
  assign n8432 = ( ~n8048 & n8050 ) | ( ~n8048 & n8059 ) | ( n8050 & n8059 ) ;
  assign n8433 = ( n8048 & ~n8060 ) | ( n8048 & n8432 ) | ( ~n8060 & n8432 ) ;
  assign n8434 = ( n8422 & n8431 ) | ( n8422 & n8433 ) | ( n8431 & n8433 ) ;
  assign n8435 = ~n5084 & n6584 ;
  assign n8436 = n2396 & n7022 ;
  assign n8437 = n2552 & ~n6588 ;
  assign n8438 = ~n2491 & n6587 ;
  assign n8439 = ( n2552 & ~n8437 ) | ( n2552 & n8438 ) | ( ~n8437 & n8438 ) ;
  assign n8440 = ( ~n8435 & n8436 ) | ( ~n8435 & n8439 ) | ( n8436 & n8439 ) ;
  assign n8441 = ( ~x11 & n8435 ) | ( ~x11 & n8440 ) | ( n8435 & n8440 ) ;
  assign n8442 = ( n8435 & n8440 ) | ( n8435 & ~n8441 ) | ( n8440 & ~n8441 ) ;
  assign n8443 = ( x11 & n8441 ) | ( x11 & ~n8442 ) | ( n8441 & ~n8442 ) ;
  assign n8444 = ( ~n8060 & n8062 ) | ( ~n8060 & n8071 ) | ( n8062 & n8071 ) ;
  assign n8445 = ( n8060 & ~n8072 ) | ( n8060 & n8444 ) | ( ~n8072 & n8444 ) ;
  assign n8446 = ( n8434 & n8443 ) | ( n8434 & n8445 ) | ( n8443 & n8445 ) ;
  assign n8447 = ~n4900 & n6584 ;
  assign n8448 = n2396 & n6587 ;
  assign n8449 = ~n2298 & n7022 ;
  assign n8450 = ~n2491 & n6588 ;
  assign n8451 = n8449 | n8450 ;
  assign n8452 = ( ~n8447 & n8448 ) | ( ~n8447 & n8451 ) | ( n8448 & n8451 ) ;
  assign n8453 = ( ~x11 & n8447 ) | ( ~x11 & n8452 ) | ( n8447 & n8452 ) ;
  assign n8454 = ( n8447 & n8452 ) | ( n8447 & ~n8453 ) | ( n8452 & ~n8453 ) ;
  assign n8455 = ( x11 & n8453 ) | ( x11 & ~n8454 ) | ( n8453 & ~n8454 ) ;
  assign n8456 = ( ~n8072 & n8074 ) | ( ~n8072 & n8083 ) | ( n8074 & n8083 ) ;
  assign n8457 = ( n8072 & ~n8084 ) | ( n8072 & n8456 ) | ( ~n8084 & n8456 ) ;
  assign n8458 = ( n8446 & n8455 ) | ( n8446 & n8457 ) | ( n8455 & n8457 ) ;
  assign n8459 = ( ~n8084 & n8093 ) | ( ~n8084 & n8095 ) | ( n8093 & n8095 ) ;
  assign n8460 = ( n8084 & ~n8096 ) | ( n8084 & n8459 ) | ( ~n8096 & n8459 ) ;
  assign n8461 = n2298 | n6587 ;
  assign n8462 = n2270 & n7022 ;
  assign n8463 = ( ~n2298 & n8461 ) | ( ~n2298 & n8462 ) | ( n8461 & n8462 ) ;
  assign n8464 = n2396 & n6588 ;
  assign n8465 = n8463 | n8464 ;
  assign n8466 = ~n4912 & n6584 ;
  assign n8467 = ( x11 & n8465 ) | ( x11 & ~n8466 ) | ( n8465 & ~n8466 ) ;
  assign n8468 = ( ~x11 & n8465 ) | ( ~x11 & n8466 ) | ( n8465 & n8466 ) ;
  assign n8469 = ( ~n8465 & n8467 ) | ( ~n8465 & n8468 ) | ( n8467 & n8468 ) ;
  assign n8470 = ( n8458 & n8460 ) | ( n8458 & n8469 ) | ( n8460 & n8469 ) ;
  assign n8471 = ( ~n8096 & n8105 ) | ( ~n8096 & n8107 ) | ( n8105 & n8107 ) ;
  assign n8472 = ( n8096 & ~n8108 ) | ( n8096 & n8471 ) | ( ~n8108 & n8471 ) ;
  assign n8473 = n4647 & n6584 ;
  assign n8474 = n2174 & n7022 ;
  assign n8475 = n2298 | n6588 ;
  assign n8476 = n2270 & n6587 ;
  assign n8477 = ( ~n2298 & n8475 ) | ( ~n2298 & n8476 ) | ( n8475 & n8476 ) ;
  assign n8478 = ( ~n8473 & n8474 ) | ( ~n8473 & n8477 ) | ( n8474 & n8477 ) ;
  assign n8479 = ( ~x11 & n8473 ) | ( ~x11 & n8478 ) | ( n8473 & n8478 ) ;
  assign n8480 = ( n8473 & n8478 ) | ( n8473 & ~n8479 ) | ( n8478 & ~n8479 ) ;
  assign n8481 = ( x11 & n8479 ) | ( x11 & ~n8480 ) | ( n8479 & ~n8480 ) ;
  assign n8482 = ( n8470 & n8472 ) | ( n8470 & n8481 ) | ( n8472 & n8481 ) ;
  assign n8483 = n4730 & n6584 ;
  assign n8484 = n2089 & n7022 ;
  assign n8485 = n2270 & ~n6588 ;
  assign n8486 = n2174 & n6587 ;
  assign n8487 = ( n2270 & ~n8485 ) | ( n2270 & n8486 ) | ( ~n8485 & n8486 ) ;
  assign n8488 = ( ~n8483 & n8484 ) | ( ~n8483 & n8487 ) | ( n8484 & n8487 ) ;
  assign n8489 = ( ~x11 & n8483 ) | ( ~x11 & n8488 ) | ( n8483 & n8488 ) ;
  assign n8490 = ( n8483 & n8488 ) | ( n8483 & ~n8489 ) | ( n8488 & ~n8489 ) ;
  assign n8491 = ( x11 & n8489 ) | ( x11 & ~n8490 ) | ( n8489 & ~n8490 ) ;
  assign n8492 = ( ~n8108 & n8110 ) | ( ~n8108 & n8119 ) | ( n8110 & n8119 ) ;
  assign n8493 = ( n8108 & ~n8120 ) | ( n8108 & n8492 ) | ( ~n8120 & n8492 ) ;
  assign n8494 = ( n8482 & n8491 ) | ( n8482 & n8493 ) | ( n8491 & n8493 ) ;
  assign n8495 = ~n4660 & n6584 ;
  assign n8496 = ~n2023 & n7022 ;
  assign n8497 = n2174 & ~n6588 ;
  assign n8498 = n2089 & n6587 ;
  assign n8499 = ( n2174 & ~n8497 ) | ( n2174 & n8498 ) | ( ~n8497 & n8498 ) ;
  assign n8500 = ( ~n8495 & n8496 ) | ( ~n8495 & n8499 ) | ( n8496 & n8499 ) ;
  assign n8501 = ( ~x11 & n8495 ) | ( ~x11 & n8500 ) | ( n8495 & n8500 ) ;
  assign n8502 = ( n8495 & n8500 ) | ( n8495 & ~n8501 ) | ( n8500 & ~n8501 ) ;
  assign n8503 = ( x11 & n8501 ) | ( x11 & ~n8502 ) | ( n8501 & ~n8502 ) ;
  assign n8504 = ( ~n8120 & n8122 ) | ( ~n8120 & n8131 ) | ( n8122 & n8131 ) ;
  assign n8505 = ( ~n8131 & n8132 ) | ( ~n8131 & n8504 ) | ( n8132 & n8504 ) ;
  assign n8506 = ( n8494 & n8503 ) | ( n8494 & ~n8505 ) | ( n8503 & ~n8505 ) ;
  assign n8507 = ~n4457 & n6584 ;
  assign n8508 = n1926 & n7022 ;
  assign n8509 = n2089 & ~n6588 ;
  assign n8510 = ~n2023 & n6587 ;
  assign n8511 = ( n2089 & ~n8509 ) | ( n2089 & n8510 ) | ( ~n8509 & n8510 ) ;
  assign n8512 = ( ~n8507 & n8508 ) | ( ~n8507 & n8511 ) | ( n8508 & n8511 ) ;
  assign n8513 = ( ~x11 & n8507 ) | ( ~x11 & n8512 ) | ( n8507 & n8512 ) ;
  assign n8514 = ( n8507 & n8512 ) | ( n8507 & ~n8513 ) | ( n8512 & ~n8513 ) ;
  assign n8515 = ( x11 & n8513 ) | ( x11 & ~n8514 ) | ( n8513 & ~n8514 ) ;
  assign n8516 = ( ~n8132 & n8134 ) | ( ~n8132 & n8143 ) | ( n8134 & n8143 ) ;
  assign n8517 = ( ~n8143 & n8144 ) | ( ~n8143 & n8516 ) | ( n8144 & n8516 ) ;
  assign n8518 = ( n8506 & n8515 ) | ( n8506 & ~n8517 ) | ( n8515 & ~n8517 ) ;
  assign n8519 = n4290 & n6584 ;
  assign n8520 = n1852 & n7022 ;
  assign n8521 = n2023 | n6588 ;
  assign n8522 = n1926 & n6587 ;
  assign n8523 = ( ~n2023 & n8521 ) | ( ~n2023 & n8522 ) | ( n8521 & n8522 ) ;
  assign n8524 = ( ~n8519 & n8520 ) | ( ~n8519 & n8523 ) | ( n8520 & n8523 ) ;
  assign n8525 = ( ~x11 & n8519 ) | ( ~x11 & n8524 ) | ( n8519 & n8524 ) ;
  assign n8526 = ( n8519 & n8524 ) | ( n8519 & ~n8525 ) | ( n8524 & ~n8525 ) ;
  assign n8527 = ( x11 & n8525 ) | ( x11 & ~n8526 ) | ( n8525 & ~n8526 ) ;
  assign n8528 = ( ~n8144 & n8146 ) | ( ~n8144 & n8155 ) | ( n8146 & n8155 ) ;
  assign n8529 = ( n8144 & ~n8156 ) | ( n8144 & n8528 ) | ( ~n8156 & n8528 ) ;
  assign n8530 = ( n8518 & n8527 ) | ( n8518 & n8529 ) | ( n8527 & n8529 ) ;
  assign n8531 = ~n4302 & n6584 ;
  assign n8532 = ~n1750 & n7022 ;
  assign n8533 = n1926 & ~n6588 ;
  assign n8534 = n1852 & n6587 ;
  assign n8535 = ( n1926 & ~n8533 ) | ( n1926 & n8534 ) | ( ~n8533 & n8534 ) ;
  assign n8536 = ( ~n8531 & n8532 ) | ( ~n8531 & n8535 ) | ( n8532 & n8535 ) ;
  assign n8537 = ( ~x11 & n8531 ) | ( ~x11 & n8536 ) | ( n8531 & n8536 ) ;
  assign n8538 = ( n8531 & n8536 ) | ( n8531 & ~n8537 ) | ( n8536 & ~n8537 ) ;
  assign n8539 = ( x11 & n8537 ) | ( x11 & ~n8538 ) | ( n8537 & ~n8538 ) ;
  assign n8540 = ( ~n8156 & n8158 ) | ( ~n8156 & n8167 ) | ( n8158 & n8167 ) ;
  assign n8541 = ( ~n8167 & n8168 ) | ( ~n8167 & n8540 ) | ( n8168 & n8540 ) ;
  assign n8542 = ( n8530 & n8539 ) | ( n8530 & ~n8541 ) | ( n8539 & ~n8541 ) ;
  assign n8543 = n4146 & n6584 ;
  assign n8544 = ~n1669 & n7022 ;
  assign n8545 = n1852 & ~n6588 ;
  assign n8546 = ~n1750 & n6587 ;
  assign n8547 = ( n1852 & ~n8545 ) | ( n1852 & n8546 ) | ( ~n8545 & n8546 ) ;
  assign n8548 = ( ~n8543 & n8544 ) | ( ~n8543 & n8547 ) | ( n8544 & n8547 ) ;
  assign n8549 = ( ~x11 & n8543 ) | ( ~x11 & n8548 ) | ( n8543 & n8548 ) ;
  assign n8550 = ( n8543 & n8548 ) | ( n8543 & ~n8549 ) | ( n8548 & ~n8549 ) ;
  assign n8551 = ( x11 & n8549 ) | ( x11 & ~n8550 ) | ( n8549 & ~n8550 ) ;
  assign n8552 = ( ~n8168 & n8170 ) | ( ~n8168 & n8179 ) | ( n8170 & n8179 ) ;
  assign n8553 = ( n8168 & ~n8180 ) | ( n8168 & n8552 ) | ( ~n8180 & n8552 ) ;
  assign n8554 = ( n8542 & n8551 ) | ( n8542 & n8553 ) | ( n8551 & n8553 ) ;
  assign n8555 = n4326 & n6584 ;
  assign n8556 = n1576 & n7022 ;
  assign n8557 = n1750 | n6588 ;
  assign n8558 = ~n1669 & n6587 ;
  assign n8559 = ( ~n1750 & n8557 ) | ( ~n1750 & n8558 ) | ( n8557 & n8558 ) ;
  assign n8560 = ( ~n8555 & n8556 ) | ( ~n8555 & n8559 ) | ( n8556 & n8559 ) ;
  assign n8561 = ( ~x11 & n8555 ) | ( ~x11 & n8560 ) | ( n8555 & n8560 ) ;
  assign n8562 = ( n8555 & n8560 ) | ( n8555 & ~n8561 ) | ( n8560 & ~n8561 ) ;
  assign n8563 = ( x11 & n8561 ) | ( x11 & ~n8562 ) | ( n8561 & ~n8562 ) ;
  assign n8564 = ( ~n8180 & n8182 ) | ( ~n8180 & n8191 ) | ( n8182 & n8191 ) ;
  assign n8565 = ( n8180 & ~n8192 ) | ( n8180 & n8564 ) | ( ~n8192 & n8564 ) ;
  assign n8566 = ( n8554 & n8563 ) | ( n8554 & n8565 ) | ( n8563 & n8565 ) ;
  assign n8567 = ( n8192 & ~n8194 ) | ( n8192 & n8203 ) | ( ~n8194 & n8203 ) ;
  assign n8568 = ( n8194 & ~n8204 ) | ( n8194 & n8567 ) | ( ~n8204 & n8567 ) ;
  assign n8569 = ~n3791 & n7296 ;
  assign n8570 = n1267 & n7299 ;
  assign n8571 = n1338 | n7300 ;
  assign n8572 = ~n1246 & n7879 ;
  assign n8573 = ( ~n1338 & n8571 ) | ( ~n1338 & n8572 ) | ( n8571 & n8572 ) ;
  assign n8574 = ( ~n8569 & n8570 ) | ( ~n8569 & n8573 ) | ( n8570 & n8573 ) ;
  assign n8575 = ( ~x8 & n8569 ) | ( ~x8 & n8574 ) | ( n8569 & n8574 ) ;
  assign n8576 = ( n8569 & n8574 ) | ( n8569 & ~n8575 ) | ( n8574 & ~n8575 ) ;
  assign n8577 = ( x8 & n8575 ) | ( x8 & ~n8576 ) | ( n8575 & ~n8576 ) ;
  assign n8578 = ( n8566 & n8568 ) | ( n8566 & n8577 ) | ( n8568 & n8577 ) ;
  assign n8579 = n3797 & n8230 ;
  assign n8580 = ~n3692 & n8225 ;
  assign n8581 = ~n3658 & n8226 ;
  assign n8582 = n8580 | n8581 ;
  assign n8583 = ( ~x5 & n8579 ) | ( ~x5 & n8582 ) | ( n8579 & n8582 ) ;
  assign n8584 = ( n8579 & n8582 ) | ( n8579 & ~n8583 ) | ( n8582 & ~n8583 ) ;
  assign n8585 = ( x5 & n8583 ) | ( x5 & ~n8584 ) | ( n8583 & ~n8584 ) ;
  assign n8586 = ( n8204 & ~n8206 ) | ( n8204 & n8215 ) | ( ~n8206 & n8215 ) ;
  assign n8587 = ( n8206 & ~n8216 ) | ( n8206 & n8586 ) | ( ~n8216 & n8586 ) ;
  assign n8588 = ( n8578 & n8585 ) | ( n8578 & n8587 ) | ( n8585 & n8587 ) ;
  assign n8589 = n6061 & n7296 ;
  assign n8590 = n3479 & n7299 ;
  assign n8591 = n3533 | n7300 ;
  assign n8592 = ~n3389 & n7879 ;
  assign n8593 = ( ~n3533 & n8591 ) | ( ~n3533 & n8592 ) | ( n8591 & n8592 ) ;
  assign n8594 = ( ~n8589 & n8590 ) | ( ~n8589 & n8593 ) | ( n8590 & n8593 ) ;
  assign n8595 = ( ~x8 & n8589 ) | ( ~x8 & n8594 ) | ( n8589 & n8594 ) ;
  assign n8596 = ( n8589 & n8594 ) | ( n8589 & ~n8595 ) | ( n8594 & ~n8595 ) ;
  assign n8597 = ( x8 & n8595 ) | ( x8 & ~n8596 ) | ( n8595 & ~n8596 ) ;
  assign n8598 = ( n3479 & n6009 ) | ( n3479 & n7296 ) | ( n6009 & n7296 ) ;
  assign n8599 = ~n3533 & n7299 ;
  assign n8600 = ~n3586 & n7300 ;
  assign n8601 = n8599 | n8600 ;
  assign n8602 = ~n3479 & n7879 ;
  assign n8603 = ( n7879 & n8601 ) | ( n7879 & ~n8602 ) | ( n8601 & ~n8602 ) ;
  assign n8604 = ( ~n6608 & n8598 ) | ( ~n6608 & n8603 ) | ( n8598 & n8603 ) ;
  assign n8605 = ~n3586 & n7878 ;
  assign n8606 = x8 & n8605 ;
  assign n8607 = ( n6009 & n6618 ) | ( n6009 & n7296 ) | ( n6618 & n7296 ) ;
  assign n8608 = ~n3533 & n7879 ;
  assign n8609 = n3586 | n7299 ;
  assign n8610 = ( ~n3586 & n8608 ) | ( ~n3586 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8611 = n8607 | n8610 ;
  assign n8612 = ( x8 & n8606 ) | ( x8 & n8611 ) | ( n8606 & n8611 ) ;
  assign n8613 = n8604 | n8612 ;
  assign n8614 = x8 & ~n8613 ;
  assign n8615 = ( n8255 & n8597 ) | ( n8255 & n8614 ) | ( n8597 & n8614 ) ;
  assign n8616 = n3389 | n7299 ;
  assign n8617 = ~n3355 & n7879 ;
  assign n8618 = ( ~n3389 & n8616 ) | ( ~n3389 & n8617 ) | ( n8616 & n8617 ) ;
  assign n8619 = n3479 & n7300 ;
  assign n8620 = n8618 | n8619 ;
  assign n8621 = ~n6104 & n7296 ;
  assign n8622 = ( x8 & n8620 ) | ( x8 & ~n8621 ) | ( n8620 & ~n8621 ) ;
  assign n8623 = ( ~x8 & n8620 ) | ( ~x8 & n8621 ) | ( n8620 & n8621 ) ;
  assign n8624 = ( ~n8620 & n8622 ) | ( ~n8620 & n8623 ) | ( n8622 & n8623 ) ;
  assign n8625 = ( n8256 & n8257 ) | ( n8256 & n8260 ) | ( n8257 & n8260 ) ;
  assign n8626 = ~n8256 & n8261 ;
  assign n8627 = ( n8256 & ~n8625 ) | ( n8256 & n8626 ) | ( ~n8625 & n8626 ) ;
  assign n8628 = ( n8615 & n8624 ) | ( n8615 & n8627 ) | ( n8624 & n8627 ) ;
  assign n8629 = ~n6154 & n7296 ;
  assign n8630 = ~n3300 & n7879 ;
  assign n8631 = n3389 | n7300 ;
  assign n8632 = ~n3355 & n7299 ;
  assign n8633 = ( ~n3389 & n8631 ) | ( ~n3389 & n8632 ) | ( n8631 & n8632 ) ;
  assign n8634 = ( ~n8629 & n8630 ) | ( ~n8629 & n8633 ) | ( n8630 & n8633 ) ;
  assign n8635 = ( ~x8 & n8629 ) | ( ~x8 & n8634 ) | ( n8629 & n8634 ) ;
  assign n8636 = ( n8629 & n8634 ) | ( n8629 & ~n8635 ) | ( n8634 & ~n8635 ) ;
  assign n8637 = ( x8 & n8635 ) | ( x8 & ~n8636 ) | ( n8635 & ~n8636 ) ;
  assign n8638 = ( n8254 & n8262 ) | ( n8254 & ~n8263 ) | ( n8262 & ~n8263 ) ;
  assign n8639 = n8263 & ~n8638 ;
  assign n8640 = ( n8628 & n8637 ) | ( n8628 & n8639 ) | ( n8637 & n8639 ) ;
  assign n8641 = n6200 & n7296 ;
  assign n8642 = ~n3300 & n7299 ;
  assign n8643 = n3355 | n7300 ;
  assign n8644 = n3239 & n7879 ;
  assign n8645 = ( ~n3355 & n8643 ) | ( ~n3355 & n8644 ) | ( n8643 & n8644 ) ;
  assign n8646 = ( ~n8641 & n8642 ) | ( ~n8641 & n8645 ) | ( n8642 & n8645 ) ;
  assign n8647 = ( ~x8 & n8641 ) | ( ~x8 & n8646 ) | ( n8641 & n8646 ) ;
  assign n8648 = ( n8641 & n8646 ) | ( n8641 & ~n8647 ) | ( n8646 & ~n8647 ) ;
  assign n8649 = ( x8 & n8647 ) | ( x8 & ~n8648 ) | ( n8647 & ~n8648 ) ;
  assign n8650 = ( n7915 & n8247 ) | ( n7915 & ~n8264 ) | ( n8247 & ~n8264 ) ;
  assign n8651 = ( n8264 & ~n8265 ) | ( n8264 & n8650 ) | ( ~n8265 & n8650 ) ;
  assign n8652 = ( n8640 & n8649 ) | ( n8640 & n8651 ) | ( n8649 & n8651 ) ;
  assign n8653 = ~n6243 & n7296 ;
  assign n8654 = n3153 & n7879 ;
  assign n8655 = n3300 | n7300 ;
  assign n8656 = n3239 & n7299 ;
  assign n8657 = ( ~n3300 & n8655 ) | ( ~n3300 & n8656 ) | ( n8655 & n8656 ) ;
  assign n8658 = ( ~n8653 & n8654 ) | ( ~n8653 & n8657 ) | ( n8654 & n8657 ) ;
  assign n8659 = ( ~x8 & n8653 ) | ( ~x8 & n8658 ) | ( n8653 & n8658 ) ;
  assign n8660 = ( n8653 & n8658 ) | ( n8653 & ~n8659 ) | ( n8658 & ~n8659 ) ;
  assign n8661 = ( x8 & n8659 ) | ( x8 & ~n8660 ) | ( n8659 & ~n8660 ) ;
  assign n8662 = ( ~n8265 & n8274 ) | ( ~n8265 & n8277 ) | ( n8274 & n8277 ) ;
  assign n8663 = ( n8265 & ~n8278 ) | ( n8265 & n8662 ) | ( ~n8278 & n8662 ) ;
  assign n8664 = ( n8652 & n8661 ) | ( n8652 & n8663 ) | ( n8661 & n8663 ) ;
  assign n8665 = ( ~n8278 & n8287 ) | ( ~n8278 & n8289 ) | ( n8287 & n8289 ) ;
  assign n8666 = ( n8278 & ~n8290 ) | ( n8278 & n8665 ) | ( ~n8290 & n8665 ) ;
  assign n8667 = n5710 & n7296 ;
  assign n8668 = n3153 & n7299 ;
  assign n8669 = n3239 & ~n7300 ;
  assign n8670 = n3078 & n7879 ;
  assign n8671 = ( n3239 & ~n8669 ) | ( n3239 & n8670 ) | ( ~n8669 & n8670 ) ;
  assign n8672 = ( ~n8667 & n8668 ) | ( ~n8667 & n8671 ) | ( n8668 & n8671 ) ;
  assign n8673 = ( ~x8 & n8667 ) | ( ~x8 & n8672 ) | ( n8667 & n8672 ) ;
  assign n8674 = ( n8667 & n8672 ) | ( n8667 & ~n8673 ) | ( n8672 & ~n8673 ) ;
  assign n8675 = ( x8 & n8673 ) | ( x8 & ~n8674 ) | ( n8673 & ~n8674 ) ;
  assign n8676 = ( n8664 & n8666 ) | ( n8664 & n8675 ) | ( n8666 & n8675 ) ;
  assign n8677 = ( ~n8290 & n8299 ) | ( ~n8290 & n8301 ) | ( n8299 & n8301 ) ;
  assign n8678 = ( n8290 & ~n8302 ) | ( n8290 & n8677 ) | ( ~n8302 & n8677 ) ;
  assign n8679 = n3078 & ~n7299 ;
  assign n8680 = ~n3046 & n7879 ;
  assign n8681 = ( n3078 & ~n8679 ) | ( n3078 & n8680 ) | ( ~n8679 & n8680 ) ;
  assign n8682 = n3153 & n7300 ;
  assign n8683 = n8681 | n8682 ;
  assign n8684 = ~n6267 & n7296 ;
  assign n8685 = ( x8 & n8683 ) | ( x8 & ~n8684 ) | ( n8683 & ~n8684 ) ;
  assign n8686 = ( ~x8 & n8683 ) | ( ~x8 & n8684 ) | ( n8683 & n8684 ) ;
  assign n8687 = ( ~n8683 & n8685 ) | ( ~n8683 & n8686 ) | ( n8685 & n8686 ) ;
  assign n8688 = ( n8676 & n8678 ) | ( n8676 & n8687 ) | ( n8678 & n8687 ) ;
  assign n8689 = ( ~n8302 & n8311 ) | ( ~n8302 & n8313 ) | ( n8311 & n8313 ) ;
  assign n8690 = ( n8302 & ~n8314 ) | ( n8302 & n8689 ) | ( ~n8314 & n8689 ) ;
  assign n8691 = n6279 & n7296 ;
  assign n8692 = ~n2965 & n7879 ;
  assign n8693 = n3078 & ~n7300 ;
  assign n8694 = ~n3046 & n7299 ;
  assign n8695 = ( n3078 & ~n8693 ) | ( n3078 & n8694 ) | ( ~n8693 & n8694 ) ;
  assign n8696 = ( ~n8691 & n8692 ) | ( ~n8691 & n8695 ) | ( n8692 & n8695 ) ;
  assign n8697 = ( ~x8 & n8691 ) | ( ~x8 & n8696 ) | ( n8691 & n8696 ) ;
  assign n8698 = ( n8691 & n8696 ) | ( n8691 & ~n8697 ) | ( n8696 & ~n8697 ) ;
  assign n8699 = ( x8 & n8697 ) | ( x8 & ~n8698 ) | ( n8697 & ~n8698 ) ;
  assign n8700 = ( n8688 & n8690 ) | ( n8688 & n8699 ) | ( n8690 & n8699 ) ;
  assign n8701 = ~n5768 & n7296 ;
  assign n8702 = ~n2910 & n7879 ;
  assign n8703 = n3046 | n7300 ;
  assign n8704 = ~n2965 & n7299 ;
  assign n8705 = ( ~n3046 & n8703 ) | ( ~n3046 & n8704 ) | ( n8703 & n8704 ) ;
  assign n8706 = ( ~n8701 & n8702 ) | ( ~n8701 & n8705 ) | ( n8702 & n8705 ) ;
  assign n8707 = ( ~x8 & n8701 ) | ( ~x8 & n8706 ) | ( n8701 & n8706 ) ;
  assign n8708 = ( n8701 & n8706 ) | ( n8701 & ~n8707 ) | ( n8706 & ~n8707 ) ;
  assign n8709 = ( x8 & n8707 ) | ( x8 & ~n8708 ) | ( n8707 & ~n8708 ) ;
  assign n8710 = ( ~n8314 & n8316 ) | ( ~n8314 & n8325 ) | ( n8316 & n8325 ) ;
  assign n8711 = ( n8314 & ~n8326 ) | ( n8314 & n8710 ) | ( ~n8326 & n8710 ) ;
  assign n8712 = ( n8700 & n8709 ) | ( n8700 & n8711 ) | ( n8709 & n8711 ) ;
  assign n8713 = n5543 & n7296 ;
  assign n8714 = ~n2910 & n7299 ;
  assign n8715 = n2965 | n7300 ;
  assign n8716 = n2843 & n7879 ;
  assign n8717 = ( ~n2965 & n8715 ) | ( ~n2965 & n8716 ) | ( n8715 & n8716 ) ;
  assign n8718 = ( ~n8713 & n8714 ) | ( ~n8713 & n8717 ) | ( n8714 & n8717 ) ;
  assign n8719 = ( ~x8 & n8713 ) | ( ~x8 & n8718 ) | ( n8713 & n8718 ) ;
  assign n8720 = ( n8713 & n8718 ) | ( n8713 & ~n8719 ) | ( n8718 & ~n8719 ) ;
  assign n8721 = ( x8 & n8719 ) | ( x8 & ~n8720 ) | ( n8719 & ~n8720 ) ;
  assign n8722 = ( ~n8326 & n8328 ) | ( ~n8326 & n8337 ) | ( n8328 & n8337 ) ;
  assign n8723 = ( n8326 & ~n8338 ) | ( n8326 & n8722 ) | ( ~n8338 & n8722 ) ;
  assign n8724 = ( n8712 & n8721 ) | ( n8712 & n8723 ) | ( n8721 & n8723 ) ;
  assign n8725 = n5791 & n7296 ;
  assign n8726 = ~n2810 & n7879 ;
  assign n8727 = n2910 | n7300 ;
  assign n8728 = n2843 & n7299 ;
  assign n8729 = ( ~n2910 & n8727 ) | ( ~n2910 & n8728 ) | ( n8727 & n8728 ) ;
  assign n8730 = ( ~n8725 & n8726 ) | ( ~n8725 & n8729 ) | ( n8726 & n8729 ) ;
  assign n8731 = ( ~x8 & n8725 ) | ( ~x8 & n8730 ) | ( n8725 & n8730 ) ;
  assign n8732 = ( n8725 & n8730 ) | ( n8725 & ~n8731 ) | ( n8730 & ~n8731 ) ;
  assign n8733 = ( x8 & n8731 ) | ( x8 & ~n8732 ) | ( n8731 & ~n8732 ) ;
  assign n8734 = ( ~n8338 & n8340 ) | ( ~n8338 & n8349 ) | ( n8340 & n8349 ) ;
  assign n8735 = ( n8338 & ~n8350 ) | ( n8338 & n8734 ) | ( ~n8350 & n8734 ) ;
  assign n8736 = ( n8724 & n8733 ) | ( n8724 & n8735 ) | ( n8733 & n8735 ) ;
  assign n8737 = ( ~n8350 & n8359 ) | ( ~n8350 & n8361 ) | ( n8359 & n8361 ) ;
  assign n8738 = ( n8350 & ~n8362 ) | ( n8350 & n8737 ) | ( ~n8362 & n8737 ) ;
  assign n8739 = ~n5586 & n7296 ;
  assign n8740 = ~n2725 & n7879 ;
  assign n8741 = n2843 & ~n7300 ;
  assign n8742 = ~n2810 & n7299 ;
  assign n8743 = ( n2843 & ~n8741 ) | ( n2843 & n8742 ) | ( ~n8741 & n8742 ) ;
  assign n8744 = ( ~n8739 & n8740 ) | ( ~n8739 & n8743 ) | ( n8740 & n8743 ) ;
  assign n8745 = ( ~x8 & n8739 ) | ( ~x8 & n8744 ) | ( n8739 & n8744 ) ;
  assign n8746 = ( n8739 & n8744 ) | ( n8739 & ~n8745 ) | ( n8744 & ~n8745 ) ;
  assign n8747 = ( x8 & n8745 ) | ( x8 & ~n8746 ) | ( n8745 & ~n8746 ) ;
  assign n8748 = ( n8736 & n8738 ) | ( n8736 & n8747 ) | ( n8738 & n8747 ) ;
  assign n8749 = ( ~n8362 & n8371 ) | ( ~n8362 & n8373 ) | ( n8371 & n8373 ) ;
  assign n8750 = ( n8362 & ~n8374 ) | ( n8362 & n8749 ) | ( ~n8374 & n8749 ) ;
  assign n8751 = n2725 | n7299 ;
  assign n8752 = n2635 & n7879 ;
  assign n8753 = ( ~n2725 & n8751 ) | ( ~n2725 & n8752 ) | ( n8751 & n8752 ) ;
  assign n8754 = ~n2810 & n7300 ;
  assign n8755 = n8753 | n8754 ;
  assign n8756 = n5232 & n7296 ;
  assign n8757 = ( x8 & n8755 ) | ( x8 & ~n8756 ) | ( n8755 & ~n8756 ) ;
  assign n8758 = ( ~x8 & n8755 ) | ( ~x8 & n8756 ) | ( n8755 & n8756 ) ;
  assign n8759 = ( ~n8755 & n8757 ) | ( ~n8755 & n8758 ) | ( n8757 & n8758 ) ;
  assign n8760 = ( n8748 & n8750 ) | ( n8748 & n8759 ) | ( n8750 & n8759 ) ;
  assign n8761 = ( ~n8374 & n8383 ) | ( ~n8374 & n8385 ) | ( n8383 & n8385 ) ;
  assign n8762 = ( n8374 & ~n8386 ) | ( n8374 & n8761 ) | ( ~n8386 & n8761 ) ;
  assign n8763 = ~n5425 & n7296 ;
  assign n8764 = n2552 & n7879 ;
  assign n8765 = n2725 | n7300 ;
  assign n8766 = n2635 & n7299 ;
  assign n8767 = ( ~n2725 & n8765 ) | ( ~n2725 & n8766 ) | ( n8765 & n8766 ) ;
  assign n8768 = ( ~n8763 & n8764 ) | ( ~n8763 & n8767 ) | ( n8764 & n8767 ) ;
  assign n8769 = ( ~x8 & n8763 ) | ( ~x8 & n8768 ) | ( n8763 & n8768 ) ;
  assign n8770 = ( n8763 & n8768 ) | ( n8763 & ~n8769 ) | ( n8768 & ~n8769 ) ;
  assign n8771 = ( x8 & n8769 ) | ( x8 & ~n8770 ) | ( n8769 & ~n8770 ) ;
  assign n8772 = ( n8760 & n8762 ) | ( n8760 & n8771 ) | ( n8762 & n8771 ) ;
  assign n8773 = ~n5270 & n7296 ;
  assign n8774 = n2552 & n7299 ;
  assign n8775 = n2635 & ~n7300 ;
  assign n8776 = ~n2491 & n7879 ;
  assign n8777 = ( n2635 & ~n8775 ) | ( n2635 & n8776 ) | ( ~n8775 & n8776 ) ;
  assign n8778 = ( ~n8773 & n8774 ) | ( ~n8773 & n8777 ) | ( n8774 & n8777 ) ;
  assign n8779 = ( ~x8 & n8773 ) | ( ~x8 & n8778 ) | ( n8773 & n8778 ) ;
  assign n8780 = ( n8773 & n8778 ) | ( n8773 & ~n8779 ) | ( n8778 & ~n8779 ) ;
  assign n8781 = ( x8 & n8779 ) | ( x8 & ~n8780 ) | ( n8779 & ~n8780 ) ;
  assign n8782 = ( ~n8386 & n8388 ) | ( ~n8386 & n8397 ) | ( n8388 & n8397 ) ;
  assign n8783 = ( n8386 & ~n8398 ) | ( n8386 & n8782 ) | ( ~n8398 & n8782 ) ;
  assign n8784 = ( n8772 & n8781 ) | ( n8772 & n8783 ) | ( n8781 & n8783 ) ;
  assign n8785 = ~n5084 & n7296 ;
  assign n8786 = n2396 & n7879 ;
  assign n8787 = n2552 & ~n7300 ;
  assign n8788 = ~n2491 & n7299 ;
  assign n8789 = ( n2552 & ~n8787 ) | ( n2552 & n8788 ) | ( ~n8787 & n8788 ) ;
  assign n8790 = ( ~n8785 & n8786 ) | ( ~n8785 & n8789 ) | ( n8786 & n8789 ) ;
  assign n8791 = ( ~x8 & n8785 ) | ( ~x8 & n8790 ) | ( n8785 & n8790 ) ;
  assign n8792 = ( n8785 & n8790 ) | ( n8785 & ~n8791 ) | ( n8790 & ~n8791 ) ;
  assign n8793 = ( x8 & n8791 ) | ( x8 & ~n8792 ) | ( n8791 & ~n8792 ) ;
  assign n8794 = ( ~n8398 & n8400 ) | ( ~n8398 & n8409 ) | ( n8400 & n8409 ) ;
  assign n8795 = ( n8398 & ~n8410 ) | ( n8398 & n8794 ) | ( ~n8410 & n8794 ) ;
  assign n8796 = ( n8784 & n8793 ) | ( n8784 & n8795 ) | ( n8793 & n8795 ) ;
  assign n8797 = ~n4900 & n7296 ;
  assign n8798 = n2396 & n7299 ;
  assign n8799 = ~n2298 & n7879 ;
  assign n8800 = ~n2491 & n7300 ;
  assign n8801 = n8799 | n8800 ;
  assign n8802 = ( ~n8797 & n8798 ) | ( ~n8797 & n8801 ) | ( n8798 & n8801 ) ;
  assign n8803 = ( ~x8 & n8797 ) | ( ~x8 & n8802 ) | ( n8797 & n8802 ) ;
  assign n8804 = ( n8797 & n8802 ) | ( n8797 & ~n8803 ) | ( n8802 & ~n8803 ) ;
  assign n8805 = ( x8 & n8803 ) | ( x8 & ~n8804 ) | ( n8803 & ~n8804 ) ;
  assign n8806 = ( ~n8410 & n8412 ) | ( ~n8410 & n8421 ) | ( n8412 & n8421 ) ;
  assign n8807 = ( n8410 & ~n8422 ) | ( n8410 & n8806 ) | ( ~n8422 & n8806 ) ;
  assign n8808 = ( n8796 & n8805 ) | ( n8796 & n8807 ) | ( n8805 & n8807 ) ;
  assign n8809 = ( ~n8422 & n8431 ) | ( ~n8422 & n8433 ) | ( n8431 & n8433 ) ;
  assign n8810 = ( n8422 & ~n8434 ) | ( n8422 & n8809 ) | ( ~n8434 & n8809 ) ;
  assign n8811 = n2298 | n7299 ;
  assign n8812 = n2270 & n7879 ;
  assign n8813 = ( ~n2298 & n8811 ) | ( ~n2298 & n8812 ) | ( n8811 & n8812 ) ;
  assign n8814 = n2396 & n7300 ;
  assign n8815 = n8813 | n8814 ;
  assign n8816 = ~n4912 & n7296 ;
  assign n8817 = ( x8 & n8815 ) | ( x8 & ~n8816 ) | ( n8815 & ~n8816 ) ;
  assign n8818 = ( ~x8 & n8815 ) | ( ~x8 & n8816 ) | ( n8815 & n8816 ) ;
  assign n8819 = ( ~n8815 & n8817 ) | ( ~n8815 & n8818 ) | ( n8817 & n8818 ) ;
  assign n8820 = ( n8808 & n8810 ) | ( n8808 & n8819 ) | ( n8810 & n8819 ) ;
  assign n8821 = ( ~n8434 & n8443 ) | ( ~n8434 & n8445 ) | ( n8443 & n8445 ) ;
  assign n8822 = ( n8434 & ~n8446 ) | ( n8434 & n8821 ) | ( ~n8446 & n8821 ) ;
  assign n8823 = n4647 & n7296 ;
  assign n8824 = n2174 & n7879 ;
  assign n8825 = n2298 | n7300 ;
  assign n8826 = n2270 & n7299 ;
  assign n8827 = ( ~n2298 & n8825 ) | ( ~n2298 & n8826 ) | ( n8825 & n8826 ) ;
  assign n8828 = ( ~n8823 & n8824 ) | ( ~n8823 & n8827 ) | ( n8824 & n8827 ) ;
  assign n8829 = ( ~x8 & n8823 ) | ( ~x8 & n8828 ) | ( n8823 & n8828 ) ;
  assign n8830 = ( n8823 & n8828 ) | ( n8823 & ~n8829 ) | ( n8828 & ~n8829 ) ;
  assign n8831 = ( x8 & n8829 ) | ( x8 & ~n8830 ) | ( n8829 & ~n8830 ) ;
  assign n8832 = ( n8820 & n8822 ) | ( n8820 & n8831 ) | ( n8822 & n8831 ) ;
  assign n8833 = ( ~n8446 & n8455 ) | ( ~n8446 & n8457 ) | ( n8455 & n8457 ) ;
  assign n8834 = ( n8446 & ~n8458 ) | ( n8446 & n8833 ) | ( ~n8458 & n8833 ) ;
  assign n8835 = n4730 & n7296 ;
  assign n8836 = n2089 & n7879 ;
  assign n8837 = n2270 & ~n7300 ;
  assign n8838 = n2174 & n7299 ;
  assign n8839 = ( n2270 & ~n8837 ) | ( n2270 & n8838 ) | ( ~n8837 & n8838 ) ;
  assign n8840 = ( ~n8835 & n8836 ) | ( ~n8835 & n8839 ) | ( n8836 & n8839 ) ;
  assign n8841 = ( ~x8 & n8835 ) | ( ~x8 & n8840 ) | ( n8835 & n8840 ) ;
  assign n8842 = ( n8835 & n8840 ) | ( n8835 & ~n8841 ) | ( n8840 & ~n8841 ) ;
  assign n8843 = ( x8 & n8841 ) | ( x8 & ~n8842 ) | ( n8841 & ~n8842 ) ;
  assign n8844 = ( n8832 & n8834 ) | ( n8832 & n8843 ) | ( n8834 & n8843 ) ;
  assign n8845 = ~n4660 & n7296 ;
  assign n8846 = ~n2023 & n7879 ;
  assign n8847 = n2174 & ~n7300 ;
  assign n8848 = n2089 & n7299 ;
  assign n8849 = ( n2174 & ~n8847 ) | ( n2174 & n8848 ) | ( ~n8847 & n8848 ) ;
  assign n8850 = ( ~n8845 & n8846 ) | ( ~n8845 & n8849 ) | ( n8846 & n8849 ) ;
  assign n8851 = ( ~x8 & n8845 ) | ( ~x8 & n8850 ) | ( n8845 & n8850 ) ;
  assign n8852 = ( n8845 & n8850 ) | ( n8845 & ~n8851 ) | ( n8850 & ~n8851 ) ;
  assign n8853 = ( x8 & n8851 ) | ( x8 & ~n8852 ) | ( n8851 & ~n8852 ) ;
  assign n8854 = ( ~n8458 & n8460 ) | ( ~n8458 & n8469 ) | ( n8460 & n8469 ) ;
  assign n8855 = ( n8458 & ~n8470 ) | ( n8458 & n8854 ) | ( ~n8470 & n8854 ) ;
  assign n8856 = ( n8844 & n8853 ) | ( n8844 & n8855 ) | ( n8853 & n8855 ) ;
  assign n8857 = ~n4457 & n7296 ;
  assign n8858 = n1926 & n7879 ;
  assign n8859 = n2089 & ~n7300 ;
  assign n8860 = ~n2023 & n7299 ;
  assign n8861 = ( n2089 & ~n8859 ) | ( n2089 & n8860 ) | ( ~n8859 & n8860 ) ;
  assign n8862 = ( ~n8857 & n8858 ) | ( ~n8857 & n8861 ) | ( n8858 & n8861 ) ;
  assign n8863 = ( ~x8 & n8857 ) | ( ~x8 & n8862 ) | ( n8857 & n8862 ) ;
  assign n8864 = ( n8857 & n8862 ) | ( n8857 & ~n8863 ) | ( n8862 & ~n8863 ) ;
  assign n8865 = ( x8 & n8863 ) | ( x8 & ~n8864 ) | ( n8863 & ~n8864 ) ;
  assign n8866 = ( ~n8470 & n8472 ) | ( ~n8470 & n8481 ) | ( n8472 & n8481 ) ;
  assign n8867 = ( n8470 & ~n8482 ) | ( n8470 & n8866 ) | ( ~n8482 & n8866 ) ;
  assign n8868 = ( n8856 & n8865 ) | ( n8856 & n8867 ) | ( n8865 & n8867 ) ;
  assign n8869 = ( ~n8482 & n8491 ) | ( ~n8482 & n8493 ) | ( n8491 & n8493 ) ;
  assign n8870 = ( n8482 & ~n8494 ) | ( n8482 & n8869 ) | ( ~n8494 & n8869 ) ;
  assign n8871 = n4290 & n7296 ;
  assign n8872 = n1852 & n7879 ;
  assign n8873 = n2023 | n7300 ;
  assign n8874 = n1926 & n7299 ;
  assign n8875 = ( ~n2023 & n8873 ) | ( ~n2023 & n8874 ) | ( n8873 & n8874 ) ;
  assign n8876 = ( ~n8871 & n8872 ) | ( ~n8871 & n8875 ) | ( n8872 & n8875 ) ;
  assign n8877 = ( ~x8 & n8871 ) | ( ~x8 & n8876 ) | ( n8871 & n8876 ) ;
  assign n8878 = ( n8871 & n8876 ) | ( n8871 & ~n8877 ) | ( n8876 & ~n8877 ) ;
  assign n8879 = ( x8 & n8877 ) | ( x8 & ~n8878 ) | ( n8877 & ~n8878 ) ;
  assign n8880 = ( n8868 & n8870 ) | ( n8868 & n8879 ) | ( n8870 & n8879 ) ;
  assign n8881 = ( n8494 & ~n8503 ) | ( n8494 & n8505 ) | ( ~n8503 & n8505 ) ;
  assign n8882 = ( ~n8494 & n8506 ) | ( ~n8494 & n8881 ) | ( n8506 & n8881 ) ;
  assign n8883 = ~n4302 & n7296 ;
  assign n8884 = ~n1750 & n7879 ;
  assign n8885 = n1926 & ~n7300 ;
  assign n8886 = n1852 & n7299 ;
  assign n8887 = ( n1926 & ~n8885 ) | ( n1926 & n8886 ) | ( ~n8885 & n8886 ) ;
  assign n8888 = ( ~n8883 & n8884 ) | ( ~n8883 & n8887 ) | ( n8884 & n8887 ) ;
  assign n8889 = ( ~x8 & n8883 ) | ( ~x8 & n8888 ) | ( n8883 & n8888 ) ;
  assign n8890 = ( n8883 & n8888 ) | ( n8883 & ~n8889 ) | ( n8888 & ~n8889 ) ;
  assign n8891 = ( x8 & n8889 ) | ( x8 & ~n8890 ) | ( n8889 & ~n8890 ) ;
  assign n8892 = ( n8880 & ~n8882 ) | ( n8880 & n8891 ) | ( ~n8882 & n8891 ) ;
  assign n8893 = ( n8506 & ~n8515 ) | ( n8506 & n8517 ) | ( ~n8515 & n8517 ) ;
  assign n8894 = ( ~n8506 & n8518 ) | ( ~n8506 & n8893 ) | ( n8518 & n8893 ) ;
  assign n8895 = n4146 & n7296 ;
  assign n8896 = ~n1669 & n7879 ;
  assign n8897 = n1852 & ~n7300 ;
  assign n8898 = ~n1750 & n7299 ;
  assign n8899 = ( n1852 & ~n8897 ) | ( n1852 & n8898 ) | ( ~n8897 & n8898 ) ;
  assign n8900 = ( ~n8895 & n8896 ) | ( ~n8895 & n8899 ) | ( n8896 & n8899 ) ;
  assign n8901 = ( ~x8 & n8895 ) | ( ~x8 & n8900 ) | ( n8895 & n8900 ) ;
  assign n8902 = ( n8895 & n8900 ) | ( n8895 & ~n8901 ) | ( n8900 & ~n8901 ) ;
  assign n8903 = ( x8 & n8901 ) | ( x8 & ~n8902 ) | ( n8901 & ~n8902 ) ;
  assign n8904 = ( n8892 & ~n8894 ) | ( n8892 & n8903 ) | ( ~n8894 & n8903 ) ;
  assign n8905 = ( ~n8518 & n8527 ) | ( ~n8518 & n8529 ) | ( n8527 & n8529 ) ;
  assign n8906 = ( n8518 & ~n8530 ) | ( n8518 & n8905 ) | ( ~n8530 & n8905 ) ;
  assign n8907 = n4326 & n7296 ;
  assign n8908 = n1576 & n7879 ;
  assign n8909 = n1750 | n7300 ;
  assign n8910 = ~n1669 & n7299 ;
  assign n8911 = ( ~n1750 & n8909 ) | ( ~n1750 & n8910 ) | ( n8909 & n8910 ) ;
  assign n8912 = ( ~n8907 & n8908 ) | ( ~n8907 & n8911 ) | ( n8908 & n8911 ) ;
  assign n8913 = ( ~x8 & n8907 ) | ( ~x8 & n8912 ) | ( n8907 & n8912 ) ;
  assign n8914 = ( n8907 & n8912 ) | ( n8907 & ~n8913 ) | ( n8912 & ~n8913 ) ;
  assign n8915 = ( x8 & n8913 ) | ( x8 & ~n8914 ) | ( n8913 & ~n8914 ) ;
  assign n8916 = ( n8904 & n8906 ) | ( n8904 & n8915 ) | ( n8906 & n8915 ) ;
  assign n8917 = ( n8530 & ~n8539 ) | ( n8530 & n8541 ) | ( ~n8539 & n8541 ) ;
  assign n8918 = ( ~n8530 & n8542 ) | ( ~n8530 & n8917 ) | ( n8542 & n8917 ) ;
  assign n8919 = ~n4159 & n7296 ;
  assign n8920 = n1458 & n7879 ;
  assign n8921 = n1669 | n7300 ;
  assign n8922 = n1576 & n7299 ;
  assign n8923 = ( ~n1669 & n8921 ) | ( ~n1669 & n8922 ) | ( n8921 & n8922 ) ;
  assign n8924 = ( ~n8919 & n8920 ) | ( ~n8919 & n8923 ) | ( n8920 & n8923 ) ;
  assign n8925 = ( ~x8 & n8919 ) | ( ~x8 & n8924 ) | ( n8919 & n8924 ) ;
  assign n8926 = ( n8919 & n8924 ) | ( n8919 & ~n8925 ) | ( n8924 & ~n8925 ) ;
  assign n8927 = ( x8 & n8925 ) | ( x8 & ~n8926 ) | ( n8925 & ~n8926 ) ;
  assign n8928 = ( n8916 & ~n8918 ) | ( n8916 & n8927 ) | ( ~n8918 & n8927 ) ;
  assign n8929 = ( ~n8542 & n8551 ) | ( ~n8542 & n8553 ) | ( n8551 & n8553 ) ;
  assign n8930 = ( n8542 & ~n8554 ) | ( n8542 & n8929 ) | ( ~n8554 & n8929 ) ;
  assign n8931 = ~n3955 & n7296 ;
  assign n8932 = ~n1338 & n7879 ;
  assign n8933 = n1458 & n7299 ;
  assign n8934 = n1576 & n7300 ;
  assign n8935 = n8933 | n8934 ;
  assign n8936 = ( ~n8931 & n8932 ) | ( ~n8931 & n8935 ) | ( n8932 & n8935 ) ;
  assign n8937 = ( ~x8 & n8931 ) | ( ~x8 & n8936 ) | ( n8931 & n8936 ) ;
  assign n8938 = ( n8931 & n8936 ) | ( n8931 & ~n8937 ) | ( n8936 & ~n8937 ) ;
  assign n8939 = ( x8 & n8937 ) | ( x8 & ~n8938 ) | ( n8937 & ~n8938 ) ;
  assign n8940 = ( n8928 & n8930 ) | ( n8928 & n8939 ) | ( n8930 & n8939 ) ;
  assign n8941 = ( ~n8554 & n8563 ) | ( ~n8554 & n8565 ) | ( n8563 & n8565 ) ;
  assign n8942 = ( n8554 & ~n8566 ) | ( n8554 & n8941 ) | ( ~n8566 & n8941 ) ;
  assign n8943 = ~n3779 & n7296 ;
  assign n8944 = n1267 & n7879 ;
  assign n8945 = n1458 & ~n7300 ;
  assign n8946 = ~n1338 & n7299 ;
  assign n8947 = ( n1458 & ~n8945 ) | ( n1458 & n8946 ) | ( ~n8945 & n8946 ) ;
  assign n8948 = ( ~n8943 & n8944 ) | ( ~n8943 & n8947 ) | ( n8944 & n8947 ) ;
  assign n8949 = ( ~x8 & n8943 ) | ( ~x8 & n8948 ) | ( n8943 & n8948 ) ;
  assign n8950 = ( n8943 & n8948 ) | ( n8943 & ~n8949 ) | ( n8948 & ~n8949 ) ;
  assign n8951 = ( x8 & n8949 ) | ( x8 & ~n8950 ) | ( n8949 & ~n8950 ) ;
  assign n8952 = ( n8940 & n8942 ) | ( n8940 & n8951 ) | ( n8942 & n8951 ) ;
  assign n8953 = ( n8566 & ~n8568 ) | ( n8566 & n8577 ) | ( ~n8568 & n8577 ) ;
  assign n8954 = ( n8568 & ~n8578 ) | ( n8568 & n8953 ) | ( ~n8578 & n8953 ) ;
  assign n8955 = n3692 & n8229 ;
  assign n8956 = ~n3658 & n8225 ;
  assign n8957 = ( n8229 & ~n8955 ) | ( n8229 & n8956 ) | ( ~n8955 & n8956 ) ;
  assign n8958 = n1290 | n8226 ;
  assign n8959 = ( ~n1290 & n8957 ) | ( ~n1290 & n8958 ) | ( n8957 & n8958 ) ;
  assign n8960 = ( ~n4182 & n8230 ) | ( ~n4182 & n8959 ) | ( n8230 & n8959 ) ;
  assign n8961 = n8959 & ~n8960 ;
  assign n8962 = ( ~x5 & n8960 ) | ( ~x5 & n8961 ) | ( n8960 & n8961 ) ;
  assign n8963 = ( n8960 & n8961 ) | ( n8960 & ~n8962 ) | ( n8961 & ~n8962 ) ;
  assign n8964 = ( x5 & n8962 ) | ( x5 & ~n8963 ) | ( n8962 & ~n8963 ) ;
  assign n8965 = ( n8952 & n8954 ) | ( n8952 & n8964 ) | ( n8954 & n8964 ) ;
  assign n8966 = x0 | x1 ;
  assign n8967 = x2 & ~n8966 ;
  assign n8968 = n36 & ~n3691 ;
  assign n8969 = ( ~n3692 & n8967 ) | ( ~n3692 & n8968 ) | ( n8967 & n8968 ) ;
  assign n8970 = x2 | n8969 ;
  assign n8971 = ( x2 & n8969 ) | ( x2 & ~n8970 ) | ( n8969 & ~n8970 ) ;
  assign n8972 = n8970 & ~n8971 ;
  assign n8973 = ~n3665 & n8230 ;
  assign n8974 = ~n1290 & n8225 ;
  assign n8975 = ~n1246 & n8226 ;
  assign n8976 = ~n3658 & n8229 ;
  assign n8977 = n8975 | n8976 ;
  assign n8978 = ( ~n8973 & n8974 ) | ( ~n8973 & n8977 ) | ( n8974 & n8977 ) ;
  assign n8979 = ( ~x5 & n8973 ) | ( ~x5 & n8978 ) | ( n8973 & n8978 ) ;
  assign n8980 = ( n8973 & n8978 ) | ( n8973 & ~n8979 ) | ( n8978 & ~n8979 ) ;
  assign n8981 = ( x5 & n8979 ) | ( x5 & ~n8980 ) | ( n8979 & ~n8980 ) ;
  assign n8982 = ( ~n8940 & n8942 ) | ( ~n8940 & n8951 ) | ( n8942 & n8951 ) ;
  assign n8983 = ( n8940 & ~n8952 ) | ( n8940 & n8982 ) | ( ~n8952 & n8982 ) ;
  assign n8984 = ( n8972 & n8981 ) | ( n8972 & n8983 ) | ( n8981 & n8983 ) ;
  assign n8985 = n6061 & n8230 ;
  assign n8986 = n3479 & n8225 ;
  assign n8987 = n3533 | n8226 ;
  assign n8988 = ~n3389 & n8229 ;
  assign n8989 = ( ~n3533 & n8987 ) | ( ~n3533 & n8988 ) | ( n8987 & n8988 ) ;
  assign n8990 = ( ~n8985 & n8986 ) | ( ~n8985 & n8989 ) | ( n8986 & n8989 ) ;
  assign n8991 = ( ~x5 & n8985 ) | ( ~x5 & n8990 ) | ( n8985 & n8990 ) ;
  assign n8992 = ( n8985 & n8990 ) | ( n8985 & ~n8991 ) | ( n8990 & ~n8991 ) ;
  assign n8993 = ( x5 & n8991 ) | ( x5 & ~n8992 ) | ( n8991 & ~n8992 ) ;
  assign n8994 = ( n3479 & n6009 ) | ( n3479 & n8230 ) | ( n6009 & n8230 ) ;
  assign n8995 = ~n3533 & n8225 ;
  assign n8996 = ~n3586 & n8226 ;
  assign n8997 = n8995 | n8996 ;
  assign n8998 = ~n3479 & n8229 ;
  assign n8999 = ( n8229 & n8997 ) | ( n8229 & ~n8998 ) | ( n8997 & ~n8998 ) ;
  assign n9000 = ( ~n6608 & n8994 ) | ( ~n6608 & n8999 ) | ( n8994 & n8999 ) ;
  assign n9001 = ~n3586 & n8228 ;
  assign n9002 = x5 & n9001 ;
  assign n9003 = ( n6009 & n6618 ) | ( n6009 & n8230 ) | ( n6618 & n8230 ) ;
  assign n9004 = ~n3533 & n8229 ;
  assign n9005 = n3586 | n8225 ;
  assign n9006 = ( ~n3586 & n9004 ) | ( ~n3586 & n9005 ) | ( n9004 & n9005 ) ;
  assign n9007 = n9003 | n9006 ;
  assign n9008 = ( x5 & n9002 ) | ( x5 & n9007 ) | ( n9002 & n9007 ) ;
  assign n9009 = n9000 | n9008 ;
  assign n9010 = x5 & ~n9009 ;
  assign n9011 = ( n8605 & n8993 ) | ( n8605 & n9010 ) | ( n8993 & n9010 ) ;
  assign n9012 = ~n3355 & n8229 ;
  assign n9013 = n3389 | n8225 ;
  assign n9014 = ( ~n3389 & n9012 ) | ( ~n3389 & n9013 ) | ( n9012 & n9013 ) ;
  assign n9015 = n3479 & ~n8226 ;
  assign n9016 = ( n3479 & n9014 ) | ( n3479 & ~n9015 ) | ( n9014 & ~n9015 ) ;
  assign n9017 = ( ~n6104 & n8230 ) | ( ~n6104 & n9016 ) | ( n8230 & n9016 ) ;
  assign n9018 = n9016 & ~n9017 ;
  assign n9019 = ( ~x5 & n9017 ) | ( ~x5 & n9018 ) | ( n9017 & n9018 ) ;
  assign n9020 = ( n9017 & n9018 ) | ( n9017 & ~n9019 ) | ( n9018 & ~n9019 ) ;
  assign n9021 = ( x5 & n9019 ) | ( x5 & ~n9020 ) | ( n9019 & ~n9020 ) ;
  assign n9022 = ( n8606 & n8607 ) | ( n8606 & n8610 ) | ( n8607 & n8610 ) ;
  assign n9023 = ~n8606 & n8611 ;
  assign n9024 = ( n8606 & ~n9022 ) | ( n8606 & n9023 ) | ( ~n9022 & n9023 ) ;
  assign n9025 = ( n9011 & n9021 ) | ( n9011 & n9024 ) | ( n9021 & n9024 ) ;
  assign n9026 = ~n6154 & n8230 ;
  assign n9027 = ~n3300 & n8229 ;
  assign n9028 = ~n3355 & n8225 ;
  assign n9029 = ~n3389 & n8226 ;
  assign n9030 = n9028 | n9029 ;
  assign n9031 = ( ~n9026 & n9027 ) | ( ~n9026 & n9030 ) | ( n9027 & n9030 ) ;
  assign n9032 = ( ~x5 & n9026 ) | ( ~x5 & n9031 ) | ( n9026 & n9031 ) ;
  assign n9033 = ( n9026 & n9031 ) | ( n9026 & ~n9032 ) | ( n9031 & ~n9032 ) ;
  assign n9034 = ( x5 & n9032 ) | ( x5 & ~n9033 ) | ( n9032 & ~n9033 ) ;
  assign n9035 = ( n8604 & n8612 ) | ( n8604 & ~n8613 ) | ( n8612 & ~n8613 ) ;
  assign n9036 = n8613 & ~n9035 ;
  assign n9037 = ( n9025 & n9034 ) | ( n9025 & n9036 ) | ( n9034 & n9036 ) ;
  assign n9038 = n6200 & n8230 ;
  assign n9039 = ~n3300 & n8225 ;
  assign n9040 = n3355 | n8226 ;
  assign n9041 = n3239 & n8229 ;
  assign n9042 = ( ~n3355 & n9040 ) | ( ~n3355 & n9041 ) | ( n9040 & n9041 ) ;
  assign n9043 = ( ~n9038 & n9039 ) | ( ~n9038 & n9042 ) | ( n9039 & n9042 ) ;
  assign n9044 = ( ~x5 & n9038 ) | ( ~x5 & n9043 ) | ( n9038 & n9043 ) ;
  assign n9045 = ( n9038 & n9043 ) | ( n9038 & ~n9044 ) | ( n9043 & ~n9044 ) ;
  assign n9046 = ( x5 & n9044 ) | ( x5 & ~n9045 ) | ( n9044 & ~n9045 ) ;
  assign n9047 = ( n8255 & n8597 ) | ( n8255 & ~n8614 ) | ( n8597 & ~n8614 ) ;
  assign n9048 = ( n8614 & ~n8615 ) | ( n8614 & n9047 ) | ( ~n8615 & n9047 ) ;
  assign n9049 = ( n9037 & n9046 ) | ( n9037 & n9048 ) | ( n9046 & n9048 ) ;
  assign n9050 = ~n6243 & n8230 ;
  assign n9051 = n3153 & n8229 ;
  assign n9052 = n3239 & n8225 ;
  assign n9053 = ~n3300 & n8226 ;
  assign n9054 = n9052 | n9053 ;
  assign n9055 = ( ~n9050 & n9051 ) | ( ~n9050 & n9054 ) | ( n9051 & n9054 ) ;
  assign n9056 = ( ~x5 & n9050 ) | ( ~x5 & n9055 ) | ( n9050 & n9055 ) ;
  assign n9057 = ( n9050 & n9055 ) | ( n9050 & ~n9056 ) | ( n9055 & ~n9056 ) ;
  assign n9058 = ( x5 & n9056 ) | ( x5 & ~n9057 ) | ( n9056 & ~n9057 ) ;
  assign n9059 = ( ~n8615 & n8624 ) | ( ~n8615 & n8627 ) | ( n8624 & n8627 ) ;
  assign n9060 = ( n8615 & ~n8628 ) | ( n8615 & n9059 ) | ( ~n8628 & n9059 ) ;
  assign n9061 = ( n9049 & n9058 ) | ( n9049 & n9060 ) | ( n9058 & n9060 ) ;
  assign n9062 = ( ~n8628 & n8637 ) | ( ~n8628 & n8639 ) | ( n8637 & n8639 ) ;
  assign n9063 = ( n8628 & ~n8640 ) | ( n8628 & n9062 ) | ( ~n8640 & n9062 ) ;
  assign n9064 = n5710 & n8230 ;
  assign n9065 = n3153 & n8225 ;
  assign n9066 = n3239 & ~n8226 ;
  assign n9067 = n3078 & n8229 ;
  assign n9068 = ( n3239 & ~n9066 ) | ( n3239 & n9067 ) | ( ~n9066 & n9067 ) ;
  assign n9069 = ( ~n9064 & n9065 ) | ( ~n9064 & n9068 ) | ( n9065 & n9068 ) ;
  assign n9070 = ( ~x5 & n9064 ) | ( ~x5 & n9069 ) | ( n9064 & n9069 ) ;
  assign n9071 = ( n9064 & n9069 ) | ( n9064 & ~n9070 ) | ( n9069 & ~n9070 ) ;
  assign n9072 = ( x5 & n9070 ) | ( x5 & ~n9071 ) | ( n9070 & ~n9071 ) ;
  assign n9073 = ( n9061 & n9063 ) | ( n9061 & n9072 ) | ( n9063 & n9072 ) ;
  assign n9074 = ( ~n8640 & n8649 ) | ( ~n8640 & n8651 ) | ( n8649 & n8651 ) ;
  assign n9075 = ( n8640 & ~n8652 ) | ( n8640 & n9074 ) | ( ~n8652 & n9074 ) ;
  assign n9076 = n3046 | n8229 ;
  assign n9077 = n3078 & n8225 ;
  assign n9078 = ( ~n3046 & n9076 ) | ( ~n3046 & n9077 ) | ( n9076 & n9077 ) ;
  assign n9079 = n3153 & ~n8226 ;
  assign n9080 = ( n3153 & n9078 ) | ( n3153 & ~n9079 ) | ( n9078 & ~n9079 ) ;
  assign n9081 = ( ~n6267 & n8230 ) | ( ~n6267 & n9080 ) | ( n8230 & n9080 ) ;
  assign n9082 = n9080 & ~n9081 ;
  assign n9083 = ( ~x5 & n9081 ) | ( ~x5 & n9082 ) | ( n9081 & n9082 ) ;
  assign n9084 = ( n9081 & n9082 ) | ( n9081 & ~n9083 ) | ( n9082 & ~n9083 ) ;
  assign n9085 = ( x5 & n9083 ) | ( x5 & ~n9084 ) | ( n9083 & ~n9084 ) ;
  assign n9086 = ( n9073 & n9075 ) | ( n9073 & n9085 ) | ( n9075 & n9085 ) ;
  assign n9087 = ( ~n8652 & n8661 ) | ( ~n8652 & n8663 ) | ( n8661 & n8663 ) ;
  assign n9088 = ( n8652 & ~n8664 ) | ( n8652 & n9087 ) | ( ~n8664 & n9087 ) ;
  assign n9089 = n6279 & n8230 ;
  assign n9090 = ~n2965 & n8229 ;
  assign n9091 = n3078 & n8226 ;
  assign n9092 = ~n3046 & n8225 ;
  assign n9093 = n9091 | n9092 ;
  assign n9094 = ( ~n9089 & n9090 ) | ( ~n9089 & n9093 ) | ( n9090 & n9093 ) ;
  assign n9095 = ( ~x5 & n9089 ) | ( ~x5 & n9094 ) | ( n9089 & n9094 ) ;
  assign n9096 = ( n9089 & n9094 ) | ( n9089 & ~n9095 ) | ( n9094 & ~n9095 ) ;
  assign n9097 = ( x5 & n9095 ) | ( x5 & ~n9096 ) | ( n9095 & ~n9096 ) ;
  assign n9098 = ( n9086 & n9088 ) | ( n9086 & n9097 ) | ( n9088 & n9097 ) ;
  assign n9099 = ~n5768 & n8230 ;
  assign n9100 = ~n2910 & n8229 ;
  assign n9101 = n3046 | n8226 ;
  assign n9102 = ~n2965 & n8225 ;
  assign n9103 = ( ~n3046 & n9101 ) | ( ~n3046 & n9102 ) | ( n9101 & n9102 ) ;
  assign n9104 = ( ~n9099 & n9100 ) | ( ~n9099 & n9103 ) | ( n9100 & n9103 ) ;
  assign n9105 = ( ~x5 & n9099 ) | ( ~x5 & n9104 ) | ( n9099 & n9104 ) ;
  assign n9106 = ( n9099 & n9104 ) | ( n9099 & ~n9105 ) | ( n9104 & ~n9105 ) ;
  assign n9107 = ( x5 & n9105 ) | ( x5 & ~n9106 ) | ( n9105 & ~n9106 ) ;
  assign n9108 = ( ~n8664 & n8666 ) | ( ~n8664 & n8675 ) | ( n8666 & n8675 ) ;
  assign n9109 = ( n8664 & ~n8676 ) | ( n8664 & n9108 ) | ( ~n8676 & n9108 ) ;
  assign n9110 = ( n9098 & n9107 ) | ( n9098 & n9109 ) | ( n9107 & n9109 ) ;
  assign n9111 = n5543 & n8230 ;
  assign n9112 = ~n2910 & n8225 ;
  assign n9113 = n2965 | n8226 ;
  assign n9114 = n2843 & n8229 ;
  assign n9115 = ( ~n2965 & n9113 ) | ( ~n2965 & n9114 ) | ( n9113 & n9114 ) ;
  assign n9116 = ( ~n9111 & n9112 ) | ( ~n9111 & n9115 ) | ( n9112 & n9115 ) ;
  assign n9117 = ( ~x5 & n9111 ) | ( ~x5 & n9116 ) | ( n9111 & n9116 ) ;
  assign n9118 = ( n9111 & n9116 ) | ( n9111 & ~n9117 ) | ( n9116 & ~n9117 ) ;
  assign n9119 = ( x5 & n9117 ) | ( x5 & ~n9118 ) | ( n9117 & ~n9118 ) ;
  assign n9120 = ( ~n8676 & n8678 ) | ( ~n8676 & n8687 ) | ( n8678 & n8687 ) ;
  assign n9121 = ( n8676 & ~n8688 ) | ( n8676 & n9120 ) | ( ~n8688 & n9120 ) ;
  assign n9122 = ( n9110 & n9119 ) | ( n9110 & n9121 ) | ( n9119 & n9121 ) ;
  assign n9123 = n5791 & n8230 ;
  assign n9124 = ~n2810 & n8229 ;
  assign n9125 = n2910 | n8226 ;
  assign n9126 = n2843 & n8225 ;
  assign n9127 = ( ~n2910 & n9125 ) | ( ~n2910 & n9126 ) | ( n9125 & n9126 ) ;
  assign n9128 = ( ~n9123 & n9124 ) | ( ~n9123 & n9127 ) | ( n9124 & n9127 ) ;
  assign n9129 = ( ~x5 & n9123 ) | ( ~x5 & n9128 ) | ( n9123 & n9128 ) ;
  assign n9130 = ( n9123 & n9128 ) | ( n9123 & ~n9129 ) | ( n9128 & ~n9129 ) ;
  assign n9131 = ( x5 & n9129 ) | ( x5 & ~n9130 ) | ( n9129 & ~n9130 ) ;
  assign n9132 = ( ~n8688 & n8690 ) | ( ~n8688 & n8699 ) | ( n8690 & n8699 ) ;
  assign n9133 = ( n8688 & ~n8700 ) | ( n8688 & n9132 ) | ( ~n8700 & n9132 ) ;
  assign n9134 = ( n9122 & n9131 ) | ( n9122 & n9133 ) | ( n9131 & n9133 ) ;
  assign n9135 = ( ~n8700 & n8709 ) | ( ~n8700 & n8711 ) | ( n8709 & n8711 ) ;
  assign n9136 = ( n8700 & ~n8712 ) | ( n8700 & n9135 ) | ( ~n8712 & n9135 ) ;
  assign n9137 = ~n5586 & n8230 ;
  assign n9138 = ~n2725 & n8229 ;
  assign n9139 = n2843 & n8226 ;
  assign n9140 = ~n2810 & n8225 ;
  assign n9141 = n9139 | n9140 ;
  assign n9142 = ( ~n9137 & n9138 ) | ( ~n9137 & n9141 ) | ( n9138 & n9141 ) ;
  assign n9143 = ( ~x5 & n9137 ) | ( ~x5 & n9142 ) | ( n9137 & n9142 ) ;
  assign n9144 = ( n9137 & n9142 ) | ( n9137 & ~n9143 ) | ( n9142 & ~n9143 ) ;
  assign n9145 = ( x5 & n9143 ) | ( x5 & ~n9144 ) | ( n9143 & ~n9144 ) ;
  assign n9146 = ( n9134 & n9136 ) | ( n9134 & n9145 ) | ( n9136 & n9145 ) ;
  assign n9147 = ( ~n8712 & n8721 ) | ( ~n8712 & n8723 ) | ( n8721 & n8723 ) ;
  assign n9148 = ( n8712 & ~n8724 ) | ( n8712 & n9147 ) | ( ~n8724 & n9147 ) ;
  assign n9149 = n2635 & ~n8229 ;
  assign n9150 = ~n2725 & n8225 ;
  assign n9151 = ( n2635 & ~n9149 ) | ( n2635 & n9150 ) | ( ~n9149 & n9150 ) ;
  assign n9152 = n2810 | n8226 ;
  assign n9153 = ( ~n2810 & n9151 ) | ( ~n2810 & n9152 ) | ( n9151 & n9152 ) ;
  assign n9154 = n5232 & n8230 ;
  assign n9155 = n9153 | n9154 ;
  assign n9156 = x5 | n9155 ;
  assign n9157 = ( x5 & n9155 ) | ( x5 & ~n9156 ) | ( n9155 & ~n9156 ) ;
  assign n9158 = n9156 & ~n9157 ;
  assign n9159 = ( n9146 & n9148 ) | ( n9146 & n9158 ) | ( n9148 & n9158 ) ;
  assign n9160 = ( ~n8724 & n8733 ) | ( ~n8724 & n8735 ) | ( n8733 & n8735 ) ;
  assign n9161 = ( n8724 & ~n8736 ) | ( n8724 & n9160 ) | ( ~n8736 & n9160 ) ;
  assign n9162 = ~n5425 & n8230 ;
  assign n9163 = n2552 & n8229 ;
  assign n9164 = ~n2725 & n8226 ;
  assign n9165 = n2635 & n8225 ;
  assign n9166 = n9164 | n9165 ;
  assign n9167 = ( ~n9162 & n9163 ) | ( ~n9162 & n9166 ) | ( n9163 & n9166 ) ;
  assign n9168 = ( ~x5 & n9162 ) | ( ~x5 & n9167 ) | ( n9162 & n9167 ) ;
  assign n9169 = ( n9162 & n9167 ) | ( n9162 & ~n9168 ) | ( n9167 & ~n9168 ) ;
  assign n9170 = ( x5 & n9168 ) | ( x5 & ~n9169 ) | ( n9168 & ~n9169 ) ;
  assign n9171 = ( n9159 & n9161 ) | ( n9159 & n9170 ) | ( n9161 & n9170 ) ;
  assign n9172 = ~n5270 & n8230 ;
  assign n9173 = n2552 & n8225 ;
  assign n9174 = n2635 & ~n8226 ;
  assign n9175 = ~n2491 & n8229 ;
  assign n9176 = ( n2635 & ~n9174 ) | ( n2635 & n9175 ) | ( ~n9174 & n9175 ) ;
  assign n9177 = ( ~n9172 & n9173 ) | ( ~n9172 & n9176 ) | ( n9173 & n9176 ) ;
  assign n9178 = ( ~x5 & n9172 ) | ( ~x5 & n9177 ) | ( n9172 & n9177 ) ;
  assign n9179 = ( n9172 & n9177 ) | ( n9172 & ~n9178 ) | ( n9177 & ~n9178 ) ;
  assign n9180 = ( x5 & n9178 ) | ( x5 & ~n9179 ) | ( n9178 & ~n9179 ) ;
  assign n9181 = ( ~n8736 & n8738 ) | ( ~n8736 & n8747 ) | ( n8738 & n8747 ) ;
  assign n9182 = ( n8736 & ~n8748 ) | ( n8736 & n9181 ) | ( ~n8748 & n9181 ) ;
  assign n9183 = ( n9171 & n9180 ) | ( n9171 & n9182 ) | ( n9180 & n9182 ) ;
  assign n9184 = ~n5084 & n8230 ;
  assign n9185 = n2396 & n8229 ;
  assign n9186 = ~n2491 & n8225 ;
  assign n9187 = n2552 & n8226 ;
  assign n9188 = n9186 | n9187 ;
  assign n9189 = ( ~n9184 & n9185 ) | ( ~n9184 & n9188 ) | ( n9185 & n9188 ) ;
  assign n9190 = ( ~x5 & n9184 ) | ( ~x5 & n9189 ) | ( n9184 & n9189 ) ;
  assign n9191 = ( n9184 & n9189 ) | ( n9184 & ~n9190 ) | ( n9189 & ~n9190 ) ;
  assign n9192 = ( x5 & n9190 ) | ( x5 & ~n9191 ) | ( n9190 & ~n9191 ) ;
  assign n9193 = ( ~n8748 & n8750 ) | ( ~n8748 & n8759 ) | ( n8750 & n8759 ) ;
  assign n9194 = ( n8748 & ~n8760 ) | ( n8748 & n9193 ) | ( ~n8760 & n9193 ) ;
  assign n9195 = ( n9183 & n9192 ) | ( n9183 & n9194 ) | ( n9192 & n9194 ) ;
  assign n9196 = ~n4900 & n8230 ;
  assign n9197 = n2396 & n8225 ;
  assign n9198 = ~n2298 & n8229 ;
  assign n9199 = ~n2491 & n8226 ;
  assign n9200 = n9198 | n9199 ;
  assign n9201 = ( ~n9196 & n9197 ) | ( ~n9196 & n9200 ) | ( n9197 & n9200 ) ;
  assign n9202 = ( ~x5 & n9196 ) | ( ~x5 & n9201 ) | ( n9196 & n9201 ) ;
  assign n9203 = ( n9196 & n9201 ) | ( n9196 & ~n9202 ) | ( n9201 & ~n9202 ) ;
  assign n9204 = ( x5 & n9202 ) | ( x5 & ~n9203 ) | ( n9202 & ~n9203 ) ;
  assign n9205 = ( ~n8760 & n8762 ) | ( ~n8760 & n8771 ) | ( n8762 & n8771 ) ;
  assign n9206 = ( n8760 & ~n8772 ) | ( n8760 & n9205 ) | ( ~n8772 & n9205 ) ;
  assign n9207 = ( n9195 & n9204 ) | ( n9195 & n9206 ) | ( n9204 & n9206 ) ;
  assign n9208 = ( ~n8772 & n8781 ) | ( ~n8772 & n8783 ) | ( n8781 & n8783 ) ;
  assign n9209 = ( n8772 & ~n8784 ) | ( n8772 & n9208 ) | ( ~n8784 & n9208 ) ;
  assign n9210 = n2270 & ~n8229 ;
  assign n9211 = ~n2298 & n8225 ;
  assign n9212 = ( n2270 & ~n9210 ) | ( n2270 & n9211 ) | ( ~n9210 & n9211 ) ;
  assign n9213 = n2396 & ~n8226 ;
  assign n9214 = ( n2396 & n9212 ) | ( n2396 & ~n9213 ) | ( n9212 & ~n9213 ) ;
  assign n9215 = ( ~n4912 & n8230 ) | ( ~n4912 & n9214 ) | ( n8230 & n9214 ) ;
  assign n9216 = n9214 & ~n9215 ;
  assign n9217 = ( ~x5 & n9215 ) | ( ~x5 & n9216 ) | ( n9215 & n9216 ) ;
  assign n9218 = ( n9215 & n9216 ) | ( n9215 & ~n9217 ) | ( n9216 & ~n9217 ) ;
  assign n9219 = ( x5 & n9217 ) | ( x5 & ~n9218 ) | ( n9217 & ~n9218 ) ;
  assign n9220 = ( n9207 & n9209 ) | ( n9207 & n9219 ) | ( n9209 & n9219 ) ;
  assign n9221 = ( ~n8784 & n8793 ) | ( ~n8784 & n8795 ) | ( n8793 & n8795 ) ;
  assign n9222 = ( n8784 & ~n8796 ) | ( n8784 & n9221 ) | ( ~n8796 & n9221 ) ;
  assign n9223 = n4647 & n8230 ;
  assign n9224 = n2174 & n8229 ;
  assign n9225 = n2298 | n8226 ;
  assign n9226 = n2270 & n8225 ;
  assign n9227 = ( ~n2298 & n9225 ) | ( ~n2298 & n9226 ) | ( n9225 & n9226 ) ;
  assign n9228 = ( ~n9223 & n9224 ) | ( ~n9223 & n9227 ) | ( n9224 & n9227 ) ;
  assign n9229 = ( ~x5 & n9223 ) | ( ~x5 & n9228 ) | ( n9223 & n9228 ) ;
  assign n9230 = ( n9223 & n9228 ) | ( n9223 & ~n9229 ) | ( n9228 & ~n9229 ) ;
  assign n9231 = ( x5 & n9229 ) | ( x5 & ~n9230 ) | ( n9229 & ~n9230 ) ;
  assign n9232 = ( n9220 & n9222 ) | ( n9220 & n9231 ) | ( n9222 & n9231 ) ;
  assign n9233 = ( ~n8796 & n8805 ) | ( ~n8796 & n8807 ) | ( n8805 & n8807 ) ;
  assign n9234 = ( n8796 & ~n8808 ) | ( n8796 & n9233 ) | ( ~n8808 & n9233 ) ;
  assign n9235 = n4730 & n8230 ;
  assign n9236 = n2089 & n8229 ;
  assign n9237 = n2270 & n8226 ;
  assign n9238 = n2174 & n8225 ;
  assign n9239 = n9237 | n9238 ;
  assign n9240 = ( ~n9235 & n9236 ) | ( ~n9235 & n9239 ) | ( n9236 & n9239 ) ;
  assign n9241 = ( ~x5 & n9235 ) | ( ~x5 & n9240 ) | ( n9235 & n9240 ) ;
  assign n9242 = ( n9235 & n9240 ) | ( n9235 & ~n9241 ) | ( n9240 & ~n9241 ) ;
  assign n9243 = ( x5 & n9241 ) | ( x5 & ~n9242 ) | ( n9241 & ~n9242 ) ;
  assign n9244 = ( n9232 & n9234 ) | ( n9232 & n9243 ) | ( n9234 & n9243 ) ;
  assign n9245 = ~n4660 & n8230 ;
  assign n9246 = ~n2023 & n8229 ;
  assign n9247 = n2174 & n8226 ;
  assign n9248 = n2089 & n8225 ;
  assign n9249 = n9247 | n9248 ;
  assign n9250 = ( ~n9245 & n9246 ) | ( ~n9245 & n9249 ) | ( n9246 & n9249 ) ;
  assign n9251 = ( ~x5 & n9245 ) | ( ~x5 & n9250 ) | ( n9245 & n9250 ) ;
  assign n9252 = ( n9245 & n9250 ) | ( n9245 & ~n9251 ) | ( n9250 & ~n9251 ) ;
  assign n9253 = ( x5 & n9251 ) | ( x5 & ~n9252 ) | ( n9251 & ~n9252 ) ;
  assign n9254 = ( ~n8808 & n8810 ) | ( ~n8808 & n8819 ) | ( n8810 & n8819 ) ;
  assign n9255 = ( n8808 & ~n8820 ) | ( n8808 & n9254 ) | ( ~n8820 & n9254 ) ;
  assign n9256 = ( n9244 & n9253 ) | ( n9244 & n9255 ) | ( n9253 & n9255 ) ;
  assign n9257 = ~n4457 & n8230 ;
  assign n9258 = n1926 & n8229 ;
  assign n9259 = ~n2023 & n8225 ;
  assign n9260 = n2089 & n8226 ;
  assign n9261 = n9259 | n9260 ;
  assign n9262 = ( ~n9257 & n9258 ) | ( ~n9257 & n9261 ) | ( n9258 & n9261 ) ;
  assign n9263 = ( ~x5 & n9257 ) | ( ~x5 & n9262 ) | ( n9257 & n9262 ) ;
  assign n9264 = ( n9257 & n9262 ) | ( n9257 & ~n9263 ) | ( n9262 & ~n9263 ) ;
  assign n9265 = ( x5 & n9263 ) | ( x5 & ~n9264 ) | ( n9263 & ~n9264 ) ;
  assign n9266 = ( ~n8820 & n8822 ) | ( ~n8820 & n8831 ) | ( n8822 & n8831 ) ;
  assign n9267 = ( n8820 & ~n8832 ) | ( n8820 & n9266 ) | ( ~n8832 & n9266 ) ;
  assign n9268 = ( n9256 & n9265 ) | ( n9256 & n9267 ) | ( n9265 & n9267 ) ;
  assign n9269 = n4290 & n8230 ;
  assign n9270 = n1852 & n8229 ;
  assign n9271 = ~n2023 & n8226 ;
  assign n9272 = n1926 & n8225 ;
  assign n9273 = n9271 | n9272 ;
  assign n9274 = ( ~n9269 & n9270 ) | ( ~n9269 & n9273 ) | ( n9270 & n9273 ) ;
  assign n9275 = ( ~x5 & n9269 ) | ( ~x5 & n9274 ) | ( n9269 & n9274 ) ;
  assign n9276 = ( n9269 & n9274 ) | ( n9269 & ~n9275 ) | ( n9274 & ~n9275 ) ;
  assign n9277 = ( x5 & n9275 ) | ( x5 & ~n9276 ) | ( n9275 & ~n9276 ) ;
  assign n9278 = ( ~n8832 & n8834 ) | ( ~n8832 & n8843 ) | ( n8834 & n8843 ) ;
  assign n9279 = ( n8832 & ~n8844 ) | ( n8832 & n9278 ) | ( ~n8844 & n9278 ) ;
  assign n9280 = ( n9268 & n9277 ) | ( n9268 & n9279 ) | ( n9277 & n9279 ) ;
  assign n9281 = ( ~n8844 & n8853 ) | ( ~n8844 & n8855 ) | ( n8853 & n8855 ) ;
  assign n9282 = ( n8844 & ~n8856 ) | ( n8844 & n9281 ) | ( ~n8856 & n9281 ) ;
  assign n9283 = ~n4302 & n8230 ;
  assign n9284 = ~n1750 & n8229 ;
  assign n9285 = n1852 & n8225 ;
  assign n9286 = n1926 & n8226 ;
  assign n9287 = n9285 | n9286 ;
  assign n9288 = ( ~n9283 & n9284 ) | ( ~n9283 & n9287 ) | ( n9284 & n9287 ) ;
  assign n9289 = ( ~x5 & n9283 ) | ( ~x5 & n9288 ) | ( n9283 & n9288 ) ;
  assign n9290 = ( n9283 & n9288 ) | ( n9283 & ~n9289 ) | ( n9288 & ~n9289 ) ;
  assign n9291 = ( x5 & n9289 ) | ( x5 & ~n9290 ) | ( n9289 & ~n9290 ) ;
  assign n9292 = ( n9280 & n9282 ) | ( n9280 & n9291 ) | ( n9282 & n9291 ) ;
  assign n9293 = ( ~n8856 & n8865 ) | ( ~n8856 & n8867 ) | ( n8865 & n8867 ) ;
  assign n9294 = ( n8856 & ~n8868 ) | ( n8856 & n9293 ) | ( ~n8868 & n9293 ) ;
  assign n9295 = n4146 & n8230 ;
  assign n9296 = ~n1669 & n8229 ;
  assign n9297 = n1852 & ~n8226 ;
  assign n9298 = ~n1750 & n8225 ;
  assign n9299 = ( n1852 & ~n9297 ) | ( n1852 & n9298 ) | ( ~n9297 & n9298 ) ;
  assign n9300 = ( ~n9295 & n9296 ) | ( ~n9295 & n9299 ) | ( n9296 & n9299 ) ;
  assign n9301 = ( ~x5 & n9295 ) | ( ~x5 & n9300 ) | ( n9295 & n9300 ) ;
  assign n9302 = ( n9295 & n9300 ) | ( n9295 & ~n9301 ) | ( n9300 & ~n9301 ) ;
  assign n9303 = ( x5 & n9301 ) | ( x5 & ~n9302 ) | ( n9301 & ~n9302 ) ;
  assign n9304 = ( n9292 & n9294 ) | ( n9292 & n9303 ) | ( n9294 & n9303 ) ;
  assign n9305 = n4326 & n8230 ;
  assign n9306 = n1576 & n8229 ;
  assign n9307 = n1750 | n8226 ;
  assign n9308 = ~n1669 & n8225 ;
  assign n9309 = ( ~n1750 & n9307 ) | ( ~n1750 & n9308 ) | ( n9307 & n9308 ) ;
  assign n9310 = ( ~n9305 & n9306 ) | ( ~n9305 & n9309 ) | ( n9306 & n9309 ) ;
  assign n9311 = ( ~x5 & n9305 ) | ( ~x5 & n9310 ) | ( n9305 & n9310 ) ;
  assign n9312 = ( n9305 & n9310 ) | ( n9305 & ~n9311 ) | ( n9310 & ~n9311 ) ;
  assign n9313 = ( x5 & n9311 ) | ( x5 & ~n9312 ) | ( n9311 & ~n9312 ) ;
  assign n9314 = ( ~n8868 & n8870 ) | ( ~n8868 & n8879 ) | ( n8870 & n8879 ) ;
  assign n9315 = ( n8868 & ~n8880 ) | ( n8868 & n9314 ) | ( ~n8880 & n9314 ) ;
  assign n9316 = ( n9304 & n9313 ) | ( n9304 & n9315 ) | ( n9313 & n9315 ) ;
  assign n9317 = ~n4159 & n8230 ;
  assign n9318 = n1458 & n8229 ;
  assign n9319 = ~n1669 & n8226 ;
  assign n9320 = n1576 & n8225 ;
  assign n9321 = n9319 | n9320 ;
  assign n9322 = ( ~n9317 & n9318 ) | ( ~n9317 & n9321 ) | ( n9318 & n9321 ) ;
  assign n9323 = ( ~x5 & n9317 ) | ( ~x5 & n9322 ) | ( n9317 & n9322 ) ;
  assign n9324 = ( n9317 & n9322 ) | ( n9317 & ~n9323 ) | ( n9322 & ~n9323 ) ;
  assign n9325 = ( x5 & n9323 ) | ( x5 & ~n9324 ) | ( n9323 & ~n9324 ) ;
  assign n9326 = ( ~n8880 & n8882 ) | ( ~n8880 & n8891 ) | ( n8882 & n8891 ) ;
  assign n9327 = ( ~n8891 & n8892 ) | ( ~n8891 & n9326 ) | ( n8892 & n9326 ) ;
  assign n9328 = ( n9316 & n9325 ) | ( n9316 & ~n9327 ) | ( n9325 & ~n9327 ) ;
  assign n9329 = ~n3955 & n8230 ;
  assign n9330 = ~n1338 & n8229 ;
  assign n9331 = n1458 & n8225 ;
  assign n9332 = n1576 & n8226 ;
  assign n9333 = n9331 | n9332 ;
  assign n9334 = ( ~n9329 & n9330 ) | ( ~n9329 & n9333 ) | ( n9330 & n9333 ) ;
  assign n9335 = ( ~x5 & n9329 ) | ( ~x5 & n9334 ) | ( n9329 & n9334 ) ;
  assign n9336 = ( n9329 & n9334 ) | ( n9329 & ~n9335 ) | ( n9334 & ~n9335 ) ;
  assign n9337 = ( x5 & n9335 ) | ( x5 & ~n9336 ) | ( n9335 & ~n9336 ) ;
  assign n9338 = ( ~n8892 & n8894 ) | ( ~n8892 & n8903 ) | ( n8894 & n8903 ) ;
  assign n9339 = ( ~n8903 & n8904 ) | ( ~n8903 & n9338 ) | ( n8904 & n9338 ) ;
  assign n9340 = ( n9328 & n9337 ) | ( n9328 & ~n9339 ) | ( n9337 & ~n9339 ) ;
  assign n9341 = ~n3779 & n8230 ;
  assign n9342 = n1267 & n8229 ;
  assign n9343 = n1458 & ~n8226 ;
  assign n9344 = ~n1338 & n8225 ;
  assign n9345 = ( n1458 & ~n9343 ) | ( n1458 & n9344 ) | ( ~n9343 & n9344 ) ;
  assign n9346 = ( ~n9341 & n9342 ) | ( ~n9341 & n9345 ) | ( n9342 & n9345 ) ;
  assign n9347 = ( ~x5 & n9341 ) | ( ~x5 & n9346 ) | ( n9341 & n9346 ) ;
  assign n9348 = ( n9341 & n9346 ) | ( n9341 & ~n9347 ) | ( n9346 & ~n9347 ) ;
  assign n9349 = ( x5 & n9347 ) | ( x5 & ~n9348 ) | ( n9347 & ~n9348 ) ;
  assign n9350 = ( ~n8904 & n8906 ) | ( ~n8904 & n8915 ) | ( n8906 & n8915 ) ;
  assign n9351 = ( n8904 & ~n8916 ) | ( n8904 & n9350 ) | ( ~n8916 & n9350 ) ;
  assign n9352 = ( n9340 & n9349 ) | ( n9340 & n9351 ) | ( n9349 & n9351 ) ;
  assign n9353 = ~n3791 & n8230 ;
  assign n9354 = n1267 & n8225 ;
  assign n9355 = n1338 | n8226 ;
  assign n9356 = ~n1246 & n8229 ;
  assign n9357 = ( ~n1338 & n9355 ) | ( ~n1338 & n9356 ) | ( n9355 & n9356 ) ;
  assign n9358 = ( ~n9353 & n9354 ) | ( ~n9353 & n9357 ) | ( n9354 & n9357 ) ;
  assign n9359 = ( ~x5 & n9353 ) | ( ~x5 & n9358 ) | ( n9353 & n9358 ) ;
  assign n9360 = ( n9353 & n9358 ) | ( n9353 & ~n9359 ) | ( n9358 & ~n9359 ) ;
  assign n9361 = ( x5 & n9359 ) | ( x5 & ~n9360 ) | ( n9359 & ~n9360 ) ;
  assign n9362 = ( ~n8916 & n8918 ) | ( ~n8916 & n8927 ) | ( n8918 & n8927 ) ;
  assign n9363 = ( ~n8927 & n8928 ) | ( ~n8927 & n9362 ) | ( n8928 & n9362 ) ;
  assign n9364 = ( n9352 & n9361 ) | ( n9352 & ~n9363 ) | ( n9361 & ~n9363 ) ;
  assign n9365 = n3621 & n8230 ;
  assign n9366 = ~n1290 & n8229 ;
  assign n9367 = ~n1246 & n8225 ;
  assign n9368 = n1267 & n8226 ;
  assign n9369 = n9367 | n9368 ;
  assign n9370 = ( ~n9365 & n9366 ) | ( ~n9365 & n9369 ) | ( n9366 & n9369 ) ;
  assign n9371 = ( ~x5 & n9365 ) | ( ~x5 & n9370 ) | ( n9365 & n9370 ) ;
  assign n9372 = ( n9365 & n9370 ) | ( n9365 & ~n9371 ) | ( n9370 & ~n9371 ) ;
  assign n9373 = ( x5 & n9371 ) | ( x5 & ~n9372 ) | ( n9371 & ~n9372 ) ;
  assign n9374 = ( ~n8928 & n8930 ) | ( ~n8928 & n8939 ) | ( n8930 & n8939 ) ;
  assign n9375 = ( n8928 & ~n8940 ) | ( n8928 & n9374 ) | ( ~n8940 & n9374 ) ;
  assign n9376 = ( n9364 & n9373 ) | ( n9364 & n9375 ) | ( n9373 & n9375 ) ;
  assign n9377 = n36 & n6200 ;
  assign n9378 = ~x0 & x1 ;
  assign n9379 = ~n3355 & n8967 ;
  assign n9380 = n35 & n3239 ;
  assign n9381 = n9379 | n9380 ;
  assign n9382 = n3300 & n9378 ;
  assign n9383 = ( n9378 & n9381 ) | ( n9378 & ~n9382 ) | ( n9381 & ~n9382 ) ;
  assign n9384 = ( ~x2 & n9377 ) | ( ~x2 & n9383 ) | ( n9377 & n9383 ) ;
  assign n9385 = ( n9377 & n9383 ) | ( n9377 & ~n9384 ) | ( n9383 & ~n9384 ) ;
  assign n9386 = ( x2 & n9384 ) | ( x2 & ~n9385 ) | ( n9384 & ~n9385 ) ;
  assign n9387 = n36 & ~n6104 ;
  assign n9388 = n35 & ~n3355 ;
  assign n9389 = ( ~x0 & n3389 ) | ( ~x0 & n8966 ) | ( n3389 & n8966 ) ;
  assign n9390 = ( ~n3389 & n9388 ) | ( ~n3389 & n9389 ) | ( n9388 & n9389 ) ;
  assign n9391 = n3479 & ~n8967 ;
  assign n9392 = ( n3479 & n9390 ) | ( n3479 & ~n9391 ) | ( n9390 & ~n9391 ) ;
  assign n9393 = ( ~x2 & n9387 ) | ( ~x2 & n9392 ) | ( n9387 & n9392 ) ;
  assign n9394 = ( n9387 & n9392 ) | ( n9387 & ~n9393 ) | ( n9392 & ~n9393 ) ;
  assign n9395 = ( x2 & n9393 ) | ( x2 & ~n9394 ) | ( n9393 & ~n9394 ) ;
  assign n9396 = ~n3533 & n8967 ;
  assign n9397 = n35 & n3389 ;
  assign n9398 = ( n35 & n9396 ) | ( n35 & ~n9397 ) | ( n9396 & ~n9397 ) ;
  assign n9399 = ~n3479 & n9378 ;
  assign n9400 = ( n9378 & n9398 ) | ( n9378 & ~n9399 ) | ( n9398 & ~n9399 ) ;
  assign n9401 = n36 & n6061 ;
  assign n9402 = n9400 | n9401 ;
  assign n9403 = x2 & ~n9402 ;
  assign n9404 = ( x0 & ~x1 ) | ( x0 & n36 ) | ( ~x1 & n36 ) ;
  assign n9405 = ( x0 & n3479 ) | ( x0 & n9404 ) | ( n3479 & n9404 ) ;
  assign n9406 = ( ~x0 & n35 ) | ( ~x0 & n8966 ) | ( n35 & n8966 ) ;
  assign n9407 = ( n3479 & n8966 ) | ( n3479 & n9406 ) | ( n8966 & n9406 ) ;
  assign n9408 = ( ~n3533 & n9405 ) | ( ~n3533 & n9407 ) | ( n9405 & n9407 ) ;
  assign n9409 = n3586 | n9408 ;
  assign n9410 = ( x2 & n9408 ) | ( x2 & ~n9409 ) | ( n9408 & ~n9409 ) ;
  assign n9411 = ( n9001 & n9402 ) | ( n9001 & n9403 ) | ( n9402 & n9403 ) ;
  assign n9412 = ( n9403 & ~n9410 ) | ( n9403 & n9411 ) | ( ~n9410 & n9411 ) ;
  assign n9413 = ( n9002 & n9003 ) | ( n9002 & n9006 ) | ( n9003 & n9006 ) ;
  assign n9414 = ~n9002 & n9007 ;
  assign n9415 = ( n9002 & ~n9413 ) | ( n9002 & n9414 ) | ( ~n9413 & n9414 ) ;
  assign n9416 = ( n9395 & n9412 ) | ( n9395 & n9415 ) | ( n9412 & n9415 ) ;
  assign n9417 = n36 & ~n6154 ;
  assign n9418 = ~n3355 & n9378 ;
  assign n9419 = ~n3389 & n8967 ;
  assign n9420 = n9418 | n9419 ;
  assign n9421 = n35 | n3300 ;
  assign n9422 = ( ~n3300 & n9420 ) | ( ~n3300 & n9421 ) | ( n9420 & n9421 ) ;
  assign n9423 = ( ~x2 & n9417 ) | ( ~x2 & n9422 ) | ( n9417 & n9422 ) ;
  assign n9424 = ( n9417 & n9422 ) | ( n9417 & ~n9423 ) | ( n9422 & ~n9423 ) ;
  assign n9425 = ( x2 & n9423 ) | ( x2 & ~n9424 ) | ( n9423 & ~n9424 ) ;
  assign n9426 = ~n9000 & n9008 ;
  assign n9427 = ( ~n9008 & n9009 ) | ( ~n9008 & n9426 ) | ( n9009 & n9426 ) ;
  assign n9428 = ( n9416 & n9425 ) | ( n9416 & n9427 ) | ( n9425 & n9427 ) ;
  assign n9429 = ( n8605 & n8993 ) | ( n8605 & ~n9010 ) | ( n8993 & ~n9010 ) ;
  assign n9430 = ( n9010 & ~n9011 ) | ( n9010 & n9429 ) | ( ~n9011 & n9429 ) ;
  assign n9431 = ( n9386 & n9428 ) | ( n9386 & n9430 ) | ( n9428 & n9430 ) ;
  assign n9432 = ( ~n9011 & n9021 ) | ( ~n9011 & n9024 ) | ( n9021 & n9024 ) ;
  assign n9433 = ( n9011 & ~n9025 ) | ( n9011 & n9432 ) | ( ~n9025 & n9432 ) ;
  assign n9434 = n36 & ~n6243 ;
  assign n9435 = n35 & n3153 ;
  assign n9436 = ( x0 & n3239 ) | ( x0 & ~n8966 ) | ( n3239 & ~n8966 ) ;
  assign n9437 = ( n3239 & n9435 ) | ( n3239 & ~n9436 ) | ( n9435 & ~n9436 ) ;
  assign n9438 = n3300 | n8967 ;
  assign n9439 = ( ~n3300 & n9437 ) | ( ~n3300 & n9438 ) | ( n9437 & n9438 ) ;
  assign n9440 = ( ~x2 & n9434 ) | ( ~x2 & n9439 ) | ( n9434 & n9439 ) ;
  assign n9441 = ( n9434 & n9439 ) | ( n9434 & ~n9440 ) | ( n9439 & ~n9440 ) ;
  assign n9442 = ( x2 & n9440 ) | ( x2 & ~n9441 ) | ( n9440 & ~n9441 ) ;
  assign n9443 = ( n9431 & n9433 ) | ( n9431 & n9442 ) | ( n9433 & n9442 ) ;
  assign n9444 = n36 & n5710 ;
  assign n9445 = n35 & n3078 ;
  assign n9446 = n3239 & n8967 ;
  assign n9447 = n9445 | n9446 ;
  assign n9448 = ~n3153 & n9378 ;
  assign n9449 = ( n9378 & n9447 ) | ( n9378 & ~n9448 ) | ( n9447 & ~n9448 ) ;
  assign n9450 = ( ~x2 & n9444 ) | ( ~x2 & n9449 ) | ( n9444 & n9449 ) ;
  assign n9451 = ( n9444 & n9449 ) | ( n9444 & ~n9450 ) | ( n9449 & ~n9450 ) ;
  assign n9452 = ( x2 & n9450 ) | ( x2 & ~n9451 ) | ( n9450 & ~n9451 ) ;
  assign n9453 = ( ~n9025 & n9034 ) | ( ~n9025 & n9036 ) | ( n9034 & n9036 ) ;
  assign n9454 = ( n9025 & ~n9037 ) | ( n9025 & n9453 ) | ( ~n9037 & n9453 ) ;
  assign n9455 = ( n9443 & n9452 ) | ( n9443 & n9454 ) | ( n9452 & n9454 ) ;
  assign n9456 = n36 & ~n6267 ;
  assign n9457 = n35 & ~n3046 ;
  assign n9458 = ( x0 & n3078 ) | ( x0 & ~n8966 ) | ( n3078 & ~n8966 ) ;
  assign n9459 = ( n3078 & n9457 ) | ( n3078 & ~n9458 ) | ( n9457 & ~n9458 ) ;
  assign n9460 = n3153 & ~n8967 ;
  assign n9461 = ( n3153 & n9459 ) | ( n3153 & ~n9460 ) | ( n9459 & ~n9460 ) ;
  assign n9462 = ( ~x2 & n9456 ) | ( ~x2 & n9461 ) | ( n9456 & n9461 ) ;
  assign n9463 = ( n9456 & n9461 ) | ( n9456 & ~n9462 ) | ( n9461 & ~n9462 ) ;
  assign n9464 = ( x2 & n9462 ) | ( x2 & ~n9463 ) | ( n9462 & ~n9463 ) ;
  assign n9465 = ( ~n9037 & n9046 ) | ( ~n9037 & n9048 ) | ( n9046 & n9048 ) ;
  assign n9466 = ( n9037 & ~n9049 ) | ( n9037 & n9465 ) | ( ~n9049 & n9465 ) ;
  assign n9467 = ( n9455 & n9464 ) | ( n9455 & n9466 ) | ( n9464 & n9466 ) ;
  assign n9468 = n36 & n6279 ;
  assign n9469 = n3078 & n8967 ;
  assign n9470 = ( x0 & n3046 ) | ( x0 & n8966 ) | ( n3046 & n8966 ) ;
  assign n9471 = ( n8966 & n9469 ) | ( n8966 & ~n9470 ) | ( n9469 & ~n9470 ) ;
  assign n9472 = n35 | n2965 ;
  assign n9473 = ( ~n2965 & n9471 ) | ( ~n2965 & n9472 ) | ( n9471 & n9472 ) ;
  assign n9474 = ( ~x2 & n9468 ) | ( ~x2 & n9473 ) | ( n9468 & n9473 ) ;
  assign n9475 = ( n9468 & n9473 ) | ( n9468 & ~n9474 ) | ( n9473 & ~n9474 ) ;
  assign n9476 = ( x2 & n9474 ) | ( x2 & ~n9475 ) | ( n9474 & ~n9475 ) ;
  assign n9477 = ( ~n9049 & n9058 ) | ( ~n9049 & n9060 ) | ( n9058 & n9060 ) ;
  assign n9478 = ( n9049 & ~n9061 ) | ( n9049 & n9477 ) | ( ~n9061 & n9477 ) ;
  assign n9479 = ( n9467 & n9476 ) | ( n9467 & n9478 ) | ( n9476 & n9478 ) ;
  assign n9480 = ( ~n9061 & n9063 ) | ( ~n9061 & n9072 ) | ( n9063 & n9072 ) ;
  assign n9481 = ( n9061 & ~n9073 ) | ( n9061 & n9480 ) | ( ~n9073 & n9480 ) ;
  assign n9482 = n36 & ~n5768 ;
  assign n9483 = ~n3046 & n8967 ;
  assign n9484 = ( x0 & n2965 ) | ( x0 & n8966 ) | ( n2965 & n8966 ) ;
  assign n9485 = ( n8966 & n9483 ) | ( n8966 & ~n9484 ) | ( n9483 & ~n9484 ) ;
  assign n9486 = n35 | n2910 ;
  assign n9487 = ( ~n2910 & n9485 ) | ( ~n2910 & n9486 ) | ( n9485 & n9486 ) ;
  assign n9488 = ( ~x2 & n9482 ) | ( ~x2 & n9487 ) | ( n9482 & n9487 ) ;
  assign n9489 = ( n9482 & n9487 ) | ( n9482 & ~n9488 ) | ( n9487 & ~n9488 ) ;
  assign n9490 = ( x2 & n9488 ) | ( x2 & ~n9489 ) | ( n9488 & ~n9489 ) ;
  assign n9491 = ( n9479 & n9481 ) | ( n9479 & n9490 ) | ( n9481 & n9490 ) ;
  assign n9492 = ( ~n9073 & n9075 ) | ( ~n9073 & n9085 ) | ( n9075 & n9085 ) ;
  assign n9493 = ( n9073 & ~n9086 ) | ( n9073 & n9492 ) | ( ~n9086 & n9492 ) ;
  assign n9494 = n36 & n5543 ;
  assign n9495 = ~n2965 & n8967 ;
  assign n9496 = n35 & n2843 ;
  assign n9497 = n9495 | n9496 ;
  assign n9498 = n2910 & n9378 ;
  assign n9499 = ( n9378 & n9497 ) | ( n9378 & ~n9498 ) | ( n9497 & ~n9498 ) ;
  assign n9500 = ( ~x2 & n9494 ) | ( ~x2 & n9499 ) | ( n9494 & n9499 ) ;
  assign n9501 = ( n9494 & n9499 ) | ( n9494 & ~n9500 ) | ( n9499 & ~n9500 ) ;
  assign n9502 = ( x2 & n9500 ) | ( x2 & ~n9501 ) | ( n9500 & ~n9501 ) ;
  assign n9503 = ( n9491 & n9493 ) | ( n9491 & n9502 ) | ( n9493 & n9502 ) ;
  assign n9504 = ( ~n9086 & n9088 ) | ( ~n9086 & n9097 ) | ( n9088 & n9097 ) ;
  assign n9505 = ( n9086 & ~n9098 ) | ( n9086 & n9504 ) | ( ~n9098 & n9504 ) ;
  assign n9506 = n36 & n5791 ;
  assign n9507 = ~n2910 & n8967 ;
  assign n9508 = ( x0 & ~n2843 ) | ( x0 & n8966 ) | ( ~n2843 & n8966 ) ;
  assign n9509 = ( n8966 & n9507 ) | ( n8966 & ~n9508 ) | ( n9507 & ~n9508 ) ;
  assign n9510 = n35 | n2810 ;
  assign n9511 = ( ~n2810 & n9509 ) | ( ~n2810 & n9510 ) | ( n9509 & n9510 ) ;
  assign n9512 = ( ~x2 & n9506 ) | ( ~x2 & n9511 ) | ( n9506 & n9511 ) ;
  assign n9513 = ( n9506 & n9511 ) | ( n9506 & ~n9512 ) | ( n9511 & ~n9512 ) ;
  assign n9514 = ( x2 & n9512 ) | ( x2 & ~n9513 ) | ( n9512 & ~n9513 ) ;
  assign n9515 = ( n9503 & n9505 ) | ( n9503 & n9514 ) | ( n9505 & n9514 ) ;
  assign n9516 = n36 & ~n5586 ;
  assign n9517 = n2843 & n8967 ;
  assign n9518 = ( x0 & n2810 ) | ( x0 & n8966 ) | ( n2810 & n8966 ) ;
  assign n9519 = ( n8966 & n9517 ) | ( n8966 & ~n9518 ) | ( n9517 & ~n9518 ) ;
  assign n9520 = n35 | n2725 ;
  assign n9521 = ( ~n2725 & n9519 ) | ( ~n2725 & n9520 ) | ( n9519 & n9520 ) ;
  assign n9522 = ( ~x2 & n9516 ) | ( ~x2 & n9521 ) | ( n9516 & n9521 ) ;
  assign n9523 = ( n9516 & n9521 ) | ( n9516 & ~n9522 ) | ( n9521 & ~n9522 ) ;
  assign n9524 = ( x2 & n9522 ) | ( x2 & ~n9523 ) | ( n9522 & ~n9523 ) ;
  assign n9525 = ( ~n9098 & n9107 ) | ( ~n9098 & n9109 ) | ( n9107 & n9109 ) ;
  assign n9526 = ( n9098 & ~n9110 ) | ( n9098 & n9525 ) | ( ~n9110 & n9525 ) ;
  assign n9527 = ( n9515 & n9524 ) | ( n9515 & n9526 ) | ( n9524 & n9526 ) ;
  assign n9528 = n36 & n5232 ;
  assign n9529 = n2810 | n8967 ;
  assign n9530 = n35 & n2635 ;
  assign n9531 = ( n9406 & ~n9520 ) | ( n9406 & n9530 ) | ( ~n9520 & n9530 ) ;
  assign n9532 = ( ~n2810 & n9529 ) | ( ~n2810 & n9531 ) | ( n9529 & n9531 ) ;
  assign n9533 = ( ~x2 & n9528 ) | ( ~x2 & n9532 ) | ( n9528 & n9532 ) ;
  assign n9534 = ( n9528 & n9532 ) | ( n9528 & ~n9533 ) | ( n9532 & ~n9533 ) ;
  assign n9535 = ( x2 & n9533 ) | ( x2 & ~n9534 ) | ( n9533 & ~n9534 ) ;
  assign n9536 = ( ~n9110 & n9119 ) | ( ~n9110 & n9121 ) | ( n9119 & n9121 ) ;
  assign n9537 = ( n9110 & ~n9122 ) | ( n9110 & n9536 ) | ( ~n9122 & n9536 ) ;
  assign n9538 = ( n9527 & n9535 ) | ( n9527 & n9537 ) | ( n9535 & n9537 ) ;
  assign n9539 = n36 & ~n5425 ;
  assign n9540 = ~n2725 & n8967 ;
  assign n9541 = ( x0 & ~n2635 ) | ( x0 & n8966 ) | ( ~n2635 & n8966 ) ;
  assign n9542 = ( n8966 & n9540 ) | ( n8966 & ~n9541 ) | ( n9540 & ~n9541 ) ;
  assign n9543 = ~n35 & n2552 ;
  assign n9544 = ( n2552 & n9542 ) | ( n2552 & ~n9543 ) | ( n9542 & ~n9543 ) ;
  assign n9545 = ( ~x2 & n9539 ) | ( ~x2 & n9544 ) | ( n9539 & n9544 ) ;
  assign n9546 = ( n9539 & n9544 ) | ( n9539 & ~n9545 ) | ( n9544 & ~n9545 ) ;
  assign n9547 = ( x2 & n9545 ) | ( x2 & ~n9546 ) | ( n9545 & ~n9546 ) ;
  assign n9548 = ( ~n9122 & n9131 ) | ( ~n9122 & n9133 ) | ( n9131 & n9133 ) ;
  assign n9549 = ( n9122 & ~n9134 ) | ( n9122 & n9548 ) | ( ~n9134 & n9548 ) ;
  assign n9550 = ( n9538 & n9547 ) | ( n9538 & n9549 ) | ( n9547 & n9549 ) ;
  assign n9551 = ( ~n9134 & n9136 ) | ( ~n9134 & n9145 ) | ( n9136 & n9145 ) ;
  assign n9552 = ( n9134 & ~n9146 ) | ( n9134 & n9551 ) | ( ~n9146 & n9551 ) ;
  assign n9553 = n36 & ~n5270 ;
  assign n9554 = n35 & ~n2491 ;
  assign n9555 = n2635 & n8967 ;
  assign n9556 = n9554 | n9555 ;
  assign n9557 = ~n2552 & n9378 ;
  assign n9558 = ( n9378 & n9556 ) | ( n9378 & ~n9557 ) | ( n9556 & ~n9557 ) ;
  assign n9559 = ( ~x2 & n9553 ) | ( ~x2 & n9558 ) | ( n9553 & n9558 ) ;
  assign n9560 = ( n9553 & n9558 ) | ( n9553 & ~n9559 ) | ( n9558 & ~n9559 ) ;
  assign n9561 = ( x2 & n9559 ) | ( x2 & ~n9560 ) | ( n9559 & ~n9560 ) ;
  assign n9562 = ( n9550 & n9552 ) | ( n9550 & n9561 ) | ( n9552 & n9561 ) ;
  assign n9563 = ( ~n9146 & n9148 ) | ( ~n9146 & n9158 ) | ( n9148 & n9158 ) ;
  assign n9564 = ( n9146 & ~n9159 ) | ( n9146 & n9563 ) | ( ~n9159 & n9563 ) ;
  assign n9565 = n36 & ~n5084 ;
  assign n9566 = ~n2491 & n9378 ;
  assign n9567 = n2552 & n8967 ;
  assign n9568 = n9566 | n9567 ;
  assign n9569 = ~n35 & n2396 ;
  assign n9570 = ( n2396 & n9568 ) | ( n2396 & ~n9569 ) | ( n9568 & ~n9569 ) ;
  assign n9571 = ( ~x2 & n9565 ) | ( ~x2 & n9570 ) | ( n9565 & n9570 ) ;
  assign n9572 = ( n9565 & n9570 ) | ( n9565 & ~n9571 ) | ( n9570 & ~n9571 ) ;
  assign n9573 = ( x2 & n9571 ) | ( x2 & ~n9572 ) | ( n9571 & ~n9572 ) ;
  assign n9574 = ( n9562 & n9564 ) | ( n9562 & n9573 ) | ( n9564 & n9573 ) ;
  assign n9575 = ( ~n9159 & n9161 ) | ( ~n9159 & n9170 ) | ( n9161 & n9170 ) ;
  assign n9576 = ( n9159 & ~n9171 ) | ( n9159 & n9575 ) | ( ~n9171 & n9575 ) ;
  assign n9577 = n36 & ~n4900 ;
  assign n9578 = n35 & ~n2298 ;
  assign n9579 = ~n2491 & n8967 ;
  assign n9580 = n9578 | n9579 ;
  assign n9581 = ~n2396 & n9378 ;
  assign n9582 = ( n9378 & n9580 ) | ( n9378 & ~n9581 ) | ( n9580 & ~n9581 ) ;
  assign n9583 = ( ~x2 & n9577 ) | ( ~x2 & n9582 ) | ( n9577 & n9582 ) ;
  assign n9584 = ( n9577 & n9582 ) | ( n9577 & ~n9583 ) | ( n9582 & ~n9583 ) ;
  assign n9585 = ( x2 & n9583 ) | ( x2 & ~n9584 ) | ( n9583 & ~n9584 ) ;
  assign n9586 = ( n9574 & n9576 ) | ( n9574 & n9585 ) | ( n9576 & n9585 ) ;
  assign n9587 = n36 & ~n4912 ;
  assign n9588 = n35 & n2270 ;
  assign n9589 = ( ~x0 & n2298 ) | ( ~x0 & n8966 ) | ( n2298 & n8966 ) ;
  assign n9590 = ( ~n2298 & n9588 ) | ( ~n2298 & n9589 ) | ( n9588 & n9589 ) ;
  assign n9591 = n2396 & ~n8967 ;
  assign n9592 = ( n2396 & n9590 ) | ( n2396 & ~n9591 ) | ( n9590 & ~n9591 ) ;
  assign n9593 = ( ~x2 & n9587 ) | ( ~x2 & n9592 ) | ( n9587 & n9592 ) ;
  assign n9594 = ( n9587 & n9592 ) | ( n9587 & ~n9593 ) | ( n9592 & ~n9593 ) ;
  assign n9595 = ( x2 & n9593 ) | ( x2 & ~n9594 ) | ( n9593 & ~n9594 ) ;
  assign n9596 = ( ~n9171 & n9180 ) | ( ~n9171 & n9182 ) | ( n9180 & n9182 ) ;
  assign n9597 = ( n9171 & ~n9183 ) | ( n9171 & n9596 ) | ( ~n9183 & n9596 ) ;
  assign n9598 = ( n9586 & n9595 ) | ( n9586 & n9597 ) | ( n9595 & n9597 ) ;
  assign n9599 = n36 & n4647 ;
  assign n9600 = ~n2298 & n8967 ;
  assign n9601 = ( x0 & ~n2270 ) | ( x0 & n8966 ) | ( ~n2270 & n8966 ) ;
  assign n9602 = ( n8966 & n9600 ) | ( n8966 & ~n9601 ) | ( n9600 & ~n9601 ) ;
  assign n9603 = ~n35 & n2174 ;
  assign n9604 = ( n2174 & n9602 ) | ( n2174 & ~n9603 ) | ( n9602 & ~n9603 ) ;
  assign n9605 = ( ~x2 & n9599 ) | ( ~x2 & n9604 ) | ( n9599 & n9604 ) ;
  assign n9606 = ( n9599 & n9604 ) | ( n9599 & ~n9605 ) | ( n9604 & ~n9605 ) ;
  assign n9607 = ( x2 & n9605 ) | ( x2 & ~n9606 ) | ( n9605 & ~n9606 ) ;
  assign n9608 = ( ~n9183 & n9192 ) | ( ~n9183 & n9194 ) | ( n9192 & n9194 ) ;
  assign n9609 = ( n9183 & ~n9195 ) | ( n9183 & n9608 ) | ( ~n9195 & n9608 ) ;
  assign n9610 = ( n9598 & n9607 ) | ( n9598 & n9609 ) | ( n9607 & n9609 ) ;
  assign n9611 = n36 & n4730 ;
  assign n9612 = n2270 & n8967 ;
  assign n9613 = ( x0 & ~n2174 ) | ( x0 & n8966 ) | ( ~n2174 & n8966 ) ;
  assign n9614 = ( n8966 & n9612 ) | ( n8966 & ~n9613 ) | ( n9612 & ~n9613 ) ;
  assign n9615 = ~n35 & n2089 ;
  assign n9616 = ( n2089 & n9614 ) | ( n2089 & ~n9615 ) | ( n9614 & ~n9615 ) ;
  assign n9617 = ( ~x2 & n9611 ) | ( ~x2 & n9616 ) | ( n9611 & n9616 ) ;
  assign n9618 = ( n9611 & n9616 ) | ( n9611 & ~n9617 ) | ( n9616 & ~n9617 ) ;
  assign n9619 = ( x2 & n9617 ) | ( x2 & ~n9618 ) | ( n9617 & ~n9618 ) ;
  assign n9620 = ( ~n9195 & n9204 ) | ( ~n9195 & n9206 ) | ( n9204 & n9206 ) ;
  assign n9621 = ( n9195 & ~n9207 ) | ( n9195 & n9620 ) | ( ~n9207 & n9620 ) ;
  assign n9622 = ( n9610 & n9619 ) | ( n9610 & n9621 ) | ( n9619 & n9621 ) ;
  assign n9623 = ( ~n9207 & n9209 ) | ( ~n9207 & n9219 ) | ( n9209 & n9219 ) ;
  assign n9624 = ( n9207 & ~n9220 ) | ( n9207 & n9623 ) | ( ~n9220 & n9623 ) ;
  assign n9625 = n36 & ~n4660 ;
  assign n9626 = n2174 & n8967 ;
  assign n9627 = ( n35 & n2089 ) | ( n35 & n9406 ) | ( n2089 & n9406 ) ;
  assign n9628 = x0 & n2023 ;
  assign n9629 = ( n9626 & n9627 ) | ( n9626 & ~n9628 ) | ( n9627 & ~n9628 ) ;
  assign n9630 = ( ~x2 & n9625 ) | ( ~x2 & n9629 ) | ( n9625 & n9629 ) ;
  assign n9631 = ( n9625 & n9629 ) | ( n9625 & ~n9630 ) | ( n9629 & ~n9630 ) ;
  assign n9632 = ( x2 & n9630 ) | ( x2 & ~n9631 ) | ( n9630 & ~n9631 ) ;
  assign n9633 = ( n9622 & n9624 ) | ( n9622 & n9632 ) | ( n9624 & n9632 ) ;
  assign n9634 = ( ~n9220 & n9222 ) | ( ~n9220 & n9231 ) | ( n9222 & n9231 ) ;
  assign n9635 = ( n9220 & ~n9232 ) | ( n9220 & n9634 ) | ( ~n9232 & n9634 ) ;
  assign n9636 = n36 & ~n4457 ;
  assign n9637 = ~n2023 & n9378 ;
  assign n9638 = n2089 & n8967 ;
  assign n9639 = n9637 | n9638 ;
  assign n9640 = ~n35 & n1926 ;
  assign n9641 = ( n1926 & n9639 ) | ( n1926 & ~n9640 ) | ( n9639 & ~n9640 ) ;
  assign n9642 = ( ~x2 & n9636 ) | ( ~x2 & n9641 ) | ( n9636 & n9641 ) ;
  assign n9643 = ( n9636 & n9641 ) | ( n9636 & ~n9642 ) | ( n9641 & ~n9642 ) ;
  assign n9644 = ( x2 & n9642 ) | ( x2 & ~n9643 ) | ( n9642 & ~n9643 ) ;
  assign n9645 = ( n9633 & n9635 ) | ( n9633 & n9644 ) | ( n9635 & n9644 ) ;
  assign n9646 = ( ~n9232 & n9234 ) | ( ~n9232 & n9243 ) | ( n9234 & n9243 ) ;
  assign n9647 = ( n9232 & ~n9244 ) | ( n9232 & n9646 ) | ( ~n9244 & n9646 ) ;
  assign n9648 = n36 & n4290 ;
  assign n9649 = ~n2023 & n8967 ;
  assign n9650 = ( x0 & ~n1926 ) | ( x0 & n8966 ) | ( ~n1926 & n8966 ) ;
  assign n9651 = ( n8966 & n9649 ) | ( n8966 & ~n9650 ) | ( n9649 & ~n9650 ) ;
  assign n9652 = ~n35 & n1852 ;
  assign n9653 = ( n1852 & n9651 ) | ( n1852 & ~n9652 ) | ( n9651 & ~n9652 ) ;
  assign n9654 = ( ~x2 & n9648 ) | ( ~x2 & n9653 ) | ( n9648 & n9653 ) ;
  assign n9655 = ( n9648 & n9653 ) | ( n9648 & ~n9654 ) | ( n9653 & ~n9654 ) ;
  assign n9656 = ( x2 & n9654 ) | ( x2 & ~n9655 ) | ( n9654 & ~n9655 ) ;
  assign n9657 = ( n9645 & n9647 ) | ( n9645 & n9656 ) | ( n9647 & n9656 ) ;
  assign n9658 = n36 & ~n4302 ;
  assign n9659 = n1852 & n9378 ;
  assign n9660 = n1926 & n8967 ;
  assign n9661 = n9659 | n9660 ;
  assign n9662 = n35 | n1750 ;
  assign n9663 = ( ~n1750 & n9661 ) | ( ~n1750 & n9662 ) | ( n9661 & n9662 ) ;
  assign n9664 = ( ~x2 & n9658 ) | ( ~x2 & n9663 ) | ( n9658 & n9663 ) ;
  assign n9665 = ( n9658 & n9663 ) | ( n9658 & ~n9664 ) | ( n9663 & ~n9664 ) ;
  assign n9666 = ( x2 & n9664 ) | ( x2 & ~n9665 ) | ( n9664 & ~n9665 ) ;
  assign n9667 = ( ~n9244 & n9253 ) | ( ~n9244 & n9255 ) | ( n9253 & n9255 ) ;
  assign n9668 = ( n9244 & ~n9256 ) | ( n9244 & n9667 ) | ( ~n9256 & n9667 ) ;
  assign n9669 = ( n9657 & n9666 ) | ( n9657 & n9668 ) | ( n9666 & n9668 ) ;
  assign n9670 = n36 & n4146 ;
  assign n9671 = n1852 & n8967 ;
  assign n9672 = ( x0 & n1750 ) | ( x0 & n8966 ) | ( n1750 & n8966 ) ;
  assign n9673 = ( n8966 & n9671 ) | ( n8966 & ~n9672 ) | ( n9671 & ~n9672 ) ;
  assign n9674 = n35 | n1669 ;
  assign n9675 = ( ~n1669 & n9673 ) | ( ~n1669 & n9674 ) | ( n9673 & n9674 ) ;
  assign n9676 = ( ~x2 & n9670 ) | ( ~x2 & n9675 ) | ( n9670 & n9675 ) ;
  assign n9677 = ( n9670 & n9675 ) | ( n9670 & ~n9676 ) | ( n9675 & ~n9676 ) ;
  assign n9678 = ( x2 & n9676 ) | ( x2 & ~n9677 ) | ( n9676 & ~n9677 ) ;
  assign n9679 = ( ~n9256 & n9265 ) | ( ~n9256 & n9267 ) | ( n9265 & n9267 ) ;
  assign n9680 = ( n9256 & ~n9268 ) | ( n9256 & n9679 ) | ( ~n9268 & n9679 ) ;
  assign n9681 = ( n9669 & n9678 ) | ( n9669 & n9680 ) | ( n9678 & n9680 ) ;
  assign n9682 = n36 & n4326 ;
  assign n9683 = ~n1750 & n8967 ;
  assign n9684 = ( x0 & n1669 ) | ( x0 & n8966 ) | ( n1669 & n8966 ) ;
  assign n9685 = ( n8966 & n9683 ) | ( n8966 & ~n9684 ) | ( n9683 & ~n9684 ) ;
  assign n9686 = ~n35 & n1576 ;
  assign n9687 = ( n1576 & n9685 ) | ( n1576 & ~n9686 ) | ( n9685 & ~n9686 ) ;
  assign n9688 = ( ~x2 & n9682 ) | ( ~x2 & n9687 ) | ( n9682 & n9687 ) ;
  assign n9689 = ( n9682 & n9687 ) | ( n9682 & ~n9688 ) | ( n9687 & ~n9688 ) ;
  assign n9690 = ( x2 & n9688 ) | ( x2 & ~n9689 ) | ( n9688 & ~n9689 ) ;
  assign n9691 = ( ~n9268 & n9277 ) | ( ~n9268 & n9279 ) | ( n9277 & n9279 ) ;
  assign n9692 = ( n9268 & ~n9280 ) | ( n9268 & n9691 ) | ( ~n9280 & n9691 ) ;
  assign n9693 = ( n9681 & n9690 ) | ( n9681 & n9692 ) | ( n9690 & n9692 ) ;
  assign n9694 = ( ~n9280 & n9282 ) | ( ~n9280 & n9291 ) | ( n9282 & n9291 ) ;
  assign n9695 = ( n9280 & ~n9292 ) | ( n9280 & n9694 ) | ( ~n9292 & n9694 ) ;
  assign n9696 = n36 & ~n4159 ;
  assign n9697 = ~n1669 & n8967 ;
  assign n9698 = n35 & ~n1458 ;
  assign n9699 = ( n35 & n9697 ) | ( n35 & ~n9698 ) | ( n9697 & ~n9698 ) ;
  assign n9700 = ~n1576 & n9378 ;
  assign n9701 = ( n9378 & n9699 ) | ( n9378 & ~n9700 ) | ( n9699 & ~n9700 ) ;
  assign n9702 = ( ~x2 & n9696 ) | ( ~x2 & n9701 ) | ( n9696 & n9701 ) ;
  assign n9703 = ( n9696 & n9701 ) | ( n9696 & ~n9702 ) | ( n9701 & ~n9702 ) ;
  assign n9704 = ( x2 & n9702 ) | ( x2 & ~n9703 ) | ( n9702 & ~n9703 ) ;
  assign n9705 = ( n9693 & n9695 ) | ( n9693 & n9704 ) | ( n9695 & n9704 ) ;
  assign n9706 = ( ~n9292 & n9294 ) | ( ~n9292 & n9303 ) | ( n9294 & n9303 ) ;
  assign n9707 = ( n9292 & ~n9304 ) | ( n9292 & n9706 ) | ( ~n9304 & n9706 ) ;
  assign n9708 = n36 & ~n3955 ;
  assign n9709 = n35 & n1338 ;
  assign n9710 = n1458 & n9378 ;
  assign n9711 = ( n35 & ~n9709 ) | ( n35 & n9710 ) | ( ~n9709 & n9710 ) ;
  assign n9712 = n1576 & ~n8967 ;
  assign n9713 = ( n1576 & n9711 ) | ( n1576 & ~n9712 ) | ( n9711 & ~n9712 ) ;
  assign n9714 = ( ~x2 & n9708 ) | ( ~x2 & n9713 ) | ( n9708 & n9713 ) ;
  assign n9715 = ( n9708 & n9713 ) | ( n9708 & ~n9714 ) | ( n9713 & ~n9714 ) ;
  assign n9716 = ( x2 & n9714 ) | ( x2 & ~n9715 ) | ( n9714 & ~n9715 ) ;
  assign n9717 = ( n9705 & n9707 ) | ( n9705 & n9716 ) | ( n9707 & n9716 ) ;
  assign n9718 = n36 & ~n3779 ;
  assign n9719 = n1458 & n8967 ;
  assign n9720 = ( x0 & n1338 ) | ( x0 & n8966 ) | ( n1338 & n8966 ) ;
  assign n9721 = ( n8966 & n9719 ) | ( n8966 & ~n9720 ) | ( n9719 & ~n9720 ) ;
  assign n9722 = ~n35 & n1267 ;
  assign n9723 = ( n1267 & n9721 ) | ( n1267 & ~n9722 ) | ( n9721 & ~n9722 ) ;
  assign n9724 = ( ~x2 & n9718 ) | ( ~x2 & n9723 ) | ( n9718 & n9723 ) ;
  assign n9725 = ( n9718 & n9723 ) | ( n9718 & ~n9724 ) | ( n9723 & ~n9724 ) ;
  assign n9726 = ( x2 & n9724 ) | ( x2 & ~n9725 ) | ( n9724 & ~n9725 ) ;
  assign n9727 = ( ~n9304 & n9313 ) | ( ~n9304 & n9315 ) | ( n9313 & n9315 ) ;
  assign n9728 = ( n9304 & ~n9316 ) | ( n9304 & n9727 ) | ( ~n9316 & n9727 ) ;
  assign n9729 = ( n9717 & n9726 ) | ( n9717 & n9728 ) | ( n9726 & n9728 ) ;
  assign n9730 = ( n9316 & ~n9325 ) | ( n9316 & n9327 ) | ( ~n9325 & n9327 ) ;
  assign n9731 = ( ~n9316 & n9328 ) | ( ~n9316 & n9730 ) | ( n9328 & n9730 ) ;
  assign n9732 = n36 & ~n3791 ;
  assign n9733 = n35 & ~n1246 ;
  assign n9734 = ~n1338 & n8967 ;
  assign n9735 = n9733 | n9734 ;
  assign n9736 = ~n1267 & n9378 ;
  assign n9737 = ( n9378 & n9735 ) | ( n9378 & ~n9736 ) | ( n9735 & ~n9736 ) ;
  assign n9738 = ( ~x2 & n9732 ) | ( ~x2 & n9737 ) | ( n9732 & n9737 ) ;
  assign n9739 = ( n9732 & n9737 ) | ( n9732 & ~n9738 ) | ( n9737 & ~n9738 ) ;
  assign n9740 = ( x2 & n9738 ) | ( x2 & ~n9739 ) | ( n9738 & ~n9739 ) ;
  assign n9741 = ( n9729 & ~n9731 ) | ( n9729 & n9740 ) | ( ~n9731 & n9740 ) ;
  assign n9742 = ( n9328 & ~n9337 ) | ( n9328 & n9339 ) | ( ~n9337 & n9339 ) ;
  assign n9743 = ( ~n9328 & n9340 ) | ( ~n9328 & n9742 ) | ( n9340 & n9742 ) ;
  assign n9744 = n36 & n3621 ;
  assign n9745 = ~n1246 & n9378 ;
  assign n9746 = n1267 & n8967 ;
  assign n9747 = n9745 | n9746 ;
  assign n9748 = n35 | n1290 ;
  assign n9749 = ( ~n1290 & n9747 ) | ( ~n1290 & n9748 ) | ( n9747 & n9748 ) ;
  assign n9750 = ( ~x2 & n9744 ) | ( ~x2 & n9749 ) | ( n9744 & n9749 ) ;
  assign n9751 = ( n9744 & n9749 ) | ( n9744 & ~n9750 ) | ( n9749 & ~n9750 ) ;
  assign n9752 = ( x2 & n9750 ) | ( x2 & ~n9751 ) | ( n9750 & ~n9751 ) ;
  assign n9753 = ( n9741 & ~n9743 ) | ( n9741 & n9752 ) | ( ~n9743 & n9752 ) ;
  assign n9754 = ( ~n9340 & n9349 ) | ( ~n9340 & n9351 ) | ( n9349 & n9351 ) ;
  assign n9755 = ( n9340 & ~n9352 ) | ( n9340 & n9754 ) | ( ~n9352 & n9754 ) ;
  assign n9756 = n36 & ~n3665 ;
  assign n9757 = n1246 & n8967 ;
  assign n9758 = n35 & ~n3658 ;
  assign n9759 = ( n8967 & ~n9757 ) | ( n8967 & n9758 ) | ( ~n9757 & n9758 ) ;
  assign n9760 = n1290 & n9378 ;
  assign n9761 = ( n9378 & n9759 ) | ( n9378 & ~n9760 ) | ( n9759 & ~n9760 ) ;
  assign n9762 = ( ~x2 & n9756 ) | ( ~x2 & n9761 ) | ( n9756 & n9761 ) ;
  assign n9763 = ( n9756 & n9761 ) | ( n9756 & ~n9762 ) | ( n9761 & ~n9762 ) ;
  assign n9764 = ( x2 & n9762 ) | ( x2 & ~n9763 ) | ( n9762 & ~n9763 ) ;
  assign n9765 = ( n9753 & n9755 ) | ( n9753 & n9764 ) | ( n9755 & n9764 ) ;
  assign n9766 = ( n9352 & ~n9361 ) | ( n9352 & n9363 ) | ( ~n9361 & n9363 ) ;
  assign n9767 = ( ~n9352 & n9364 ) | ( ~n9352 & n9766 ) | ( n9364 & n9766 ) ;
  assign n9768 = n36 & ~n4182 ;
  assign n9769 = n35 & ~n3692 ;
  assign n9770 = ( ~x0 & n3658 ) | ( ~x0 & n8966 ) | ( n3658 & n8966 ) ;
  assign n9771 = ( ~n3658 & n9769 ) | ( ~n3658 & n9770 ) | ( n9769 & n9770 ) ;
  assign n9772 = n1290 | n8967 ;
  assign n9773 = ( ~n1290 & n9771 ) | ( ~n1290 & n9772 ) | ( n9771 & n9772 ) ;
  assign n9774 = ( ~x2 & n9768 ) | ( ~x2 & n9773 ) | ( n9768 & n9773 ) ;
  assign n9775 = ( n9768 & n9773 ) | ( n9768 & ~n9774 ) | ( n9773 & ~n9774 ) ;
  assign n9776 = ( x2 & n9774 ) | ( x2 & ~n9775 ) | ( n9774 & ~n9775 ) ;
  assign n9777 = ( n9765 & ~n9767 ) | ( n9765 & n9776 ) | ( ~n9767 & n9776 ) ;
  assign n9778 = ( ~n9364 & n9373 ) | ( ~n9364 & n9375 ) | ( n9373 & n9375 ) ;
  assign n9779 = ( n9364 & ~n9376 ) | ( n9364 & n9778 ) | ( ~n9376 & n9778 ) ;
  assign n9780 = n36 & n3797 ;
  assign n9781 = ~n3692 & n9378 ;
  assign n9782 = ~n3658 & n8967 ;
  assign n9783 = n9781 | n9782 ;
  assign n9784 = ( ~x2 & n9780 ) | ( ~x2 & n9783 ) | ( n9780 & n9783 ) ;
  assign n9785 = ( n9780 & n9783 ) | ( n9780 & ~n9784 ) | ( n9783 & ~n9784 ) ;
  assign n9786 = ( x2 & n9784 ) | ( x2 & ~n9785 ) | ( n9784 & ~n9785 ) ;
  assign n9787 = ( n9777 & n9779 ) | ( n9777 & n9786 ) | ( n9779 & n9786 ) ;
  assign n9788 = ( n8972 & ~n8981 ) | ( n8972 & n8983 ) | ( ~n8981 & n8983 ) ;
  assign n9789 = ( n8981 & ~n8984 ) | ( n8981 & n9788 ) | ( ~n8984 & n9788 ) ;
  assign n9790 = ( n9376 & n9787 ) | ( n9376 & n9789 ) | ( n9787 & n9789 ) ;
  assign n9791 = ( n8952 & ~n8954 ) | ( n8952 & n8964 ) | ( ~n8954 & n8964 ) ;
  assign n9792 = ( n8954 & ~n8965 ) | ( n8954 & n9791 ) | ( ~n8965 & n9791 ) ;
  assign n9793 = ( n8984 & n9790 ) | ( n8984 & n9792 ) | ( n9790 & n9792 ) ;
  assign n9794 = ( n8578 & ~n8585 ) | ( n8578 & n8587 ) | ( ~n8585 & n8587 ) ;
  assign n9795 = ( n8585 & ~n8588 ) | ( n8585 & n9794 ) | ( ~n8588 & n9794 ) ;
  assign n9796 = ( n8965 & n9793 ) | ( n8965 & n9795 ) | ( n9793 & n9795 ) ;
  assign n9797 = ( n8216 & n8235 ) | ( n8216 & n8237 ) | ( n8235 & n8237 ) ;
  assign n9798 = ( n8237 & n8238 ) | ( n8237 & ~n9797 ) | ( n8238 & ~n9797 ) ;
  assign n9799 = ( n8588 & n9796 ) | ( n8588 & ~n9798 ) | ( n9796 & ~n9798 ) ;
  assign n9800 = ( n7886 & ~n7895 ) | ( n7886 & n7897 ) | ( ~n7895 & n7897 ) ;
  assign n9801 = ( n7895 & ~n7898 ) | ( n7895 & n9800 ) | ( ~n7898 & n9800 ) ;
  assign n9802 = ( n8238 & n9799 ) | ( n8238 & n9801 ) | ( n9799 & n9801 ) ;
  assign n9803 = ( n7580 & n7587 ) | ( n7580 & n7589 ) | ( n7587 & n7589 ) ;
  assign n9804 = ( n7589 & n7590 ) | ( n7589 & ~n9803 ) | ( n7590 & ~n9803 ) ;
  assign n9805 = ( n7898 & n9802 ) | ( n7898 & ~n9804 ) | ( n9802 & ~n9804 ) ;
  assign n9806 = ( ~n7289 & n7306 ) | ( ~n7289 & n7308 ) | ( n7306 & n7308 ) ;
  assign n9807 = ( n7289 & ~n7309 ) | ( n7289 & n9806 ) | ( ~n7309 & n9806 ) ;
  assign n9808 = ( n7590 & n9805 ) | ( n7590 & n9807 ) | ( n9805 & n9807 ) ;
  assign n9809 = ( n7029 & ~n7038 ) | ( n7029 & n7040 ) | ( ~n7038 & n7040 ) ;
  assign n9810 = ( n7038 & ~n7041 ) | ( n7038 & n9809 ) | ( ~n7041 & n9809 ) ;
  assign n9811 = ( n7309 & n9808 ) | ( n7309 & n9810 ) | ( n9808 & n9810 ) ;
  assign n9812 = ( n6797 & ~n6804 ) | ( n6797 & n6806 ) | ( ~n6804 & n6806 ) ;
  assign n9813 = ( n6804 & ~n6807 ) | ( n6804 & n9812 ) | ( ~n6807 & n9812 ) ;
  assign n9814 = ( n7041 & n9811 ) | ( n7041 & n9813 ) | ( n9811 & n9813 ) ;
  assign n9815 = ( n6577 & ~n6594 ) | ( n6577 & n6596 ) | ( ~n6594 & n6596 ) ;
  assign n9816 = ( n6594 & ~n6597 ) | ( n6594 & n9815 ) | ( ~n6597 & n9815 ) ;
  assign n9817 = ( n6807 & n9814 ) | ( n6807 & n9816 ) | ( n9814 & n9816 ) ;
  assign n9818 = ( n6471 & ~n6480 ) | ( n6471 & n6482 ) | ( ~n6480 & n6482 ) ;
  assign n9819 = ( n6480 & ~n6483 ) | ( n6480 & n9818 ) | ( ~n6483 & n9818 ) ;
  assign n9820 = ( n6597 & n9817 ) | ( n6597 & n9819 ) | ( n9817 & n9819 ) ;
  assign n9821 = ( n6366 & ~n6373 ) | ( n6366 & n6375 ) | ( ~n6373 & n6375 ) ;
  assign n9822 = ( n6373 & ~n6376 ) | ( n6373 & n9821 ) | ( ~n6376 & n9821 ) ;
  assign n9823 = ( n6483 & n9820 ) | ( n6483 & n9822 ) | ( n9820 & n9822 ) ;
  assign n9824 = ( ~n5959 & n5976 ) | ( ~n5959 & n5978 ) | ( n5976 & n5978 ) ;
  assign n9825 = ( n5959 & ~n5979 ) | ( n5959 & n9824 ) | ( ~n5979 & n9824 ) ;
  assign n9826 = ( n6376 & n9823 ) | ( n6376 & n9825 ) | ( n9823 & n9825 ) ;
  assign n9827 = ( n5866 & n5875 ) | ( n5866 & n5877 ) | ( n5875 & n5877 ) ;
  assign n9828 = ( n5877 & n5878 ) | ( n5877 & ~n9827 ) | ( n5878 & ~n9827 ) ;
  assign n9829 = ( n5979 & n9826 ) | ( n5979 & ~n9828 ) | ( n9826 & ~n9828 ) ;
  assign n9830 = ( n5661 & ~n5663 ) | ( n5661 & n5672 ) | ( ~n5663 & n5672 ) ;
  assign n9831 = ( n5663 & ~n5673 ) | ( n5663 & n9830 ) | ( ~n5673 & n9830 ) ;
  assign n9832 = ( n5878 & n9829 ) | ( n5878 & n9831 ) | ( n9829 & n9831 ) ;
  assign n9833 = ( n5497 & n5513 ) | ( n5497 & n5515 ) | ( n5513 & n5515 ) ;
  assign n9834 = ( n5515 & n5516 ) | ( n5515 & ~n9833 ) | ( n5516 & ~n9833 ) ;
  assign n9835 = ( n5673 & n9832 ) | ( n5673 & ~n9834 ) | ( n9832 & ~n9834 ) ;
  assign n9836 = ( n5405 & ~n5414 ) | ( n5405 & n5416 ) | ( ~n5414 & n5416 ) ;
  assign n9837 = ( n5414 & ~n5417 ) | ( n5414 & n9836 ) | ( ~n5417 & n9836 ) ;
  assign n9838 = ( n5516 & n9835 ) | ( n5516 & n9837 ) | ( n9835 & n9837 ) ;
  assign n9839 = ( ~n5336 & n5338 ) | ( ~n5336 & n5345 ) | ( n5338 & n5345 ) ;
  assign n9840 = ( n5336 & ~n5346 ) | ( n5336 & n9839 ) | ( ~n5346 & n9839 ) ;
  assign n9841 = ( n5417 & n9838 ) | ( n5417 & n9840 ) | ( n9838 & n9840 ) ;
  assign n9842 = ( n4963 & n4979 ) | ( n4963 & n4981 ) | ( n4979 & n4981 ) ;
  assign n9843 = ( n4981 & n4982 ) | ( n4981 & ~n9842 ) | ( n4982 & ~n9842 ) ;
  assign n9844 = ( n5346 & n9841 ) | ( n5346 & ~n9843 ) | ( n9841 & ~n9843 ) ;
  assign n9845 = ( n4801 & ~n4810 ) | ( n4801 & n4824 ) | ( ~n4810 & n4824 ) ;
  assign n9846 = ( n4810 & ~n4825 ) | ( n4810 & n9845 ) | ( ~n4825 & n9845 ) ;
  assign n9847 = ( n4982 & n9844 ) | ( n4982 & n9846 ) | ( n9844 & n9846 ) ;
  assign n9848 = ~n3692 & n4792 ;
  assign n9849 = ~n3658 & n4709 ;
  assign n9850 = n9848 | n9849 ;
  assign n9851 = n3797 & n4713 ;
  assign n9852 = n9850 | n9851 ;
  assign n9853 = ( ~n4690 & n4692 ) | ( ~n4690 & n4701 ) | ( n4692 & n4701 ) ;
  assign n9854 = ( ~n4701 & n4702 ) | ( ~n4701 & n9853 ) | ( n4702 & n9853 ) ;
  assign n9855 = n4822 & ~n9854 ;
  assign n9856 = n4822 & n9854 ;
  assign n9857 = ( n9854 & n9855 ) | ( n9854 & ~n9856 ) | ( n9855 & ~n9856 ) ;
  assign n9858 = ( x23 & n9852 ) | ( x23 & ~n9857 ) | ( n9852 & ~n9857 ) ;
  assign n9859 = ( ~x23 & n9852 ) | ( ~x23 & n9857 ) | ( n9852 & n9857 ) ;
  assign n9860 = ( ~n9852 & n9858 ) | ( ~n9852 & n9859 ) | ( n9858 & n9859 ) ;
  assign n9861 = ( n4825 & n9847 ) | ( n4825 & ~n9860 ) | ( n9847 & ~n9860 ) ;
  assign n9862 = ( n4702 & ~n4718 ) | ( n4702 & n4720 ) | ( ~n4718 & n4720 ) ;
  assign n9863 = ( n4718 & ~n4721 ) | ( n4718 & n9862 ) | ( ~n4721 & n9862 ) ;
  assign n9864 = ( n4822 & ~n9854 ) | ( n4822 & n9860 ) | ( ~n9854 & n9860 ) ;
  assign n9865 = ( n9861 & n9863 ) | ( n9861 & n9864 ) | ( n9863 & n9864 ) ;
  assign n9866 = ( n4373 & ~n4382 ) | ( n4373 & n4384 ) | ( ~n4382 & n4384 ) ;
  assign n9867 = ( n4382 & ~n4385 ) | ( n4382 & n9866 ) | ( ~n4385 & n9866 ) ;
  assign n9868 = ( n4721 & n9865 ) | ( n4721 & n9867 ) | ( n9865 & n9867 ) ;
  assign n9869 = ( n4341 & ~n4343 ) | ( n4341 & n4351 ) | ( ~n4343 & n4351 ) ;
  assign n9870 = ( n4343 & ~n4352 ) | ( n4343 & n9869 ) | ( ~n4352 & n9869 ) ;
  assign n9871 = ( n4385 & n9868 ) | ( n4385 & n9870 ) | ( n9868 & n9870 ) ;
  assign n9872 = ( n4207 & ~n4216 ) | ( n4207 & n4218 ) | ( ~n4216 & n4218 ) ;
  assign n9873 = ( n4216 & ~n4219 ) | ( n4216 & n9872 ) | ( ~n4219 & n9872 ) ;
  assign n9874 = ( n4352 & n9871 ) | ( n4352 & n9873 ) | ( n9871 & n9873 ) ;
  assign n9875 = ( n4177 & ~n4179 ) | ( n4177 & n4191 ) | ( ~n4179 & n4191 ) ;
  assign n9876 = ( ~n4177 & n4192 ) | ( ~n4177 & n9875 ) | ( n4192 & n9875 ) ;
  assign n9877 = ( n4219 & n9874 ) | ( n4219 & n9876 ) | ( n9874 & n9876 ) ;
  assign n9878 = ( n3794 & ~n3795 ) | ( n3794 & n3808 ) | ( ~n3795 & n3808 ) ;
  assign n9879 = ( n3795 & ~n3809 ) | ( n3795 & n9878 ) | ( ~n3809 & n9878 ) ;
  assign n9880 = ( ~n4192 & n9877 ) | ( ~n4192 & n9879 ) | ( n9877 & n9879 ) ;
  assign n9881 = ( ~n3707 & n3809 ) | ( ~n3707 & n9880 ) | ( n3809 & n9880 ) ;
  assign n9882 = ( n3707 & n3809 ) | ( n3707 & n9880 ) | ( n3809 & n9880 ) ;
  assign n9883 = ( n3707 & n9881 ) | ( n3707 & ~n9882 ) | ( n9881 & ~n9882 ) ;
  assign n9884 = n607 & ~n9883 ;
  assign n9885 = n366 | n1168 ;
  assign n9886 = ( ~n1218 & n5049 ) | ( ~n1218 & n6025 ) | ( n5049 & n6025 ) ;
  assign n9887 = n1218 | n9886 ;
  assign n9888 = n2353 | n2412 ;
  assign n9889 = n450 | n796 ;
  assign n9890 = n540 | n956 ;
  assign n9891 = n2683 | n9890 ;
  assign n9892 = ( ~n9888 & n9889 ) | ( ~n9888 & n9891 ) | ( n9889 & n9891 ) ;
  assign n9893 = n9888 | n9892 ;
  assign n9894 = ( n312 & ~n382 ) | ( n312 & n463 ) | ( ~n382 & n463 ) ;
  assign n9895 = n382 | n1835 ;
  assign n9896 = ( n378 & ~n9894 ) | ( n378 & n9895 ) | ( ~n9894 & n9895 ) ;
  assign n9897 = n9894 | n9896 ;
  assign n9898 = ( n95 & ~n9893 ) | ( n95 & n9897 ) | ( ~n9893 & n9897 ) ;
  assign n9899 = n9893 | n9898 ;
  assign n9900 = ( ~n9885 & n9887 ) | ( ~n9885 & n9899 ) | ( n9887 & n9899 ) ;
  assign n9901 = n9885 | n9900 ;
  assign n9902 = ( x29 & n744 ) | ( x29 & ~n9901 ) | ( n744 & ~n9901 ) ;
  assign n9903 = ( x29 & ~n744 ) | ( x29 & n9901 ) | ( ~n744 & n9901 ) ;
  assign n9904 = ( ~x29 & n9902 ) | ( ~x29 & n9903 ) | ( n9902 & n9903 ) ;
  assign n9905 = n1250 & ~n3658 ;
  assign n9906 = n607 & n1290 ;
  assign n9907 = ( n607 & n9905 ) | ( n607 & ~n9906 ) | ( n9905 & ~n9906 ) ;
  assign n9908 = n1248 & ~n4182 ;
  assign n9909 = n9907 | n9908 ;
  assign n9910 = ( n3625 & n9904 ) | ( n3625 & n9909 ) | ( n9904 & n9909 ) ;
  assign n9911 = ( n3625 & ~n9904 ) | ( n3625 & n9909 ) | ( ~n9904 & n9909 ) ;
  assign n9912 = ( n9904 & ~n9910 ) | ( n9904 & n9911 ) | ( ~n9910 & n9911 ) ;
  assign n9913 = ( ~n3628 & n3667 ) | ( ~n3628 & n3707 ) | ( n3667 & n3707 ) ;
  assign n9914 = ( n9881 & n9912 ) | ( n9881 & n9913 ) | ( n9912 & n9913 ) ;
  assign n9915 = ( ~n9881 & n9912 ) | ( ~n9881 & n9913 ) | ( n9912 & n9913 ) ;
  assign n9916 = ( n9881 & ~n9914 ) | ( n9881 & n9915 ) | ( ~n9914 & n9915 ) ;
  assign n9917 = n1250 & n9916 ;
  assign n9918 = n9884 | n9917 ;
  assign n9919 = ( n1001 & ~n1235 ) | ( n1001 & n3081 ) | ( ~n1235 & n3081 ) ;
  assign n9920 = n1235 | n9919 ;
  assign n9921 = ( n1213 & n1226 ) | ( n1213 & ~n9920 ) | ( n1226 & ~n9920 ) ;
  assign n9922 = n9920 | n9921 ;
  assign n9923 = ( ~n3651 & n3685 ) | ( ~n3651 & n9922 ) | ( n3685 & n9922 ) ;
  assign n9924 = ( n3651 & ~n5138 ) | ( n3651 & n9923 ) | ( ~n5138 & n9923 ) ;
  assign n9925 = n5138 | n9924 ;
  assign n9926 = ~n95 & n375 ;
  assign n9927 = ( ~n1434 & n9925 ) | ( ~n1434 & n9926 ) | ( n9925 & n9926 ) ;
  assign n9928 = ~n9925 & n9927 ;
  assign n9929 = n1250 & ~n3692 ;
  assign n9930 = n1248 & n3797 ;
  assign n9931 = n9929 | n9930 ;
  assign n9932 = ( ~n9902 & n9928 ) | ( ~n9902 & n9931 ) | ( n9928 & n9931 ) ;
  assign n9933 = ( n9928 & n9931 ) | ( n9928 & ~n9932 ) | ( n9931 & ~n9932 ) ;
  assign n9934 = ( n9902 & n9932 ) | ( n9902 & ~n9933 ) | ( n9932 & ~n9933 ) ;
  assign n9935 = ( n9910 & n9914 ) | ( n9910 & ~n9934 ) | ( n9914 & ~n9934 ) ;
  assign n9936 = ( n9910 & ~n9914 ) | ( n9910 & n9934 ) | ( ~n9914 & n9934 ) ;
  assign n9937 = ( ~n9910 & n9935 ) | ( ~n9910 & n9936 ) | ( n9935 & n9936 ) ;
  assign n9938 = n606 & n9937 ;
  assign n9939 = ( n606 & n9918 ) | ( n606 & ~n9938 ) | ( n9918 & ~n9938 ) ;
  assign n9940 = ( n9877 & n9879 ) | ( n9877 & ~n9880 ) | ( n9879 & ~n9880 ) ;
  assign n9941 = ( n4192 & n9880 ) | ( n4192 & ~n9940 ) | ( n9880 & ~n9940 ) ;
  assign n9942 = ( n4219 & ~n9874 ) | ( n4219 & n9876 ) | ( ~n9874 & n9876 ) ;
  assign n9943 = ( n9874 & ~n9877 ) | ( n9874 & n9942 ) | ( ~n9877 & n9942 ) ;
  assign n9944 = ( n4352 & ~n9871 ) | ( n4352 & n9873 ) | ( ~n9871 & n9873 ) ;
  assign n9945 = ( n9871 & ~n9874 ) | ( n9871 & n9944 ) | ( ~n9874 & n9944 ) ;
  assign n9946 = ( n4385 & ~n9868 ) | ( n4385 & n9870 ) | ( ~n9868 & n9870 ) ;
  assign n9947 = ( n9868 & ~n9871 ) | ( n9868 & n9946 ) | ( ~n9871 & n9946 ) ;
  assign n9948 = ( n4721 & ~n9865 ) | ( n4721 & n9867 ) | ( ~n9865 & n9867 ) ;
  assign n9949 = ( n9865 & ~n9868 ) | ( n9865 & n9948 ) | ( ~n9868 & n9948 ) ;
  assign n9950 = ( ~n9861 & n9863 ) | ( ~n9861 & n9864 ) | ( n9863 & n9864 ) ;
  assign n9951 = ( n9861 & ~n9865 ) | ( n9861 & n9950 ) | ( ~n9865 & n9950 ) ;
  assign n9952 = ( n4825 & ~n9847 ) | ( n4825 & n9860 ) | ( ~n9847 & n9860 ) ;
  assign n9953 = ( ~n4825 & n9861 ) | ( ~n4825 & n9952 ) | ( n9861 & n9952 ) ;
  assign n9954 = ( n4982 & ~n9844 ) | ( n4982 & n9846 ) | ( ~n9844 & n9846 ) ;
  assign n9955 = ( n9844 & ~n9847 ) | ( n9844 & n9954 ) | ( ~n9847 & n9954 ) ;
  assign n9956 = ( n5346 & ~n9841 ) | ( n5346 & n9843 ) | ( ~n9841 & n9843 ) ;
  assign n9957 = ( ~n5346 & n9844 ) | ( ~n5346 & n9956 ) | ( n9844 & n9956 ) ;
  assign n9958 = ( n5417 & ~n9838 ) | ( n5417 & n9840 ) | ( ~n9838 & n9840 ) ;
  assign n9959 = ( n9838 & ~n9841 ) | ( n9838 & n9958 ) | ( ~n9841 & n9958 ) ;
  assign n9960 = ( n5516 & ~n9835 ) | ( n5516 & n9837 ) | ( ~n9835 & n9837 ) ;
  assign n9961 = ( n9835 & ~n9838 ) | ( n9835 & n9960 ) | ( ~n9838 & n9960 ) ;
  assign n9962 = ( n5673 & ~n9832 ) | ( n5673 & n9834 ) | ( ~n9832 & n9834 ) ;
  assign n9963 = ( ~n5673 & n9835 ) | ( ~n5673 & n9962 ) | ( n9835 & n9962 ) ;
  assign n9964 = ( n5878 & ~n9829 ) | ( n5878 & n9831 ) | ( ~n9829 & n9831 ) ;
  assign n9965 = ( n9829 & ~n9832 ) | ( n9829 & n9964 ) | ( ~n9832 & n9964 ) ;
  assign n9966 = ( n5979 & ~n9826 ) | ( n5979 & n9828 ) | ( ~n9826 & n9828 ) ;
  assign n9967 = ( ~n5979 & n9829 ) | ( ~n5979 & n9966 ) | ( n9829 & n9966 ) ;
  assign n9968 = ( n6376 & ~n9823 ) | ( n6376 & n9825 ) | ( ~n9823 & n9825 ) ;
  assign n9969 = ( n9823 & ~n9826 ) | ( n9823 & n9968 ) | ( ~n9826 & n9968 ) ;
  assign n9970 = ( n6483 & ~n9820 ) | ( n6483 & n9822 ) | ( ~n9820 & n9822 ) ;
  assign n9971 = ( n9820 & ~n9823 ) | ( n9820 & n9970 ) | ( ~n9823 & n9970 ) ;
  assign n9972 = ( n6597 & ~n9817 ) | ( n6597 & n9819 ) | ( ~n9817 & n9819 ) ;
  assign n9973 = ( n9817 & ~n9820 ) | ( n9817 & n9972 ) | ( ~n9820 & n9972 ) ;
  assign n9974 = ( n6807 & ~n9814 ) | ( n6807 & n9816 ) | ( ~n9814 & n9816 ) ;
  assign n9975 = ( n9814 & ~n9817 ) | ( n9814 & n9974 ) | ( ~n9817 & n9974 ) ;
  assign n9976 = ( n7041 & ~n9811 ) | ( n7041 & n9813 ) | ( ~n9811 & n9813 ) ;
  assign n9977 = ( n9811 & ~n9814 ) | ( n9811 & n9976 ) | ( ~n9814 & n9976 ) ;
  assign n9978 = ( n7309 & ~n9808 ) | ( n7309 & n9810 ) | ( ~n9808 & n9810 ) ;
  assign n9979 = ( n9808 & ~n9811 ) | ( n9808 & n9978 ) | ( ~n9811 & n9978 ) ;
  assign n9980 = ( n7590 & ~n9805 ) | ( n7590 & n9807 ) | ( ~n9805 & n9807 ) ;
  assign n9981 = ( n9805 & ~n9808 ) | ( n9805 & n9980 ) | ( ~n9808 & n9980 ) ;
  assign n9982 = ( n7898 & ~n9802 ) | ( n7898 & n9804 ) | ( ~n9802 & n9804 ) ;
  assign n9983 = ( ~n7898 & n9805 ) | ( ~n7898 & n9982 ) | ( n9805 & n9982 ) ;
  assign n9984 = ( n8238 & ~n9799 ) | ( n8238 & n9801 ) | ( ~n9799 & n9801 ) ;
  assign n9985 = ( n9799 & ~n9802 ) | ( n9799 & n9984 ) | ( ~n9802 & n9984 ) ;
  assign n9986 = ( n8588 & ~n9796 ) | ( n8588 & n9798 ) | ( ~n9796 & n9798 ) ;
  assign n9987 = ( ~n8588 & n9799 ) | ( ~n8588 & n9986 ) | ( n9799 & n9986 ) ;
  assign n9988 = ( n8965 & ~n9793 ) | ( n8965 & n9795 ) | ( ~n9793 & n9795 ) ;
  assign n9989 = ( n9793 & ~n9796 ) | ( n9793 & n9988 ) | ( ~n9796 & n9988 ) ;
  assign n9990 = ( n8984 & ~n9790 ) | ( n8984 & n9792 ) | ( ~n9790 & n9792 ) ;
  assign n9991 = ( n9790 & ~n9793 ) | ( n9790 & n9990 ) | ( ~n9793 & n9990 ) ;
  assign n9992 = ( n9376 & ~n9787 ) | ( n9376 & n9789 ) | ( ~n9787 & n9789 ) ;
  assign n9993 = ( n9787 & ~n9790 ) | ( n9787 & n9992 ) | ( ~n9790 & n9992 ) ;
  assign n9994 = ( ~n9777 & n9779 ) | ( ~n9777 & n9786 ) | ( n9779 & n9786 ) ;
  assign n9995 = ( n9777 & ~n9787 ) | ( n9777 & n9994 ) | ( ~n9787 & n9994 ) ;
  assign n9996 = ( ~n9765 & n9767 ) | ( ~n9765 & n9776 ) | ( n9767 & n9776 ) ;
  assign n9997 = ( ~n9776 & n9777 ) | ( ~n9776 & n9996 ) | ( n9777 & n9996 ) ;
  assign n9998 = ( ~n9753 & n9755 ) | ( ~n9753 & n9764 ) | ( n9755 & n9764 ) ;
  assign n9999 = ( n9753 & ~n9765 ) | ( n9753 & n9998 ) | ( ~n9765 & n9998 ) ;
  assign n10000 = ( ~n9741 & n9743 ) | ( ~n9741 & n9752 ) | ( n9743 & n9752 ) ;
  assign n10001 = ( ~n9752 & n9753 ) | ( ~n9752 & n10000 ) | ( n9753 & n10000 ) ;
  assign n10002 = ( ~n9729 & n9731 ) | ( ~n9729 & n9740 ) | ( n9731 & n9740 ) ;
  assign n10003 = ( ~n9740 & n9741 ) | ( ~n9740 & n10002 ) | ( n9741 & n10002 ) ;
  assign n10004 = ( n9999 & ~n10001 ) | ( n9999 & n10003 ) | ( ~n10001 & n10003 ) ;
  assign n10005 = ~n9999 & n10004 ;
  assign n10006 = n10001 | n10005 ;
  assign n10007 = ( n9997 & ~n9999 ) | ( n9997 & n10006 ) | ( ~n9999 & n10006 ) ;
  assign n10008 = ( ~n9995 & n9997 ) | ( ~n9995 & n10007 ) | ( n9997 & n10007 ) ;
  assign n10009 = ( n9993 & n9995 ) | ( n9993 & ~n10008 ) | ( n9995 & ~n10008 ) ;
  assign n10010 = ( n9991 & n9993 ) | ( n9991 & n10009 ) | ( n9993 & n10009 ) ;
  assign n10011 = ( n9989 & n9991 ) | ( n9989 & n10010 ) | ( n9991 & n10010 ) ;
  assign n10012 = ( ~n9987 & n9989 ) | ( ~n9987 & n10011 ) | ( n9989 & n10011 ) ;
  assign n10013 = ( n9985 & ~n9987 ) | ( n9985 & n10012 ) | ( ~n9987 & n10012 ) ;
  assign n10014 = ( ~n9983 & n9985 ) | ( ~n9983 & n10013 ) | ( n9985 & n10013 ) ;
  assign n10015 = ( n9981 & ~n9983 ) | ( n9981 & n10014 ) | ( ~n9983 & n10014 ) ;
  assign n10016 = ( n9979 & n9981 ) | ( n9979 & n10015 ) | ( n9981 & n10015 ) ;
  assign n10017 = ( n9977 & n9979 ) | ( n9977 & n10016 ) | ( n9979 & n10016 ) ;
  assign n10018 = ( n9975 & n9977 ) | ( n9975 & n10017 ) | ( n9977 & n10017 ) ;
  assign n10019 = ( n9973 & n9975 ) | ( n9973 & n10018 ) | ( n9975 & n10018 ) ;
  assign n10020 = ( n9971 & n9973 ) | ( n9971 & n10019 ) | ( n9973 & n10019 ) ;
  assign n10021 = ( n9969 & n9971 ) | ( n9969 & n10020 ) | ( n9971 & n10020 ) ;
  assign n10022 = ( ~n9967 & n9969 ) | ( ~n9967 & n10021 ) | ( n9969 & n10021 ) ;
  assign n10023 = ( n9965 & ~n9967 ) | ( n9965 & n10022 ) | ( ~n9967 & n10022 ) ;
  assign n10024 = ( ~n9963 & n9965 ) | ( ~n9963 & n10023 ) | ( n9965 & n10023 ) ;
  assign n10025 = ( n9961 & ~n9963 ) | ( n9961 & n10024 ) | ( ~n9963 & n10024 ) ;
  assign n10026 = ( n9959 & n9961 ) | ( n9959 & n10025 ) | ( n9961 & n10025 ) ;
  assign n10027 = ( ~n9957 & n9959 ) | ( ~n9957 & n10026 ) | ( n9959 & n10026 ) ;
  assign n10028 = ( n9955 & ~n9957 ) | ( n9955 & n10027 ) | ( ~n9957 & n10027 ) ;
  assign n10029 = ( ~n9953 & n9955 ) | ( ~n9953 & n10028 ) | ( n9955 & n10028 ) ;
  assign n10030 = ( n9951 & ~n9953 ) | ( n9951 & n10029 ) | ( ~n9953 & n10029 ) ;
  assign n10031 = ( n9949 & n9951 ) | ( n9949 & n10030 ) | ( n9951 & n10030 ) ;
  assign n10032 = ( n9947 & n9949 ) | ( n9947 & n10031 ) | ( n9949 & n10031 ) ;
  assign n10033 = ( n9945 & n9947 ) | ( n9945 & n10032 ) | ( n9947 & n10032 ) ;
  assign n10034 = ( n9943 & n9945 ) | ( n9943 & n10033 ) | ( n9945 & n10033 ) ;
  assign n10035 = ( ~n9941 & n9943 ) | ( ~n9941 & n10034 ) | ( n9943 & n10034 ) ;
  assign n10036 = ( n9883 & n9941 ) | ( n9883 & ~n10035 ) | ( n9941 & ~n10035 ) ;
  assign n10037 = ( n9883 & ~n9916 ) | ( n9883 & n10036 ) | ( ~n9916 & n10036 ) ;
  assign n10038 = ( ~n9916 & n9937 ) | ( ~n9916 & n10037 ) | ( n9937 & n10037 ) ;
  assign n10039 = ( n9916 & ~n9937 ) | ( n9916 & n10037 ) | ( ~n9937 & n10037 ) ;
  assign n10040 = ( ~n10037 & n10038 ) | ( ~n10037 & n10039 ) | ( n10038 & n10039 ) ;
  assign n10041 = n1248 & n10040 ;
  assign n10042 = n9939 | n10041 ;
  assign n10043 = ( n311 & n605 ) | ( n311 & n10042 ) | ( n605 & n10042 ) ;
  assign n10044 = n1254 | n1870 ;
  assign n10045 = ( n72 & n129 ) | ( n72 & n160 ) | ( n129 & n160 ) ;
  assign n10046 = n55 | n10045 ;
  assign n10047 = ( n3679 & ~n10044 ) | ( n3679 & n10046 ) | ( ~n10044 & n10046 ) ;
  assign n10048 = n10044 | n10047 ;
  assign n10049 = ( n1230 & n3655 ) | ( n1230 & n9897 ) | ( n3655 & n9897 ) ;
  assign n10050 = ( n1230 & n10048 ) | ( n1230 & ~n10049 ) | ( n10048 & ~n10049 ) ;
  assign n10051 = ~n10048 & n10050 ;
  assign n10052 = n9928 & ~n10051 ;
  assign n10053 = n9928 & n10051 ;
  assign n10054 = ( n10051 & n10052 ) | ( n10051 & ~n10053 ) | ( n10052 & ~n10053 ) ;
  assign n10055 = ( n9932 & n9935 ) | ( n9932 & ~n10054 ) | ( n9935 & ~n10054 ) ;
  assign n10056 = ( n9932 & ~n9935 ) | ( n9932 & n10054 ) | ( ~n9935 & n10054 ) ;
  assign n10057 = ( ~n9932 & n10055 ) | ( ~n9932 & n10056 ) | ( n10055 & n10056 ) ;
  assign n10058 = n606 & n10057 ;
  assign n10059 = ( n607 & n1250 ) | ( n607 & ~n9937 ) | ( n1250 & ~n9937 ) ;
  assign n10060 = ( n9917 & ~n9937 ) | ( n9917 & n10059 ) | ( ~n9937 & n10059 ) ;
  assign n10061 = ( n606 & ~n10058 ) | ( n606 & n10060 ) | ( ~n10058 & n10060 ) ;
  assign n10062 = ( n9937 & n10038 ) | ( n9937 & n10057 ) | ( n10038 & n10057 ) ;
  assign n10063 = ( ~n9937 & n10038 ) | ( ~n9937 & n10057 ) | ( n10038 & n10057 ) ;
  assign n10064 = ( n9937 & ~n10062 ) | ( n9937 & n10063 ) | ( ~n10062 & n10063 ) ;
  assign n10065 = n1248 & ~n10064 ;
  assign n10066 = n10061 | n10065 ;
  assign n10067 = ( ~n462 & n10043 ) | ( ~n462 & n10066 ) | ( n10043 & n10066 ) ;
  assign n10068 = ( n462 & n10043 ) | ( n462 & n10066 ) | ( n10043 & n10066 ) ;
  assign n10069 = ( n462 & n10067 ) | ( n462 & ~n10068 ) | ( n10067 & ~n10068 ) ;
  assign n10070 = n3162 | n3731 ;
  assign n10071 = ( n295 & n691 ) | ( n295 & ~n916 ) | ( n691 & ~n916 ) ;
  assign n10072 = n916 | n10071 ;
  assign n10073 = n2126 | n3747 ;
  assign n10074 = ( n913 & n1257 ) | ( n913 & ~n2126 ) | ( n1257 & ~n2126 ) ;
  assign n10075 = ( ~n10072 & n10073 ) | ( ~n10072 & n10074 ) | ( n10073 & n10074 ) ;
  assign n10076 = n10072 | n10075 ;
  assign n10077 = ( n3873 & ~n10070 ) | ( n3873 & n10076 ) | ( ~n10070 & n10076 ) ;
  assign n10078 = n10070 | n10077 ;
  assign n10079 = n422 | n513 ;
  assign n10080 = ( n153 & n969 ) | ( n153 & ~n10079 ) | ( n969 & ~n10079 ) ;
  assign n10081 = n10079 | n10080 ;
  assign n10082 = n51 | n316 ;
  assign n10083 = n254 | n10082 ;
  assign n10084 = ( n2975 & n9890 ) | ( n2975 & ~n10083 ) | ( n9890 & ~n10083 ) ;
  assign n10085 = n10083 | n10084 ;
  assign n10086 = n5015 | n10085 ;
  assign n10087 = n2791 | n2929 ;
  assign n10088 = n81 | n824 ;
  assign n10089 = ( n2484 & n6206 ) | ( n2484 & ~n10088 ) | ( n6206 & ~n10088 ) ;
  assign n10090 = n10088 | n10089 ;
  assign n10091 = ( n4426 & ~n10087 ) | ( n4426 & n10090 ) | ( ~n10087 & n10090 ) ;
  assign n10092 = n10087 | n10091 ;
  assign n10093 = ( ~n10081 & n10086 ) | ( ~n10081 & n10092 ) | ( n10086 & n10092 ) ;
  assign n10094 = n10081 | n10093 ;
  assign n10095 = n4486 | n10094 ;
  assign n10096 = n287 | n1351 ;
  assign n10097 = ( n57 & n102 ) | ( n57 & n145 ) | ( n102 & n145 ) ;
  assign n10098 = n990 | n10097 ;
  assign n10099 = n1487 | n2033 ;
  assign n10100 = n3390 | n10099 ;
  assign n10101 = ( ~n10096 & n10098 ) | ( ~n10096 & n10100 ) | ( n10098 & n10100 ) ;
  assign n10102 = n10096 | n10101 ;
  assign n10103 = n246 | n3902 ;
  assign n10104 = ( n5573 & ~n10102 ) | ( n5573 & n10103 ) | ( ~n10102 & n10103 ) ;
  assign n10105 = n10102 | n10104 ;
  assign n10106 = ( ~n10078 & n10095 ) | ( ~n10078 & n10105 ) | ( n10095 & n10105 ) ;
  assign n10107 = n10078 | n10106 ;
  assign n10108 = n1526 | n2207 ;
  assign n10109 = ( n57 & n66 ) | ( n57 & n73 ) | ( n66 & n73 ) ;
  assign n10110 = ( n66 & n129 ) | ( n66 & n160 ) | ( n129 & n160 ) ;
  assign n10111 = ( n1721 & n10109 ) | ( n1721 & ~n10110 ) | ( n10109 & ~n10110 ) ;
  assign n10112 = n368 | n641 ;
  assign n10113 = n512 | n10112 ;
  assign n10114 = ( n10110 & ~n10111 ) | ( n10110 & n10113 ) | ( ~n10111 & n10113 ) ;
  assign n10115 = n10111 | n10114 ;
  assign n10116 = n110 | n146 ;
  assign n10117 = ( ~n10108 & n10115 ) | ( ~n10108 & n10116 ) | ( n10115 & n10116 ) ;
  assign n10118 = n10108 | n10117 ;
  assign n10119 = n690 | n3520 ;
  assign n10120 = n440 | n838 ;
  assign n10121 = ( n4069 & n4873 ) | ( n4069 & ~n10120 ) | ( n4873 & ~n10120 ) ;
  assign n10122 = n10120 | n10121 ;
  assign n10123 = n337 | n353 ;
  assign n10124 = ( n433 & n609 ) | ( n433 & ~n10123 ) | ( n609 & ~n10123 ) ;
  assign n10125 = n10123 | n10124 ;
  assign n10126 = ( ~n10119 & n10122 ) | ( ~n10119 & n10125 ) | ( n10122 & n10125 ) ;
  assign n10127 = n10119 | n10126 ;
  assign n10128 = ( n4537 & ~n5750 ) | ( n4537 & n10127 ) | ( ~n5750 & n10127 ) ;
  assign n10129 = n239 | n492 ;
  assign n10130 = n719 | n1208 ;
  assign n10131 = ( n1059 & ~n10129 ) | ( n1059 & n10130 ) | ( ~n10129 & n10130 ) ;
  assign n10132 = n10129 | n10131 ;
  assign n10133 = ( n5750 & ~n10128 ) | ( n5750 & n10132 ) | ( ~n10128 & n10132 ) ;
  assign n10134 = n10128 | n10133 ;
  assign n10135 = ( ~n4890 & n10118 ) | ( ~n4890 & n10134 ) | ( n10118 & n10134 ) ;
  assign n10136 = ( n73 & n80 ) | ( n73 & n136 ) | ( n80 & n136 ) ;
  assign n10137 = n379 | n10136 ;
  assign n10138 = ( n59 & n145 ) | ( n59 & n166 ) | ( n145 & n166 ) ;
  assign n10139 = n132 | n10138 ;
  assign n10140 = n45 | n514 ;
  assign n10141 = n928 | n10140 ;
  assign n10142 = ( ~n10137 & n10139 ) | ( ~n10137 & n10141 ) | ( n10139 & n10141 ) ;
  assign n10143 = n10137 | n10142 ;
  assign n10144 = n2011 | n2071 ;
  assign n10145 = ( n2232 & n2467 ) | ( n2232 & ~n10144 ) | ( n2467 & ~n10144 ) ;
  assign n10146 = n10144 | n10145 ;
  assign n10147 = ( n1963 & ~n10143 ) | ( n1963 & n10146 ) | ( ~n10143 & n10146 ) ;
  assign n10148 = n10143 | n10147 ;
  assign n10149 = ( n66 & n84 ) | ( n66 & n119 ) | ( n84 & n119 ) ;
  assign n10150 = ( n549 & n732 ) | ( n549 & ~n10149 ) | ( n732 & ~n10149 ) ;
  assign n10151 = n10149 | n10150 ;
  assign n10152 = n138 | n1436 ;
  assign n10153 = ( n6175 & ~n10151 ) | ( n6175 & n10152 ) | ( ~n10151 & n10152 ) ;
  assign n10154 = n10151 | n10153 ;
  assign n10155 = n292 | n1494 ;
  assign n10156 = ( n3997 & n6092 ) | ( n3997 & ~n10155 ) | ( n6092 & ~n10155 ) ;
  assign n10157 = n10155 | n10156 ;
  assign n10158 = ( n548 & ~n10154 ) | ( n548 & n10157 ) | ( ~n10154 & n10157 ) ;
  assign n10159 = n10154 | n10158 ;
  assign n10160 = ( ~n10118 & n10148 ) | ( ~n10118 & n10159 ) | ( n10148 & n10159 ) ;
  assign n10161 = ( ~n4890 & n10135 ) | ( ~n4890 & n10160 ) | ( n10135 & n10160 ) ;
  assign n10162 = n4890 | n10161 ;
  assign n10163 = ( x23 & n4712 ) | ( x23 & n4792 ) | ( n4712 & n4792 ) ;
  assign n10164 = n4712 | n4792 ;
  assign n10165 = x22 | n10164 ;
  assign n10166 = ~n10163 & n10165 ;
  assign n10167 = ( n10107 & n10162 ) | ( n10107 & ~n10166 ) | ( n10162 & ~n10166 ) ;
  assign n10168 = n607 | n9941 ;
  assign n10169 = n1250 & ~n9883 ;
  assign n10170 = ( ~n9941 & n10168 ) | ( ~n9941 & n10169 ) | ( n10168 & n10169 ) ;
  assign n10171 = n606 & ~n9916 ;
  assign n10172 = ( n606 & n10170 ) | ( n606 & ~n10171 ) | ( n10170 & ~n10171 ) ;
  assign n10173 = ( n9883 & n9916 ) | ( n9883 & n10036 ) | ( n9916 & n10036 ) ;
  assign n10174 = ( n9916 & n10037 ) | ( n9916 & ~n10173 ) | ( n10037 & ~n10173 ) ;
  assign n10175 = n1248 & n10174 ;
  assign n10176 = n10172 | n10175 ;
  assign n10177 = ( n311 & n10167 ) | ( n311 & n10176 ) | ( n10167 & n10176 ) ;
  assign n10178 = ( n59 & n98 ) | ( n59 & n328 ) | ( n98 & n328 ) ;
  assign n10179 = ( n290 & n746 ) | ( n290 & ~n10178 ) | ( n746 & ~n10178 ) ;
  assign n10180 = n10178 | n10179 ;
  assign n10181 = n234 | n655 ;
  assign n10182 = n1693 | n3828 ;
  assign n10183 = ( n847 & ~n10181 ) | ( n847 & n10182 ) | ( ~n10181 & n10182 ) ;
  assign n10184 = n10181 | n10183 ;
  assign n10185 = ( n4488 & ~n10180 ) | ( n4488 & n10184 ) | ( ~n10180 & n10184 ) ;
  assign n10186 = n10180 | n10185 ;
  assign n10187 = ~n1171 & n1742 ;
  assign n10188 = n1048 | n1237 ;
  assign n10189 = n302 | n10188 ;
  assign n10190 = ( n807 & n10187 ) | ( n807 & n10189 ) | ( n10187 & n10189 ) ;
  assign n10191 = n10187 & ~n10190 ;
  assign n10192 = ( n3428 & ~n10186 ) | ( n3428 & n10191 ) | ( ~n10186 & n10191 ) ;
  assign n10193 = n1658 | n3378 ;
  assign n10194 = n3351 | n10193 ;
  assign n10195 = n79 | n338 ;
  assign n10196 = ( n483 & n1225 ) | ( n483 & ~n10195 ) | ( n1225 & ~n10195 ) ;
  assign n10197 = n10195 | n10196 ;
  assign n10198 = ( n4510 & ~n10193 ) | ( n4510 & n10197 ) | ( ~n10193 & n10197 ) ;
  assign n10199 = ( n781 & n2353 ) | ( n781 & ~n10198 ) | ( n2353 & ~n10198 ) ;
  assign n10200 = n10198 | n10199 ;
  assign n10201 = n300 | n1110 ;
  assign n10202 = ( ~n54 & n73 ) | ( ~n54 & n166 ) | ( n73 & n166 ) ;
  assign n10203 = n174 | n312 ;
  assign n10204 = ( n479 & n662 ) | ( n479 & ~n10203 ) | ( n662 & ~n10203 ) ;
  assign n10205 = n10203 | n10204 ;
  assign n10206 = ( ~n10201 & n10202 ) | ( ~n10201 & n10205 ) | ( n10202 & n10205 ) ;
  assign n10207 = n10201 | n10206 ;
  assign n10208 = ( ~n10194 & n10200 ) | ( ~n10194 & n10207 ) | ( n10200 & n10207 ) ;
  assign n10209 = n10194 | n10208 ;
  assign n10210 = ( n10094 & n10191 ) | ( n10094 & n10209 ) | ( n10191 & n10209 ) ;
  assign n10211 = ( n3428 & n10192 ) | ( n3428 & ~n10210 ) | ( n10192 & ~n10210 ) ;
  assign n10212 = ~n3428 & n10211 ;
  assign n10213 = n609 | n2945 ;
  assign n10214 = n1680 | n1716 ;
  assign n10215 = n686 | n1690 ;
  assign n10216 = ( ~n10213 & n10214 ) | ( ~n10213 & n10215 ) | ( n10214 & n10215 ) ;
  assign n10217 = n10213 | n10216 ;
  assign n10218 = ( n64 & n97 ) | ( n64 & n122 ) | ( n97 & n122 ) ;
  assign n10219 = n2827 | n5002 ;
  assign n10220 = n10218 | n10219 ;
  assign n10221 = ( n1332 & n3415 ) | ( n1332 & ~n10220 ) | ( n3415 & ~n10220 ) ;
  assign n10222 = n10220 | n10221 ;
  assign n10223 = ( n2392 & ~n10217 ) | ( n2392 & n10222 ) | ( ~n10217 & n10222 ) ;
  assign n10224 = n10217 | n10223 ;
  assign n10225 = ( n1113 & n1892 ) | ( n1113 & ~n2078 ) | ( n1892 & ~n2078 ) ;
  assign n10226 = n2078 | n10225 ;
  assign n10227 = n2124 | n3584 ;
  assign n10228 = n445 | n4100 ;
  assign n10229 = n234 | n394 ;
  assign n10230 = ( n1078 & n1790 ) | ( n1078 & ~n10229 ) | ( n1790 & ~n10229 ) ;
  assign n10231 = n10229 | n10230 ;
  assign n10232 = ( n465 & ~n977 ) | ( n465 & n1637 ) | ( ~n977 & n1637 ) ;
  assign n10233 = n977 | n10232 ;
  assign n10234 = ( ~n10228 & n10231 ) | ( ~n10228 & n10233 ) | ( n10231 & n10233 ) ;
  assign n10235 = n10228 | n10234 ;
  assign n10236 = ( ~n10226 & n10227 ) | ( ~n10226 & n10235 ) | ( n10227 & n10235 ) ;
  assign n10237 = n10226 | n10236 ;
  assign n10238 = ( n2677 & n10224 ) | ( n2677 & ~n10237 ) | ( n10224 & ~n10237 ) ;
  assign n10239 = ~n10224 & n10238 ;
  assign n10240 = ( n4966 & n4967 ) | ( n4966 & ~n5397 ) | ( n4967 & ~n5397 ) ;
  assign n10241 = ( n4970 & ~n4972 ) | ( n4970 & n5398 ) | ( ~n4972 & n5398 ) ;
  assign n10242 = ( ~x20 & n10240 ) | ( ~x20 & n10241 ) | ( n10240 & n10241 ) ;
  assign n10243 = ( n10212 & n10239 ) | ( n10212 & n10242 ) | ( n10239 & n10242 ) ;
  assign n10244 = n79 | n347 ;
  assign n10245 = ( n80 & n149 ) | ( n80 & n160 ) | ( n149 & n160 ) ;
  assign n10246 = ( n131 & n185 ) | ( n131 & ~n10245 ) | ( n185 & ~n10245 ) ;
  assign n10247 = n10245 | n10246 ;
  assign n10248 = ( n762 & ~n10244 ) | ( n762 & n10247 ) | ( ~n10244 & n10247 ) ;
  assign n10249 = n10244 | n10248 ;
  assign n10250 = n732 | n749 ;
  assign n10251 = n889 | n10250 ;
  assign n10252 = n103 | n352 ;
  assign n10253 = ( n206 & n625 ) | ( n206 & ~n10252 ) | ( n625 & ~n10252 ) ;
  assign n10254 = n10252 | n10253 ;
  assign n10255 = n2661 | n2726 ;
  assign n10256 = ( ~n10251 & n10254 ) | ( ~n10251 & n10255 ) | ( n10254 & n10255 ) ;
  assign n10257 = n10251 | n10256 ;
  assign n10258 = n192 | n367 ;
  assign n10259 = n810 | n10258 ;
  assign n10260 = ( ~n10249 & n10257 ) | ( ~n10249 & n10259 ) | ( n10257 & n10259 ) ;
  assign n10261 = n10249 | n10260 ;
  assign n10262 = n2520 | n3538 ;
  assign n10263 = ( n3769 & ~n10261 ) | ( n3769 & n10262 ) | ( ~n10261 & n10262 ) ;
  assign n10264 = n10261 | n10263 ;
  assign n10265 = n607 & n9947 ;
  assign n10266 = n1250 & n9945 ;
  assign n10267 = n10265 | n10266 ;
  assign n10268 = n606 & ~n9943 ;
  assign n10269 = ( n606 & n10267 ) | ( n606 & ~n10268 ) | ( n10267 & ~n10268 ) ;
  assign n10270 = ( n9943 & ~n9945 ) | ( n9943 & n10033 ) | ( ~n9945 & n10033 ) ;
  assign n10271 = ( n9945 & ~n10034 ) | ( n9945 & n10270 ) | ( ~n10034 & n10270 ) ;
  assign n10272 = n1248 & n10271 ;
  assign n10273 = n10269 | n10272 ;
  assign n10274 = ( n10243 & n10264 ) | ( n10243 & n10273 ) | ( n10264 & n10273 ) ;
  assign n10275 = ( n10107 & n10243 ) | ( n10107 & ~n10274 ) | ( n10243 & ~n10274 ) ;
  assign n10276 = ( n10107 & n10162 ) | ( n10107 & n10166 ) | ( n10162 & n10166 ) ;
  assign n10277 = ( n10166 & n10167 ) | ( n10166 & ~n10276 ) | ( n10167 & ~n10276 ) ;
  assign n10278 = n607 & n9943 ;
  assign n10279 = n1250 & ~n9941 ;
  assign n10280 = n10278 | n10279 ;
  assign n10281 = n606 & n9883 ;
  assign n10282 = ( n606 & n10280 ) | ( n606 & ~n10281 ) | ( n10280 & ~n10281 ) ;
  assign n10283 = ( n9883 & n9941 ) | ( n9883 & ~n10036 ) | ( n9941 & ~n10036 ) ;
  assign n10284 = ( n10035 & n10036 ) | ( n10035 & ~n10283 ) | ( n10036 & ~n10283 ) ;
  assign n10285 = n1248 & n10284 ;
  assign n10286 = n10282 | n10285 ;
  assign n10287 = ( n10275 & n10277 ) | ( n10275 & ~n10286 ) | ( n10277 & ~n10286 ) ;
  assign n10288 = ( ~n311 & n10167 ) | ( ~n311 & n10176 ) | ( n10167 & n10176 ) ;
  assign n10289 = ( n311 & ~n10177 ) | ( n311 & n10288 ) | ( ~n10177 & n10288 ) ;
  assign n10290 = n197 | n540 ;
  assign n10291 = ( n455 & n463 ) | ( n455 & ~n10290 ) | ( n463 & ~n10290 ) ;
  assign n10292 = n10290 | n10291 ;
  assign n10293 = n1213 | n1420 ;
  assign n10294 = n406 | n10293 ;
  assign n10295 = ( n1288 & n10292 ) | ( n1288 & ~n10294 ) | ( n10292 & ~n10294 ) ;
  assign n10296 = ~n10292 & n10295 ;
  assign n10297 = n9928 & n10296 ;
  assign n10298 = n9928 | n10296 ;
  assign n10299 = ~n10297 & n10298 ;
  assign n10300 = ( n10052 & n10055 ) | ( n10052 & ~n10299 ) | ( n10055 & ~n10299 ) ;
  assign n10301 = ( n10052 & ~n10055 ) | ( n10052 & n10299 ) | ( ~n10055 & n10299 ) ;
  assign n10302 = ( ~n10052 & n10300 ) | ( ~n10052 & n10301 ) | ( n10300 & n10301 ) ;
  assign n10303 = ( n10057 & n10062 ) | ( n10057 & n10302 ) | ( n10062 & n10302 ) ;
  assign n10304 = ( ~n10057 & n10062 ) | ( ~n10057 & n10302 ) | ( n10062 & n10302 ) ;
  assign n10305 = ( n10057 & ~n10303 ) | ( n10057 & n10304 ) | ( ~n10303 & n10304 ) ;
  assign n10306 = n3800 & ~n10305 ;
  assign n10307 = n3799 & ~n10302 ;
  assign n10308 = n3700 & ~n9937 ;
  assign n10309 = n3802 & ~n10057 ;
  assign n10310 = n10308 | n10309 ;
  assign n10311 = ( ~n10306 & n10307 ) | ( ~n10306 & n10310 ) | ( n10307 & n10310 ) ;
  assign n10312 = ( ~x29 & n10306 ) | ( ~x29 & n10311 ) | ( n10306 & n10311 ) ;
  assign n10313 = ( n10306 & n10311 ) | ( n10306 & ~n10312 ) | ( n10311 & ~n10312 ) ;
  assign n10314 = ( x29 & n10312 ) | ( x29 & ~n10313 ) | ( n10312 & ~n10313 ) ;
  assign n10315 = ( ~n10287 & n10289 ) | ( ~n10287 & n10314 ) | ( n10289 & n10314 ) ;
  assign n10316 = ( n311 & ~n605 ) | ( n311 & n10042 ) | ( ~n605 & n10042 ) ;
  assign n10317 = ( n605 & ~n10043 ) | ( n605 & n10316 ) | ( ~n10043 & n10316 ) ;
  assign n10318 = ( n10177 & n10315 ) | ( n10177 & n10317 ) | ( n10315 & n10317 ) ;
  assign n10319 = n851 | n3711 ;
  assign n10320 = ( ~n1560 & n2543 ) | ( ~n1560 & n2943 ) | ( n2543 & n2943 ) ;
  assign n10321 = ( n1560 & ~n6091 ) | ( n1560 & n10320 ) | ( ~n6091 & n10320 ) ;
  assign n10322 = n6091 | n10321 ;
  assign n10323 = ( ~n3757 & n10264 ) | ( ~n3757 & n10322 ) | ( n10264 & n10322 ) ;
  assign n10324 = n1620 | n2029 ;
  assign n10325 = ( n320 & n1169 ) | ( n320 & ~n1547 ) | ( n1169 & ~n1547 ) ;
  assign n10326 = n1547 | n10325 ;
  assign n10327 = n317 | n956 ;
  assign n10328 = n890 | n10327 ;
  assign n10329 = ( n4410 & ~n10326 ) | ( n4410 & n10328 ) | ( ~n10326 & n10328 ) ;
  assign n10330 = n10326 | n10329 ;
  assign n10331 = ( n4065 & ~n10324 ) | ( n4065 & n10330 ) | ( ~n10324 & n10330 ) ;
  assign n10332 = n10324 | n10331 ;
  assign n10333 = n1079 | n1720 ;
  assign n10334 = n489 | n839 ;
  assign n10335 = n226 | n362 ;
  assign n10336 = ( n1511 & ~n10334 ) | ( n1511 & n10335 ) | ( ~n10334 & n10335 ) ;
  assign n10337 = n10334 | n10336 ;
  assign n10338 = ( ~n6109 & n10333 ) | ( ~n6109 & n10337 ) | ( n10333 & n10337 ) ;
  assign n10339 = ( n2181 & n6109 ) | ( n2181 & ~n10338 ) | ( n6109 & ~n10338 ) ;
  assign n10340 = n10338 | n10339 ;
  assign n10341 = ( ~n10322 & n10332 ) | ( ~n10322 & n10340 ) | ( n10332 & n10340 ) ;
  assign n10342 = ( ~n3757 & n10323 ) | ( ~n3757 & n10341 ) | ( n10323 & n10341 ) ;
  assign n10343 = n3757 | n10342 ;
  assign n10344 = ( n3639 & ~n10319 ) | ( n3639 & n10343 ) | ( ~n10319 & n10343 ) ;
  assign n10345 = n10319 | n10344 ;
  assign n10346 = ( ~n10297 & n10300 ) | ( ~n10297 & n10345 ) | ( n10300 & n10345 ) ;
  assign n10347 = ( n10302 & n10303 ) | ( n10302 & ~n10346 ) | ( n10303 & ~n10346 ) ;
  assign n10348 = n10346 & ~n10347 ;
  assign n10349 = n3800 & n10348 ;
  assign n10350 = n3700 & ~n10302 ;
  assign n10351 = n3799 | n10350 ;
  assign n10352 = ( n3802 & ~n10349 ) | ( n3802 & n10351 ) | ( ~n10349 & n10351 ) ;
  assign n10353 = ( ~x29 & n10349 ) | ( ~x29 & n10352 ) | ( n10349 & n10352 ) ;
  assign n10354 = ( n10349 & n10352 ) | ( n10349 & ~n10353 ) | ( n10352 & ~n10353 ) ;
  assign n10355 = ( x29 & n10353 ) | ( x29 & ~n10354 ) | ( n10353 & ~n10354 ) ;
  assign n10356 = ( ~n10069 & n10318 ) | ( ~n10069 & n10355 ) | ( n10318 & n10355 ) ;
  assign n10357 = ( n10069 & n10318 ) | ( n10069 & n10355 ) | ( n10318 & n10355 ) ;
  assign n10358 = ( n10069 & n10356 ) | ( n10069 & ~n10357 ) | ( n10356 & ~n10357 ) ;
  assign n10359 = ( n10177 & ~n10315 ) | ( n10177 & n10317 ) | ( ~n10315 & n10317 ) ;
  assign n10360 = ( n10315 & ~n10318 ) | ( n10315 & n10359 ) | ( ~n10318 & n10359 ) ;
  assign n10361 = ( ~n10302 & n10303 ) | ( ~n10302 & n10346 ) | ( n10303 & n10346 ) ;
  assign n10362 = ( ~n10303 & n10347 ) | ( ~n10303 & n10361 ) | ( n10347 & n10361 ) ;
  assign n10363 = n3800 & n10362 ;
  assign n10364 = n3799 & n10346 ;
  assign n10365 = n3700 & ~n10057 ;
  assign n10366 = n3802 & ~n10302 ;
  assign n10367 = n10365 | n10366 ;
  assign n10368 = ( ~n10363 & n10364 ) | ( ~n10363 & n10367 ) | ( n10364 & n10367 ) ;
  assign n10369 = ( ~x29 & n10363 ) | ( ~x29 & n10368 ) | ( n10363 & n10368 ) ;
  assign n10370 = ( n10363 & n10368 ) | ( n10363 & ~n10369 ) | ( n10368 & ~n10369 ) ;
  assign n10371 = ( x29 & n10369 ) | ( x29 & ~n10370 ) | ( n10369 & ~n10370 ) ;
  assign n10372 = ( n38 & n10360 ) | ( n38 & n10371 ) | ( n10360 & n10371 ) ;
  assign n10373 = n3800 & n10040 ;
  assign n10374 = n3799 & ~n9937 ;
  assign n10375 = n3700 & ~n9883 ;
  assign n10376 = n3802 & n9916 ;
  assign n10377 = n10375 | n10376 ;
  assign n10378 = ( ~n10373 & n10374 ) | ( ~n10373 & n10377 ) | ( n10374 & n10377 ) ;
  assign n10379 = ( ~x29 & n10373 ) | ( ~x29 & n10378 ) | ( n10373 & n10378 ) ;
  assign n10380 = ( n10373 & n10378 ) | ( n10373 & ~n10379 ) | ( n10378 & ~n10379 ) ;
  assign n10381 = ( x29 & n10379 ) | ( x29 & ~n10380 ) | ( n10379 & ~n10380 ) ;
  assign n10382 = ( n10107 & ~n10243 ) | ( n10107 & n10274 ) | ( ~n10243 & n10274 ) ;
  assign n10383 = ( ~n10107 & n10275 ) | ( ~n10107 & n10382 ) | ( n10275 & n10382 ) ;
  assign n10384 = n607 & n9945 ;
  assign n10385 = n1250 & n9943 ;
  assign n10386 = n10384 | n10385 ;
  assign n10387 = n606 & n9941 ;
  assign n10388 = ( n606 & n10386 ) | ( n606 & ~n10387 ) | ( n10386 & ~n10387 ) ;
  assign n10389 = ( n9941 & ~n9943 ) | ( n9941 & n10034 ) | ( ~n9943 & n10034 ) ;
  assign n10390 = ( ~n10034 & n10035 ) | ( ~n10034 & n10389 ) | ( n10035 & n10389 ) ;
  assign n10391 = n1248 & n10390 ;
  assign n10392 = ( n1248 & n10388 ) | ( n1248 & ~n10391 ) | ( n10388 & ~n10391 ) ;
  assign n10393 = ( n10381 & n10383 ) | ( n10381 & n10392 ) | ( n10383 & n10392 ) ;
  assign n10394 = ( n10275 & n10277 ) | ( n10275 & n10286 ) | ( n10277 & n10286 ) ;
  assign n10395 = ( n10286 & n10287 ) | ( n10286 & ~n10394 ) | ( n10287 & ~n10394 ) ;
  assign n10396 = n3800 & ~n10064 ;
  assign n10397 = n3799 & ~n10057 ;
  assign n10398 = n3700 & n9916 ;
  assign n10399 = n3802 & ~n9937 ;
  assign n10400 = n10398 | n10399 ;
  assign n10401 = ( ~n10396 & n10397 ) | ( ~n10396 & n10400 ) | ( n10397 & n10400 ) ;
  assign n10402 = ( ~x29 & n10396 ) | ( ~x29 & n10401 ) | ( n10396 & n10401 ) ;
  assign n10403 = ( n10396 & n10401 ) | ( n10396 & ~n10402 ) | ( n10401 & ~n10402 ) ;
  assign n10404 = ( x29 & n10402 ) | ( x29 & ~n10403 ) | ( n10402 & ~n10403 ) ;
  assign n10405 = ( n10393 & n10395 ) | ( n10393 & n10404 ) | ( n10395 & n10404 ) ;
  assign n10406 = n4195 | n10346 ;
  assign n10407 = ( n4200 & n4202 ) | ( n4200 & n10406 ) | ( n4202 & n10406 ) ;
  assign n10408 = n4201 | n4345 ;
  assign n10409 = ( x26 & n10407 ) | ( x26 & ~n10408 ) | ( n10407 & ~n10408 ) ;
  assign n10410 = ( ~x26 & n10407 ) | ( ~x26 & n10408 ) | ( n10407 & n10408 ) ;
  assign n10411 = ( ~n10407 & n10409 ) | ( ~n10407 & n10410 ) | ( n10409 & n10410 ) ;
  assign n10412 = ( n10289 & n10314 ) | ( n10289 & ~n10315 ) | ( n10314 & ~n10315 ) ;
  assign n10413 = ( n10287 & n10315 ) | ( n10287 & ~n10412 ) | ( n10315 & ~n10412 ) ;
  assign n10414 = ( n10405 & n10411 ) | ( n10405 & ~n10413 ) | ( n10411 & ~n10413 ) ;
  assign n10415 = ( n83 & n98 ) | ( n83 & n100 ) | ( n98 & n100 ) ;
  assign n10416 = ( ~n78 & n97 ) | ( ~n78 & n122 ) | ( n97 & n122 ) ;
  assign n10417 = n10415 | n10416 ;
  assign n10418 = ( n44 & n73 ) | ( n44 & n98 ) | ( n73 & n98 ) ;
  assign n10419 = ( n217 & n444 ) | ( n217 & ~n10418 ) | ( n444 & ~n10418 ) ;
  assign n10420 = n10418 | n10419 ;
  assign n10421 = ( n3485 & ~n10417 ) | ( n3485 & n10420 ) | ( ~n10417 & n10420 ) ;
  assign n10422 = ( n1565 & n10417 ) | ( n1565 & ~n10421 ) | ( n10417 & ~n10421 ) ;
  assign n10423 = n10421 | n10422 ;
  assign n10424 = n1323 | n1929 ;
  assign n10425 = ( n712 & n2726 ) | ( n712 & ~n10424 ) | ( n2726 & ~n10424 ) ;
  assign n10426 = n10424 | n10425 ;
  assign n10427 = ( n2869 & ~n10423 ) | ( n2869 & n10426 ) | ( ~n10423 & n10426 ) ;
  assign n10428 = n10423 | n10427 ;
  assign n10429 = ( n150 & ~n1754 ) | ( n150 & n2883 ) | ( ~n1754 & n2883 ) ;
  assign n10430 = n1754 | n10429 ;
  assign n10431 = n745 | n1092 ;
  assign n10432 = n686 | n931 ;
  assign n10433 = ( n2292 & n10431 ) | ( n2292 & ~n10432 ) | ( n10431 & ~n10432 ) ;
  assign n10434 = ( n2878 & n10432 ) | ( n2878 & ~n10433 ) | ( n10432 & ~n10433 ) ;
  assign n10435 = n10433 | n10434 ;
  assign n10436 = n266 | n332 ;
  assign n10437 = n1171 | n10436 ;
  assign n10438 = n1174 | n1473 ;
  assign n10439 = n230 | n824 ;
  assign n10440 = ( n697 & n4503 ) | ( n697 & ~n10439 ) | ( n4503 & ~n10439 ) ;
  assign n10441 = n10439 | n10440 ;
  assign n10442 = ( ~n10437 & n10438 ) | ( ~n10437 & n10441 ) | ( n10438 & n10441 ) ;
  assign n10443 = n10437 | n10442 ;
  assign n10444 = ( ~n10430 & n10435 ) | ( ~n10430 & n10443 ) | ( n10435 & n10443 ) ;
  assign n10445 = n10430 | n10444 ;
  assign n10446 = ( n5131 & n10428 ) | ( n5131 & ~n10445 ) | ( n10428 & ~n10445 ) ;
  assign n10447 = ~n10428 & n10446 ;
  assign n10448 = n607 & n9951 ;
  assign n10449 = n1250 & n9949 ;
  assign n10450 = n10448 | n10449 ;
  assign n10451 = n606 & ~n9947 ;
  assign n10452 = ( n606 & n10450 ) | ( n606 & ~n10451 ) | ( n10450 & ~n10451 ) ;
  assign n10453 = ( n9947 & ~n9949 ) | ( n9947 & n10031 ) | ( ~n9949 & n10031 ) ;
  assign n10454 = ( n9949 & ~n10032 ) | ( n9949 & n10453 ) | ( ~n10032 & n10453 ) ;
  assign n10455 = n1248 & n10454 ;
  assign n10456 = n10452 | n10455 ;
  assign n10457 = ( n10212 & ~n10447 ) | ( n10212 & n10456 ) | ( ~n10447 & n10456 ) ;
  assign n10458 = ( n10212 & n10239 ) | ( n10212 & ~n10242 ) | ( n10239 & ~n10242 ) ;
  assign n10459 = ( n10242 & ~n10243 ) | ( n10242 & n10458 ) | ( ~n10243 & n10458 ) ;
  assign n10460 = n607 & n9949 ;
  assign n10461 = n1250 & n9947 ;
  assign n10462 = n10460 | n10461 ;
  assign n10463 = n606 & ~n9945 ;
  assign n10464 = ( n606 & n10462 ) | ( n606 & ~n10463 ) | ( n10462 & ~n10463 ) ;
  assign n10465 = ( n9945 & ~n9947 ) | ( n9945 & n10032 ) | ( ~n9947 & n10032 ) ;
  assign n10466 = ( n9947 & ~n10033 ) | ( n9947 & n10465 ) | ( ~n10033 & n10465 ) ;
  assign n10467 = n1248 & n10466 ;
  assign n10468 = n10464 | n10467 ;
  assign n10469 = ( n10457 & ~n10459 ) | ( n10457 & n10468 ) | ( ~n10459 & n10468 ) ;
  assign n10470 = ( ~n10243 & n10264 ) | ( ~n10243 & n10273 ) | ( n10264 & n10273 ) ;
  assign n10471 = ( n10243 & ~n10274 ) | ( n10243 & n10470 ) | ( ~n10274 & n10470 ) ;
  assign n10472 = n3800 & n10174 ;
  assign n10473 = n3799 & n9916 ;
  assign n10474 = n3700 | n9941 ;
  assign n10475 = n3802 & ~n9883 ;
  assign n10476 = ( ~n9941 & n10474 ) | ( ~n9941 & n10475 ) | ( n10474 & n10475 ) ;
  assign n10477 = ( ~n10472 & n10473 ) | ( ~n10472 & n10476 ) | ( n10473 & n10476 ) ;
  assign n10478 = ( ~x29 & n10472 ) | ( ~x29 & n10477 ) | ( n10472 & n10477 ) ;
  assign n10479 = ( n10472 & n10477 ) | ( n10472 & ~n10478 ) | ( n10477 & ~n10478 ) ;
  assign n10480 = ( x29 & n10478 ) | ( x29 & ~n10479 ) | ( n10478 & ~n10479 ) ;
  assign n10481 = ( n10469 & n10471 ) | ( n10469 & n10480 ) | ( n10471 & n10480 ) ;
  assign n10482 = ( n10381 & ~n10383 ) | ( n10381 & n10392 ) | ( ~n10383 & n10392 ) ;
  assign n10483 = ( n10383 & ~n10393 ) | ( n10383 & n10482 ) | ( ~n10393 & n10482 ) ;
  assign n10484 = n4202 & n10362 ;
  assign n10485 = n4201 & n10346 ;
  assign n10486 = n4200 & ~n10057 ;
  assign n10487 = n4345 & ~n10302 ;
  assign n10488 = n10486 | n10487 ;
  assign n10489 = ( ~n10484 & n10485 ) | ( ~n10484 & n10488 ) | ( n10485 & n10488 ) ;
  assign n10490 = ( ~x26 & n10484 ) | ( ~x26 & n10489 ) | ( n10484 & n10489 ) ;
  assign n10491 = ( n10484 & n10489 ) | ( n10484 & ~n10490 ) | ( n10489 & ~n10490 ) ;
  assign n10492 = ( x26 & n10490 ) | ( x26 & ~n10491 ) | ( n10490 & ~n10491 ) ;
  assign n10493 = ( n10481 & n10483 ) | ( n10481 & n10492 ) | ( n10483 & n10492 ) ;
  assign n10494 = ( n10393 & ~n10395 ) | ( n10393 & n10404 ) | ( ~n10395 & n10404 ) ;
  assign n10495 = ( n10395 & ~n10405 ) | ( n10395 & n10494 ) | ( ~n10405 & n10494 ) ;
  assign n10496 = n4202 & n10348 ;
  assign n10497 = n4345 & n10346 ;
  assign n10498 = n4200 & ~n10302 ;
  assign n10499 = n4201 | n10498 ;
  assign n10500 = ( ~n10496 & n10497 ) | ( ~n10496 & n10499 ) | ( n10497 & n10499 ) ;
  assign n10501 = ( ~x26 & n10496 ) | ( ~x26 & n10500 ) | ( n10496 & n10500 ) ;
  assign n10502 = ( n10496 & n10500 ) | ( n10496 & ~n10501 ) | ( n10500 & ~n10501 ) ;
  assign n10503 = ( x26 & n10501 ) | ( x26 & ~n10502 ) | ( n10501 & ~n10502 ) ;
  assign n10504 = ( n10493 & n10495 ) | ( n10493 & n10503 ) | ( n10495 & n10503 ) ;
  assign n10505 = n2407 | n3328 ;
  assign n10506 = ( n73 & n84 ) | ( n73 & n122 ) | ( n84 & n122 ) ;
  assign n10507 = ( n177 & n435 ) | ( n177 & ~n10506 ) | ( n435 & ~n10506 ) ;
  assign n10508 = n10506 | n10507 ;
  assign n10509 = ( n5201 & ~n10505 ) | ( n5201 & n10508 ) | ( ~n10505 & n10508 ) ;
  assign n10510 = n10505 | n10509 ;
  assign n10511 = ( ~n3237 & n4024 ) | ( ~n3237 & n10510 ) | ( n4024 & n10510 ) ;
  assign n10512 = n566 | n675 ;
  assign n10513 = ( n995 & n1376 ) | ( n995 & ~n10512 ) | ( n1376 & ~n10512 ) ;
  assign n10514 = n10512 | n10513 ;
  assign n10515 = ( ~n2398 & n3568 ) | ( ~n2398 & n10514 ) | ( n3568 & n10514 ) ;
  assign n10516 = ~n10514 & n10515 ;
  assign n10517 = n299 | n1366 ;
  assign n10518 = n684 | n884 ;
  assign n10519 = n10517 | n10518 ;
  assign n10520 = n1027 | n1225 ;
  assign n10521 = n1235 | n1940 ;
  assign n10522 = ( n288 & n1488 ) | ( n288 & ~n10521 ) | ( n1488 & ~n10521 ) ;
  assign n10523 = n10521 | n10522 ;
  assign n10524 = ( ~n10519 & n10520 ) | ( ~n10519 & n10523 ) | ( n10520 & n10523 ) ;
  assign n10525 = n10519 | n10524 ;
  assign n10526 = ( n10510 & n10516 ) | ( n10510 & ~n10525 ) | ( n10516 & ~n10525 ) ;
  assign n10527 = ( n3237 & ~n10511 ) | ( n3237 & n10526 ) | ( ~n10511 & n10526 ) ;
  assign n10528 = ~n3237 & n10527 ;
  assign n10529 = ( x17 & n5507 ) | ( x17 & n5666 ) | ( n5507 & n5666 ) ;
  assign n10530 = n5507 | n5666 ;
  assign n10531 = x16 | n10530 ;
  assign n10532 = ~n10529 & n10531 ;
  assign n10533 = ( n775 & n952 ) | ( n775 & ~n3034 ) | ( n952 & ~n3034 ) ;
  assign n10534 = n3034 | n10533 ;
  assign n10535 = n943 | n2628 ;
  assign n10536 = n466 | n2443 ;
  assign n10537 = n81 | n576 ;
  assign n10538 = n153 | n549 ;
  assign n10539 = ( n1003 & ~n10537 ) | ( n1003 & n10538 ) | ( ~n10537 & n10538 ) ;
  assign n10540 = n10537 | n10539 ;
  assign n10541 = ( ~n10535 & n10536 ) | ( ~n10535 & n10540 ) | ( n10536 & n10540 ) ;
  assign n10542 = n10535 | n10541 ;
  assign n10543 = ( n10113 & ~n10534 ) | ( n10113 & n10542 ) | ( ~n10534 & n10542 ) ;
  assign n10544 = n6087 | n10543 ;
  assign n10545 = ( n10186 & n10534 ) | ( n10186 & ~n10544 ) | ( n10534 & ~n10544 ) ;
  assign n10546 = n10544 | n10545 ;
  assign n10547 = ( n624 & ~n4860 ) | ( n624 & n10546 ) | ( ~n4860 & n10546 ) ;
  assign n10548 = ( n3426 & n4860 ) | ( n3426 & ~n10547 ) | ( n4860 & ~n10547 ) ;
  assign n10549 = n10547 | n10548 ;
  assign n10550 = ( n10528 & n10532 ) | ( n10528 & ~n10549 ) | ( n10532 & ~n10549 ) ;
  assign n10551 = n607 & ~n9953 ;
  assign n10552 = n1250 & n9951 ;
  assign n10553 = n10551 | n10552 ;
  assign n10554 = n606 & ~n9949 ;
  assign n10555 = ( n606 & n10553 ) | ( n606 & ~n10554 ) | ( n10553 & ~n10554 ) ;
  assign n10556 = ( n9949 & ~n9951 ) | ( n9949 & n10030 ) | ( ~n9951 & n10030 ) ;
  assign n10557 = ( n9951 & ~n10031 ) | ( n9951 & n10556 ) | ( ~n10031 & n10556 ) ;
  assign n10558 = n1248 & n10557 ;
  assign n10559 = n10555 | n10558 ;
  assign n10560 = ( n10212 & ~n10550 ) | ( n10212 & n10559 ) | ( ~n10550 & n10559 ) ;
  assign n10561 = n607 & n9959 ;
  assign n10562 = n1250 & ~n9957 ;
  assign n10563 = n10561 | n10562 ;
  assign n10564 = n606 & ~n9955 ;
  assign n10565 = ( n606 & n10563 ) | ( n606 & ~n10564 ) | ( n10563 & ~n10564 ) ;
  assign n10566 = ( ~n9955 & n9957 ) | ( ~n9955 & n10027 ) | ( n9957 & n10027 ) ;
  assign n10567 = ( ~n10027 & n10028 ) | ( ~n10027 & n10566 ) | ( n10028 & n10566 ) ;
  assign n10568 = n1248 & ~n10567 ;
  assign n10569 = n10565 | n10568 ;
  assign n10570 = ( n262 & n3484 ) | ( n262 & ~n10134 ) | ( n3484 & ~n10134 ) ;
  assign n10571 = n10134 | n10570 ;
  assign n10572 = n712 | n10218 ;
  assign n10573 = n449 | n540 ;
  assign n10574 = n512 | n10573 ;
  assign n10575 = ( n819 & ~n10572 ) | ( n819 & n10574 ) | ( ~n10572 & n10574 ) ;
  assign n10576 = n10572 | n10575 ;
  assign n10577 = ( ~n3556 & n10571 ) | ( ~n3556 & n10576 ) | ( n10571 & n10576 ) ;
  assign n10578 = ( n100 & n102 ) | ( n100 & n136 ) | ( n102 & n136 ) ;
  assign n10579 = ( n83 & n84 ) | ( n83 & n109 ) | ( n84 & n109 ) ;
  assign n10580 = n215 | n10579 ;
  assign n10581 = ( n346 & ~n10578 ) | ( n346 & n10580 ) | ( ~n10578 & n10580 ) ;
  assign n10582 = n10578 | n10581 ;
  assign n10583 = n991 | n3317 ;
  assign n10584 = ( n625 & n961 ) | ( n625 & ~n991 ) | ( n961 & ~n991 ) ;
  assign n10585 = ( ~n10582 & n10583 ) | ( ~n10582 & n10584 ) | ( n10583 & n10584 ) ;
  assign n10586 = n10582 | n10585 ;
  assign n10587 = ( n50 & n64 ) | ( n50 & n149 ) | ( n64 & n149 ) ;
  assign n10588 = ( n485 & n2302 ) | ( n485 & ~n10587 ) | ( n2302 & ~n10587 ) ;
  assign n10589 = n10587 | n10588 ;
  assign n10590 = n2628 | n3303 ;
  assign n10591 = ( n2882 & ~n10589 ) | ( n2882 & n10590 ) | ( ~n10589 & n10590 ) ;
  assign n10592 = n10589 | n10591 ;
  assign n10593 = ( ~n10576 & n10586 ) | ( ~n10576 & n10592 ) | ( n10586 & n10592 ) ;
  assign n10594 = ( ~n3556 & n10577 ) | ( ~n3556 & n10593 ) | ( n10577 & n10593 ) ;
  assign n10595 = n3556 | n10594 ;
  assign n10596 = ( n153 & n331 ) | ( n153 & ~n5074 ) | ( n331 & ~n5074 ) ;
  assign n10597 = n5074 | n10596 ;
  assign n10598 = n195 | n5208 ;
  assign n10599 = n492 | n764 ;
  assign n10600 = n1001 | n1031 ;
  assign n10601 = ( ~n524 & n957 ) | ( ~n524 & n10600 ) | ( n957 & n10600 ) ;
  assign n10602 = ( n524 & ~n10599 ) | ( n524 & n10601 ) | ( ~n10599 & n10601 ) ;
  assign n10603 = n10599 | n10602 ;
  assign n10604 = n1171 | n1185 ;
  assign n10605 = ( ~n10598 & n10603 ) | ( ~n10598 & n10604 ) | ( n10603 & n10604 ) ;
  assign n10606 = n10598 | n10605 ;
  assign n10607 = ( n2213 & ~n3529 ) | ( n2213 & n10606 ) | ( ~n3529 & n10606 ) ;
  assign n10608 = n1542 | n10607 ;
  assign n10609 = ( n3529 & ~n10597 ) | ( n3529 & n10608 ) | ( ~n10597 & n10608 ) ;
  assign n10610 = n10597 | n10609 ;
  assign n10611 = ( n48 & n75 ) | ( n48 & n98 ) | ( n75 & n98 ) ;
  assign n10612 = n104 | n10611 ;
  assign n10613 = n112 | n921 ;
  assign n10614 = ( n136 & n149 ) | ( n136 & n152 ) | ( n149 & n152 ) ;
  assign n10615 = ( ~n10612 & n10613 ) | ( ~n10612 & n10614 ) | ( n10613 & n10614 ) ;
  assign n10616 = n10612 | n10615 ;
  assign n10617 = n1810 | n3970 ;
  assign n10618 = n1346 | n1556 ;
  assign n10619 = n230 | n1082 ;
  assign n10620 = ( n690 & ~n1793 ) | ( n690 & n10619 ) | ( ~n1793 & n10619 ) ;
  assign n10621 = ( n1793 & ~n10618 ) | ( n1793 & n10620 ) | ( ~n10618 & n10620 ) ;
  assign n10622 = n10618 | n10621 ;
  assign n10623 = ( ~n10616 & n10617 ) | ( ~n10616 & n10622 ) | ( n10617 & n10622 ) ;
  assign n10624 = n10616 | n10623 ;
  assign n10625 = n2776 & ~n6234 ;
  assign n10626 = n175 | n2256 ;
  assign n10627 = n4588 | n10626 ;
  assign n10628 = ( n2737 & n4523 ) | ( n2737 & ~n10627 ) | ( n4523 & ~n10627 ) ;
  assign n10629 = n10627 | n10628 ;
  assign n10630 = ( n10624 & n10625 ) | ( n10624 & ~n10629 ) | ( n10625 & ~n10629 ) ;
  assign n10631 = ~n10624 & n10630 ;
  assign n10632 = n10610 & ~n10631 ;
  assign n10633 = n10610 & n10631 ;
  assign n10634 = ( n10631 & n10632 ) | ( n10631 & ~n10633 ) | ( n10632 & ~n10633 ) ;
  assign n10635 = n5969 | n6464 ;
  assign n10636 = n5965 | n10635 ;
  assign n10637 = n5966 | n10636 ;
  assign n10638 = ( ~x14 & n10634 ) | ( ~x14 & n10637 ) | ( n10634 & n10637 ) ;
  assign n10639 = ( n10634 & n10637 ) | ( n10634 & ~n10638 ) | ( n10637 & ~n10638 ) ;
  assign n10640 = ( x14 & n10638 ) | ( x14 & ~n10639 ) | ( n10638 & ~n10639 ) ;
  assign n10641 = ( ~n10610 & n10631 ) | ( ~n10610 & n10640 ) | ( n10631 & n10640 ) ;
  assign n10642 = ( n10569 & ~n10595 ) | ( n10569 & n10641 ) | ( ~n10595 & n10641 ) ;
  assign n10643 = ( n10528 & n10569 ) | ( n10528 & ~n10642 ) | ( n10569 & ~n10642 ) ;
  assign n10644 = ( n10528 & n10532 ) | ( n10528 & n10549 ) | ( n10532 & n10549 ) ;
  assign n10645 = ( n10549 & n10550 ) | ( n10549 & ~n10644 ) | ( n10550 & ~n10644 ) ;
  assign n10646 = n607 & n9955 ;
  assign n10647 = n1250 & ~n9953 ;
  assign n10648 = n10646 | n10647 ;
  assign n10649 = n606 & ~n9951 ;
  assign n10650 = ( n606 & n10648 ) | ( n606 & ~n10649 ) | ( n10648 & ~n10649 ) ;
  assign n10651 = ( ~n9951 & n9953 ) | ( ~n9951 & n10029 ) | ( n9953 & n10029 ) ;
  assign n10652 = ( ~n10029 & n10030 ) | ( ~n10029 & n10651 ) | ( n10030 & n10651 ) ;
  assign n10653 = n1248 & ~n10652 ;
  assign n10654 = n10650 | n10653 ;
  assign n10655 = ( n10643 & n10645 ) | ( n10643 & n10654 ) | ( n10645 & n10654 ) ;
  assign n10656 = ( n10212 & n10559 ) | ( n10212 & ~n10560 ) | ( n10559 & ~n10560 ) ;
  assign n10657 = ( n10550 & n10560 ) | ( n10550 & ~n10656 ) | ( n10560 & ~n10656 ) ;
  assign n10658 = n3800 & n10271 ;
  assign n10659 = n3799 & n9943 ;
  assign n10660 = n3700 & n9947 ;
  assign n10661 = n3802 & n9945 ;
  assign n10662 = n10660 | n10661 ;
  assign n10663 = ( ~n10658 & n10659 ) | ( ~n10658 & n10662 ) | ( n10659 & n10662 ) ;
  assign n10664 = ( ~x29 & n10658 ) | ( ~x29 & n10663 ) | ( n10658 & n10663 ) ;
  assign n10665 = ( n10658 & n10663 ) | ( n10658 & ~n10664 ) | ( n10663 & ~n10664 ) ;
  assign n10666 = ( x29 & n10664 ) | ( x29 & ~n10665 ) | ( n10664 & ~n10665 ) ;
  assign n10667 = ( n10655 & ~n10657 ) | ( n10655 & n10666 ) | ( ~n10657 & n10666 ) ;
  assign n10668 = ( n10212 & n10447 ) | ( n10212 & n10456 ) | ( n10447 & n10456 ) ;
  assign n10669 = ( n10447 & n10457 ) | ( n10447 & ~n10668 ) | ( n10457 & ~n10668 ) ;
  assign n10670 = ( n10560 & n10667 ) | ( n10560 & ~n10669 ) | ( n10667 & ~n10669 ) ;
  assign n10671 = ( n10457 & n10459 ) | ( n10457 & n10468 ) | ( n10459 & n10468 ) ;
  assign n10672 = ( n10459 & n10469 ) | ( n10459 & ~n10671 ) | ( n10469 & ~n10671 ) ;
  assign n10673 = n3800 & n10284 ;
  assign n10674 = n3799 & ~n9883 ;
  assign n10675 = n3700 & n9943 ;
  assign n10676 = n3802 & ~n9941 ;
  assign n10677 = n10675 | n10676 ;
  assign n10678 = ( ~n10673 & n10674 ) | ( ~n10673 & n10677 ) | ( n10674 & n10677 ) ;
  assign n10679 = ( ~x29 & n10673 ) | ( ~x29 & n10678 ) | ( n10673 & n10678 ) ;
  assign n10680 = ( n10673 & n10678 ) | ( n10673 & ~n10679 ) | ( n10678 & ~n10679 ) ;
  assign n10681 = ( x29 & n10679 ) | ( x29 & ~n10680 ) | ( n10679 & ~n10680 ) ;
  assign n10682 = ( n10670 & ~n10672 ) | ( n10670 & n10681 ) | ( ~n10672 & n10681 ) ;
  assign n10683 = ( ~n10469 & n10471 ) | ( ~n10469 & n10480 ) | ( n10471 & n10480 ) ;
  assign n10684 = ( n10469 & ~n10481 ) | ( n10469 & n10683 ) | ( ~n10481 & n10683 ) ;
  assign n10685 = n4202 & ~n10305 ;
  assign n10686 = n4201 & ~n10302 ;
  assign n10687 = n4200 & ~n9937 ;
  assign n10688 = n4345 & ~n10057 ;
  assign n10689 = n10687 | n10688 ;
  assign n10690 = ( ~n10685 & n10686 ) | ( ~n10685 & n10689 ) | ( n10686 & n10689 ) ;
  assign n10691 = ( ~x26 & n10685 ) | ( ~x26 & n10690 ) | ( n10685 & n10690 ) ;
  assign n10692 = ( n10685 & n10690 ) | ( n10685 & ~n10691 ) | ( n10690 & ~n10691 ) ;
  assign n10693 = ( x26 & n10691 ) | ( x26 & ~n10692 ) | ( n10691 & ~n10692 ) ;
  assign n10694 = ( n10682 & n10684 ) | ( n10682 & n10693 ) | ( n10684 & n10693 ) ;
  assign n10695 = ( n10481 & ~n10483 ) | ( n10481 & n10492 ) | ( ~n10483 & n10492 ) ;
  assign n10696 = ( n10483 & ~n10493 ) | ( n10483 & n10695 ) | ( ~n10493 & n10695 ) ;
  assign n10697 = ( x20 & ~x23 ) | ( x20 & n10165 ) | ( ~x23 & n10165 ) ;
  assign n10698 = ( ~x23 & n4704 ) | ( ~x23 & n10697 ) | ( n4704 & n10697 ) ;
  assign n10699 = ( n10694 & n10696 ) | ( n10694 & n10698 ) | ( n10696 & n10698 ) ;
  assign n10700 = n4202 & n10040 ;
  assign n10701 = n4201 & ~n9937 ;
  assign n10702 = n4200 & ~n9883 ;
  assign n10703 = n4345 & n9916 ;
  assign n10704 = n10702 | n10703 ;
  assign n10705 = ( ~n10700 & n10701 ) | ( ~n10700 & n10704 ) | ( n10701 & n10704 ) ;
  assign n10706 = ( ~x26 & n10700 ) | ( ~x26 & n10705 ) | ( n10700 & n10705 ) ;
  assign n10707 = ( n10700 & n10705 ) | ( n10700 & ~n10706 ) | ( n10705 & ~n10706 ) ;
  assign n10708 = ( x26 & n10706 ) | ( x26 & ~n10707 ) | ( n10706 & ~n10707 ) ;
  assign n10709 = ( n10560 & n10667 ) | ( n10560 & n10669 ) | ( n10667 & n10669 ) ;
  assign n10710 = ( n10669 & n10670 ) | ( n10669 & ~n10709 ) | ( n10670 & ~n10709 ) ;
  assign n10711 = n3800 & ~n10390 ;
  assign n10712 = n3799 & ~n9941 ;
  assign n10713 = n3700 & n9945 ;
  assign n10714 = n3802 & n9943 ;
  assign n10715 = n10713 | n10714 ;
  assign n10716 = ( ~n10711 & n10712 ) | ( ~n10711 & n10715 ) | ( n10712 & n10715 ) ;
  assign n10717 = ( ~x29 & n10711 ) | ( ~x29 & n10716 ) | ( n10711 & n10716 ) ;
  assign n10718 = ( n10711 & n10716 ) | ( n10711 & ~n10717 ) | ( n10716 & ~n10717 ) ;
  assign n10719 = ( x29 & n10717 ) | ( x29 & ~n10718 ) | ( n10717 & ~n10718 ) ;
  assign n10720 = ( n10708 & ~n10710 ) | ( n10708 & n10719 ) | ( ~n10710 & n10719 ) ;
  assign n10721 = ( ~n10670 & n10672 ) | ( ~n10670 & n10681 ) | ( n10672 & n10681 ) ;
  assign n10722 = ( ~n10681 & n10682 ) | ( ~n10681 & n10721 ) | ( n10682 & n10721 ) ;
  assign n10723 = n4202 & ~n10064 ;
  assign n10724 = n4201 & ~n10057 ;
  assign n10725 = n4200 & n9916 ;
  assign n10726 = n4345 & ~n9937 ;
  assign n10727 = n10725 | n10726 ;
  assign n10728 = ( ~n10723 & n10724 ) | ( ~n10723 & n10727 ) | ( n10724 & n10727 ) ;
  assign n10729 = ( ~x26 & n10723 ) | ( ~x26 & n10728 ) | ( n10723 & n10728 ) ;
  assign n10730 = ( n10723 & n10728 ) | ( n10723 & ~n10729 ) | ( n10728 & ~n10729 ) ;
  assign n10731 = ( x26 & n10729 ) | ( x26 & ~n10730 ) | ( n10729 & ~n10730 ) ;
  assign n10732 = ( n10720 & ~n10722 ) | ( n10720 & n10731 ) | ( ~n10722 & n10731 ) ;
  assign n10733 = ( ~n10682 & n10684 ) | ( ~n10682 & n10693 ) | ( n10684 & n10693 ) ;
  assign n10734 = ( n10682 & ~n10694 ) | ( n10682 & n10733 ) | ( ~n10694 & n10733 ) ;
  assign n10735 = n4709 & ~n10346 ;
  assign n10736 = ( n4709 & n10164 ) | ( n4709 & ~n10735 ) | ( n10164 & ~n10735 ) ;
  assign n10737 = ( ~x23 & n4713 ) | ( ~x23 & n10736 ) | ( n4713 & n10736 ) ;
  assign n10738 = ( n4713 & n10736 ) | ( n4713 & ~n10737 ) | ( n10736 & ~n10737 ) ;
  assign n10739 = ( x23 & n10737 ) | ( x23 & ~n10738 ) | ( n10737 & ~n10738 ) ;
  assign n10740 = ( n10732 & n10734 ) | ( n10732 & n10739 ) | ( n10734 & n10739 ) ;
  assign n10741 = ( n10569 & n10595 ) | ( n10569 & n10641 ) | ( n10595 & n10641 ) ;
  assign n10742 = ( n10528 & n10641 ) | ( n10528 & ~n10741 ) | ( n10641 & ~n10741 ) ;
  assign n10743 = ( ~n10528 & n10643 ) | ( ~n10528 & n10742 ) | ( n10643 & n10742 ) ;
  assign n10744 = n607 & ~n9957 ;
  assign n10745 = n1250 & n9955 ;
  assign n10746 = n10744 | n10745 ;
  assign n10747 = n606 & n9953 ;
  assign n10748 = ( n606 & n10746 ) | ( n606 & ~n10747 ) | ( n10746 & ~n10747 ) ;
  assign n10749 = ( n9953 & ~n9955 ) | ( n9953 & n10028 ) | ( ~n9955 & n10028 ) ;
  assign n10750 = ( ~n10028 & n10029 ) | ( ~n10028 & n10749 ) | ( n10029 & n10749 ) ;
  assign n10751 = n1248 & ~n10750 ;
  assign n10752 = n10748 | n10751 ;
  assign n10753 = n3800 & n10454 ;
  assign n10754 = n3799 & n9947 ;
  assign n10755 = n3700 & n9951 ;
  assign n10756 = n3802 & n9949 ;
  assign n10757 = n10755 | n10756 ;
  assign n10758 = ( ~n10753 & n10754 ) | ( ~n10753 & n10757 ) | ( n10754 & n10757 ) ;
  assign n10759 = ( ~x29 & n10753 ) | ( ~x29 & n10758 ) | ( n10753 & n10758 ) ;
  assign n10760 = ( n10753 & n10758 ) | ( n10753 & ~n10759 ) | ( n10758 & ~n10759 ) ;
  assign n10761 = ( x29 & n10759 ) | ( x29 & ~n10760 ) | ( n10759 & ~n10760 ) ;
  assign n10762 = ( ~n10743 & n10752 ) | ( ~n10743 & n10761 ) | ( n10752 & n10761 ) ;
  assign n10763 = n3800 & n10466 ;
  assign n10764 = n3799 & n9945 ;
  assign n10765 = n3700 & n9949 ;
  assign n10766 = n3802 & n9947 ;
  assign n10767 = n10765 | n10766 ;
  assign n10768 = ( ~n10763 & n10764 ) | ( ~n10763 & n10767 ) | ( n10764 & n10767 ) ;
  assign n10769 = ( ~x29 & n10763 ) | ( ~x29 & n10768 ) | ( n10763 & n10768 ) ;
  assign n10770 = ( n10763 & n10768 ) | ( n10763 & ~n10769 ) | ( n10768 & ~n10769 ) ;
  assign n10771 = ( x29 & n10769 ) | ( x29 & ~n10770 ) | ( n10769 & ~n10770 ) ;
  assign n10772 = ( n10643 & ~n10645 ) | ( n10643 & n10654 ) | ( ~n10645 & n10654 ) ;
  assign n10773 = ( n10645 & ~n10655 ) | ( n10645 & n10772 ) | ( ~n10655 & n10772 ) ;
  assign n10774 = ( n10762 & n10771 ) | ( n10762 & n10773 ) | ( n10771 & n10773 ) ;
  assign n10775 = ( n10655 & n10657 ) | ( n10655 & n10666 ) | ( n10657 & n10666 ) ;
  assign n10776 = ( n10657 & n10667 ) | ( n10657 & ~n10775 ) | ( n10667 & ~n10775 ) ;
  assign n10777 = n4202 & n10174 ;
  assign n10778 = n4201 & n9916 ;
  assign n10779 = n4200 | n9941 ;
  assign n10780 = n4345 & ~n9883 ;
  assign n10781 = ( ~n9941 & n10779 ) | ( ~n9941 & n10780 ) | ( n10779 & n10780 ) ;
  assign n10782 = ( ~n10777 & n10778 ) | ( ~n10777 & n10781 ) | ( n10778 & n10781 ) ;
  assign n10783 = ( ~x26 & n10777 ) | ( ~x26 & n10782 ) | ( n10777 & n10782 ) ;
  assign n10784 = ( n10777 & n10782 ) | ( n10777 & ~n10783 ) | ( n10782 & ~n10783 ) ;
  assign n10785 = ( x26 & n10783 ) | ( x26 & ~n10784 ) | ( n10783 & ~n10784 ) ;
  assign n10786 = ( n10774 & ~n10776 ) | ( n10774 & n10785 ) | ( ~n10776 & n10785 ) ;
  assign n10787 = ( n10708 & n10710 ) | ( n10708 & n10719 ) | ( n10710 & n10719 ) ;
  assign n10788 = ( n10710 & n10720 ) | ( n10710 & ~n10787 ) | ( n10720 & ~n10787 ) ;
  assign n10789 = n4713 & n10362 ;
  assign n10790 = n4712 & n10346 ;
  assign n10791 = n4709 & ~n10057 ;
  assign n10792 = n4792 & ~n10302 ;
  assign n10793 = n10791 | n10792 ;
  assign n10794 = ( ~n10789 & n10790 ) | ( ~n10789 & n10793 ) | ( n10790 & n10793 ) ;
  assign n10795 = ( ~x23 & n10789 ) | ( ~x23 & n10794 ) | ( n10789 & n10794 ) ;
  assign n10796 = ( n10789 & n10794 ) | ( n10789 & ~n10795 ) | ( n10794 & ~n10795 ) ;
  assign n10797 = ( x23 & n10795 ) | ( x23 & ~n10796 ) | ( n10795 & ~n10796 ) ;
  assign n10798 = ( n10786 & ~n10788 ) | ( n10786 & n10797 ) | ( ~n10788 & n10797 ) ;
  assign n10799 = ( n10720 & n10722 ) | ( n10720 & n10731 ) | ( n10722 & n10731 ) ;
  assign n10800 = ( n10722 & n10732 ) | ( n10722 & ~n10799 ) | ( n10732 & ~n10799 ) ;
  assign n10801 = n4713 & n10348 ;
  assign n10802 = n4792 & n10346 ;
  assign n10803 = n4709 & ~n10302 ;
  assign n10804 = n4712 | n10803 ;
  assign n10805 = ( ~n10801 & n10802 ) | ( ~n10801 & n10804 ) | ( n10802 & n10804 ) ;
  assign n10806 = ( ~x23 & n10801 ) | ( ~x23 & n10805 ) | ( n10801 & n10805 ) ;
  assign n10807 = ( n10801 & n10805 ) | ( n10801 & ~n10806 ) | ( n10805 & ~n10806 ) ;
  assign n10808 = ( x23 & n10806 ) | ( x23 & ~n10807 ) | ( n10806 & ~n10807 ) ;
  assign n10809 = ( n10798 & ~n10800 ) | ( n10798 & n10808 ) | ( ~n10800 & n10808 ) ;
  assign n10810 = n384 | n1914 ;
  assign n10811 = n2238 | n10810 ;
  assign n10812 = n1550 | n10811 ;
  assign n10813 = n440 | n960 ;
  assign n10814 = n217 | n360 ;
  assign n10815 = ( n3930 & ~n10813 ) | ( n3930 & n10814 ) | ( ~n10813 & n10814 ) ;
  assign n10816 = n10813 | n10815 ;
  assign n10817 = n92 | n176 ;
  assign n10818 = ( n239 & n873 ) | ( n239 & ~n10817 ) | ( n873 & ~n10817 ) ;
  assign n10819 = n10817 | n10818 ;
  assign n10820 = n292 | n1460 ;
  assign n10821 = ( n2077 & ~n10819 ) | ( n2077 & n10820 ) | ( ~n10819 & n10820 ) ;
  assign n10822 = n10819 | n10821 ;
  assign n10823 = ( n487 & ~n10816 ) | ( n487 & n10822 ) | ( ~n10816 & n10822 ) ;
  assign n10824 = n10816 | n10823 ;
  assign n10825 = ( n828 & ~n10812 ) | ( n828 & n10824 ) | ( ~n10812 & n10824 ) ;
  assign n10826 = n10812 | n10825 ;
  assign n10827 = n208 | n450 ;
  assign n10828 = n153 | n851 ;
  assign n10829 = ( n136 & n145 ) | ( n136 & n166 ) | ( n145 & n166 ) ;
  assign n10830 = ( n1824 & ~n10828 ) | ( n1824 & n10829 ) | ( ~n10828 & n10829 ) ;
  assign n10831 = n10828 | n10830 ;
  assign n10832 = ( n66 & n122 ) | ( n66 & n152 ) | ( n122 & n152 ) ;
  assign n10833 = ( n348 & n885 ) | ( n348 & ~n10832 ) | ( n885 & ~n10832 ) ;
  assign n10834 = n10832 | n10833 ;
  assign n10835 = ( ~n10827 & n10831 ) | ( ~n10827 & n10834 ) | ( n10831 & n10834 ) ;
  assign n10836 = n2126 | n2791 ;
  assign n10837 = n499 | n1172 ;
  assign n10838 = n732 | n1237 ;
  assign n10839 = n146 | n300 ;
  assign n10840 = ( n4059 & ~n10838 ) | ( n4059 & n10839 ) | ( ~n10838 & n10839 ) ;
  assign n10841 = n10838 | n10840 ;
  assign n10842 = ( ~n10836 & n10837 ) | ( ~n10836 & n10841 ) | ( n10837 & n10841 ) ;
  assign n10843 = n10836 | n10842 ;
  assign n10844 = ( n10827 & ~n10835 ) | ( n10827 & n10843 ) | ( ~n10835 & n10843 ) ;
  assign n10845 = n10835 | n10844 ;
  assign n10846 = n1790 | n4397 ;
  assign n10847 = n792 | n10846 ;
  assign n10848 = ( ~n3814 & n10845 ) | ( ~n3814 & n10847 ) | ( n10845 & n10847 ) ;
  assign n10849 = ( n3044 & n3194 ) | ( n3044 & ~n3814 ) | ( n3194 & ~n3814 ) ;
  assign n10850 = n3814 | n10849 ;
  assign n10851 = ( ~n10826 & n10848 ) | ( ~n10826 & n10850 ) | ( n10848 & n10850 ) ;
  assign n10852 = n10826 | n10851 ;
  assign n10853 = n607 & ~n9963 ;
  assign n10854 = n1250 & n9961 ;
  assign n10855 = n10853 | n10854 ;
  assign n10856 = n606 & ~n9959 ;
  assign n10857 = ( n606 & n10855 ) | ( n606 & ~n10856 ) | ( n10855 & ~n10856 ) ;
  assign n10858 = ( n9959 & ~n9961 ) | ( n9959 & n10025 ) | ( ~n9961 & n10025 ) ;
  assign n10859 = ( n9961 & ~n10026 ) | ( n9961 & n10858 ) | ( ~n10026 & n10858 ) ;
  assign n10860 = n1248 & n10859 ;
  assign n10861 = n10857 | n10860 ;
  assign n10862 = ( ~n10610 & n10852 ) | ( ~n10610 & n10861 ) | ( n10852 & n10861 ) ;
  assign n10863 = n607 & n9961 ;
  assign n10864 = n1250 & n9959 ;
  assign n10865 = n10863 | n10864 ;
  assign n10866 = n606 & n9957 ;
  assign n10867 = ( n606 & n10865 ) | ( n606 & ~n10866 ) | ( n10865 & ~n10866 ) ;
  assign n10868 = ( n9957 & ~n9959 ) | ( n9957 & n10026 ) | ( ~n9959 & n10026 ) ;
  assign n10869 = ( ~n10026 & n10027 ) | ( ~n10026 & n10868 ) | ( n10027 & n10868 ) ;
  assign n10870 = n1248 & ~n10869 ;
  assign n10871 = n10867 | n10870 ;
  assign n10872 = ( n10640 & n10862 ) | ( n10640 & n10871 ) | ( n10862 & n10871 ) ;
  assign n10873 = ( n10595 & n10642 ) | ( n10595 & ~n10741 ) | ( n10642 & ~n10741 ) ;
  assign n10874 = n3800 & n10557 ;
  assign n10875 = n3799 & n9949 ;
  assign n10876 = n3700 & ~n9953 ;
  assign n10877 = n3802 & n9951 ;
  assign n10878 = n10876 | n10877 ;
  assign n10879 = ( ~n10874 & n10875 ) | ( ~n10874 & n10878 ) | ( n10875 & n10878 ) ;
  assign n10880 = ( ~x29 & n10874 ) | ( ~x29 & n10879 ) | ( n10874 & n10879 ) ;
  assign n10881 = ( n10874 & n10879 ) | ( n10874 & ~n10880 ) | ( n10879 & ~n10880 ) ;
  assign n10882 = ( x29 & n10880 ) | ( x29 & ~n10881 ) | ( n10880 & ~n10881 ) ;
  assign n10883 = ( n10872 & n10873 ) | ( n10872 & n10882 ) | ( n10873 & n10882 ) ;
  assign n10884 = ( n10752 & n10761 ) | ( n10752 & ~n10762 ) | ( n10761 & ~n10762 ) ;
  assign n10885 = ( n10743 & n10762 ) | ( n10743 & ~n10884 ) | ( n10762 & ~n10884 ) ;
  assign n10886 = n4202 & ~n10390 ;
  assign n10887 = n4201 & ~n9941 ;
  assign n10888 = n4200 & n9945 ;
  assign n10889 = n4345 & n9943 ;
  assign n10890 = n10888 | n10889 ;
  assign n10891 = ( ~n10886 & n10887 ) | ( ~n10886 & n10890 ) | ( n10887 & n10890 ) ;
  assign n10892 = ( ~x26 & n10886 ) | ( ~x26 & n10891 ) | ( n10886 & n10891 ) ;
  assign n10893 = ( n10886 & n10891 ) | ( n10886 & ~n10892 ) | ( n10891 & ~n10892 ) ;
  assign n10894 = ( x26 & n10892 ) | ( x26 & ~n10893 ) | ( n10892 & ~n10893 ) ;
  assign n10895 = ( n10883 & ~n10885 ) | ( n10883 & n10894 ) | ( ~n10885 & n10894 ) ;
  assign n10896 = n4202 & n10284 ;
  assign n10897 = n4201 & ~n9883 ;
  assign n10898 = n4200 & n9943 ;
  assign n10899 = n4345 & ~n9941 ;
  assign n10900 = n10898 | n10899 ;
  assign n10901 = ( ~n10896 & n10897 ) | ( ~n10896 & n10900 ) | ( n10897 & n10900 ) ;
  assign n10902 = ( ~x26 & n10896 ) | ( ~x26 & n10901 ) | ( n10896 & n10901 ) ;
  assign n10903 = ( n10896 & n10901 ) | ( n10896 & ~n10902 ) | ( n10901 & ~n10902 ) ;
  assign n10904 = ( x26 & n10902 ) | ( x26 & ~n10903 ) | ( n10902 & ~n10903 ) ;
  assign n10905 = ( ~n10762 & n10771 ) | ( ~n10762 & n10773 ) | ( n10771 & n10773 ) ;
  assign n10906 = ( n10762 & ~n10774 ) | ( n10762 & n10905 ) | ( ~n10774 & n10905 ) ;
  assign n10907 = ( n10895 & n10904 ) | ( n10895 & n10906 ) | ( n10904 & n10906 ) ;
  assign n10908 = ( n10774 & n10776 ) | ( n10774 & n10785 ) | ( n10776 & n10785 ) ;
  assign n10909 = ( n10776 & n10786 ) | ( n10776 & ~n10908 ) | ( n10786 & ~n10908 ) ;
  assign n10910 = n4713 & ~n10305 ;
  assign n10911 = n4712 & ~n10302 ;
  assign n10912 = n4709 & ~n9937 ;
  assign n10913 = n4792 & ~n10057 ;
  assign n10914 = n10912 | n10913 ;
  assign n10915 = ( ~n10910 & n10911 ) | ( ~n10910 & n10914 ) | ( n10911 & n10914 ) ;
  assign n10916 = ( ~x23 & n10910 ) | ( ~x23 & n10915 ) | ( n10910 & n10915 ) ;
  assign n10917 = ( n10910 & n10915 ) | ( n10910 & ~n10916 ) | ( n10915 & ~n10916 ) ;
  assign n10918 = ( x23 & n10916 ) | ( x23 & ~n10917 ) | ( n10916 & ~n10917 ) ;
  assign n10919 = ( n10907 & ~n10909 ) | ( n10907 & n10918 ) | ( ~n10909 & n10918 ) ;
  assign n10920 = ( n10786 & n10788 ) | ( n10786 & n10797 ) | ( n10788 & n10797 ) ;
  assign n10921 = ( n10788 & n10798 ) | ( n10788 & ~n10920 ) | ( n10798 & ~n10920 ) ;
  assign n10922 = ( n10242 & n10919 ) | ( n10242 & ~n10921 ) | ( n10919 & ~n10921 ) ;
  assign n10923 = n607 & n9965 ;
  assign n10924 = n1250 & ~n9963 ;
  assign n10925 = n10923 | n10924 ;
  assign n10926 = n606 & ~n9961 ;
  assign n10927 = ( n606 & n10925 ) | ( n606 & ~n10926 ) | ( n10925 & ~n10926 ) ;
  assign n10928 = ( ~n9961 & n9963 ) | ( ~n9961 & n10024 ) | ( n9963 & n10024 ) ;
  assign n10929 = ( ~n10024 & n10025 ) | ( ~n10024 & n10928 ) | ( n10025 & n10928 ) ;
  assign n10930 = n1248 & ~n10929 ;
  assign n10931 = n10927 | n10930 ;
  assign n10932 = n253 | n433 ;
  assign n10933 = n685 | n10932 ;
  assign n10934 = n1235 | n4509 ;
  assign n10935 = ( n4420 & ~n10933 ) | ( n4420 & n10934 ) | ( ~n10933 & n10934 ) ;
  assign n10936 = n10933 | n10935 ;
  assign n10937 = n176 | n947 ;
  assign n10938 = ( ~n653 & n1902 ) | ( ~n653 & n5049 ) | ( n1902 & n5049 ) ;
  assign n10939 = ( n653 & ~n10937 ) | ( n653 & n10938 ) | ( ~n10937 & n10938 ) ;
  assign n10940 = n10937 | n10939 ;
  assign n10941 = n362 | n1460 ;
  assign n10942 = n701 | n10941 ;
  assign n10943 = n241 | n576 ;
  assign n10944 = ( n150 & n1169 ) | ( n150 & ~n10943 ) | ( n1169 & ~n10943 ) ;
  assign n10945 = n10943 | n10944 ;
  assign n10946 = ( n2935 & n10942 ) | ( n2935 & ~n10945 ) | ( n10942 & ~n10945 ) ;
  assign n10947 = n120 | n529 ;
  assign n10948 = ( n54 & n78 ) | ( n54 & ~n80 ) | ( n78 & ~n80 ) ;
  assign n10949 = ( n2347 & n10947 ) | ( n2347 & n10948 ) | ( n10947 & n10948 ) ;
  assign n10950 = n1220 | n2576 ;
  assign n10951 = ( n48 & n72 ) | ( n48 & n98 ) | ( n72 & n98 ) ;
  assign n10952 = ( ~n3127 & n10950 ) | ( ~n3127 & n10951 ) | ( n10950 & n10951 ) ;
  assign n10953 = n3127 | n10952 ;
  assign n10954 = ( n10948 & n10949 ) | ( n10948 & ~n10953 ) | ( n10949 & ~n10953 ) ;
  assign n10955 = ~n10949 & n10954 ;
  assign n10956 = ( ~n10945 & n10946 ) | ( ~n10945 & n10955 ) | ( n10946 & n10955 ) ;
  assign n10957 = ~n10946 & n10956 ;
  assign n10958 = ( n10936 & ~n10940 ) | ( n10936 & n10957 ) | ( ~n10940 & n10957 ) ;
  assign n10959 = ~n10936 & n10958 ;
  assign n10960 = ( n1017 & n5701 ) | ( n1017 & n10959 ) | ( n5701 & n10959 ) ;
  assign n10961 = n10959 & ~n10960 ;
  assign n10962 = n1707 | n2245 ;
  assign n10963 = n1509 | n4510 ;
  assign n10964 = n692 | n2067 ;
  assign n10965 = n167 | n536 ;
  assign n10966 = n952 | n2215 ;
  assign n10967 = ( n262 & n525 ) | ( n262 & ~n10966 ) | ( n525 & ~n10966 ) ;
  assign n10968 = n10966 | n10967 ;
  assign n10969 = ( ~n10964 & n10965 ) | ( ~n10964 & n10968 ) | ( n10965 & n10968 ) ;
  assign n10970 = n10964 | n10969 ;
  assign n10971 = ( n3184 & ~n10963 ) | ( n3184 & n10970 ) | ( ~n10963 & n10970 ) ;
  assign n10972 = n10963 | n10971 ;
  assign n10973 = n295 | n447 ;
  assign n10974 = ( ~n764 & n2182 ) | ( ~n764 & n3128 ) | ( n2182 & n3128 ) ;
  assign n10975 = ( n764 & ~n10973 ) | ( n764 & n10974 ) | ( ~n10973 & n10974 ) ;
  assign n10976 = n10973 | n10975 ;
  assign n10977 = ( n250 & n10972 ) | ( n250 & ~n10976 ) | ( n10972 & ~n10976 ) ;
  assign n10978 = ~n10972 & n10977 ;
  assign n10979 = ( ~n5575 & n10962 ) | ( ~n5575 & n10978 ) | ( n10962 & n10978 ) ;
  assign n10980 = ~n10962 & n10979 ;
  assign n10981 = n10961 | n10980 ;
  assign n10982 = ( n10961 & n10980 ) | ( n10961 & ~n10981 ) | ( n10980 & ~n10981 ) ;
  assign n10983 = n10981 & ~n10982 ;
  assign n10984 = n6587 | n7022 ;
  assign n10985 = n6583 | n10984 ;
  assign n10986 = n6584 | n10985 ;
  assign n10987 = ( ~x11 & n10983 ) | ( ~x11 & n10986 ) | ( n10983 & n10986 ) ;
  assign n10988 = ( n10983 & n10986 ) | ( n10983 & ~n10987 ) | ( n10986 & ~n10987 ) ;
  assign n10989 = ( x11 & n10987 ) | ( x11 & ~n10988 ) | ( n10987 & ~n10988 ) ;
  assign n10990 = ( n10961 & n10980 ) | ( n10961 & ~n10989 ) | ( n10980 & ~n10989 ) ;
  assign n10991 = ( n10610 & ~n10931 ) | ( n10610 & n10990 ) | ( ~n10931 & n10990 ) ;
  assign n10992 = n607 & n9971 ;
  assign n10993 = n1250 & n9969 ;
  assign n10994 = n10992 | n10993 ;
  assign n10995 = n606 & n9967 ;
  assign n10996 = ( n606 & n10994 ) | ( n606 & ~n10995 ) | ( n10994 & ~n10995 ) ;
  assign n10997 = ( n9967 & ~n9969 ) | ( n9967 & n10021 ) | ( ~n9969 & n10021 ) ;
  assign n10998 = ( ~n10021 & n10022 ) | ( ~n10021 & n10997 ) | ( n10022 & n10997 ) ;
  assign n10999 = n1248 & ~n10998 ;
  assign n11000 = n10996 | n10999 ;
  assign n11001 = n101 | n1595 ;
  assign n11002 = n890 | n11001 ;
  assign n11003 = n320 | n1430 ;
  assign n11004 = ( n1512 & n2504 ) | ( n1512 & ~n11003 ) | ( n2504 & ~n11003 ) ;
  assign n11005 = ( n549 & n1313 ) | ( n549 & ~n11003 ) | ( n1313 & ~n11003 ) ;
  assign n11006 = n11003 | n11005 ;
  assign n11007 = ( ~n11002 & n11004 ) | ( ~n11002 & n11006 ) | ( n11004 & n11006 ) ;
  assign n11008 = n11002 | n11007 ;
  assign n11009 = n1578 | n11008 ;
  assign n11010 = n969 | n1463 ;
  assign n11011 = n590 | n1341 ;
  assign n11012 = n764 | n11011 ;
  assign n11013 = n172 | n384 ;
  assign n11014 = n1174 | n1626 ;
  assign n11015 = n2914 | n11014 ;
  assign n11016 = ( ~n11012 & n11013 ) | ( ~n11012 & n11015 ) | ( n11013 & n11015 ) ;
  assign n11017 = ( n4032 & ~n11012 ) | ( n4032 & n11016 ) | ( ~n11012 & n11016 ) ;
  assign n11018 = n11012 | n11017 ;
  assign n11019 = ( ~n11009 & n11010 ) | ( ~n11009 & n11018 ) | ( n11010 & n11018 ) ;
  assign n11020 = n11009 | n11019 ;
  assign n11021 = n3210 | n10118 ;
  assign n11022 = n1790 | n2982 ;
  assign n11023 = n164 | n294 ;
  assign n11024 = n795 | n11023 ;
  assign n11025 = n2308 | n4436 ;
  assign n11026 = ( n837 & n1751 ) | ( n837 & ~n2308 ) | ( n1751 & ~n2308 ) ;
  assign n11027 = ( ~n11024 & n11025 ) | ( ~n11024 & n11026 ) | ( n11025 & n11026 ) ;
  assign n11028 = n11024 | n11027 ;
  assign n11029 = ( n1131 & ~n11022 ) | ( n1131 & n11028 ) | ( ~n11022 & n11028 ) ;
  assign n11030 = n11022 | n11029 ;
  assign n11031 = ( ~n11020 & n11021 ) | ( ~n11020 & n11030 ) | ( n11021 & n11030 ) ;
  assign n11032 = n11020 | n11031 ;
  assign n11033 = ( n72 & n116 ) | ( n72 & n166 ) | ( n116 & n166 ) ;
  assign n11034 = ( n202 & n1096 ) | ( n202 & ~n11033 ) | ( n1096 & ~n11033 ) ;
  assign n11035 = n11033 | n11034 ;
  assign n11036 = n1881 | n5017 ;
  assign n11037 = n167 | n274 ;
  assign n11038 = n810 | n11037 ;
  assign n11039 = ( ~n11035 & n11036 ) | ( ~n11035 & n11038 ) | ( n11036 & n11038 ) ;
  assign n11040 = n11035 | n11039 ;
  assign n11041 = ( n64 & n145 ) | ( n64 & n719 ) | ( n145 & n719 ) ;
  assign n11042 = ( n433 & n1082 ) | ( n433 & ~n11041 ) | ( n1082 & ~n11041 ) ;
  assign n11043 = n11041 | n11042 ;
  assign n11044 = ( n1320 & n2576 ) | ( n1320 & ~n2663 ) | ( n2576 & ~n2663 ) ;
  assign n11045 = n2663 | n11044 ;
  assign n11046 = ( n2952 & n11043 ) | ( n2952 & ~n11045 ) | ( n11043 & ~n11045 ) ;
  assign n11047 = ~n11043 & n11046 ;
  assign n11048 = n2671 | n2829 ;
  assign n11049 = n757 | n866 ;
  assign n11050 = n225 | n299 ;
  assign n11051 = n888 | n11050 ;
  assign n11052 = ( n66 & n80 ) | ( n66 & n145 ) | ( n80 & n145 ) ;
  assign n11053 = n320 | n11052 ;
  assign n11054 = ( n317 & ~n11051 ) | ( n317 & n11053 ) | ( ~n11051 & n11053 ) ;
  assign n11055 = n11051 | n11054 ;
  assign n11056 = ( ~n11048 & n11049 ) | ( ~n11048 & n11055 ) | ( n11049 & n11055 ) ;
  assign n11057 = n11048 | n11056 ;
  assign n11058 = ( n11040 & n11047 ) | ( n11040 & ~n11057 ) | ( n11047 & ~n11057 ) ;
  assign n11059 = ~n11040 & n11058 ;
  assign n11060 = ( n940 & n2230 ) | ( n940 & n11059 ) | ( n2230 & n11059 ) ;
  assign n11061 = n11059 & ~n11060 ;
  assign n11062 = n11032 & ~n11061 ;
  assign n11063 = n11032 & n11061 ;
  assign n11064 = ( n11061 & n11062 ) | ( n11061 & ~n11063 ) | ( n11062 & ~n11063 ) ;
  assign n11065 = n7299 | n7879 ;
  assign n11066 = n7295 | n11065 ;
  assign n11067 = n7296 | n11066 ;
  assign n11068 = ( ~x8 & n11064 ) | ( ~x8 & n11067 ) | ( n11064 & n11067 ) ;
  assign n11069 = ( n11064 & n11067 ) | ( n11064 & ~n11068 ) | ( n11067 & ~n11068 ) ;
  assign n11070 = ( x8 & n11068 ) | ( x8 & ~n11069 ) | ( n11068 & ~n11069 ) ;
  assign n11071 = ( ~n11032 & n11061 ) | ( ~n11032 & n11070 ) | ( n11061 & n11070 ) ;
  assign n11072 = ( n10961 & n11000 ) | ( n10961 & ~n11071 ) | ( n11000 & ~n11071 ) ;
  assign n11073 = n446 | n1133 ;
  assign n11074 = n544 | n1870 ;
  assign n11075 = n10201 | n11074 ;
  assign n11076 = n5056 | n11075 ;
  assign n11077 = ( n4987 & ~n11073 ) | ( n4987 & n11076 ) | ( ~n11073 & n11076 ) ;
  assign n11078 = n11073 | n11077 ;
  assign n11079 = n353 | n1692 ;
  assign n11080 = n1306 | n11079 ;
  assign n11081 = n4638 | n11080 ;
  assign n11082 = n332 | n346 ;
  assign n11083 = n277 | n294 ;
  assign n11084 = ( n206 & n661 ) | ( n206 & ~n11083 ) | ( n661 & ~n11083 ) ;
  assign n11085 = n11083 | n11084 ;
  assign n11086 = ( n2619 & ~n10810 ) | ( n2619 & n11085 ) | ( ~n10810 & n11085 ) ;
  assign n11087 = ( n1378 & n10810 ) | ( n1378 & ~n11086 ) | ( n10810 & ~n11086 ) ;
  assign n11088 = n11086 | n11087 ;
  assign n11089 = ( ~n11080 & n11082 ) | ( ~n11080 & n11088 ) | ( n11082 & n11088 ) ;
  assign n11090 = ( ~n11078 & n11081 ) | ( ~n11078 & n11089 ) | ( n11081 & n11089 ) ;
  assign n11091 = n117 | n764 ;
  assign n11092 = ( n653 & n888 ) | ( n653 & ~n11091 ) | ( n888 & ~n11091 ) ;
  assign n11093 = n11091 | n11092 ;
  assign n11094 = ( n1163 & n1351 ) | ( n1163 & ~n11093 ) | ( n1351 & ~n11093 ) ;
  assign n11095 = n11093 | n11094 ;
  assign n11096 = n171 | n254 ;
  assign n11097 = ( n549 & n878 ) | ( n549 & ~n11096 ) | ( n878 & ~n11096 ) ;
  assign n11098 = n11096 | n11097 ;
  assign n11099 = ( ~n2409 & n2892 ) | ( ~n2409 & n11098 ) | ( n2892 & n11098 ) ;
  assign n11100 = ~n11098 & n11099 ;
  assign n11101 = n163 | n985 ;
  assign n11102 = ( n995 & n1838 ) | ( n995 & ~n11101 ) | ( n1838 & ~n11101 ) ;
  assign n11103 = n11101 | n11102 ;
  assign n11104 = n2412 | n2443 ;
  assign n11105 = n773 | n1494 ;
  assign n11106 = ( n1369 & ~n11104 ) | ( n1369 & n11105 ) | ( ~n11104 & n11105 ) ;
  assign n11107 = n11104 | n11106 ;
  assign n11108 = ( n3444 & ~n11103 ) | ( n3444 & n11107 ) | ( ~n11103 & n11107 ) ;
  assign n11109 = n11103 | n11108 ;
  assign n11110 = ( n11095 & n11100 ) | ( n11095 & ~n11109 ) | ( n11100 & ~n11109 ) ;
  assign n11111 = ~n11095 & n11110 ;
  assign n11112 = ( ~n11078 & n11090 ) | ( ~n11078 & n11111 ) | ( n11090 & n11111 ) ;
  assign n11113 = ~n11090 & n11112 ;
  assign n11114 = ( n10961 & n11072 ) | ( n10961 & ~n11113 ) | ( n11072 & ~n11113 ) ;
  assign n11115 = n607 & ~n9967 ;
  assign n11116 = n1250 & n9965 ;
  assign n11117 = n11115 | n11116 ;
  assign n11118 = n606 & n9963 ;
  assign n11119 = ( n606 & n11117 ) | ( n606 & ~n11118 ) | ( n11117 & ~n11118 ) ;
  assign n11120 = ( n9963 & ~n9965 ) | ( n9963 & n10023 ) | ( ~n9965 & n10023 ) ;
  assign n11121 = ( ~n10023 & n10024 ) | ( ~n10023 & n11120 ) | ( n10024 & n11120 ) ;
  assign n11122 = n1248 & ~n11121 ;
  assign n11123 = n11119 | n11122 ;
  assign n11124 = ( ~n10989 & n11114 ) | ( ~n10989 & n11123 ) | ( n11114 & n11123 ) ;
  assign n11125 = ( n10610 & n10931 ) | ( n10610 & n10990 ) | ( n10931 & n10990 ) ;
  assign n11126 = ( n10931 & n10991 ) | ( n10931 & ~n11125 ) | ( n10991 & ~n11125 ) ;
  assign n11127 = n3800 & ~n10567 ;
  assign n11128 = n3799 & n9955 ;
  assign n11129 = n3700 & n9959 ;
  assign n11130 = n3802 & ~n9957 ;
  assign n11131 = n11129 | n11130 ;
  assign n11132 = ( ~n11127 & n11128 ) | ( ~n11127 & n11131 ) | ( n11128 & n11131 ) ;
  assign n11133 = ( ~x29 & n11127 ) | ( ~x29 & n11132 ) | ( n11127 & n11132 ) ;
  assign n11134 = ( n11127 & n11132 ) | ( n11127 & ~n11133 ) | ( n11132 & ~n11133 ) ;
  assign n11135 = ( x29 & n11133 ) | ( x29 & ~n11134 ) | ( n11133 & ~n11134 ) ;
  assign n11136 = ( n11124 & n11126 ) | ( n11124 & n11135 ) | ( n11126 & n11135 ) ;
  assign n11137 = ( n10852 & n10861 ) | ( n10852 & ~n10862 ) | ( n10861 & ~n10862 ) ;
  assign n11138 = ( n10610 & n10862 ) | ( n10610 & ~n11137 ) | ( n10862 & ~n11137 ) ;
  assign n11139 = ( n10991 & ~n11136 ) | ( n10991 & n11138 ) | ( ~n11136 & n11138 ) ;
  assign n11140 = ( ~n10640 & n10862 ) | ( ~n10640 & n10871 ) | ( n10862 & n10871 ) ;
  assign n11141 = ( n10640 & ~n10872 ) | ( n10640 & n11140 ) | ( ~n10872 & n11140 ) ;
  assign n11142 = n3800 & ~n10652 ;
  assign n11143 = n3799 & n9951 ;
  assign n11144 = n3700 & n9955 ;
  assign n11145 = n3802 & ~n9953 ;
  assign n11146 = n11144 | n11145 ;
  assign n11147 = ( ~n11142 & n11143 ) | ( ~n11142 & n11146 ) | ( n11143 & n11146 ) ;
  assign n11148 = ( ~x29 & n11142 ) | ( ~x29 & n11147 ) | ( n11142 & n11147 ) ;
  assign n11149 = ( n11142 & n11147 ) | ( n11142 & ~n11148 ) | ( n11147 & ~n11148 ) ;
  assign n11150 = ( x29 & n11148 ) | ( x29 & ~n11149 ) | ( n11148 & ~n11149 ) ;
  assign n11151 = ( ~n11139 & n11141 ) | ( ~n11139 & n11150 ) | ( n11141 & n11150 ) ;
  assign n11152 = ( ~n10872 & n10873 ) | ( ~n10872 & n10882 ) | ( n10873 & n10882 ) ;
  assign n11153 = ( n10872 & ~n10883 ) | ( n10872 & n11152 ) | ( ~n10883 & n11152 ) ;
  assign n11154 = n4202 & n10271 ;
  assign n11155 = n4201 & n9943 ;
  assign n11156 = n4200 & n9947 ;
  assign n11157 = n4345 & n9945 ;
  assign n11158 = n11156 | n11157 ;
  assign n11159 = ( ~n11154 & n11155 ) | ( ~n11154 & n11158 ) | ( n11155 & n11158 ) ;
  assign n11160 = ( ~x26 & n11154 ) | ( ~x26 & n11159 ) | ( n11154 & n11159 ) ;
  assign n11161 = ( n11154 & n11159 ) | ( n11154 & ~n11160 ) | ( n11159 & ~n11160 ) ;
  assign n11162 = ( x26 & n11160 ) | ( x26 & ~n11161 ) | ( n11160 & ~n11161 ) ;
  assign n11163 = ( n11151 & n11153 ) | ( n11151 & n11162 ) | ( n11153 & n11162 ) ;
  assign n11164 = ( ~n10883 & n10885 ) | ( ~n10883 & n10894 ) | ( n10885 & n10894 ) ;
  assign n11165 = ( ~n10894 & n10895 ) | ( ~n10894 & n11164 ) | ( n10895 & n11164 ) ;
  assign n11166 = n4713 & n10040 ;
  assign n11167 = n4712 & ~n9937 ;
  assign n11168 = n4709 & ~n9883 ;
  assign n11169 = n4792 & n9916 ;
  assign n11170 = n11168 | n11169 ;
  assign n11171 = ( ~n11166 & n11167 ) | ( ~n11166 & n11170 ) | ( n11167 & n11170 ) ;
  assign n11172 = ( ~x23 & n11166 ) | ( ~x23 & n11171 ) | ( n11166 & n11171 ) ;
  assign n11173 = ( n11166 & n11171 ) | ( n11166 & ~n11172 ) | ( n11171 & ~n11172 ) ;
  assign n11174 = ( x23 & n11172 ) | ( x23 & ~n11173 ) | ( n11172 & ~n11173 ) ;
  assign n11175 = ( n11163 & ~n11165 ) | ( n11163 & n11174 ) | ( ~n11165 & n11174 ) ;
  assign n11176 = ( ~n10895 & n10904 ) | ( ~n10895 & n10906 ) | ( n10904 & n10906 ) ;
  assign n11177 = ( n10895 & ~n10907 ) | ( n10895 & n11176 ) | ( ~n10907 & n11176 ) ;
  assign n11178 = n4713 & ~n10064 ;
  assign n11179 = n4712 & ~n10057 ;
  assign n11180 = n4709 & n9916 ;
  assign n11181 = n4792 & ~n9937 ;
  assign n11182 = n11180 | n11181 ;
  assign n11183 = ( ~n11178 & n11179 ) | ( ~n11178 & n11182 ) | ( n11179 & n11182 ) ;
  assign n11184 = ( ~x23 & n11178 ) | ( ~x23 & n11183 ) | ( n11178 & n11183 ) ;
  assign n11185 = ( n11178 & n11183 ) | ( n11178 & ~n11184 ) | ( n11183 & ~n11184 ) ;
  assign n11186 = ( x23 & n11184 ) | ( x23 & ~n11185 ) | ( n11184 & ~n11185 ) ;
  assign n11187 = ( n11175 & n11177 ) | ( n11175 & n11186 ) | ( n11177 & n11186 ) ;
  assign n11188 = ( ~n10907 & n10909 ) | ( ~n10907 & n10918 ) | ( n10909 & n10918 ) ;
  assign n11189 = ( ~n10918 & n10919 ) | ( ~n10918 & n11188 ) | ( n10919 & n11188 ) ;
  assign n11190 = n4972 | n5398 ;
  assign n11191 = ~n4973 & n10346 ;
  assign n11192 = ( n10346 & n11190 ) | ( n10346 & ~n11191 ) | ( n11190 & ~n11191 ) ;
  assign n11193 = ( ~x20 & n4974 ) | ( ~x20 & n11192 ) | ( n4974 & n11192 ) ;
  assign n11194 = ( n4974 & n11192 ) | ( n4974 & ~n11193 ) | ( n11192 & ~n11193 ) ;
  assign n11195 = ( x20 & n11193 ) | ( x20 & ~n11194 ) | ( n11193 & ~n11194 ) ;
  assign n11196 = ( n11187 & ~n11189 ) | ( n11187 & n11195 ) | ( ~n11189 & n11195 ) ;
  assign n11197 = ( ~n10991 & n11136 ) | ( ~n10991 & n11138 ) | ( n11136 & n11138 ) ;
  assign n11198 = ( ~n11138 & n11139 ) | ( ~n11138 & n11197 ) | ( n11139 & n11197 ) ;
  assign n11199 = n3800 & ~n10750 ;
  assign n11200 = n3799 & ~n9953 ;
  assign n11201 = n3700 & ~n9957 ;
  assign n11202 = n3802 & n9955 ;
  assign n11203 = n11201 | n11202 ;
  assign n11204 = ( ~n11199 & n11200 ) | ( ~n11199 & n11203 ) | ( n11200 & n11203 ) ;
  assign n11205 = ( ~x29 & n11199 ) | ( ~x29 & n11204 ) | ( n11199 & n11204 ) ;
  assign n11206 = ( n11199 & n11204 ) | ( n11199 & ~n11205 ) | ( n11204 & ~n11205 ) ;
  assign n11207 = ( x29 & n11205 ) | ( x29 & ~n11206 ) | ( n11205 & ~n11206 ) ;
  assign n11208 = n4202 & n10454 ;
  assign n11209 = n4201 & n9947 ;
  assign n11210 = n4200 & n9951 ;
  assign n11211 = n4345 & n9949 ;
  assign n11212 = n11210 | n11211 ;
  assign n11213 = ( ~n11208 & n11209 ) | ( ~n11208 & n11212 ) | ( n11209 & n11212 ) ;
  assign n11214 = ( ~x26 & n11208 ) | ( ~x26 & n11213 ) | ( n11208 & n11213 ) ;
  assign n11215 = ( n11208 & n11213 ) | ( n11208 & ~n11214 ) | ( n11213 & ~n11214 ) ;
  assign n11216 = ( x26 & n11214 ) | ( x26 & ~n11215 ) | ( n11214 & ~n11215 ) ;
  assign n11217 = ( n11198 & n11207 ) | ( n11198 & n11216 ) | ( n11207 & n11216 ) ;
  assign n11218 = ( n11141 & n11150 ) | ( n11141 & ~n11151 ) | ( n11150 & ~n11151 ) ;
  assign n11219 = ( n11139 & n11151 ) | ( n11139 & ~n11218 ) | ( n11151 & ~n11218 ) ;
  assign n11220 = n4202 & n10466 ;
  assign n11221 = n4201 & n9945 ;
  assign n11222 = n4200 & n9949 ;
  assign n11223 = n4345 & n9947 ;
  assign n11224 = n11222 | n11223 ;
  assign n11225 = ( ~n11220 & n11221 ) | ( ~n11220 & n11224 ) | ( n11221 & n11224 ) ;
  assign n11226 = ( ~x26 & n11220 ) | ( ~x26 & n11225 ) | ( n11220 & n11225 ) ;
  assign n11227 = ( n11220 & n11225 ) | ( n11220 & ~n11226 ) | ( n11225 & ~n11226 ) ;
  assign n11228 = ( x26 & n11226 ) | ( x26 & ~n11227 ) | ( n11226 & ~n11227 ) ;
  assign n11229 = ( n11217 & ~n11219 ) | ( n11217 & n11228 ) | ( ~n11219 & n11228 ) ;
  assign n11230 = ( n11151 & ~n11153 ) | ( n11151 & n11162 ) | ( ~n11153 & n11162 ) ;
  assign n11231 = ( n11153 & ~n11163 ) | ( n11153 & n11230 ) | ( ~n11163 & n11230 ) ;
  assign n11232 = n4713 & n10174 ;
  assign n11233 = n4712 & n9916 ;
  assign n11234 = n4792 | n9883 ;
  assign n11235 = n4709 & ~n9941 ;
  assign n11236 = ( ~n9883 & n11234 ) | ( ~n9883 & n11235 ) | ( n11234 & n11235 ) ;
  assign n11237 = ( ~n11232 & n11233 ) | ( ~n11232 & n11236 ) | ( n11233 & n11236 ) ;
  assign n11238 = ( ~x23 & n11232 ) | ( ~x23 & n11237 ) | ( n11232 & n11237 ) ;
  assign n11239 = ( n11232 & n11237 ) | ( n11232 & ~n11238 ) | ( n11237 & ~n11238 ) ;
  assign n11240 = ( x23 & n11238 ) | ( x23 & ~n11239 ) | ( n11238 & ~n11239 ) ;
  assign n11241 = ( n11229 & n11231 ) | ( n11229 & n11240 ) | ( n11231 & n11240 ) ;
  assign n11242 = ( ~n11163 & n11165 ) | ( ~n11163 & n11174 ) | ( n11165 & n11174 ) ;
  assign n11243 = ( ~n11174 & n11175 ) | ( ~n11174 & n11242 ) | ( n11175 & n11242 ) ;
  assign n11244 = n4974 & n10362 ;
  assign n11245 = n5398 & n10346 ;
  assign n11246 = n4973 & ~n10057 ;
  assign n11247 = n4972 & ~n10302 ;
  assign n11248 = n11246 | n11247 ;
  assign n11249 = ( ~n11244 & n11245 ) | ( ~n11244 & n11248 ) | ( n11245 & n11248 ) ;
  assign n11250 = ( ~x20 & n11244 ) | ( ~x20 & n11249 ) | ( n11244 & n11249 ) ;
  assign n11251 = ( n11244 & n11249 ) | ( n11244 & ~n11250 ) | ( n11249 & ~n11250 ) ;
  assign n11252 = ( x20 & n11250 ) | ( x20 & ~n11251 ) | ( n11250 & ~n11251 ) ;
  assign n11253 = ( n11241 & ~n11243 ) | ( n11241 & n11252 ) | ( ~n11243 & n11252 ) ;
  assign n11254 = n4974 & n10348 ;
  assign n11255 = n4972 & n10346 ;
  assign n11256 = n4973 & ~n10302 ;
  assign n11257 = n5398 | n11256 ;
  assign n11258 = ( ~n11254 & n11255 ) | ( ~n11254 & n11257 ) | ( n11255 & n11257 ) ;
  assign n11259 = ( ~x20 & n11254 ) | ( ~x20 & n11258 ) | ( n11254 & n11258 ) ;
  assign n11260 = ( n11254 & n11258 ) | ( n11254 & ~n11259 ) | ( n11258 & ~n11259 ) ;
  assign n11261 = ( x20 & n11259 ) | ( x20 & ~n11260 ) | ( n11259 & ~n11260 ) ;
  assign n11262 = ( ~n11175 & n11177 ) | ( ~n11175 & n11186 ) | ( n11177 & n11186 ) ;
  assign n11263 = ( n11175 & ~n11187 ) | ( n11175 & n11262 ) | ( ~n11187 & n11262 ) ;
  assign n11264 = ( n11253 & n11261 ) | ( n11253 & n11263 ) | ( n11261 & n11263 ) ;
  assign n11265 = ( ~n10961 & n11072 ) | ( ~n10961 & n11113 ) | ( n11072 & n11113 ) ;
  assign n11266 = ( ~n11072 & n11114 ) | ( ~n11072 & n11265 ) | ( n11114 & n11265 ) ;
  assign n11267 = n607 & n9969 ;
  assign n11268 = n1250 & ~n9967 ;
  assign n11269 = n11267 | n11268 ;
  assign n11270 = n606 & ~n9965 ;
  assign n11271 = ( n606 & n11269 ) | ( n606 & ~n11270 ) | ( n11269 & ~n11270 ) ;
  assign n11272 = ( ~n9965 & n9967 ) | ( ~n9965 & n10022 ) | ( n9967 & n10022 ) ;
  assign n11273 = ( ~n10022 & n10023 ) | ( ~n10022 & n11272 ) | ( n10023 & n11272 ) ;
  assign n11274 = n1248 & ~n11273 ;
  assign n11275 = n11271 | n11274 ;
  assign n11276 = n3800 & n10859 ;
  assign n11277 = n3799 & n9959 ;
  assign n11278 = n3700 & ~n9963 ;
  assign n11279 = n3802 & n9961 ;
  assign n11280 = n11278 | n11279 ;
  assign n11281 = ( ~n11276 & n11277 ) | ( ~n11276 & n11280 ) | ( n11277 & n11280 ) ;
  assign n11282 = ( ~x29 & n11276 ) | ( ~x29 & n11281 ) | ( n11276 & n11281 ) ;
  assign n11283 = ( n11276 & n11281 ) | ( n11276 & ~n11282 ) | ( n11281 & ~n11282 ) ;
  assign n11284 = ( x29 & n11282 ) | ( x29 & ~n11283 ) | ( n11282 & ~n11283 ) ;
  assign n11285 = ( ~n11266 & n11275 ) | ( ~n11266 & n11284 ) | ( n11275 & n11284 ) ;
  assign n11286 = ( n10989 & ~n11114 ) | ( n10989 & n11123 ) | ( ~n11114 & n11123 ) ;
  assign n11287 = ( ~n11123 & n11124 ) | ( ~n11123 & n11286 ) | ( n11124 & n11286 ) ;
  assign n11288 = n3800 & ~n10869 ;
  assign n11289 = n3799 & ~n9957 ;
  assign n11290 = n3700 & n9961 ;
  assign n11291 = n3802 & n9959 ;
  assign n11292 = n11290 | n11291 ;
  assign n11293 = ( ~n11288 & n11289 ) | ( ~n11288 & n11292 ) | ( n11289 & n11292 ) ;
  assign n11294 = ( ~x29 & n11288 ) | ( ~x29 & n11293 ) | ( n11288 & n11293 ) ;
  assign n11295 = ( n11288 & n11293 ) | ( n11288 & ~n11294 ) | ( n11293 & ~n11294 ) ;
  assign n11296 = ( x29 & n11294 ) | ( x29 & ~n11295 ) | ( n11294 & ~n11295 ) ;
  assign n11297 = ( n11285 & ~n11287 ) | ( n11285 & n11296 ) | ( ~n11287 & n11296 ) ;
  assign n11298 = ( n11124 & ~n11126 ) | ( n11124 & n11135 ) | ( ~n11126 & n11135 ) ;
  assign n11299 = ( n11126 & ~n11136 ) | ( n11126 & n11298 ) | ( ~n11136 & n11298 ) ;
  assign n11300 = n4202 & n10557 ;
  assign n11301 = n4201 & n9949 ;
  assign n11302 = n4200 & ~n9953 ;
  assign n11303 = n4345 & n9951 ;
  assign n11304 = n11302 | n11303 ;
  assign n11305 = ( ~n11300 & n11301 ) | ( ~n11300 & n11304 ) | ( n11301 & n11304 ) ;
  assign n11306 = ( ~x26 & n11300 ) | ( ~x26 & n11305 ) | ( n11300 & n11305 ) ;
  assign n11307 = ( n11300 & n11305 ) | ( n11300 & ~n11306 ) | ( n11305 & ~n11306 ) ;
  assign n11308 = ( x26 & n11306 ) | ( x26 & ~n11307 ) | ( n11306 & ~n11307 ) ;
  assign n11309 = ( n11297 & n11299 ) | ( n11297 & n11308 ) | ( n11299 & n11308 ) ;
  assign n11310 = ( n11198 & ~n11207 ) | ( n11198 & n11216 ) | ( ~n11207 & n11216 ) ;
  assign n11311 = ( n11207 & ~n11217 ) | ( n11207 & n11310 ) | ( ~n11217 & n11310 ) ;
  assign n11312 = n4713 & ~n10390 ;
  assign n11313 = n4712 & ~n9941 ;
  assign n11314 = n4709 & n9945 ;
  assign n11315 = n4792 & n9943 ;
  assign n11316 = n11314 | n11315 ;
  assign n11317 = ( ~n11312 & n11313 ) | ( ~n11312 & n11316 ) | ( n11313 & n11316 ) ;
  assign n11318 = ( ~x23 & n11312 ) | ( ~x23 & n11317 ) | ( n11312 & n11317 ) ;
  assign n11319 = ( n11312 & n11317 ) | ( n11312 & ~n11318 ) | ( n11317 & ~n11318 ) ;
  assign n11320 = ( x23 & n11318 ) | ( x23 & ~n11319 ) | ( n11318 & ~n11319 ) ;
  assign n11321 = ( n11309 & n11311 ) | ( n11309 & n11320 ) | ( n11311 & n11320 ) ;
  assign n11322 = ( ~n11217 & n11219 ) | ( ~n11217 & n11228 ) | ( n11219 & n11228 ) ;
  assign n11323 = ( ~n11228 & n11229 ) | ( ~n11228 & n11322 ) | ( n11229 & n11322 ) ;
  assign n11324 = n4713 & n10284 ;
  assign n11325 = n4712 & ~n9883 ;
  assign n11326 = n4709 & n9943 ;
  assign n11327 = n4792 & ~n9941 ;
  assign n11328 = n11326 | n11327 ;
  assign n11329 = ( ~n11324 & n11325 ) | ( ~n11324 & n11328 ) | ( n11325 & n11328 ) ;
  assign n11330 = ( ~x23 & n11324 ) | ( ~x23 & n11329 ) | ( n11324 & n11329 ) ;
  assign n11331 = ( n11324 & n11329 ) | ( n11324 & ~n11330 ) | ( n11329 & ~n11330 ) ;
  assign n11332 = ( x23 & n11330 ) | ( x23 & ~n11331 ) | ( n11330 & ~n11331 ) ;
  assign n11333 = ( n11321 & ~n11323 ) | ( n11321 & n11332 ) | ( ~n11323 & n11332 ) ;
  assign n11334 = ( n11229 & ~n11231 ) | ( n11229 & n11240 ) | ( ~n11231 & n11240 ) ;
  assign n11335 = ( n11231 & ~n11241 ) | ( n11231 & n11334 ) | ( ~n11241 & n11334 ) ;
  assign n11336 = n4974 & ~n10305 ;
  assign n11337 = n5398 & ~n10302 ;
  assign n11338 = n4973 & ~n9937 ;
  assign n11339 = n4972 & ~n10057 ;
  assign n11340 = n11338 | n11339 ;
  assign n11341 = ( ~n11336 & n11337 ) | ( ~n11336 & n11340 ) | ( n11337 & n11340 ) ;
  assign n11342 = ( ~x20 & n11336 ) | ( ~x20 & n11341 ) | ( n11336 & n11341 ) ;
  assign n11343 = ( n11336 & n11341 ) | ( n11336 & ~n11342 ) | ( n11341 & ~n11342 ) ;
  assign n11344 = ( x20 & n11342 ) | ( x20 & ~n11343 ) | ( n11342 & ~n11343 ) ;
  assign n11345 = ( n11333 & n11335 ) | ( n11333 & n11344 ) | ( n11335 & n11344 ) ;
  assign n11346 = ( ~n11241 & n11243 ) | ( ~n11241 & n11252 ) | ( n11243 & n11252 ) ;
  assign n11347 = ( ~n11252 & n11253 ) | ( ~n11252 & n11346 ) | ( n11253 & n11346 ) ;
  assign n11348 = n5499 & ~n10530 ;
  assign n11349 = ( ~x17 & n10531 ) | ( ~x17 & n11348 ) | ( n10531 & n11348 ) ;
  assign n11350 = ( n11345 & ~n11347 ) | ( n11345 & n11349 ) | ( ~n11347 & n11349 ) ;
  assign n11351 = ( x0 & ~x2 ) | ( x0 & n9378 ) | ( ~x2 & n9378 ) ;
  assign n11352 = ~n3878 & n10955 ;
  assign n11353 = n238 | n2798 ;
  assign n11354 = ( n1680 & n3733 ) | ( n1680 & ~n11353 ) | ( n3733 & ~n11353 ) ;
  assign n11355 = n11353 | n11354 ;
  assign n11356 = n3397 | n4106 ;
  assign n11357 = n1728 | n3105 ;
  assign n11358 = n10626 | n11357 ;
  assign n11359 = n2207 | n2680 ;
  assign n11360 = n945 | n11359 ;
  assign n11361 = n789 | n1593 ;
  assign n11362 = n115 | n290 ;
  assign n11363 = ( n613 & n1096 ) | ( n613 & ~n11362 ) | ( n1096 & ~n11362 ) ;
  assign n11364 = n11362 | n11363 ;
  assign n11365 = ( n262 & n505 ) | ( n262 & ~n775 ) | ( n505 & ~n775 ) ;
  assign n11366 = n775 | n11365 ;
  assign n11367 = ( ~n11361 & n11364 ) | ( ~n11361 & n11366 ) | ( n11364 & n11366 ) ;
  assign n11368 = n11361 | n11367 ;
  assign n11369 = ( n1355 & ~n11360 ) | ( n1355 & n11368 ) | ( ~n11360 & n11368 ) ;
  assign n11370 = n11360 | n11369 ;
  assign n11371 = ( ~n11356 & n11358 ) | ( ~n11356 & n11370 ) | ( n11358 & n11370 ) ;
  assign n11372 = n11356 | n11371 ;
  assign n11373 = n185 | n1005 ;
  assign n11374 = ( n1692 & n11098 ) | ( n1692 & ~n11373 ) | ( n11098 & ~n11373 ) ;
  assign n11375 = n11373 | n11374 ;
  assign n11376 = ( ~n11355 & n11372 ) | ( ~n11355 & n11375 ) | ( n11372 & n11375 ) ;
  assign n11377 = n11355 | n11376 ;
  assign n11378 = n745 | n1710 ;
  assign n11379 = ( n3404 & n3841 ) | ( n3404 & ~n11378 ) | ( n3841 & ~n11378 ) ;
  assign n11380 = n11378 | n11379 ;
  assign n11381 = n5678 | n6094 ;
  assign n11382 = n277 | n886 ;
  assign n11383 = ( n1312 & n4100 ) | ( n1312 & ~n11382 ) | ( n4100 & ~n11382 ) ;
  assign n11384 = n11382 | n11383 ;
  assign n11385 = ( ~n11380 & n11381 ) | ( ~n11380 & n11384 ) | ( n11381 & n11384 ) ;
  assign n11386 = n11380 | n11385 ;
  assign n11387 = ( n11352 & n11377 ) | ( n11352 & n11386 ) | ( n11377 & n11386 ) ;
  assign n11388 = n11352 & ~n11387 ;
  assign n11389 = n8225 | n8229 ;
  assign n11390 = x4 | n11389 ;
  assign n11391 = x4 & n8218 ;
  assign n11392 = ( ~x5 & n11390 ) | ( ~x5 & n11391 ) | ( n11390 & n11391 ) ;
  assign n11393 = ( n11351 & n11388 ) | ( n11351 & n11392 ) | ( n11388 & n11392 ) ;
  assign n11394 = n607 & n9977 ;
  assign n11395 = n1250 & n9975 ;
  assign n11396 = n11394 | n11395 ;
  assign n11397 = n606 & ~n9973 ;
  assign n11398 = ( n606 & n11396 ) | ( n606 & ~n11397 ) | ( n11396 & ~n11397 ) ;
  assign n11399 = ( n9973 & ~n9975 ) | ( n9973 & n10018 ) | ( ~n9975 & n10018 ) ;
  assign n11400 = ( n9975 & ~n10019 ) | ( n9975 & n11399 ) | ( ~n10019 & n11399 ) ;
  assign n11401 = n1248 & n11400 ;
  assign n11402 = n11398 | n11401 ;
  assign n11403 = ( n11032 & n11393 ) | ( n11032 & ~n11402 ) | ( n11393 & ~n11402 ) ;
  assign n11404 = n577 | n1694 ;
  assign n11405 = n2966 | n11404 ;
  assign n11406 = n1110 | n2181 ;
  assign n11407 = n519 | n11406 ;
  assign n11408 = n1413 | n11407 ;
  assign n11409 = n138 | n294 ;
  assign n11410 = ( n41 & ~n78 ) | ( n41 & n149 ) | ( ~n78 & n149 ) ;
  assign n11411 = n215 | n11410 ;
  assign n11412 = ( n1692 & ~n11409 ) | ( n1692 & n11411 ) | ( ~n11409 & n11411 ) ;
  assign n11413 = n11409 | n11412 ;
  assign n11414 = ( n1394 & ~n5099 ) | ( n1394 & n11413 ) | ( ~n5099 & n11413 ) ;
  assign n11415 = ( n5099 & n11051 ) | ( n5099 & ~n11414 ) | ( n11051 & ~n11414 ) ;
  assign n11416 = n11414 | n11415 ;
  assign n11417 = ( ~n11405 & n11408 ) | ( ~n11405 & n11416 ) | ( n11408 & n11416 ) ;
  assign n11418 = n11405 | n11417 ;
  assign n11419 = ( ~n2755 & n2907 ) | ( ~n2755 & n11418 ) | ( n2907 & n11418 ) ;
  assign n11420 = ~n11418 & n11419 ;
  assign n11421 = ( n11032 & n11403 ) | ( n11032 & n11420 ) | ( n11403 & n11420 ) ;
  assign n11422 = n607 & n9973 ;
  assign n11423 = n1250 & n9971 ;
  assign n11424 = n11422 | n11423 ;
  assign n11425 = n606 & ~n9969 ;
  assign n11426 = ( n606 & n11424 ) | ( n606 & ~n11425 ) | ( n11424 & ~n11425 ) ;
  assign n11427 = ( n9969 & ~n9971 ) | ( n9969 & n10020 ) | ( ~n9971 & n10020 ) ;
  assign n11428 = ( n9971 & ~n10021 ) | ( n9971 & n11427 ) | ( ~n10021 & n11427 ) ;
  assign n11429 = n1248 & n11428 ;
  assign n11430 = n11426 | n11429 ;
  assign n11431 = ( n11070 & ~n11421 ) | ( n11070 & n11430 ) | ( ~n11421 & n11430 ) ;
  assign n11432 = ( n10961 & n11000 ) | ( n10961 & ~n11072 ) | ( n11000 & ~n11072 ) ;
  assign n11433 = ( n11071 & n11072 ) | ( n11071 & ~n11432 ) | ( n11072 & ~n11432 ) ;
  assign n11434 = n3800 & ~n10929 ;
  assign n11435 = n3799 & n9961 ;
  assign n11436 = n3700 & n9965 ;
  assign n11437 = n3802 & ~n9963 ;
  assign n11438 = n11436 | n11437 ;
  assign n11439 = ( ~n11434 & n11435 ) | ( ~n11434 & n11438 ) | ( n11435 & n11438 ) ;
  assign n11440 = ( ~x29 & n11434 ) | ( ~x29 & n11439 ) | ( n11434 & n11439 ) ;
  assign n11441 = ( n11434 & n11439 ) | ( n11434 & ~n11440 ) | ( n11439 & ~n11440 ) ;
  assign n11442 = ( x29 & n11440 ) | ( x29 & ~n11441 ) | ( n11440 & ~n11441 ) ;
  assign n11443 = ( n11431 & ~n11433 ) | ( n11431 & n11442 ) | ( ~n11433 & n11442 ) ;
  assign n11444 = ( n11275 & n11284 ) | ( n11275 & ~n11285 ) | ( n11284 & ~n11285 ) ;
  assign n11445 = ( n11266 & n11285 ) | ( n11266 & ~n11444 ) | ( n11285 & ~n11444 ) ;
  assign n11446 = n4202 & ~n10750 ;
  assign n11447 = n4201 & ~n9953 ;
  assign n11448 = n4200 & ~n9957 ;
  assign n11449 = n4345 & n9955 ;
  assign n11450 = n11448 | n11449 ;
  assign n11451 = ( ~n11446 & n11447 ) | ( ~n11446 & n11450 ) | ( n11447 & n11450 ) ;
  assign n11452 = ( ~x26 & n11446 ) | ( ~x26 & n11451 ) | ( n11446 & n11451 ) ;
  assign n11453 = ( n11446 & n11451 ) | ( n11446 & ~n11452 ) | ( n11451 & ~n11452 ) ;
  assign n11454 = ( x26 & n11452 ) | ( x26 & ~n11453 ) | ( n11452 & ~n11453 ) ;
  assign n11455 = ( n11443 & ~n11445 ) | ( n11443 & n11454 ) | ( ~n11445 & n11454 ) ;
  assign n11456 = n4202 & ~n10652 ;
  assign n11457 = n4201 & n9951 ;
  assign n11458 = n4200 & n9955 ;
  assign n11459 = n4345 & ~n9953 ;
  assign n11460 = n11458 | n11459 ;
  assign n11461 = ( ~n11456 & n11457 ) | ( ~n11456 & n11460 ) | ( n11457 & n11460 ) ;
  assign n11462 = ( ~x26 & n11456 ) | ( ~x26 & n11461 ) | ( n11456 & n11461 ) ;
  assign n11463 = ( n11456 & n11461 ) | ( n11456 & ~n11462 ) | ( n11461 & ~n11462 ) ;
  assign n11464 = ( x26 & n11462 ) | ( x26 & ~n11463 ) | ( n11462 & ~n11463 ) ;
  assign n11465 = ( ~n11285 & n11287 ) | ( ~n11285 & n11296 ) | ( n11287 & n11296 ) ;
  assign n11466 = ( ~n11296 & n11297 ) | ( ~n11296 & n11465 ) | ( n11297 & n11465 ) ;
  assign n11467 = ( n11455 & n11464 ) | ( n11455 & ~n11466 ) | ( n11464 & ~n11466 ) ;
  assign n11468 = ( n11297 & ~n11299 ) | ( n11297 & n11308 ) | ( ~n11299 & n11308 ) ;
  assign n11469 = ( n11299 & ~n11309 ) | ( n11299 & n11468 ) | ( ~n11309 & n11468 ) ;
  assign n11470 = n4713 & n10271 ;
  assign n11471 = n4712 & n9943 ;
  assign n11472 = n4709 & n9947 ;
  assign n11473 = n4792 & n9945 ;
  assign n11474 = n11472 | n11473 ;
  assign n11475 = ( ~n11470 & n11471 ) | ( ~n11470 & n11474 ) | ( n11471 & n11474 ) ;
  assign n11476 = ( ~x23 & n11470 ) | ( ~x23 & n11475 ) | ( n11470 & n11475 ) ;
  assign n11477 = ( n11470 & n11475 ) | ( n11470 & ~n11476 ) | ( n11475 & ~n11476 ) ;
  assign n11478 = ( x23 & n11476 ) | ( x23 & ~n11477 ) | ( n11476 & ~n11477 ) ;
  assign n11479 = ( n11467 & n11469 ) | ( n11467 & n11478 ) | ( n11469 & n11478 ) ;
  assign n11480 = ( n11309 & ~n11311 ) | ( n11309 & n11320 ) | ( ~n11311 & n11320 ) ;
  assign n11481 = ( n11311 & ~n11321 ) | ( n11311 & n11480 ) | ( ~n11321 & n11480 ) ;
  assign n11482 = n4974 & n10040 ;
  assign n11483 = n5398 & ~n9937 ;
  assign n11484 = n4973 & ~n9883 ;
  assign n11485 = n4972 & n9916 ;
  assign n11486 = n11484 | n11485 ;
  assign n11487 = ( ~n11482 & n11483 ) | ( ~n11482 & n11486 ) | ( n11483 & n11486 ) ;
  assign n11488 = ( ~x20 & n11482 ) | ( ~x20 & n11487 ) | ( n11482 & n11487 ) ;
  assign n11489 = ( n11482 & n11487 ) | ( n11482 & ~n11488 ) | ( n11487 & ~n11488 ) ;
  assign n11490 = ( x20 & n11488 ) | ( x20 & ~n11489 ) | ( n11488 & ~n11489 ) ;
  assign n11491 = ( n11479 & n11481 ) | ( n11479 & n11490 ) | ( n11481 & n11490 ) ;
  assign n11492 = ( ~n11321 & n11323 ) | ( ~n11321 & n11332 ) | ( n11323 & n11332 ) ;
  assign n11493 = ( ~n11332 & n11333 ) | ( ~n11332 & n11492 ) | ( n11333 & n11492 ) ;
  assign n11494 = n4974 & ~n10064 ;
  assign n11495 = n5398 & ~n10057 ;
  assign n11496 = n4973 & n9916 ;
  assign n11497 = n4972 & ~n9937 ;
  assign n11498 = n11496 | n11497 ;
  assign n11499 = ( ~n11494 & n11495 ) | ( ~n11494 & n11498 ) | ( n11495 & n11498 ) ;
  assign n11500 = ( ~x20 & n11494 ) | ( ~x20 & n11499 ) | ( n11494 & n11499 ) ;
  assign n11501 = ( n11494 & n11499 ) | ( n11494 & ~n11500 ) | ( n11499 & ~n11500 ) ;
  assign n11502 = ( x20 & n11500 ) | ( x20 & ~n11501 ) | ( n11500 & ~n11501 ) ;
  assign n11503 = ( n11491 & ~n11493 ) | ( n11491 & n11502 ) | ( ~n11493 & n11502 ) ;
  assign n11504 = ( n11333 & ~n11335 ) | ( n11333 & n11344 ) | ( ~n11335 & n11344 ) ;
  assign n11505 = ( n11335 & ~n11345 ) | ( n11335 & n11504 ) | ( ~n11345 & n11504 ) ;
  assign n11506 = n5504 & ~n10346 ;
  assign n11507 = ( n5504 & n10530 ) | ( n5504 & ~n11506 ) | ( n10530 & ~n11506 ) ;
  assign n11508 = ( ~x17 & n5508 ) | ( ~x17 & n11507 ) | ( n5508 & n11507 ) ;
  assign n11509 = ( n5508 & n11507 ) | ( n5508 & ~n11508 ) | ( n11507 & ~n11508 ) ;
  assign n11510 = ( x17 & n11508 ) | ( x17 & ~n11509 ) | ( n11508 & ~n11509 ) ;
  assign n11511 = ( n11503 & n11505 ) | ( n11503 & n11510 ) | ( n11505 & n11510 ) ;
  assign n11512 = n262 | n2442 ;
  assign n11513 = n241 | n337 ;
  assign n11514 = ( n942 & n3131 ) | ( n942 & ~n5185 ) | ( n3131 & ~n5185 ) ;
  assign n11515 = n5185 | n11514 ;
  assign n11516 = ( n445 & ~n11513 ) | ( n445 & n11515 ) | ( ~n11513 & n11515 ) ;
  assign n11517 = n11513 | n11516 ;
  assign n11518 = ( ~n231 & n293 ) | ( ~n231 & n1032 ) | ( n293 & n1032 ) ;
  assign n11519 = n231 | n11518 ;
  assign n11520 = n567 | n1082 ;
  assign n11521 = n207 | n11520 ;
  assign n11522 = ( ~n718 & n11519 ) | ( ~n718 & n11521 ) | ( n11519 & n11521 ) ;
  assign n11523 = n718 | n11522 ;
  assign n11524 = ( n1732 & n2321 ) | ( n1732 & ~n3351 ) | ( n2321 & ~n3351 ) ;
  assign n11525 = n3351 | n11524 ;
  assign n11526 = ( n3885 & ~n11523 ) | ( n3885 & n11525 ) | ( ~n11523 & n11525 ) ;
  assign n11527 = n11523 | n11526 ;
  assign n11528 = ( n2723 & ~n11517 ) | ( n2723 & n11527 ) | ( ~n11517 & n11527 ) ;
  assign n11529 = n11517 | n11528 ;
  assign n11530 = ( n746 & n886 ) | ( n746 & ~n2671 ) | ( n886 & ~n2671 ) ;
  assign n11531 = n2671 | n11530 ;
  assign n11532 = ( ~n11512 & n11529 ) | ( ~n11512 & n11531 ) | ( n11529 & n11531 ) ;
  assign n11533 = n11512 | n11532 ;
  assign n11534 = ~n807 & n3568 ;
  assign n11535 = n514 | n719 ;
  assign n11536 = ( n2708 & n11534 ) | ( n2708 & n11535 ) | ( n11534 & n11535 ) ;
  assign n11537 = n11534 & ~n11536 ;
  assign n11538 = ( n10428 & ~n11533 ) | ( n10428 & n11537 ) | ( ~n11533 & n11537 ) ;
  assign n11539 = n361 | n1116 ;
  assign n11540 = ( n64 & n83 ) | ( n64 & n116 ) | ( n83 & n116 ) ;
  assign n11541 = n609 | n11540 ;
  assign n11542 = ( n6110 & n11539 ) | ( n6110 & ~n11541 ) | ( n11539 & ~n11541 ) ;
  assign n11543 = ( n199 & n11541 ) | ( n199 & ~n11542 ) | ( n11541 & ~n11542 ) ;
  assign n11544 = n11542 | n11543 ;
  assign n11545 = n132 | n233 ;
  assign n11546 = n1313 | n11545 ;
  assign n11547 = n751 | n11098 ;
  assign n11548 = ( n101 & n641 ) | ( n101 & ~n1792 ) | ( n641 & ~n1792 ) ;
  assign n11549 = n1792 | n11548 ;
  assign n11550 = ( ~n11546 & n11547 ) | ( ~n11546 & n11549 ) | ( n11547 & n11549 ) ;
  assign n11551 = n11546 | n11550 ;
  assign n11552 = ( n11537 & n11544 ) | ( n11537 & n11551 ) | ( n11544 & n11551 ) ;
  assign n11553 = ( n10428 & n11538 ) | ( n10428 & ~n11552 ) | ( n11538 & ~n11552 ) ;
  assign n11554 = ~n10428 & n11553 ;
  assign n11555 = n607 & n9985 ;
  assign n11556 = n1250 & ~n9983 ;
  assign n11557 = n11555 | n11556 ;
  assign n11558 = n606 & ~n9981 ;
  assign n11559 = ( n606 & n11557 ) | ( n606 & ~n11558 ) | ( n11557 & ~n11558 ) ;
  assign n11560 = ( ~n9981 & n9983 ) | ( ~n9981 & n10014 ) | ( n9983 & n10014 ) ;
  assign n11561 = ( ~n10014 & n10015 ) | ( ~n10014 & n11560 ) | ( n10015 & n11560 ) ;
  assign n11562 = n1248 & ~n11561 ;
  assign n11563 = n11559 | n11562 ;
  assign n11564 = ( n11351 & ~n11554 ) | ( n11351 & n11563 ) | ( ~n11554 & n11563 ) ;
  assign n11565 = n466 | n851 ;
  assign n11566 = n519 | n11565 ;
  assign n11567 = ( n913 & n2328 ) | ( n913 & ~n11566 ) | ( n2328 & ~n11566 ) ;
  assign n11568 = n11566 | n11567 ;
  assign n11569 = ( n314 & ~n1757 ) | ( n314 & n2870 ) | ( ~n1757 & n2870 ) ;
  assign n11570 = n1757 | n11569 ;
  assign n11571 = ( n729 & ~n11568 ) | ( n729 & n11570 ) | ( ~n11568 & n11570 ) ;
  assign n11572 = n11568 | n11571 ;
  assign n11573 = n4397 | n10181 ;
  assign n11574 = n2636 | n2846 ;
  assign n11575 = ( n10254 & ~n11573 ) | ( n10254 & n11574 ) | ( ~n11573 & n11574 ) ;
  assign n11576 = n11573 | n11575 ;
  assign n11577 = ( ~n11377 & n11572 ) | ( ~n11377 & n11576 ) | ( n11572 & n11576 ) ;
  assign n11578 = n455 | n1589 ;
  assign n11579 = n10120 | n11578 ;
  assign n11580 = ( n11377 & ~n11577 ) | ( n11377 & n11579 ) | ( ~n11577 & n11579 ) ;
  assign n11581 = n11577 | n11580 ;
  assign n11582 = ( n11351 & n11564 ) | ( n11351 & n11581 ) | ( n11564 & n11581 ) ;
  assign n11583 = n627 | n835 ;
  assign n11584 = n1626 | n2827 ;
  assign n11585 = n2967 & ~n3168 ;
  assign n11586 = ( n4418 & n10613 ) | ( n4418 & n11585 ) | ( n10613 & n11585 ) ;
  assign n11587 = n11585 & ~n11586 ;
  assign n11588 = n120 | n641 ;
  assign n11589 = ( n447 & n586 ) | ( n447 & ~n11588 ) | ( n586 & ~n11588 ) ;
  assign n11590 = n11588 | n11589 ;
  assign n11591 = ( n11584 & n11587 ) | ( n11584 & ~n11590 ) | ( n11587 & ~n11590 ) ;
  assign n11592 = ~n11584 & n11591 ;
  assign n11593 = ( n627 & ~n3554 ) | ( n627 & n11592 ) | ( ~n3554 & n11592 ) ;
  assign n11594 = ( n532 & n11583 ) | ( n532 & n11593 ) | ( n11583 & n11593 ) ;
  assign n11595 = ( ~n3869 & n11593 ) | ( ~n3869 & n11594 ) | ( n11593 & n11594 ) ;
  assign n11596 = ~n11594 & n11595 ;
  assign n11597 = ( n11351 & n11582 ) | ( n11351 & ~n11596 ) | ( n11582 & ~n11596 ) ;
  assign n11598 = ( n11351 & ~n11388 ) | ( n11351 & n11392 ) | ( ~n11388 & n11392 ) ;
  assign n11599 = ( n11388 & ~n11393 ) | ( n11388 & n11598 ) | ( ~n11393 & n11598 ) ;
  assign n11600 = n607 & n9979 ;
  assign n11601 = n1250 & n9977 ;
  assign n11602 = n11600 | n11601 ;
  assign n11603 = n606 & ~n9975 ;
  assign n11604 = ( n606 & n11602 ) | ( n606 & ~n11603 ) | ( n11602 & ~n11603 ) ;
  assign n11605 = ( n9975 & ~n9977 ) | ( n9975 & n10017 ) | ( ~n9977 & n10017 ) ;
  assign n11606 = ( n9977 & ~n10018 ) | ( n9977 & n11605 ) | ( ~n10018 & n11605 ) ;
  assign n11607 = n1248 & n11606 ;
  assign n11608 = n11604 | n11607 ;
  assign n11609 = ( n11597 & ~n11599 ) | ( n11597 & n11608 ) | ( ~n11599 & n11608 ) ;
  assign n11610 = ( ~n11032 & n11393 ) | ( ~n11032 & n11402 ) | ( n11393 & n11402 ) ;
  assign n11611 = ( ~n11393 & n11403 ) | ( ~n11393 & n11610 ) | ( n11403 & n11610 ) ;
  assign n11612 = n3800 & ~n10998 ;
  assign n11613 = n3799 & ~n9967 ;
  assign n11614 = n3700 & n9971 ;
  assign n11615 = n3802 & n9969 ;
  assign n11616 = n11614 | n11615 ;
  assign n11617 = ( ~n11612 & n11613 ) | ( ~n11612 & n11616 ) | ( n11613 & n11616 ) ;
  assign n11618 = ( ~x29 & n11612 ) | ( ~x29 & n11617 ) | ( n11612 & n11617 ) ;
  assign n11619 = ( n11612 & n11617 ) | ( n11612 & ~n11618 ) | ( n11617 & ~n11618 ) ;
  assign n11620 = ( x29 & n11618 ) | ( x29 & ~n11619 ) | ( n11618 & ~n11619 ) ;
  assign n11621 = ( n11609 & n11611 ) | ( n11609 & n11620 ) | ( n11611 & n11620 ) ;
  assign n11622 = ( n11402 & n11420 ) | ( n11402 & ~n11610 ) | ( n11420 & ~n11610 ) ;
  assign n11623 = ( n11403 & ~n11421 ) | ( n11403 & n11622 ) | ( ~n11421 & n11622 ) ;
  assign n11624 = n607 & n9975 ;
  assign n11625 = n1250 & n9973 ;
  assign n11626 = n11624 | n11625 ;
  assign n11627 = n606 & ~n9971 ;
  assign n11628 = ( n606 & n11626 ) | ( n606 & ~n11627 ) | ( n11626 & ~n11627 ) ;
  assign n11629 = ( n9971 & ~n9973 ) | ( n9971 & n10019 ) | ( ~n9973 & n10019 ) ;
  assign n11630 = ( n9973 & ~n10020 ) | ( n9973 & n11629 ) | ( ~n10020 & n11629 ) ;
  assign n11631 = n1248 & n11630 ;
  assign n11632 = n11628 | n11631 ;
  assign n11633 = ( n11621 & ~n11623 ) | ( n11621 & n11632 ) | ( ~n11623 & n11632 ) ;
  assign n11634 = n3800 & ~n11121 ;
  assign n11635 = n3799 & ~n9963 ;
  assign n11636 = n3700 & ~n9967 ;
  assign n11637 = n3802 & n9965 ;
  assign n11638 = n11636 | n11637 ;
  assign n11639 = ( ~n11634 & n11635 ) | ( ~n11634 & n11638 ) | ( n11635 & n11638 ) ;
  assign n11640 = ( ~x29 & n11634 ) | ( ~x29 & n11639 ) | ( n11634 & n11639 ) ;
  assign n11641 = ( n11634 & n11639 ) | ( n11634 & ~n11640 ) | ( n11639 & ~n11640 ) ;
  assign n11642 = ( x29 & n11640 ) | ( x29 & ~n11641 ) | ( n11640 & ~n11641 ) ;
  assign n11643 = ( n11070 & n11430 ) | ( n11070 & ~n11431 ) | ( n11430 & ~n11431 ) ;
  assign n11644 = ( n11421 & n11431 ) | ( n11421 & ~n11643 ) | ( n11431 & ~n11643 ) ;
  assign n11645 = ( n11633 & n11642 ) | ( n11633 & ~n11644 ) | ( n11642 & ~n11644 ) ;
  assign n11646 = ( ~n11431 & n11433 ) | ( ~n11431 & n11442 ) | ( n11433 & n11442 ) ;
  assign n11647 = ( ~n11442 & n11443 ) | ( ~n11442 & n11646 ) | ( n11443 & n11646 ) ;
  assign n11648 = n4202 & ~n10567 ;
  assign n11649 = n4201 & n9955 ;
  assign n11650 = n4200 & n9959 ;
  assign n11651 = n4345 & ~n9957 ;
  assign n11652 = n11650 | n11651 ;
  assign n11653 = ( ~n11648 & n11649 ) | ( ~n11648 & n11652 ) | ( n11649 & n11652 ) ;
  assign n11654 = ( ~x26 & n11648 ) | ( ~x26 & n11653 ) | ( n11648 & n11653 ) ;
  assign n11655 = ( n11648 & n11653 ) | ( n11648 & ~n11654 ) | ( n11653 & ~n11654 ) ;
  assign n11656 = ( x26 & n11654 ) | ( x26 & ~n11655 ) | ( n11654 & ~n11655 ) ;
  assign n11657 = ( n11645 & ~n11647 ) | ( n11645 & n11656 ) | ( ~n11647 & n11656 ) ;
  assign n11658 = ( ~n11443 & n11445 ) | ( ~n11443 & n11454 ) | ( n11445 & n11454 ) ;
  assign n11659 = ( ~n11454 & n11455 ) | ( ~n11454 & n11658 ) | ( n11455 & n11658 ) ;
  assign n11660 = n4713 & n10454 ;
  assign n11661 = n4712 & n9947 ;
  assign n11662 = n4709 & n9951 ;
  assign n11663 = n4792 & n9949 ;
  assign n11664 = n11662 | n11663 ;
  assign n11665 = ( ~n11660 & n11661 ) | ( ~n11660 & n11664 ) | ( n11661 & n11664 ) ;
  assign n11666 = ( ~x23 & n11660 ) | ( ~x23 & n11665 ) | ( n11660 & n11665 ) ;
  assign n11667 = ( n11660 & n11665 ) | ( n11660 & ~n11666 ) | ( n11665 & ~n11666 ) ;
  assign n11668 = ( x23 & n11666 ) | ( x23 & ~n11667 ) | ( n11666 & ~n11667 ) ;
  assign n11669 = ( n11657 & ~n11659 ) | ( n11657 & n11668 ) | ( ~n11659 & n11668 ) ;
  assign n11670 = ( n11455 & ~n11464 ) | ( n11455 & n11466 ) | ( ~n11464 & n11466 ) ;
  assign n11671 = ( ~n11455 & n11467 ) | ( ~n11455 & n11670 ) | ( n11467 & n11670 ) ;
  assign n11672 = n4713 & n10466 ;
  assign n11673 = n4712 & n9945 ;
  assign n11674 = n4709 & n9949 ;
  assign n11675 = n4792 & n9947 ;
  assign n11676 = n11674 | n11675 ;
  assign n11677 = ( ~n11672 & n11673 ) | ( ~n11672 & n11676 ) | ( n11673 & n11676 ) ;
  assign n11678 = ( ~x23 & n11672 ) | ( ~x23 & n11677 ) | ( n11672 & n11677 ) ;
  assign n11679 = ( n11672 & n11677 ) | ( n11672 & ~n11678 ) | ( n11677 & ~n11678 ) ;
  assign n11680 = ( x23 & n11678 ) | ( x23 & ~n11679 ) | ( n11678 & ~n11679 ) ;
  assign n11681 = ( n11669 & ~n11671 ) | ( n11669 & n11680 ) | ( ~n11671 & n11680 ) ;
  assign n11682 = ( n11467 & ~n11469 ) | ( n11467 & n11478 ) | ( ~n11469 & n11478 ) ;
  assign n11683 = ( n11469 & ~n11479 ) | ( n11469 & n11682 ) | ( ~n11479 & n11682 ) ;
  assign n11684 = n4974 & n10174 ;
  assign n11685 = n5398 & n9916 ;
  assign n11686 = n4972 | n9883 ;
  assign n11687 = n4973 & ~n9941 ;
  assign n11688 = ( ~n9883 & n11686 ) | ( ~n9883 & n11687 ) | ( n11686 & n11687 ) ;
  assign n11689 = ( ~n11684 & n11685 ) | ( ~n11684 & n11688 ) | ( n11685 & n11688 ) ;
  assign n11690 = ( ~x20 & n11684 ) | ( ~x20 & n11689 ) | ( n11684 & n11689 ) ;
  assign n11691 = ( n11684 & n11689 ) | ( n11684 & ~n11690 ) | ( n11689 & ~n11690 ) ;
  assign n11692 = ( x20 & n11690 ) | ( x20 & ~n11691 ) | ( n11690 & ~n11691 ) ;
  assign n11693 = ( n11681 & n11683 ) | ( n11681 & n11692 ) | ( n11683 & n11692 ) ;
  assign n11694 = ( n11479 & ~n11481 ) | ( n11479 & n11490 ) | ( ~n11481 & n11490 ) ;
  assign n11695 = ( n11481 & ~n11491 ) | ( n11481 & n11694 ) | ( ~n11491 & n11694 ) ;
  assign n11696 = n5508 & n10362 ;
  assign n11697 = n5507 & n10346 ;
  assign n11698 = n5504 & ~n10057 ;
  assign n11699 = n5666 & ~n10302 ;
  assign n11700 = n11698 | n11699 ;
  assign n11701 = ( ~n11696 & n11697 ) | ( ~n11696 & n11700 ) | ( n11697 & n11700 ) ;
  assign n11702 = ( ~x17 & n11696 ) | ( ~x17 & n11701 ) | ( n11696 & n11701 ) ;
  assign n11703 = ( n11696 & n11701 ) | ( n11696 & ~n11702 ) | ( n11701 & ~n11702 ) ;
  assign n11704 = ( x17 & n11702 ) | ( x17 & ~n11703 ) | ( n11702 & ~n11703 ) ;
  assign n11705 = ( n11693 & n11695 ) | ( n11693 & n11704 ) | ( n11695 & n11704 ) ;
  assign n11706 = n5508 & n10348 ;
  assign n11707 = n5666 & n10346 ;
  assign n11708 = n5504 & ~n10302 ;
  assign n11709 = n5507 | n11708 ;
  assign n11710 = ( ~n11706 & n11707 ) | ( ~n11706 & n11709 ) | ( n11707 & n11709 ) ;
  assign n11711 = ( ~x17 & n11706 ) | ( ~x17 & n11710 ) | ( n11706 & n11710 ) ;
  assign n11712 = ( n11706 & n11710 ) | ( n11706 & ~n11711 ) | ( n11710 & ~n11711 ) ;
  assign n11713 = ( x17 & n11711 ) | ( x17 & ~n11712 ) | ( n11711 & ~n11712 ) ;
  assign n11714 = ( ~n11491 & n11493 ) | ( ~n11491 & n11502 ) | ( n11493 & n11502 ) ;
  assign n11715 = ( ~n11502 & n11503 ) | ( ~n11502 & n11714 ) | ( n11503 & n11714 ) ;
  assign n11716 = ( n11705 & n11713 ) | ( n11705 & ~n11715 ) | ( n11713 & ~n11715 ) ;
  assign n11717 = ( n11621 & n11623 ) | ( n11621 & n11632 ) | ( n11623 & n11632 ) ;
  assign n11718 = ( n11623 & n11633 ) | ( n11623 & ~n11717 ) | ( n11633 & ~n11717 ) ;
  assign n11719 = n3800 & ~n11273 ;
  assign n11720 = n3799 & n9965 ;
  assign n11721 = n3700 & n9969 ;
  assign n11722 = n3802 & ~n9967 ;
  assign n11723 = n11721 | n11722 ;
  assign n11724 = ( ~n11719 & n11720 ) | ( ~n11719 & n11723 ) | ( n11720 & n11723 ) ;
  assign n11725 = ( ~x29 & n11719 ) | ( ~x29 & n11724 ) | ( n11719 & n11724 ) ;
  assign n11726 = ( n11719 & n11724 ) | ( n11719 & ~n11725 ) | ( n11724 & ~n11725 ) ;
  assign n11727 = ( x29 & n11725 ) | ( x29 & ~n11726 ) | ( n11725 & ~n11726 ) ;
  assign n11728 = n4202 & n10859 ;
  assign n11729 = n4201 & n9959 ;
  assign n11730 = n4200 & ~n9963 ;
  assign n11731 = n4345 & n9961 ;
  assign n11732 = n11730 | n11731 ;
  assign n11733 = ( ~n11728 & n11729 ) | ( ~n11728 & n11732 ) | ( n11729 & n11732 ) ;
  assign n11734 = ( ~x26 & n11728 ) | ( ~x26 & n11733 ) | ( n11728 & n11733 ) ;
  assign n11735 = ( n11728 & n11733 ) | ( n11728 & ~n11734 ) | ( n11733 & ~n11734 ) ;
  assign n11736 = ( x26 & n11734 ) | ( x26 & ~n11735 ) | ( n11734 & ~n11735 ) ;
  assign n11737 = ( ~n11718 & n11727 ) | ( ~n11718 & n11736 ) | ( n11727 & n11736 ) ;
  assign n11738 = ( n11633 & ~n11642 ) | ( n11633 & n11644 ) | ( ~n11642 & n11644 ) ;
  assign n11739 = ( ~n11633 & n11645 ) | ( ~n11633 & n11738 ) | ( n11645 & n11738 ) ;
  assign n11740 = n4202 & ~n10869 ;
  assign n11741 = n4201 & ~n9957 ;
  assign n11742 = n4200 & n9961 ;
  assign n11743 = n4345 & n9959 ;
  assign n11744 = n11742 | n11743 ;
  assign n11745 = ( ~n11740 & n11741 ) | ( ~n11740 & n11744 ) | ( n11741 & n11744 ) ;
  assign n11746 = ( ~x26 & n11740 ) | ( ~x26 & n11745 ) | ( n11740 & n11745 ) ;
  assign n11747 = ( n11740 & n11745 ) | ( n11740 & ~n11746 ) | ( n11745 & ~n11746 ) ;
  assign n11748 = ( x26 & n11746 ) | ( x26 & ~n11747 ) | ( n11746 & ~n11747 ) ;
  assign n11749 = ( n11737 & ~n11739 ) | ( n11737 & n11748 ) | ( ~n11739 & n11748 ) ;
  assign n11750 = ( ~n11645 & n11647 ) | ( ~n11645 & n11656 ) | ( n11647 & n11656 ) ;
  assign n11751 = ( ~n11656 & n11657 ) | ( ~n11656 & n11750 ) | ( n11657 & n11750 ) ;
  assign n11752 = n4713 & n10557 ;
  assign n11753 = n4712 & n9949 ;
  assign n11754 = n4709 & ~n9953 ;
  assign n11755 = n4792 & n9951 ;
  assign n11756 = n11754 | n11755 ;
  assign n11757 = ( ~n11752 & n11753 ) | ( ~n11752 & n11756 ) | ( n11753 & n11756 ) ;
  assign n11758 = ( ~x23 & n11752 ) | ( ~x23 & n11757 ) | ( n11752 & n11757 ) ;
  assign n11759 = ( n11752 & n11757 ) | ( n11752 & ~n11758 ) | ( n11757 & ~n11758 ) ;
  assign n11760 = ( x23 & n11758 ) | ( x23 & ~n11759 ) | ( n11758 & ~n11759 ) ;
  assign n11761 = ( n11749 & ~n11751 ) | ( n11749 & n11760 ) | ( ~n11751 & n11760 ) ;
  assign n11762 = ( ~n11657 & n11659 ) | ( ~n11657 & n11668 ) | ( n11659 & n11668 ) ;
  assign n11763 = ( ~n11668 & n11669 ) | ( ~n11668 & n11762 ) | ( n11669 & n11762 ) ;
  assign n11764 = n4974 & ~n10390 ;
  assign n11765 = n5398 & ~n9941 ;
  assign n11766 = n4973 & n9945 ;
  assign n11767 = n4972 & n9943 ;
  assign n11768 = n11766 | n11767 ;
  assign n11769 = ( ~n11764 & n11765 ) | ( ~n11764 & n11768 ) | ( n11765 & n11768 ) ;
  assign n11770 = ( ~x20 & n11764 ) | ( ~x20 & n11769 ) | ( n11764 & n11769 ) ;
  assign n11771 = ( n11764 & n11769 ) | ( n11764 & ~n11770 ) | ( n11769 & ~n11770 ) ;
  assign n11772 = ( x20 & n11770 ) | ( x20 & ~n11771 ) | ( n11770 & ~n11771 ) ;
  assign n11773 = ( n11761 & ~n11763 ) | ( n11761 & n11772 ) | ( ~n11763 & n11772 ) ;
  assign n11774 = ( ~n11669 & n11671 ) | ( ~n11669 & n11680 ) | ( n11671 & n11680 ) ;
  assign n11775 = ( ~n11680 & n11681 ) | ( ~n11680 & n11774 ) | ( n11681 & n11774 ) ;
  assign n11776 = n4974 & n10284 ;
  assign n11777 = n5398 & ~n9883 ;
  assign n11778 = n4973 & n9943 ;
  assign n11779 = n4972 & ~n9941 ;
  assign n11780 = n11778 | n11779 ;
  assign n11781 = ( ~n11776 & n11777 ) | ( ~n11776 & n11780 ) | ( n11777 & n11780 ) ;
  assign n11782 = ( ~x20 & n11776 ) | ( ~x20 & n11781 ) | ( n11776 & n11781 ) ;
  assign n11783 = ( n11776 & n11781 ) | ( n11776 & ~n11782 ) | ( n11781 & ~n11782 ) ;
  assign n11784 = ( x20 & n11782 ) | ( x20 & ~n11783 ) | ( n11782 & ~n11783 ) ;
  assign n11785 = ( n11773 & ~n11775 ) | ( n11773 & n11784 ) | ( ~n11775 & n11784 ) ;
  assign n11786 = ( n11681 & ~n11683 ) | ( n11681 & n11692 ) | ( ~n11683 & n11692 ) ;
  assign n11787 = ( n11683 & ~n11693 ) | ( n11683 & n11786 ) | ( ~n11693 & n11786 ) ;
  assign n11788 = n5508 & ~n10305 ;
  assign n11789 = n5507 & ~n10302 ;
  assign n11790 = n5504 & ~n9937 ;
  assign n11791 = n5666 & ~n10057 ;
  assign n11792 = n11790 | n11791 ;
  assign n11793 = ( ~n11788 & n11789 ) | ( ~n11788 & n11792 ) | ( n11789 & n11792 ) ;
  assign n11794 = ( ~x17 & n11788 ) | ( ~x17 & n11793 ) | ( n11788 & n11793 ) ;
  assign n11795 = ( n11788 & n11793 ) | ( n11788 & ~n11794 ) | ( n11793 & ~n11794 ) ;
  assign n11796 = ( x17 & n11794 ) | ( x17 & ~n11795 ) | ( n11794 & ~n11795 ) ;
  assign n11797 = ( n11785 & n11787 ) | ( n11785 & n11796 ) | ( n11787 & n11796 ) ;
  assign n11798 = x14 | n10637 ;
  assign n11799 = ( x14 & n10637 ) | ( x14 & ~n11798 ) | ( n10637 & ~n11798 ) ;
  assign n11800 = n11798 & ~n11799 ;
  assign n11801 = ( n11693 & ~n11695 ) | ( n11693 & n11704 ) | ( ~n11695 & n11704 ) ;
  assign n11802 = ( n11695 & ~n11705 ) | ( n11695 & n11801 ) | ( ~n11705 & n11801 ) ;
  assign n11803 = ( n11797 & n11800 ) | ( n11797 & n11802 ) | ( n11800 & n11802 ) ;
  assign n11804 = n10001 & ~n10003 ;
  assign n11805 = ~n10001 & n10003 ;
  assign n11806 = ( n1248 & n11804 ) | ( n1248 & n11805 ) | ( n11804 & n11805 ) ;
  assign n11807 = ( n606 & ~n10001 ) | ( n606 & n11806 ) | ( ~n10001 & n11806 ) ;
  assign n11808 = ( n1250 & ~n10003 ) | ( n1250 & n11806 ) | ( ~n10003 & n11806 ) ;
  assign n11809 = n11807 | n11808 ;
  assign n11810 = n195 | n873 ;
  assign n11811 = n1129 | n11810 ;
  assign n11812 = ( ~n54 & n100 ) | ( ~n54 & n102 ) | ( n100 & n102 ) ;
  assign n11813 = n1059 | n11812 ;
  assign n11814 = ( n2251 & ~n11811 ) | ( n2251 & n11813 ) | ( ~n11811 & n11813 ) ;
  assign n11815 = n11811 | n11814 ;
  assign n11816 = n151 | n233 ;
  assign n11817 = n1278 | n4548 ;
  assign n11818 = ( n11815 & n11816 ) | ( n11815 & ~n11817 ) | ( n11816 & ~n11817 ) ;
  assign n11819 = n1347 | n1435 ;
  assign n11820 = n5527 | n11819 ;
  assign n11821 = n949 | n1204 ;
  assign n11822 = n689 | n786 ;
  assign n11823 = ( n265 & n810 ) | ( n265 & ~n11822 ) | ( n810 & ~n11822 ) ;
  assign n11824 = n11822 | n11823 ;
  assign n11825 = ( n466 & n2071 ) | ( n466 & ~n11824 ) | ( n2071 & ~n11824 ) ;
  assign n11826 = n11824 | n11825 ;
  assign n11827 = ( ~n11820 & n11821 ) | ( ~n11820 & n11826 ) | ( n11821 & n11826 ) ;
  assign n11828 = n11820 | n11827 ;
  assign n11829 = ( n11817 & ~n11818 ) | ( n11817 & n11828 ) | ( ~n11818 & n11828 ) ;
  assign n11830 = n11818 | n11829 ;
  assign n11831 = n3298 & ~n6073 ;
  assign n11832 = n904 | n2467 ;
  assign n11833 = n583 | n2918 ;
  assign n11834 = ( n1032 & ~n11832 ) | ( n1032 & n11833 ) | ( ~n11832 & n11833 ) ;
  assign n11835 = ( n338 & n11832 ) | ( n338 & ~n11834 ) | ( n11832 & ~n11834 ) ;
  assign n11836 = n11834 | n11835 ;
  assign n11837 = n509 | n3024 ;
  assign n11838 = ( n3000 & ~n3059 ) | ( n3000 & n11837 ) | ( ~n3059 & n11837 ) ;
  assign n11839 = n3059 | n11838 ;
  assign n11840 = ( ~n6073 & n11836 ) | ( ~n6073 & n11839 ) | ( n11836 & n11839 ) ;
  assign n11841 = ( n11830 & n11831 ) | ( n11830 & ~n11840 ) | ( n11831 & ~n11840 ) ;
  assign n11842 = ~n11830 & n11841 ;
  assign n11843 = n11809 & ~n11842 ;
  assign n11844 = n718 | n3761 ;
  assign n11845 = n11544 | n11844 ;
  assign n11846 = n1024 | n1860 ;
  assign n11847 = n110 | n120 ;
  assign n11848 = n329 | n338 ;
  assign n11849 = ( n762 & n783 ) | ( n762 & ~n11848 ) | ( n783 & ~n11848 ) ;
  assign n11850 = n11848 | n11849 ;
  assign n11851 = ( n922 & ~n11847 ) | ( n922 & n11850 ) | ( ~n11847 & n11850 ) ;
  assign n11852 = n11847 | n11851 ;
  assign n11853 = ( n2362 & ~n11846 ) | ( n2362 & n11852 ) | ( ~n11846 & n11852 ) ;
  assign n11854 = n11846 | n11853 ;
  assign n11855 = ( ~n78 & n109 ) | ( ~n78 & n129 ) | ( n109 & n129 ) ;
  assign n11856 = ( n1556 & ~n1581 ) | ( n1556 & n11855 ) | ( ~n1581 & n11855 ) ;
  assign n11857 = n1581 | n11856 ;
  assign n11858 = ( ~n11844 & n11854 ) | ( ~n11844 & n11857 ) | ( n11854 & n11857 ) ;
  assign n11859 = ( ~n10148 & n11845 ) | ( ~n10148 & n11858 ) | ( n11845 & n11858 ) ;
  assign n11860 = ( ~n10148 & n11111 ) | ( ~n10148 & n11859 ) | ( n11111 & n11859 ) ;
  assign n11861 = ~n11859 & n11860 ;
  assign n11862 = n607 & ~n10003 ;
  assign n11863 = n1250 & ~n10001 ;
  assign n11864 = n11862 | n11863 ;
  assign n11865 = n606 & ~n9999 ;
  assign n11866 = ( n606 & n11864 ) | ( n606 & ~n11865 ) | ( n11864 & ~n11865 ) ;
  assign n11867 = n9999 & n11805 ;
  assign n11868 = ( n9999 & n10005 ) | ( n9999 & ~n11867 ) | ( n10005 & ~n11867 ) ;
  assign n11869 = n1248 & n11868 ;
  assign n11870 = n11866 | n11869 ;
  assign n11871 = ( n11843 & ~n11861 ) | ( n11843 & n11870 ) | ( ~n11861 & n11870 ) ;
  assign n11872 = n1193 | n3470 ;
  assign n11873 = n105 | n318 ;
  assign n11874 = n1887 | n11873 ;
  assign n11875 = n4117 | n5190 ;
  assign n11876 = ( n66 & n102 ) | ( n66 & n145 ) | ( n102 & n145 ) ;
  assign n11877 = ( n514 & n587 ) | ( n514 & ~n11876 ) | ( n587 & ~n11876 ) ;
  assign n11878 = n11876 | n11877 ;
  assign n11879 = ( ~n11874 & n11875 ) | ( ~n11874 & n11878 ) | ( n11875 & n11878 ) ;
  assign n11880 = n11874 | n11879 ;
  assign n11881 = ( n6165 & ~n11872 ) | ( n6165 & n11880 ) | ( ~n11872 & n11880 ) ;
  assign n11882 = n11872 | n11881 ;
  assign n11883 = ( n1076 & ~n4112 ) | ( n1076 & n11882 ) | ( ~n4112 & n11882 ) ;
  assign n11884 = ( n621 & n4112 ) | ( n621 & ~n11883 ) | ( n4112 & ~n11883 ) ;
  assign n11885 = n11883 | n11884 ;
  assign n11886 = n607 & ~n10001 ;
  assign n11887 = n1250 & n9999 ;
  assign n11888 = n11886 | n11887 ;
  assign n11889 = n606 & n9997 ;
  assign n11890 = ( n606 & n11888 ) | ( n606 & ~n11889 ) | ( n11888 & ~n11889 ) ;
  assign n11891 = ( n9997 & n9999 ) | ( n9997 & n10006 ) | ( n9999 & n10006 ) ;
  assign n11892 = ( n9999 & n10007 ) | ( n9999 & ~n11891 ) | ( n10007 & ~n11891 ) ;
  assign n11893 = n1248 & n11892 ;
  assign n11894 = n11890 | n11893 ;
  assign n11895 = ( n11871 & n11885 ) | ( n11871 & n11894 ) | ( n11885 & n11894 ) ;
  assign n11896 = n1237 | n4069 ;
  assign n11897 = n177 | n262 ;
  assign n11898 = ( n220 & n11896 ) | ( n220 & ~n11897 ) | ( n11896 & ~n11897 ) ;
  assign n11899 = ~n11896 & n11898 ;
  assign n11900 = n582 | n1967 ;
  assign n11901 = n10520 | n11900 ;
  assign n11902 = n135 | n885 ;
  assign n11903 = ( n1588 & n4255 ) | ( n1588 & ~n11902 ) | ( n4255 & ~n11902 ) ;
  assign n11904 = n11902 | n11903 ;
  assign n11905 = n567 | n591 ;
  assign n11906 = ( n581 & n856 ) | ( n581 & ~n11905 ) | ( n856 & ~n11905 ) ;
  assign n11907 = n11905 | n11906 ;
  assign n11908 = ( n969 & n3646 ) | ( n969 & ~n11907 ) | ( n3646 & ~n11907 ) ;
  assign n11909 = n11907 | n11908 ;
  assign n11910 = ( ~n11901 & n11904 ) | ( ~n11901 & n11909 ) | ( n11904 & n11909 ) ;
  assign n11911 = n11901 | n11910 ;
  assign n11912 = ( n11078 & n11899 ) | ( n11078 & n11911 ) | ( n11899 & n11911 ) ;
  assign n11913 = n11899 & ~n11912 ;
  assign n11914 = ~n3180 & n11913 ;
  assign n11915 = n147 | n2661 ;
  assign n11916 = ( n1131 & n1802 ) | ( n1131 & ~n11915 ) | ( n1802 & ~n11915 ) ;
  assign n11917 = n11915 | n11916 ;
  assign n11918 = ( n64 & n109 ) | ( n64 & n255 ) | ( n109 & n255 ) ;
  assign n11919 = ( n238 & n713 ) | ( n238 & ~n11918 ) | ( n713 & ~n11918 ) ;
  assign n11920 = n11918 | n11919 ;
  assign n11921 = n212 | n991 ;
  assign n11922 = n2188 | n11921 ;
  assign n11923 = n11920 | n11922 ;
  assign n11924 = ( n4888 & ~n11917 ) | ( n4888 & n11923 ) | ( ~n11917 & n11923 ) ;
  assign n11925 = ( n11914 & n11917 ) | ( n11914 & n11924 ) | ( n11917 & n11924 ) ;
  assign n11926 = ( ~n805 & n11914 ) | ( ~n805 & n11925 ) | ( n11914 & n11925 ) ;
  assign n11927 = ~n11925 & n11926 ;
  assign n11928 = n607 & n9999 ;
  assign n11929 = n1250 & ~n9997 ;
  assign n11930 = n11928 | n11929 ;
  assign n11931 = n606 & ~n9995 ;
  assign n11932 = ( n606 & n11930 ) | ( n606 & ~n11931 ) | ( n11930 & ~n11931 ) ;
  assign n11933 = ( n9995 & ~n9997 ) | ( n9995 & n10007 ) | ( ~n9997 & n10007 ) ;
  assign n11934 = ( ~n10007 & n10008 ) | ( ~n10007 & n11933 ) | ( n10008 & n11933 ) ;
  assign n11935 = n1248 & n11934 ;
  assign n11936 = n11932 | n11935 ;
  assign n11937 = ( n11895 & ~n11927 ) | ( n11895 & n11936 ) | ( ~n11927 & n11936 ) ;
  assign n11938 = n679 | n1460 ;
  assign n11939 = n492 | n888 ;
  assign n11940 = ( n968 & ~n2011 ) | ( n968 & n2357 ) | ( ~n2011 & n2357 ) ;
  assign n11941 = ( n2011 & ~n11939 ) | ( n2011 & n11940 ) | ( ~n11939 & n11940 ) ;
  assign n11942 = n11939 | n11941 ;
  assign n11943 = ( ~n258 & n536 ) | ( ~n258 & n851 ) | ( n536 & n851 ) ;
  assign n11944 = n258 | n11943 ;
  assign n11945 = ( ~n11938 & n11942 ) | ( ~n11938 & n11944 ) | ( n11942 & n11944 ) ;
  assign n11946 = n11938 | n11945 ;
  assign n11947 = ( n2771 & ~n10332 ) | ( n2771 & n11946 ) | ( ~n10332 & n11946 ) ;
  assign n11948 = ( n3729 & ~n10332 ) | ( n3729 & n11947 ) | ( ~n10332 & n11947 ) ;
  assign n11949 = n192 | n488 ;
  assign n11950 = ( ~n54 & n302 ) | ( ~n54 & n3141 ) | ( n302 & n3141 ) ;
  assign n11951 = n930 | n11950 ;
  assign n11952 = ( n3741 & ~n11949 ) | ( n3741 & n11951 ) | ( ~n11949 & n11951 ) ;
  assign n11953 = n11949 | n11952 ;
  assign n11954 = ~n2343 & n11047 ;
  assign n11955 = n1589 | n1914 ;
  assign n11956 = n1312 | n2798 ;
  assign n11957 = ( n648 & n2214 ) | ( n648 & ~n3339 ) | ( n2214 & ~n3339 ) ;
  assign n11958 = n3339 | n11957 ;
  assign n11959 = ( ~n11955 & n11956 ) | ( ~n11955 & n11958 ) | ( n11956 & n11958 ) ;
  assign n11960 = n11955 | n11959 ;
  assign n11961 = ( n11953 & n11954 ) | ( n11953 & ~n11960 ) | ( n11954 & ~n11960 ) ;
  assign n11962 = ~n11953 & n11961 ;
  assign n11963 = ( ~n10332 & n11948 ) | ( ~n10332 & n11962 ) | ( n11948 & n11962 ) ;
  assign n11964 = ~n11948 & n11963 ;
  assign n11965 = n607 & ~n9997 ;
  assign n11966 = n1250 & n9995 ;
  assign n11967 = n11965 | n11966 ;
  assign n11968 = n606 & ~n9993 ;
  assign n11969 = ( n606 & n11967 ) | ( n606 & ~n11968 ) | ( n11967 & ~n11968 ) ;
  assign n11970 = ( n9993 & n9995 ) | ( n9993 & ~n10009 ) | ( n9995 & ~n10009 ) ;
  assign n11971 = ( n10008 & n10009 ) | ( n10008 & ~n11970 ) | ( n10009 & ~n11970 ) ;
  assign n11972 = n1248 & ~n11971 ;
  assign n11973 = n11969 | n11972 ;
  assign n11974 = ( n11937 & ~n11964 ) | ( n11937 & n11973 ) | ( ~n11964 & n11973 ) ;
  assign n11975 = ( n41 & n48 ) | ( n41 & n145 ) | ( n48 & n145 ) ;
  assign n11976 = n293 | n11975 ;
  assign n11977 = n2428 | n11976 ;
  assign n11978 = n662 | n792 ;
  assign n11979 = ( n192 & n4397 ) | ( n192 & ~n11978 ) | ( n4397 & ~n11978 ) ;
  assign n11980 = n11978 | n11979 ;
  assign n11981 = ( n48 & n57 ) | ( n48 & n60 ) | ( n57 & n60 ) ;
  assign n11982 = ( n316 & n492 ) | ( n316 & ~n777 ) | ( n492 & ~n777 ) ;
  assign n11983 = ( n550 & ~n777 ) | ( n550 & n921 ) | ( ~n777 & n921 ) ;
  assign n11984 = n777 | n11983 ;
  assign n11985 = ( ~n11981 & n11982 ) | ( ~n11981 & n11984 ) | ( n11982 & n11984 ) ;
  assign n11986 = n11981 | n11985 ;
  assign n11987 = ( ~n11977 & n11980 ) | ( ~n11977 & n11986 ) | ( n11980 & n11986 ) ;
  assign n11988 = n11977 | n11987 ;
  assign n11989 = ( n4078 & n6143 ) | ( n4078 & ~n11988 ) | ( n6143 & ~n11988 ) ;
  assign n11990 = n11988 | n11989 ;
  assign n11991 = n359 | n6217 ;
  assign n11992 = n5152 | n11002 ;
  assign n11993 = n208 | n1363 ;
  assign n11994 = ( n129 & n136 ) | ( n129 & n152 ) | ( n136 & n152 ) ;
  assign n11995 = ( n416 & ~n11993 ) | ( n416 & n11994 ) | ( ~n11993 & n11994 ) ;
  assign n11996 = n11993 | n11995 ;
  assign n11997 = n1510 | n3131 ;
  assign n11998 = n10600 | n11997 ;
  assign n11999 = ( n336 & ~n11996 ) | ( n336 & n11998 ) | ( ~n11996 & n11998 ) ;
  assign n12000 = n11996 | n11999 ;
  assign n12001 = n371 | n1093 ;
  assign n12002 = ( ~n11992 & n12000 ) | ( ~n11992 & n12001 ) | ( n12000 & n12001 ) ;
  assign n12003 = n11992 | n12002 ;
  assign n12004 = n11991 | n12003 ;
  assign n12005 = ( n482 & n760 ) | ( n482 & ~n862 ) | ( n760 & ~n862 ) ;
  assign n12006 = n862 | n12005 ;
  assign n12007 = n980 | n1808 ;
  assign n12008 = ( n10843 & ~n12006 ) | ( n10843 & n12007 ) | ( ~n12006 & n12007 ) ;
  assign n12009 = n12006 | n12008 ;
  assign n12010 = n3961 | n10619 ;
  assign n12011 = n1235 | n2846 ;
  assign n12012 = n266 | n746 ;
  assign n12013 = ( n586 & n2349 ) | ( n586 & ~n12012 ) | ( n2349 & ~n12012 ) ;
  assign n12014 = n12012 | n12013 ;
  assign n12015 = ( ~n12010 & n12011 ) | ( ~n12010 & n12014 ) | ( n12011 & n12014 ) ;
  assign n12016 = n12010 | n12015 ;
  assign n12017 = ( ~n11991 & n12009 ) | ( ~n11991 & n12016 ) | ( n12009 & n12016 ) ;
  assign n12018 = ( ~n11990 & n12004 ) | ( ~n11990 & n12017 ) | ( n12004 & n12017 ) ;
  assign n12019 = n11990 | n12018 ;
  assign n12020 = n607 & n9995 ;
  assign n12021 = n1250 & n9993 ;
  assign n12022 = n12020 | n12021 ;
  assign n12023 = n606 & ~n9991 ;
  assign n12024 = ( n606 & n12022 ) | ( n606 & ~n12023 ) | ( n12022 & ~n12023 ) ;
  assign n12025 = ( n9991 & n9993 ) | ( n9991 & ~n10009 ) | ( n9993 & ~n10009 ) ;
  assign n12026 = ( n10009 & ~n10010 ) | ( n10009 & n12025 ) | ( ~n10010 & n12025 ) ;
  assign n12027 = n1248 & n12026 ;
  assign n12028 = n12024 | n12027 ;
  assign n12029 = ( n11974 & n12019 ) | ( n11974 & n12028 ) | ( n12019 & n12028 ) ;
  assign n12030 = ( ~n128 & n3945 ) | ( ~n128 & n4136 ) | ( n3945 & n4136 ) ;
  assign n12031 = n1543 | n2361 ;
  assign n12032 = ( n4494 & n11826 ) | ( n4494 & ~n12031 ) | ( n11826 & ~n12031 ) ;
  assign n12033 = n12031 | n12032 ;
  assign n12034 = n55 | n186 ;
  assign n12035 = ( n759 & n1027 ) | ( n759 & ~n12034 ) | ( n1027 & ~n12034 ) ;
  assign n12036 = n12034 | n12035 ;
  assign n12037 = n318 | n782 ;
  assign n12038 = ( n1093 & ~n2523 ) | ( n1093 & n12037 ) | ( ~n2523 & n12037 ) ;
  assign n12039 = ( n2523 & ~n12036 ) | ( n2523 & n12038 ) | ( ~n12036 & n12038 ) ;
  assign n12040 = n12036 | n12039 ;
  assign n12041 = ( ~n4136 & n12033 ) | ( ~n4136 & n12040 ) | ( n12033 & n12040 ) ;
  assign n12042 = ( ~n128 & n12030 ) | ( ~n128 & n12041 ) | ( n12030 & n12041 ) ;
  assign n12043 = n128 | n12042 ;
  assign n12044 = n607 & n9993 ;
  assign n12045 = n1250 & n9991 ;
  assign n12046 = n12044 | n12045 ;
  assign n12047 = n606 & ~n9989 ;
  assign n12048 = ( n606 & n12046 ) | ( n606 & ~n12047 ) | ( n12046 & ~n12047 ) ;
  assign n12049 = ( n9989 & n9991 ) | ( n9989 & ~n10010 ) | ( n9991 & ~n10010 ) ;
  assign n12050 = ( n10010 & ~n10011 ) | ( n10010 & n12049 ) | ( ~n10011 & n12049 ) ;
  assign n12051 = n1248 & n12050 ;
  assign n12052 = n12048 | n12051 ;
  assign n12053 = ( n12029 & n12043 ) | ( n12029 & n12052 ) | ( n12043 & n12052 ) ;
  assign n12054 = n2523 | n4510 ;
  assign n12055 = ( n613 & n876 ) | ( n613 & ~n2077 ) | ( n876 & ~n2077 ) ;
  assign n12056 = n2077 | n12055 ;
  assign n12057 = n150 | n205 ;
  assign n12058 = ( ~n333 & n1096 ) | ( ~n333 & n12057 ) | ( n1096 & n12057 ) ;
  assign n12059 = ( n333 & n1057 ) | ( n333 & ~n2558 ) | ( n1057 & ~n2558 ) ;
  assign n12060 = n2558 | n12059 ;
  assign n12061 = ( ~n12056 & n12058 ) | ( ~n12056 & n12060 ) | ( n12058 & n12060 ) ;
  assign n12062 = n12056 | n12061 ;
  assign n12063 = ( n3403 & ~n12054 ) | ( n3403 & n12062 ) | ( ~n12054 & n12062 ) ;
  assign n12064 = n12054 | n12063 ;
  assign n12065 = ( ~n2697 & n3366 ) | ( ~n2697 & n11533 ) | ( n3366 & n11533 ) ;
  assign n12066 = ( n2697 & ~n12064 ) | ( n2697 & n12065 ) | ( ~n12064 & n12065 ) ;
  assign n12067 = n12064 | n12066 ;
  assign n12068 = n607 & n9991 ;
  assign n12069 = n1250 & n9989 ;
  assign n12070 = n12068 | n12069 ;
  assign n12071 = n606 & n9987 ;
  assign n12072 = ( n606 & n12070 ) | ( n606 & ~n12071 ) | ( n12070 & ~n12071 ) ;
  assign n12073 = ( n9987 & ~n9989 ) | ( n9987 & n10011 ) | ( ~n9989 & n10011 ) ;
  assign n12074 = ( ~n10011 & n10012 ) | ( ~n10011 & n12073 ) | ( n10012 & n12073 ) ;
  assign n12075 = n1248 & ~n12074 ;
  assign n12076 = n12072 | n12075 ;
  assign n12077 = ( n12053 & n12067 ) | ( n12053 & n12076 ) | ( n12067 & n12076 ) ;
  assign n12078 = ( n1091 & ~n1850 ) | ( n1091 & n2116 ) | ( ~n1850 & n2116 ) ;
  assign n12079 = n3522 | n3997 ;
  assign n12080 = n3291 | n12079 ;
  assign n12081 = n1693 | n2205 ;
  assign n12082 = n1401 | n1595 ;
  assign n12083 = n55 | n517 ;
  assign n12084 = ( n185 & n783 ) | ( n185 & ~n12083 ) | ( n783 & ~n12083 ) ;
  assign n12085 = n12083 | n12084 ;
  assign n12086 = ( ~n12081 & n12082 ) | ( ~n12081 & n12085 ) | ( n12082 & n12085 ) ;
  assign n12087 = n12081 | n12086 ;
  assign n12088 = ( n3571 & ~n12080 ) | ( n3571 & n12087 ) | ( ~n12080 & n12087 ) ;
  assign n12089 = n12080 | n12088 ;
  assign n12090 = ( ~n1091 & n5740 ) | ( ~n1091 & n12089 ) | ( n5740 & n12089 ) ;
  assign n12091 = ( ~n1850 & n12078 ) | ( ~n1850 & n12090 ) | ( n12078 & n12090 ) ;
  assign n12092 = n1850 | n12091 ;
  assign n12093 = n607 & n9989 ;
  assign n12094 = n1250 & ~n9987 ;
  assign n12095 = n12093 | n12094 ;
  assign n12096 = n606 & ~n9985 ;
  assign n12097 = ( n606 & n12095 ) | ( n606 & ~n12096 ) | ( n12095 & ~n12096 ) ;
  assign n12098 = ( ~n9985 & n9987 ) | ( ~n9985 & n10012 ) | ( n9987 & n10012 ) ;
  assign n12099 = ( ~n10012 & n10013 ) | ( ~n10012 & n12098 ) | ( n10013 & n12098 ) ;
  assign n12100 = n1248 & ~n12099 ;
  assign n12101 = n12097 | n12100 ;
  assign n12102 = ( n12077 & n12092 ) | ( n12077 & n12101 ) | ( n12092 & n12101 ) ;
  assign n12103 = n133 | n1621 ;
  assign n12104 = ( n98 & n145 ) | ( n98 & n149 ) | ( n145 & n149 ) ;
  assign n12105 = n174 | n12104 ;
  assign n12106 = ( n3544 & ~n12103 ) | ( n3544 & n12105 ) | ( ~n12103 & n12105 ) ;
  assign n12107 = n12103 | n12106 ;
  assign n12108 = ( ~n1877 & n4860 ) | ( ~n1877 & n12107 ) | ( n4860 & n12107 ) ;
  assign n12109 = n1056 | n3569 ;
  assign n12110 = n1473 | n1533 ;
  assign n12111 = ( n3139 & ~n12109 ) | ( n3139 & n12110 ) | ( ~n12109 & n12110 ) ;
  assign n12112 = n12109 | n12111 ;
  assign n12113 = ( n4072 & n10940 ) | ( n4072 & ~n12112 ) | ( n10940 & ~n12112 ) ;
  assign n12114 = n12112 | n12113 ;
  assign n12115 = n225 | n549 ;
  assign n12116 = n922 | n12115 ;
  assign n12117 = n582 | n795 ;
  assign n12118 = ( n3710 & ~n12116 ) | ( n3710 & n12117 ) | ( ~n12116 & n12117 ) ;
  assign n12119 = n12116 | n12118 ;
  assign n12120 = ( ~n12107 & n12114 ) | ( ~n12107 & n12119 ) | ( n12114 & n12119 ) ;
  assign n12121 = ( ~n1877 & n12108 ) | ( ~n1877 & n12120 ) | ( n12108 & n12120 ) ;
  assign n12122 = n1877 | n12121 ;
  assign n12123 = n607 & ~n9987 ;
  assign n12124 = n1250 & n9985 ;
  assign n12125 = n12123 | n12124 ;
  assign n12126 = n606 & n9983 ;
  assign n12127 = ( n606 & n12125 ) | ( n606 & ~n12126 ) | ( n12125 & ~n12126 ) ;
  assign n12128 = ( n9983 & ~n9985 ) | ( n9983 & n10013 ) | ( ~n9985 & n10013 ) ;
  assign n12129 = ( ~n10013 & n10014 ) | ( ~n10013 & n12128 ) | ( n10014 & n12128 ) ;
  assign n12130 = n1248 & ~n12129 ;
  assign n12131 = n12127 | n12130 ;
  assign n12132 = ( n12102 & n12122 ) | ( n12102 & n12131 ) | ( n12122 & n12131 ) ;
  assign n12133 = ( ~n11351 & n11554 ) | ( ~n11351 & n11563 ) | ( n11554 & n11563 ) ;
  assign n12134 = ( ~n11563 & n11564 ) | ( ~n11563 & n12133 ) | ( n11564 & n12133 ) ;
  assign n12135 = n3800 & n11606 ;
  assign n12136 = n3799 & n9975 ;
  assign n12137 = n3700 & n9979 ;
  assign n12138 = n3802 & n9977 ;
  assign n12139 = n12137 | n12138 ;
  assign n12140 = ( ~n12135 & n12136 ) | ( ~n12135 & n12139 ) | ( n12136 & n12139 ) ;
  assign n12141 = ( ~x29 & n12135 ) | ( ~x29 & n12140 ) | ( n12135 & n12140 ) ;
  assign n12142 = ( n12135 & n12140 ) | ( n12135 & ~n12141 ) | ( n12140 & ~n12141 ) ;
  assign n12143 = ( x29 & n12141 ) | ( x29 & ~n12142 ) | ( n12141 & ~n12142 ) ;
  assign n12144 = ( n12132 & ~n12134 ) | ( n12132 & n12143 ) | ( ~n12134 & n12143 ) ;
  assign n12145 = ( ~n11351 & n11564 ) | ( ~n11351 & n11581 ) | ( n11564 & n11581 ) ;
  assign n12146 = ( n11351 & ~n11582 ) | ( n11351 & n12145 ) | ( ~n11582 & n12145 ) ;
  assign n12147 = n607 & ~n9983 ;
  assign n12148 = n1250 & n9981 ;
  assign n12149 = n12147 | n12148 ;
  assign n12150 = n606 & ~n9979 ;
  assign n12151 = ( n606 & n12149 ) | ( n606 & ~n12150 ) | ( n12149 & ~n12150 ) ;
  assign n12152 = ( n9979 & ~n9981 ) | ( n9979 & n10015 ) | ( ~n9981 & n10015 ) ;
  assign n12153 = ( n9981 & ~n10016 ) | ( n9981 & n12152 ) | ( ~n10016 & n12152 ) ;
  assign n12154 = n1248 & n12153 ;
  assign n12155 = n12151 | n12154 ;
  assign n12156 = ( n12144 & n12146 ) | ( n12144 & n12155 ) | ( n12146 & n12155 ) ;
  assign n12157 = ( ~n11351 & n11582 ) | ( ~n11351 & n11596 ) | ( n11582 & n11596 ) ;
  assign n12158 = ( ~n11582 & n11597 ) | ( ~n11582 & n12157 ) | ( n11597 & n12157 ) ;
  assign n12159 = n607 & n9981 ;
  assign n12160 = n1250 & n9979 ;
  assign n12161 = n12159 | n12160 ;
  assign n12162 = n606 & ~n9977 ;
  assign n12163 = ( n606 & n12161 ) | ( n606 & ~n12162 ) | ( n12161 & ~n12162 ) ;
  assign n12164 = ( n9977 & ~n9979 ) | ( n9977 & n10016 ) | ( ~n9979 & n10016 ) ;
  assign n12165 = ( n9979 & ~n10017 ) | ( n9979 & n12164 ) | ( ~n10017 & n12164 ) ;
  assign n12166 = n1248 & n12165 ;
  assign n12167 = n12163 | n12166 ;
  assign n12168 = ( n12156 & ~n12158 ) | ( n12156 & n12167 ) | ( ~n12158 & n12167 ) ;
  assign n12169 = ( ~n11597 & n11599 ) | ( ~n11597 & n11608 ) | ( n11599 & n11608 ) ;
  assign n12170 = ( ~n11608 & n11609 ) | ( ~n11608 & n12169 ) | ( n11609 & n12169 ) ;
  assign n12171 = n3800 & n11428 ;
  assign n12172 = n3799 & n9969 ;
  assign n12173 = n3700 & n9973 ;
  assign n12174 = n3802 & n9971 ;
  assign n12175 = n12173 | n12174 ;
  assign n12176 = ( ~n12171 & n12172 ) | ( ~n12171 & n12175 ) | ( n12172 & n12175 ) ;
  assign n12177 = ( ~x29 & n12171 ) | ( ~x29 & n12176 ) | ( n12171 & n12176 ) ;
  assign n12178 = ( n12171 & n12176 ) | ( n12171 & ~n12177 ) | ( n12176 & ~n12177 ) ;
  assign n12179 = ( x29 & n12177 ) | ( x29 & ~n12178 ) | ( n12177 & ~n12178 ) ;
  assign n12180 = ( n12168 & ~n12170 ) | ( n12168 & n12179 ) | ( ~n12170 & n12179 ) ;
  assign n12181 = ( n11609 & ~n11611 ) | ( n11609 & n11620 ) | ( ~n11611 & n11620 ) ;
  assign n12182 = ( n11611 & ~n11621 ) | ( n11611 & n12181 ) | ( ~n11621 & n12181 ) ;
  assign n12183 = n4202 & ~n10929 ;
  assign n12184 = n4201 & n9961 ;
  assign n12185 = n4200 & n9965 ;
  assign n12186 = n4345 & ~n9963 ;
  assign n12187 = n12185 | n12186 ;
  assign n12188 = ( ~n12183 & n12184 ) | ( ~n12183 & n12187 ) | ( n12184 & n12187 ) ;
  assign n12189 = ( ~x26 & n12183 ) | ( ~x26 & n12188 ) | ( n12183 & n12188 ) ;
  assign n12190 = ( n12183 & n12188 ) | ( n12183 & ~n12189 ) | ( n12188 & ~n12189 ) ;
  assign n12191 = ( x26 & n12189 ) | ( x26 & ~n12190 ) | ( n12189 & ~n12190 ) ;
  assign n12192 = ( n12180 & n12182 ) | ( n12180 & n12191 ) | ( n12182 & n12191 ) ;
  assign n12193 = ( n11727 & n11736 ) | ( n11727 & ~n11737 ) | ( n11736 & ~n11737 ) ;
  assign n12194 = ( n11718 & n11737 ) | ( n11718 & ~n12193 ) | ( n11737 & ~n12193 ) ;
  assign n12195 = n4713 & ~n10750 ;
  assign n12196 = n4712 & ~n9953 ;
  assign n12197 = n4709 & ~n9957 ;
  assign n12198 = n4792 & n9955 ;
  assign n12199 = n12197 | n12198 ;
  assign n12200 = ( ~n12195 & n12196 ) | ( ~n12195 & n12199 ) | ( n12196 & n12199 ) ;
  assign n12201 = ( ~x23 & n12195 ) | ( ~x23 & n12200 ) | ( n12195 & n12200 ) ;
  assign n12202 = ( n12195 & n12200 ) | ( n12195 & ~n12201 ) | ( n12200 & ~n12201 ) ;
  assign n12203 = ( x23 & n12201 ) | ( x23 & ~n12202 ) | ( n12201 & ~n12202 ) ;
  assign n12204 = ( n12192 & ~n12194 ) | ( n12192 & n12203 ) | ( ~n12194 & n12203 ) ;
  assign n12205 = ( ~n11737 & n11739 ) | ( ~n11737 & n11748 ) | ( n11739 & n11748 ) ;
  assign n12206 = ( ~n11748 & n11749 ) | ( ~n11748 & n12205 ) | ( n11749 & n12205 ) ;
  assign n12207 = n4713 & ~n10652 ;
  assign n12208 = n4712 & n9951 ;
  assign n12209 = n4709 & n9955 ;
  assign n12210 = n4792 & ~n9953 ;
  assign n12211 = n12209 | n12210 ;
  assign n12212 = ( ~n12207 & n12208 ) | ( ~n12207 & n12211 ) | ( n12208 & n12211 ) ;
  assign n12213 = ( ~x23 & n12207 ) | ( ~x23 & n12212 ) | ( n12207 & n12212 ) ;
  assign n12214 = ( n12207 & n12212 ) | ( n12207 & ~n12213 ) | ( n12212 & ~n12213 ) ;
  assign n12215 = ( x23 & n12213 ) | ( x23 & ~n12214 ) | ( n12213 & ~n12214 ) ;
  assign n12216 = ( n12204 & ~n12206 ) | ( n12204 & n12215 ) | ( ~n12206 & n12215 ) ;
  assign n12217 = ( ~n11749 & n11751 ) | ( ~n11749 & n11760 ) | ( n11751 & n11760 ) ;
  assign n12218 = ( ~n11760 & n11761 ) | ( ~n11760 & n12217 ) | ( n11761 & n12217 ) ;
  assign n12219 = n4974 & n10271 ;
  assign n12220 = n5398 & n9943 ;
  assign n12221 = n4973 & n9947 ;
  assign n12222 = n4972 & n9945 ;
  assign n12223 = n12221 | n12222 ;
  assign n12224 = ( ~n12219 & n12220 ) | ( ~n12219 & n12223 ) | ( n12220 & n12223 ) ;
  assign n12225 = ( ~x20 & n12219 ) | ( ~x20 & n12224 ) | ( n12219 & n12224 ) ;
  assign n12226 = ( n12219 & n12224 ) | ( n12219 & ~n12225 ) | ( n12224 & ~n12225 ) ;
  assign n12227 = ( x20 & n12225 ) | ( x20 & ~n12226 ) | ( n12225 & ~n12226 ) ;
  assign n12228 = ( n12216 & ~n12218 ) | ( n12216 & n12227 ) | ( ~n12218 & n12227 ) ;
  assign n12229 = ( ~n11761 & n11763 ) | ( ~n11761 & n11772 ) | ( n11763 & n11772 ) ;
  assign n12230 = ( ~n11772 & n11773 ) | ( ~n11772 & n12229 ) | ( n11773 & n12229 ) ;
  assign n12231 = n5508 & n10040 ;
  assign n12232 = n5507 & ~n9937 ;
  assign n12233 = n5504 & ~n9883 ;
  assign n12234 = n5666 & n9916 ;
  assign n12235 = n12233 | n12234 ;
  assign n12236 = ( ~n12231 & n12232 ) | ( ~n12231 & n12235 ) | ( n12232 & n12235 ) ;
  assign n12237 = ( ~x17 & n12231 ) | ( ~x17 & n12236 ) | ( n12231 & n12236 ) ;
  assign n12238 = ( n12231 & n12236 ) | ( n12231 & ~n12237 ) | ( n12236 & ~n12237 ) ;
  assign n12239 = ( x17 & n12237 ) | ( x17 & ~n12238 ) | ( n12237 & ~n12238 ) ;
  assign n12240 = ( n12228 & ~n12230 ) | ( n12228 & n12239 ) | ( ~n12230 & n12239 ) ;
  assign n12241 = ( ~n11773 & n11775 ) | ( ~n11773 & n11784 ) | ( n11775 & n11784 ) ;
  assign n12242 = ( ~n11784 & n11785 ) | ( ~n11784 & n12241 ) | ( n11785 & n12241 ) ;
  assign n12243 = n5508 & ~n10064 ;
  assign n12244 = n5507 & ~n10057 ;
  assign n12245 = n5504 & n9916 ;
  assign n12246 = n5666 & ~n9937 ;
  assign n12247 = n12245 | n12246 ;
  assign n12248 = ( ~n12243 & n12244 ) | ( ~n12243 & n12247 ) | ( n12244 & n12247 ) ;
  assign n12249 = ( ~x17 & n12243 ) | ( ~x17 & n12248 ) | ( n12243 & n12248 ) ;
  assign n12250 = ( n12243 & n12248 ) | ( n12243 & ~n12249 ) | ( n12248 & ~n12249 ) ;
  assign n12251 = ( x17 & n12249 ) | ( x17 & ~n12250 ) | ( n12249 & ~n12250 ) ;
  assign n12252 = ( n12240 & ~n12242 ) | ( n12240 & n12251 ) | ( ~n12242 & n12251 ) ;
  assign n12253 = ( n11785 & ~n11787 ) | ( n11785 & n11796 ) | ( ~n11787 & n11796 ) ;
  assign n12254 = ( n11787 & ~n11797 ) | ( n11787 & n12253 ) | ( ~n11797 & n12253 ) ;
  assign n12255 = ~n5970 & n10346 ;
  assign n12256 = ( n10346 & n10635 ) | ( n10346 & ~n12255 ) | ( n10635 & ~n12255 ) ;
  assign n12257 = ( ~x14 & n5966 ) | ( ~x14 & n12256 ) | ( n5966 & n12256 ) ;
  assign n12258 = ( n5966 & n12256 ) | ( n5966 & ~n12257 ) | ( n12256 & ~n12257 ) ;
  assign n12259 = ( x14 & n12257 ) | ( x14 & ~n12258 ) | ( n12257 & ~n12258 ) ;
  assign n12260 = ( n12252 & n12254 ) | ( n12252 & n12259 ) | ( n12254 & n12259 ) ;
  assign n12261 = ( ~n12156 & n12158 ) | ( ~n12156 & n12167 ) | ( n12158 & n12167 ) ;
  assign n12262 = ( ~n12167 & n12168 ) | ( ~n12167 & n12261 ) | ( n12168 & n12261 ) ;
  assign n12263 = n3800 & n11630 ;
  assign n12264 = n3799 & n9971 ;
  assign n12265 = n3700 & n9975 ;
  assign n12266 = n3802 & n9973 ;
  assign n12267 = n12265 | n12266 ;
  assign n12268 = ( ~n12263 & n12264 ) | ( ~n12263 & n12267 ) | ( n12264 & n12267 ) ;
  assign n12269 = ( ~x29 & n12263 ) | ( ~x29 & n12268 ) | ( n12263 & n12268 ) ;
  assign n12270 = ( n12263 & n12268 ) | ( n12263 & ~n12269 ) | ( n12268 & ~n12269 ) ;
  assign n12271 = ( x29 & n12269 ) | ( x29 & ~n12270 ) | ( n12269 & ~n12270 ) ;
  assign n12272 = n4202 & ~n11273 ;
  assign n12273 = n4201 & n9965 ;
  assign n12274 = n4200 & n9969 ;
  assign n12275 = n4345 & ~n9967 ;
  assign n12276 = n12274 | n12275 ;
  assign n12277 = ( ~n12272 & n12273 ) | ( ~n12272 & n12276 ) | ( n12273 & n12276 ) ;
  assign n12278 = ( ~x26 & n12272 ) | ( ~x26 & n12277 ) | ( n12272 & n12277 ) ;
  assign n12279 = ( n12272 & n12277 ) | ( n12272 & ~n12278 ) | ( n12277 & ~n12278 ) ;
  assign n12280 = ( x26 & n12278 ) | ( x26 & ~n12279 ) | ( n12278 & ~n12279 ) ;
  assign n12281 = ( ~n12262 & n12271 ) | ( ~n12262 & n12280 ) | ( n12271 & n12280 ) ;
  assign n12282 = n4202 & ~n11121 ;
  assign n12283 = n4201 & ~n9963 ;
  assign n12284 = n4200 & ~n9967 ;
  assign n12285 = n4345 & n9965 ;
  assign n12286 = n12284 | n12285 ;
  assign n12287 = ( ~n12282 & n12283 ) | ( ~n12282 & n12286 ) | ( n12283 & n12286 ) ;
  assign n12288 = ( ~x26 & n12282 ) | ( ~x26 & n12287 ) | ( n12282 & n12287 ) ;
  assign n12289 = ( n12282 & n12287 ) | ( n12282 & ~n12288 ) | ( n12287 & ~n12288 ) ;
  assign n12290 = ( x26 & n12288 ) | ( x26 & ~n12289 ) | ( n12288 & ~n12289 ) ;
  assign n12291 = ( ~n12168 & n12170 ) | ( ~n12168 & n12179 ) | ( n12170 & n12179 ) ;
  assign n12292 = ( ~n12179 & n12180 ) | ( ~n12179 & n12291 ) | ( n12180 & n12291 ) ;
  assign n12293 = ( n12281 & n12290 ) | ( n12281 & ~n12292 ) | ( n12290 & ~n12292 ) ;
  assign n12294 = ( n12180 & ~n12182 ) | ( n12180 & n12191 ) | ( ~n12182 & n12191 ) ;
  assign n12295 = ( n12182 & ~n12192 ) | ( n12182 & n12294 ) | ( ~n12192 & n12294 ) ;
  assign n12296 = n4713 & ~n10567 ;
  assign n12297 = n4712 & n9955 ;
  assign n12298 = n4709 & n9959 ;
  assign n12299 = n4792 & ~n9957 ;
  assign n12300 = n12298 | n12299 ;
  assign n12301 = ( ~n12296 & n12297 ) | ( ~n12296 & n12300 ) | ( n12297 & n12300 ) ;
  assign n12302 = ( ~x23 & n12296 ) | ( ~x23 & n12301 ) | ( n12296 & n12301 ) ;
  assign n12303 = ( n12296 & n12301 ) | ( n12296 & ~n12302 ) | ( n12301 & ~n12302 ) ;
  assign n12304 = ( x23 & n12302 ) | ( x23 & ~n12303 ) | ( n12302 & ~n12303 ) ;
  assign n12305 = ( n12293 & n12295 ) | ( n12293 & n12304 ) | ( n12295 & n12304 ) ;
  assign n12306 = ( ~n12192 & n12194 ) | ( ~n12192 & n12203 ) | ( n12194 & n12203 ) ;
  assign n12307 = ( ~n12203 & n12204 ) | ( ~n12203 & n12306 ) | ( n12204 & n12306 ) ;
  assign n12308 = n4974 & n10454 ;
  assign n12309 = n5398 & n9947 ;
  assign n12310 = n4973 & n9951 ;
  assign n12311 = n4972 & n9949 ;
  assign n12312 = n12310 | n12311 ;
  assign n12313 = ( ~n12308 & n12309 ) | ( ~n12308 & n12312 ) | ( n12309 & n12312 ) ;
  assign n12314 = ( ~x20 & n12308 ) | ( ~x20 & n12313 ) | ( n12308 & n12313 ) ;
  assign n12315 = ( n12308 & n12313 ) | ( n12308 & ~n12314 ) | ( n12313 & ~n12314 ) ;
  assign n12316 = ( x20 & n12314 ) | ( x20 & ~n12315 ) | ( n12314 & ~n12315 ) ;
  assign n12317 = ( n12305 & ~n12307 ) | ( n12305 & n12316 ) | ( ~n12307 & n12316 ) ;
  assign n12318 = ( ~n12204 & n12206 ) | ( ~n12204 & n12215 ) | ( n12206 & n12215 ) ;
  assign n12319 = ( ~n12215 & n12216 ) | ( ~n12215 & n12318 ) | ( n12216 & n12318 ) ;
  assign n12320 = n4974 & n10466 ;
  assign n12321 = n5398 & n9945 ;
  assign n12322 = n4973 & n9949 ;
  assign n12323 = n4972 & n9947 ;
  assign n12324 = n12322 | n12323 ;
  assign n12325 = ( ~n12320 & n12321 ) | ( ~n12320 & n12324 ) | ( n12321 & n12324 ) ;
  assign n12326 = ( ~x20 & n12320 ) | ( ~x20 & n12325 ) | ( n12320 & n12325 ) ;
  assign n12327 = ( n12320 & n12325 ) | ( n12320 & ~n12326 ) | ( n12325 & ~n12326 ) ;
  assign n12328 = ( x20 & n12326 ) | ( x20 & ~n12327 ) | ( n12326 & ~n12327 ) ;
  assign n12329 = ( n12317 & ~n12319 ) | ( n12317 & n12328 ) | ( ~n12319 & n12328 ) ;
  assign n12330 = ( ~n12216 & n12218 ) | ( ~n12216 & n12227 ) | ( n12218 & n12227 ) ;
  assign n12331 = ( ~n12227 & n12228 ) | ( ~n12227 & n12330 ) | ( n12228 & n12330 ) ;
  assign n12332 = n5508 & n10174 ;
  assign n12333 = n5507 & n9916 ;
  assign n12334 = n5666 | n9883 ;
  assign n12335 = n5504 & ~n9941 ;
  assign n12336 = ( ~n9883 & n12334 ) | ( ~n9883 & n12335 ) | ( n12334 & n12335 ) ;
  assign n12337 = ( ~n12332 & n12333 ) | ( ~n12332 & n12336 ) | ( n12333 & n12336 ) ;
  assign n12338 = ( ~x17 & n12332 ) | ( ~x17 & n12337 ) | ( n12332 & n12337 ) ;
  assign n12339 = ( n12332 & n12337 ) | ( n12332 & ~n12338 ) | ( n12337 & ~n12338 ) ;
  assign n12340 = ( x17 & n12338 ) | ( x17 & ~n12339 ) | ( n12338 & ~n12339 ) ;
  assign n12341 = ( n12329 & ~n12331 ) | ( n12329 & n12340 ) | ( ~n12331 & n12340 ) ;
  assign n12342 = ( ~n12228 & n12230 ) | ( ~n12228 & n12239 ) | ( n12230 & n12239 ) ;
  assign n12343 = ( ~n12239 & n12240 ) | ( ~n12239 & n12342 ) | ( n12240 & n12342 ) ;
  assign n12344 = n5966 & n10362 ;
  assign n12345 = n6464 & n10346 ;
  assign n12346 = n5970 & ~n10057 ;
  assign n12347 = n5969 & ~n10302 ;
  assign n12348 = n12346 | n12347 ;
  assign n12349 = ( ~n12344 & n12345 ) | ( ~n12344 & n12348 ) | ( n12345 & n12348 ) ;
  assign n12350 = ( ~x14 & n12344 ) | ( ~x14 & n12349 ) | ( n12344 & n12349 ) ;
  assign n12351 = ( n12344 & n12349 ) | ( n12344 & ~n12350 ) | ( n12349 & ~n12350 ) ;
  assign n12352 = ( x14 & n12350 ) | ( x14 & ~n12351 ) | ( n12350 & ~n12351 ) ;
  assign n12353 = ( n12341 & ~n12343 ) | ( n12341 & n12352 ) | ( ~n12343 & n12352 ) ;
  assign n12354 = n5966 & n10348 ;
  assign n12355 = n5969 & n10346 ;
  assign n12356 = n5970 & ~n10302 ;
  assign n12357 = n6464 | n12356 ;
  assign n12358 = ( ~n12354 & n12355 ) | ( ~n12354 & n12357 ) | ( n12355 & n12357 ) ;
  assign n12359 = ( ~x14 & n12354 ) | ( ~x14 & n12358 ) | ( n12354 & n12358 ) ;
  assign n12360 = ( n12354 & n12358 ) | ( n12354 & ~n12359 ) | ( n12358 & ~n12359 ) ;
  assign n12361 = ( x14 & n12359 ) | ( x14 & ~n12360 ) | ( n12359 & ~n12360 ) ;
  assign n12362 = ( ~n12240 & n12242 ) | ( ~n12240 & n12251 ) | ( n12242 & n12251 ) ;
  assign n12363 = ( ~n12251 & n12252 ) | ( ~n12251 & n12362 ) | ( n12252 & n12362 ) ;
  assign n12364 = ( n12353 & n12361 ) | ( n12353 & ~n12363 ) | ( n12361 & ~n12363 ) ;
  assign n12365 = ( ~n12144 & n12146 ) | ( ~n12144 & n12155 ) | ( n12146 & n12155 ) ;
  assign n12366 = ( n12144 & ~n12156 ) | ( n12144 & n12365 ) | ( ~n12156 & n12365 ) ;
  assign n12367 = n3800 & n11400 ;
  assign n12368 = n3799 & n9973 ;
  assign n12369 = n3700 & n9977 ;
  assign n12370 = n3802 & n9975 ;
  assign n12371 = n12369 | n12370 ;
  assign n12372 = ( ~n12367 & n12368 ) | ( ~n12367 & n12371 ) | ( n12368 & n12371 ) ;
  assign n12373 = ( ~x29 & n12367 ) | ( ~x29 & n12372 ) | ( n12367 & n12372 ) ;
  assign n12374 = ( n12367 & n12372 ) | ( n12367 & ~n12373 ) | ( n12372 & ~n12373 ) ;
  assign n12375 = ( x29 & n12373 ) | ( x29 & ~n12374 ) | ( n12373 & ~n12374 ) ;
  assign n12376 = n4202 & ~n10998 ;
  assign n12377 = n4201 & ~n9967 ;
  assign n12378 = n4200 & n9971 ;
  assign n12379 = n4345 & n9969 ;
  assign n12380 = n12378 | n12379 ;
  assign n12381 = ( ~n12376 & n12377 ) | ( ~n12376 & n12380 ) | ( n12377 & n12380 ) ;
  assign n12382 = ( ~x26 & n12376 ) | ( ~x26 & n12381 ) | ( n12376 & n12381 ) ;
  assign n12383 = ( n12376 & n12381 ) | ( n12376 & ~n12382 ) | ( n12381 & ~n12382 ) ;
  assign n12384 = ( x26 & n12382 ) | ( x26 & ~n12383 ) | ( n12382 & ~n12383 ) ;
  assign n12385 = ( n12366 & n12375 ) | ( n12366 & n12384 ) | ( n12375 & n12384 ) ;
  assign n12386 = ( n12271 & n12280 ) | ( n12271 & ~n12281 ) | ( n12280 & ~n12281 ) ;
  assign n12387 = ( n12262 & n12281 ) | ( n12262 & ~n12386 ) | ( n12281 & ~n12386 ) ;
  assign n12388 = n4713 & n10859 ;
  assign n12389 = n4712 & n9959 ;
  assign n12390 = n4709 & ~n9963 ;
  assign n12391 = n4792 & n9961 ;
  assign n12392 = n12390 | n12391 ;
  assign n12393 = ( ~n12388 & n12389 ) | ( ~n12388 & n12392 ) | ( n12389 & n12392 ) ;
  assign n12394 = ( ~x23 & n12388 ) | ( ~x23 & n12393 ) | ( n12388 & n12393 ) ;
  assign n12395 = ( n12388 & n12393 ) | ( n12388 & ~n12394 ) | ( n12393 & ~n12394 ) ;
  assign n12396 = ( x23 & n12394 ) | ( x23 & ~n12395 ) | ( n12394 & ~n12395 ) ;
  assign n12397 = ( n12385 & ~n12387 ) | ( n12385 & n12396 ) | ( ~n12387 & n12396 ) ;
  assign n12398 = ( n12281 & ~n12290 ) | ( n12281 & n12292 ) | ( ~n12290 & n12292 ) ;
  assign n12399 = ( ~n12281 & n12293 ) | ( ~n12281 & n12398 ) | ( n12293 & n12398 ) ;
  assign n12400 = n4713 & ~n10869 ;
  assign n12401 = n4712 & ~n9957 ;
  assign n12402 = n4709 & n9961 ;
  assign n12403 = n4792 & n9959 ;
  assign n12404 = n12402 | n12403 ;
  assign n12405 = ( ~n12400 & n12401 ) | ( ~n12400 & n12404 ) | ( n12401 & n12404 ) ;
  assign n12406 = ( ~x23 & n12400 ) | ( ~x23 & n12405 ) | ( n12400 & n12405 ) ;
  assign n12407 = ( n12400 & n12405 ) | ( n12400 & ~n12406 ) | ( n12405 & ~n12406 ) ;
  assign n12408 = ( x23 & n12406 ) | ( x23 & ~n12407 ) | ( n12406 & ~n12407 ) ;
  assign n12409 = ( n12397 & ~n12399 ) | ( n12397 & n12408 ) | ( ~n12399 & n12408 ) ;
  assign n12410 = ( n12293 & ~n12295 ) | ( n12293 & n12304 ) | ( ~n12295 & n12304 ) ;
  assign n12411 = ( n12295 & ~n12305 ) | ( n12295 & n12410 ) | ( ~n12305 & n12410 ) ;
  assign n12412 = n4974 & n10557 ;
  assign n12413 = n5398 & n9949 ;
  assign n12414 = n4973 & ~n9953 ;
  assign n12415 = n4972 & n9951 ;
  assign n12416 = n12414 | n12415 ;
  assign n12417 = ( ~n12412 & n12413 ) | ( ~n12412 & n12416 ) | ( n12413 & n12416 ) ;
  assign n12418 = ( ~x20 & n12412 ) | ( ~x20 & n12417 ) | ( n12412 & n12417 ) ;
  assign n12419 = ( n12412 & n12417 ) | ( n12412 & ~n12418 ) | ( n12417 & ~n12418 ) ;
  assign n12420 = ( x20 & n12418 ) | ( x20 & ~n12419 ) | ( n12418 & ~n12419 ) ;
  assign n12421 = ( n12409 & n12411 ) | ( n12409 & n12420 ) | ( n12411 & n12420 ) ;
  assign n12422 = ( ~n12305 & n12307 ) | ( ~n12305 & n12316 ) | ( n12307 & n12316 ) ;
  assign n12423 = ( ~n12316 & n12317 ) | ( ~n12316 & n12422 ) | ( n12317 & n12422 ) ;
  assign n12424 = n5508 & ~n10390 ;
  assign n12425 = n5507 & ~n9941 ;
  assign n12426 = n5504 & n9945 ;
  assign n12427 = n5666 & n9943 ;
  assign n12428 = n12426 | n12427 ;
  assign n12429 = ( ~n12424 & n12425 ) | ( ~n12424 & n12428 ) | ( n12425 & n12428 ) ;
  assign n12430 = ( ~x17 & n12424 ) | ( ~x17 & n12429 ) | ( n12424 & n12429 ) ;
  assign n12431 = ( n12424 & n12429 ) | ( n12424 & ~n12430 ) | ( n12429 & ~n12430 ) ;
  assign n12432 = ( x17 & n12430 ) | ( x17 & ~n12431 ) | ( n12430 & ~n12431 ) ;
  assign n12433 = ( n12421 & ~n12423 ) | ( n12421 & n12432 ) | ( ~n12423 & n12432 ) ;
  assign n12434 = ( ~n12317 & n12319 ) | ( ~n12317 & n12328 ) | ( n12319 & n12328 ) ;
  assign n12435 = ( ~n12328 & n12329 ) | ( ~n12328 & n12434 ) | ( n12329 & n12434 ) ;
  assign n12436 = n5508 & n10284 ;
  assign n12437 = n5507 & ~n9883 ;
  assign n12438 = n5504 & n9943 ;
  assign n12439 = n5666 & ~n9941 ;
  assign n12440 = n12438 | n12439 ;
  assign n12441 = ( ~n12436 & n12437 ) | ( ~n12436 & n12440 ) | ( n12437 & n12440 ) ;
  assign n12442 = ( ~x17 & n12436 ) | ( ~x17 & n12441 ) | ( n12436 & n12441 ) ;
  assign n12443 = ( n12436 & n12441 ) | ( n12436 & ~n12442 ) | ( n12441 & ~n12442 ) ;
  assign n12444 = ( x17 & n12442 ) | ( x17 & ~n12443 ) | ( n12442 & ~n12443 ) ;
  assign n12445 = ( n12433 & ~n12435 ) | ( n12433 & n12444 ) | ( ~n12435 & n12444 ) ;
  assign n12446 = ( ~n12329 & n12331 ) | ( ~n12329 & n12340 ) | ( n12331 & n12340 ) ;
  assign n12447 = ( ~n12340 & n12341 ) | ( ~n12340 & n12446 ) | ( n12341 & n12446 ) ;
  assign n12448 = n5966 & ~n10305 ;
  assign n12449 = n6464 & ~n10302 ;
  assign n12450 = n5970 & ~n9937 ;
  assign n12451 = n5969 & ~n10057 ;
  assign n12452 = n12450 | n12451 ;
  assign n12453 = ( ~n12448 & n12449 ) | ( ~n12448 & n12452 ) | ( n12449 & n12452 ) ;
  assign n12454 = ( ~x14 & n12448 ) | ( ~x14 & n12453 ) | ( n12448 & n12453 ) ;
  assign n12455 = ( n12448 & n12453 ) | ( n12448 & ~n12454 ) | ( n12453 & ~n12454 ) ;
  assign n12456 = ( x14 & n12454 ) | ( x14 & ~n12455 ) | ( n12454 & ~n12455 ) ;
  assign n12457 = ( n12445 & ~n12447 ) | ( n12445 & n12456 ) | ( ~n12447 & n12456 ) ;
  assign n12458 = x11 | n10986 ;
  assign n12459 = ( x11 & n10986 ) | ( x11 & ~n12458 ) | ( n10986 & ~n12458 ) ;
  assign n12460 = n12458 & ~n12459 ;
  assign n12461 = ( ~n12341 & n12343 ) | ( ~n12341 & n12352 ) | ( n12343 & n12352 ) ;
  assign n12462 = ( ~n12352 & n12353 ) | ( ~n12352 & n12461 ) | ( n12353 & n12461 ) ;
  assign n12463 = ( n12457 & n12460 ) | ( n12457 & ~n12462 ) | ( n12460 & ~n12462 ) ;
  assign n12464 = ( n58 & n96 ) | ( n58 & ~n10003 ) | ( n96 & ~n10003 ) ;
  assign n12465 = n3800 & n11892 ;
  assign n12466 = n3799 & ~n9997 ;
  assign n12467 = n3700 & ~n10001 ;
  assign n12468 = n3802 & n9999 ;
  assign n12469 = n12467 | n12468 ;
  assign n12470 = ( ~n12465 & n12466 ) | ( ~n12465 & n12469 ) | ( n12466 & n12469 ) ;
  assign n12471 = ( ~x29 & n12465 ) | ( ~x29 & n12470 ) | ( n12465 & n12470 ) ;
  assign n12472 = ( n12465 & n12470 ) | ( n12465 & ~n12471 ) | ( n12470 & ~n12471 ) ;
  assign n12473 = ( x29 & n12471 ) | ( x29 & ~n12472 ) | ( n12471 & ~n12472 ) ;
  assign n12474 = n3700 & ~n10003 ;
  assign n12475 = n3802 & ~n10001 ;
  assign n12476 = n12474 | n12475 ;
  assign n12477 = n3799 & ~n9999 ;
  assign n12478 = ( n3799 & n12476 ) | ( n3799 & ~n12477 ) | ( n12476 & ~n12477 ) ;
  assign n12479 = n3800 & n11868 ;
  assign n12480 = n12478 | n12479 ;
  assign n12481 = n3697 & ~n10003 ;
  assign n12482 = x29 & n12481 ;
  assign n12483 = ( n3800 & n11804 ) | ( n3800 & n11805 ) | ( n11804 & n11805 ) ;
  assign n12484 = n3802 | n10003 ;
  assign n12485 = n3799 & ~n10001 ;
  assign n12486 = ( ~n10003 & n12484 ) | ( ~n10003 & n12485 ) | ( n12484 & n12485 ) ;
  assign n12487 = ( ~n12482 & n12483 ) | ( ~n12482 & n12486 ) | ( n12483 & n12486 ) ;
  assign n12488 = ( x29 & n12482 ) | ( x29 & n12487 ) | ( n12482 & n12487 ) ;
  assign n12489 = n12480 | n12488 ;
  assign n12490 = x29 & ~n12489 ;
  assign n12491 = ( n12464 & n12473 ) | ( n12464 & n12490 ) | ( n12473 & n12490 ) ;
  assign n12492 = n3800 & n11934 ;
  assign n12493 = n3799 & n9995 ;
  assign n12494 = n3700 & n9999 ;
  assign n12495 = n3802 & ~n9997 ;
  assign n12496 = n12494 | n12495 ;
  assign n12497 = ( ~n12492 & n12493 ) | ( ~n12492 & n12496 ) | ( n12493 & n12496 ) ;
  assign n12498 = ( ~x29 & n12492 ) | ( ~x29 & n12497 ) | ( n12492 & n12497 ) ;
  assign n12499 = ( n12492 & n12497 ) | ( n12492 & ~n12498 ) | ( n12497 & ~n12498 ) ;
  assign n12500 = ( x29 & n12498 ) | ( x29 & ~n12499 ) | ( n12498 & ~n12499 ) ;
  assign n12501 = n11809 & n11842 ;
  assign n12502 = ( n11842 & n11843 ) | ( n11842 & ~n12501 ) | ( n11843 & ~n12501 ) ;
  assign n12503 = ( n12491 & n12500 ) | ( n12491 & ~n12502 ) | ( n12500 & ~n12502 ) ;
  assign n12504 = n3800 & ~n11971 ;
  assign n12505 = n3799 & n9993 ;
  assign n12506 = n3700 & ~n9997 ;
  assign n12507 = n3802 & n9995 ;
  assign n12508 = n12506 | n12507 ;
  assign n12509 = ( ~n12504 & n12505 ) | ( ~n12504 & n12508 ) | ( n12505 & n12508 ) ;
  assign n12510 = ( ~x29 & n12504 ) | ( ~x29 & n12509 ) | ( n12504 & n12509 ) ;
  assign n12511 = ( n12504 & n12509 ) | ( n12504 & ~n12510 ) | ( n12509 & ~n12510 ) ;
  assign n12512 = ( x29 & n12510 ) | ( x29 & ~n12511 ) | ( n12510 & ~n12511 ) ;
  assign n12513 = ( ~n11843 & n11861 ) | ( ~n11843 & n11870 ) | ( n11861 & n11870 ) ;
  assign n12514 = ( ~n11870 & n11871 ) | ( ~n11870 & n12513 ) | ( n11871 & n12513 ) ;
  assign n12515 = ( n12503 & n12512 ) | ( n12503 & ~n12514 ) | ( n12512 & ~n12514 ) ;
  assign n12516 = n3800 & n12026 ;
  assign n12517 = n3799 & n9991 ;
  assign n12518 = n3700 & n9995 ;
  assign n12519 = n3802 & n9993 ;
  assign n12520 = n12518 | n12519 ;
  assign n12521 = ( ~n12516 & n12517 ) | ( ~n12516 & n12520 ) | ( n12517 & n12520 ) ;
  assign n12522 = ( ~x29 & n12516 ) | ( ~x29 & n12521 ) | ( n12516 & n12521 ) ;
  assign n12523 = ( n12516 & n12521 ) | ( n12516 & ~n12522 ) | ( n12521 & ~n12522 ) ;
  assign n12524 = ( x29 & n12522 ) | ( x29 & ~n12523 ) | ( n12522 & ~n12523 ) ;
  assign n12525 = ( ~n11871 & n11885 ) | ( ~n11871 & n11894 ) | ( n11885 & n11894 ) ;
  assign n12526 = ( n11871 & ~n11895 ) | ( n11871 & n12525 ) | ( ~n11895 & n12525 ) ;
  assign n12527 = ( n12515 & n12524 ) | ( n12515 & n12526 ) | ( n12524 & n12526 ) ;
  assign n12528 = n3800 & n12050 ;
  assign n12529 = n3799 & n9989 ;
  assign n12530 = n3700 & n9993 ;
  assign n12531 = n3802 & n9991 ;
  assign n12532 = n12530 | n12531 ;
  assign n12533 = ( ~n12528 & n12529 ) | ( ~n12528 & n12532 ) | ( n12529 & n12532 ) ;
  assign n12534 = ( ~x29 & n12528 ) | ( ~x29 & n12533 ) | ( n12528 & n12533 ) ;
  assign n12535 = ( n12528 & n12533 ) | ( n12528 & ~n12534 ) | ( n12533 & ~n12534 ) ;
  assign n12536 = ( x29 & n12534 ) | ( x29 & ~n12535 ) | ( n12534 & ~n12535 ) ;
  assign n12537 = ( ~n11895 & n11927 ) | ( ~n11895 & n11936 ) | ( n11927 & n11936 ) ;
  assign n12538 = ( ~n11936 & n11937 ) | ( ~n11936 & n12537 ) | ( n11937 & n12537 ) ;
  assign n12539 = ( n12527 & n12536 ) | ( n12527 & ~n12538 ) | ( n12536 & ~n12538 ) ;
  assign n12540 = n3800 & ~n12074 ;
  assign n12541 = n3799 & ~n9987 ;
  assign n12542 = n3700 & n9991 ;
  assign n12543 = n3802 & n9989 ;
  assign n12544 = n12542 | n12543 ;
  assign n12545 = ( ~n12540 & n12541 ) | ( ~n12540 & n12544 ) | ( n12541 & n12544 ) ;
  assign n12546 = ( ~x29 & n12540 ) | ( ~x29 & n12545 ) | ( n12540 & n12545 ) ;
  assign n12547 = ( n12540 & n12545 ) | ( n12540 & ~n12546 ) | ( n12545 & ~n12546 ) ;
  assign n12548 = ( x29 & n12546 ) | ( x29 & ~n12547 ) | ( n12546 & ~n12547 ) ;
  assign n12549 = ( ~n11937 & n11964 ) | ( ~n11937 & n11973 ) | ( n11964 & n11973 ) ;
  assign n12550 = ( ~n11973 & n11974 ) | ( ~n11973 & n12549 ) | ( n11974 & n12549 ) ;
  assign n12551 = ( n12539 & n12548 ) | ( n12539 & ~n12550 ) | ( n12548 & ~n12550 ) ;
  assign n12552 = n3800 & ~n12099 ;
  assign n12553 = n3799 & n9985 ;
  assign n12554 = n3700 & n9989 ;
  assign n12555 = n3802 & ~n9987 ;
  assign n12556 = n12554 | n12555 ;
  assign n12557 = ( ~n12552 & n12553 ) | ( ~n12552 & n12556 ) | ( n12553 & n12556 ) ;
  assign n12558 = ( ~x29 & n12552 ) | ( ~x29 & n12557 ) | ( n12552 & n12557 ) ;
  assign n12559 = ( n12552 & n12557 ) | ( n12552 & ~n12558 ) | ( n12557 & ~n12558 ) ;
  assign n12560 = ( x29 & n12558 ) | ( x29 & ~n12559 ) | ( n12558 & ~n12559 ) ;
  assign n12561 = ( ~n11974 & n12019 ) | ( ~n11974 & n12028 ) | ( n12019 & n12028 ) ;
  assign n12562 = ( n11974 & ~n12029 ) | ( n11974 & n12561 ) | ( ~n12029 & n12561 ) ;
  assign n12563 = ( n12551 & n12560 ) | ( n12551 & n12562 ) | ( n12560 & n12562 ) ;
  assign n12564 = n3800 & ~n12129 ;
  assign n12565 = n3799 & ~n9983 ;
  assign n12566 = n3700 & ~n9987 ;
  assign n12567 = n3802 & n9985 ;
  assign n12568 = n12566 | n12567 ;
  assign n12569 = ( ~n12564 & n12565 ) | ( ~n12564 & n12568 ) | ( n12565 & n12568 ) ;
  assign n12570 = ( ~x29 & n12564 ) | ( ~x29 & n12569 ) | ( n12564 & n12569 ) ;
  assign n12571 = ( n12564 & n12569 ) | ( n12564 & ~n12570 ) | ( n12569 & ~n12570 ) ;
  assign n12572 = ( x29 & n12570 ) | ( x29 & ~n12571 ) | ( n12570 & ~n12571 ) ;
  assign n12573 = ( ~n12029 & n12043 ) | ( ~n12029 & n12052 ) | ( n12043 & n12052 ) ;
  assign n12574 = ( n12029 & ~n12053 ) | ( n12029 & n12573 ) | ( ~n12053 & n12573 ) ;
  assign n12575 = ( n12563 & n12572 ) | ( n12563 & n12574 ) | ( n12572 & n12574 ) ;
  assign n12576 = n3800 & ~n11561 ;
  assign n12577 = n3799 & n9981 ;
  assign n12578 = n3700 & n9985 ;
  assign n12579 = n3802 & ~n9983 ;
  assign n12580 = n12578 | n12579 ;
  assign n12581 = ( ~n12576 & n12577 ) | ( ~n12576 & n12580 ) | ( n12577 & n12580 ) ;
  assign n12582 = ( ~x29 & n12576 ) | ( ~x29 & n12581 ) | ( n12576 & n12581 ) ;
  assign n12583 = ( n12576 & n12581 ) | ( n12576 & ~n12582 ) | ( n12581 & ~n12582 ) ;
  assign n12584 = ( x29 & n12582 ) | ( x29 & ~n12583 ) | ( n12582 & ~n12583 ) ;
  assign n12585 = ( ~n12053 & n12067 ) | ( ~n12053 & n12076 ) | ( n12067 & n12076 ) ;
  assign n12586 = ( n12053 & ~n12077 ) | ( n12053 & n12585 ) | ( ~n12077 & n12585 ) ;
  assign n12587 = ( n12575 & n12584 ) | ( n12575 & n12586 ) | ( n12584 & n12586 ) ;
  assign n12588 = n3800 & n12153 ;
  assign n12589 = n3799 & n9979 ;
  assign n12590 = n3700 & ~n9983 ;
  assign n12591 = n3802 & n9981 ;
  assign n12592 = n12590 | n12591 ;
  assign n12593 = ( ~n12588 & n12589 ) | ( ~n12588 & n12592 ) | ( n12589 & n12592 ) ;
  assign n12594 = ( ~x29 & n12588 ) | ( ~x29 & n12593 ) | ( n12588 & n12593 ) ;
  assign n12595 = ( n12588 & n12593 ) | ( n12588 & ~n12594 ) | ( n12593 & ~n12594 ) ;
  assign n12596 = ( x29 & n12594 ) | ( x29 & ~n12595 ) | ( n12594 & ~n12595 ) ;
  assign n12597 = ( ~n12077 & n12092 ) | ( ~n12077 & n12101 ) | ( n12092 & n12101 ) ;
  assign n12598 = ( n12077 & ~n12102 ) | ( n12077 & n12597 ) | ( ~n12102 & n12597 ) ;
  assign n12599 = ( n12587 & n12596 ) | ( n12587 & n12598 ) | ( n12596 & n12598 ) ;
  assign n12600 = n3800 & n12165 ;
  assign n12601 = n3799 & n9977 ;
  assign n12602 = n3700 & n9981 ;
  assign n12603 = n3802 & n9979 ;
  assign n12604 = n12602 | n12603 ;
  assign n12605 = ( ~n12600 & n12601 ) | ( ~n12600 & n12604 ) | ( n12601 & n12604 ) ;
  assign n12606 = ( ~x29 & n12600 ) | ( ~x29 & n12605 ) | ( n12600 & n12605 ) ;
  assign n12607 = ( n12600 & n12605 ) | ( n12600 & ~n12606 ) | ( n12605 & ~n12606 ) ;
  assign n12608 = ( x29 & n12606 ) | ( x29 & ~n12607 ) | ( n12606 & ~n12607 ) ;
  assign n12609 = ( ~n12102 & n12122 ) | ( ~n12102 & n12131 ) | ( n12122 & n12131 ) ;
  assign n12610 = ( n12102 & ~n12132 ) | ( n12102 & n12609 ) | ( ~n12132 & n12609 ) ;
  assign n12611 = ( n12599 & n12608 ) | ( n12599 & n12610 ) | ( n12608 & n12610 ) ;
  assign n12612 = ( ~n12132 & n12134 ) | ( ~n12132 & n12143 ) | ( n12134 & n12143 ) ;
  assign n12613 = ( ~n12143 & n12144 ) | ( ~n12143 & n12612 ) | ( n12144 & n12612 ) ;
  assign n12614 = n4202 & n11428 ;
  assign n12615 = n4201 & n9969 ;
  assign n12616 = n4200 & n9973 ;
  assign n12617 = n4345 & n9971 ;
  assign n12618 = n12616 | n12617 ;
  assign n12619 = ( ~n12614 & n12615 ) | ( ~n12614 & n12618 ) | ( n12615 & n12618 ) ;
  assign n12620 = ( ~x26 & n12614 ) | ( ~x26 & n12619 ) | ( n12614 & n12619 ) ;
  assign n12621 = ( n12614 & n12619 ) | ( n12614 & ~n12620 ) | ( n12619 & ~n12620 ) ;
  assign n12622 = ( x26 & n12620 ) | ( x26 & ~n12621 ) | ( n12620 & ~n12621 ) ;
  assign n12623 = ( n12611 & ~n12613 ) | ( n12611 & n12622 ) | ( ~n12613 & n12622 ) ;
  assign n12624 = ( n12366 & ~n12375 ) | ( n12366 & n12384 ) | ( ~n12375 & n12384 ) ;
  assign n12625 = ( n12375 & ~n12385 ) | ( n12375 & n12624 ) | ( ~n12385 & n12624 ) ;
  assign n12626 = n4713 & ~n10929 ;
  assign n12627 = n4712 & n9961 ;
  assign n12628 = n4709 & n9965 ;
  assign n12629 = n4792 & ~n9963 ;
  assign n12630 = n12628 | n12629 ;
  assign n12631 = ( ~n12626 & n12627 ) | ( ~n12626 & n12630 ) | ( n12627 & n12630 ) ;
  assign n12632 = ( ~x23 & n12626 ) | ( ~x23 & n12631 ) | ( n12626 & n12631 ) ;
  assign n12633 = ( n12626 & n12631 ) | ( n12626 & ~n12632 ) | ( n12631 & ~n12632 ) ;
  assign n12634 = ( x23 & n12632 ) | ( x23 & ~n12633 ) | ( n12632 & ~n12633 ) ;
  assign n12635 = ( n12623 & n12625 ) | ( n12623 & n12634 ) | ( n12625 & n12634 ) ;
  assign n12636 = ( ~n12385 & n12387 ) | ( ~n12385 & n12396 ) | ( n12387 & n12396 ) ;
  assign n12637 = ( ~n12396 & n12397 ) | ( ~n12396 & n12636 ) | ( n12397 & n12636 ) ;
  assign n12638 = n4974 & ~n10750 ;
  assign n12639 = n5398 & ~n9953 ;
  assign n12640 = n4973 & ~n9957 ;
  assign n12641 = n4972 & n9955 ;
  assign n12642 = n12640 | n12641 ;
  assign n12643 = ( ~n12638 & n12639 ) | ( ~n12638 & n12642 ) | ( n12639 & n12642 ) ;
  assign n12644 = ( ~x20 & n12638 ) | ( ~x20 & n12643 ) | ( n12638 & n12643 ) ;
  assign n12645 = ( n12638 & n12643 ) | ( n12638 & ~n12644 ) | ( n12643 & ~n12644 ) ;
  assign n12646 = ( x20 & n12644 ) | ( x20 & ~n12645 ) | ( n12644 & ~n12645 ) ;
  assign n12647 = ( n12635 & ~n12637 ) | ( n12635 & n12646 ) | ( ~n12637 & n12646 ) ;
  assign n12648 = ( ~n12397 & n12399 ) | ( ~n12397 & n12408 ) | ( n12399 & n12408 ) ;
  assign n12649 = ( ~n12408 & n12409 ) | ( ~n12408 & n12648 ) | ( n12409 & n12648 ) ;
  assign n12650 = n4974 & ~n10652 ;
  assign n12651 = n5398 & n9951 ;
  assign n12652 = n4973 & n9955 ;
  assign n12653 = n4972 & ~n9953 ;
  assign n12654 = n12652 | n12653 ;
  assign n12655 = ( ~n12650 & n12651 ) | ( ~n12650 & n12654 ) | ( n12651 & n12654 ) ;
  assign n12656 = ( ~x20 & n12650 ) | ( ~x20 & n12655 ) | ( n12650 & n12655 ) ;
  assign n12657 = ( n12650 & n12655 ) | ( n12650 & ~n12656 ) | ( n12655 & ~n12656 ) ;
  assign n12658 = ( x20 & n12656 ) | ( x20 & ~n12657 ) | ( n12656 & ~n12657 ) ;
  assign n12659 = ( n12647 & ~n12649 ) | ( n12647 & n12658 ) | ( ~n12649 & n12658 ) ;
  assign n12660 = ( n12409 & ~n12411 ) | ( n12409 & n12420 ) | ( ~n12411 & n12420 ) ;
  assign n12661 = ( n12411 & ~n12421 ) | ( n12411 & n12660 ) | ( ~n12421 & n12660 ) ;
  assign n12662 = n5508 & n10271 ;
  assign n12663 = n5507 & n9943 ;
  assign n12664 = n5504 & n9947 ;
  assign n12665 = n5666 & n9945 ;
  assign n12666 = n12664 | n12665 ;
  assign n12667 = ( ~n12662 & n12663 ) | ( ~n12662 & n12666 ) | ( n12663 & n12666 ) ;
  assign n12668 = ( ~x17 & n12662 ) | ( ~x17 & n12667 ) | ( n12662 & n12667 ) ;
  assign n12669 = ( n12662 & n12667 ) | ( n12662 & ~n12668 ) | ( n12667 & ~n12668 ) ;
  assign n12670 = ( x17 & n12668 ) | ( x17 & ~n12669 ) | ( n12668 & ~n12669 ) ;
  assign n12671 = ( n12659 & n12661 ) | ( n12659 & n12670 ) | ( n12661 & n12670 ) ;
  assign n12672 = ( ~n12421 & n12423 ) | ( ~n12421 & n12432 ) | ( n12423 & n12432 ) ;
  assign n12673 = ( ~n12432 & n12433 ) | ( ~n12432 & n12672 ) | ( n12433 & n12672 ) ;
  assign n12674 = n5966 & n10040 ;
  assign n12675 = n6464 & ~n9937 ;
  assign n12676 = n5970 & ~n9883 ;
  assign n12677 = n5969 & n9916 ;
  assign n12678 = n12676 | n12677 ;
  assign n12679 = ( ~n12674 & n12675 ) | ( ~n12674 & n12678 ) | ( n12675 & n12678 ) ;
  assign n12680 = ( ~x14 & n12674 ) | ( ~x14 & n12679 ) | ( n12674 & n12679 ) ;
  assign n12681 = ( n12674 & n12679 ) | ( n12674 & ~n12680 ) | ( n12679 & ~n12680 ) ;
  assign n12682 = ( x14 & n12680 ) | ( x14 & ~n12681 ) | ( n12680 & ~n12681 ) ;
  assign n12683 = ( n12671 & ~n12673 ) | ( n12671 & n12682 ) | ( ~n12673 & n12682 ) ;
  assign n12684 = ( ~n12433 & n12435 ) | ( ~n12433 & n12444 ) | ( n12435 & n12444 ) ;
  assign n12685 = ( ~n12444 & n12445 ) | ( ~n12444 & n12684 ) | ( n12445 & n12684 ) ;
  assign n12686 = n5966 & ~n10064 ;
  assign n12687 = n6464 & ~n10057 ;
  assign n12688 = n5970 & n9916 ;
  assign n12689 = n5969 & ~n9937 ;
  assign n12690 = n12688 | n12689 ;
  assign n12691 = ( ~n12686 & n12687 ) | ( ~n12686 & n12690 ) | ( n12687 & n12690 ) ;
  assign n12692 = ( ~x14 & n12686 ) | ( ~x14 & n12691 ) | ( n12686 & n12691 ) ;
  assign n12693 = ( n12686 & n12691 ) | ( n12686 & ~n12692 ) | ( n12691 & ~n12692 ) ;
  assign n12694 = ( x14 & n12692 ) | ( x14 & ~n12693 ) | ( n12692 & ~n12693 ) ;
  assign n12695 = ( n12683 & ~n12685 ) | ( n12683 & n12694 ) | ( ~n12685 & n12694 ) ;
  assign n12696 = ( ~n12445 & n12447 ) | ( ~n12445 & n12456 ) | ( n12447 & n12456 ) ;
  assign n12697 = ( ~n12456 & n12457 ) | ( ~n12456 & n12696 ) | ( n12457 & n12696 ) ;
  assign n12698 = ~n6588 & n10346 ;
  assign n12699 = ( n10346 & n10984 ) | ( n10346 & ~n12698 ) | ( n10984 & ~n12698 ) ;
  assign n12700 = ( ~x11 & n6584 ) | ( ~x11 & n12699 ) | ( n6584 & n12699 ) ;
  assign n12701 = ( n6584 & n12699 ) | ( n6584 & ~n12700 ) | ( n12699 & ~n12700 ) ;
  assign n12702 = ( x11 & n12700 ) | ( x11 & ~n12701 ) | ( n12700 & ~n12701 ) ;
  assign n12703 = ( n12695 & ~n12697 ) | ( n12695 & n12702 ) | ( ~n12697 & n12702 ) ;
  assign n12704 = n4202 & n11892 ;
  assign n12705 = n4201 & ~n9997 ;
  assign n12706 = n4200 & ~n10001 ;
  assign n12707 = n4345 & n9999 ;
  assign n12708 = n12706 | n12707 ;
  assign n12709 = ( ~n12704 & n12705 ) | ( ~n12704 & n12708 ) | ( n12705 & n12708 ) ;
  assign n12710 = ( ~x26 & n12704 ) | ( ~x26 & n12709 ) | ( n12704 & n12709 ) ;
  assign n12711 = ( n12704 & n12709 ) | ( n12704 & ~n12710 ) | ( n12709 & ~n12710 ) ;
  assign n12712 = ( x26 & n12710 ) | ( x26 & ~n12711 ) | ( n12710 & ~n12711 ) ;
  assign n12713 = n4200 & ~n10003 ;
  assign n12714 = n4345 & ~n10001 ;
  assign n12715 = n12713 | n12714 ;
  assign n12716 = n4201 & ~n9999 ;
  assign n12717 = ( n4201 & n12715 ) | ( n4201 & ~n12716 ) | ( n12715 & ~n12716 ) ;
  assign n12718 = n4202 & n11868 ;
  assign n12719 = n12717 | n12718 ;
  assign n12720 = n4195 & ~n10003 ;
  assign n12721 = x26 & n12720 ;
  assign n12722 = ( n4202 & n11804 ) | ( n4202 & n11805 ) | ( n11804 & n11805 ) ;
  assign n12723 = n4345 & ~n10003 ;
  assign n12724 = n4201 & ~n10001 ;
  assign n12725 = n12723 | n12724 ;
  assign n12726 = ( ~n12721 & n12722 ) | ( ~n12721 & n12725 ) | ( n12722 & n12725 ) ;
  assign n12727 = ( x26 & n12721 ) | ( x26 & n12726 ) | ( n12721 & n12726 ) ;
  assign n12728 = n12719 | n12727 ;
  assign n12729 = x26 & ~n12728 ;
  assign n12730 = ( n12481 & n12712 ) | ( n12481 & n12729 ) | ( n12712 & n12729 ) ;
  assign n12731 = n4202 & n11934 ;
  assign n12732 = n4201 & n9995 ;
  assign n12733 = n4200 & n9999 ;
  assign n12734 = n4345 & ~n9997 ;
  assign n12735 = n12733 | n12734 ;
  assign n12736 = ( ~n12731 & n12732 ) | ( ~n12731 & n12735 ) | ( n12732 & n12735 ) ;
  assign n12737 = ( ~x26 & n12731 ) | ( ~x26 & n12736 ) | ( n12731 & n12736 ) ;
  assign n12738 = ( n12731 & n12736 ) | ( n12731 & ~n12737 ) | ( n12736 & ~n12737 ) ;
  assign n12739 = ( x26 & n12737 ) | ( x26 & ~n12738 ) | ( n12737 & ~n12738 ) ;
  assign n12740 = ( n12483 & n12486 ) | ( n12483 & ~n12487 ) | ( n12486 & ~n12487 ) ;
  assign n12741 = ( n12482 & n12487 ) | ( n12482 & ~n12740 ) | ( n12487 & ~n12740 ) ;
  assign n12742 = ( n12730 & n12739 ) | ( n12730 & n12741 ) | ( n12739 & n12741 ) ;
  assign n12743 = n4202 & ~n11971 ;
  assign n12744 = n4201 & n9993 ;
  assign n12745 = n4200 & ~n9997 ;
  assign n12746 = n4345 & n9995 ;
  assign n12747 = n12745 | n12746 ;
  assign n12748 = ( ~n12743 & n12744 ) | ( ~n12743 & n12747 ) | ( n12744 & n12747 ) ;
  assign n12749 = ( ~x26 & n12743 ) | ( ~x26 & n12748 ) | ( n12743 & n12748 ) ;
  assign n12750 = ( n12743 & n12748 ) | ( n12743 & ~n12749 ) | ( n12748 & ~n12749 ) ;
  assign n12751 = ( x26 & n12749 ) | ( x26 & ~n12750 ) | ( n12749 & ~n12750 ) ;
  assign n12752 = ( n12480 & n12488 ) | ( n12480 & ~n12489 ) | ( n12488 & ~n12489 ) ;
  assign n12753 = n12489 & ~n12752 ;
  assign n12754 = ( n12742 & n12751 ) | ( n12742 & n12753 ) | ( n12751 & n12753 ) ;
  assign n12755 = n4202 & n12026 ;
  assign n12756 = n4201 & n9991 ;
  assign n12757 = n4200 & n9995 ;
  assign n12758 = n4345 & n9993 ;
  assign n12759 = n12757 | n12758 ;
  assign n12760 = ( ~n12755 & n12756 ) | ( ~n12755 & n12759 ) | ( n12756 & n12759 ) ;
  assign n12761 = ( ~x26 & n12755 ) | ( ~x26 & n12760 ) | ( n12755 & n12760 ) ;
  assign n12762 = ( n12755 & n12760 ) | ( n12755 & ~n12761 ) | ( n12760 & ~n12761 ) ;
  assign n12763 = ( x26 & n12761 ) | ( x26 & ~n12762 ) | ( n12761 & ~n12762 ) ;
  assign n12764 = ( n12464 & n12473 ) | ( n12464 & ~n12490 ) | ( n12473 & ~n12490 ) ;
  assign n12765 = ( n12490 & ~n12491 ) | ( n12490 & n12764 ) | ( ~n12491 & n12764 ) ;
  assign n12766 = ( n12754 & n12763 ) | ( n12754 & n12765 ) | ( n12763 & n12765 ) ;
  assign n12767 = n4202 & n12050 ;
  assign n12768 = n4201 & n9989 ;
  assign n12769 = n4200 & n9993 ;
  assign n12770 = n4345 & n9991 ;
  assign n12771 = n12769 | n12770 ;
  assign n12772 = ( ~n12767 & n12768 ) | ( ~n12767 & n12771 ) | ( n12768 & n12771 ) ;
  assign n12773 = ( ~x26 & n12767 ) | ( ~x26 & n12772 ) | ( n12767 & n12772 ) ;
  assign n12774 = ( n12767 & n12772 ) | ( n12767 & ~n12773 ) | ( n12772 & ~n12773 ) ;
  assign n12775 = ( x26 & n12773 ) | ( x26 & ~n12774 ) | ( n12773 & ~n12774 ) ;
  assign n12776 = ( n12491 & ~n12500 ) | ( n12491 & n12502 ) | ( ~n12500 & n12502 ) ;
  assign n12777 = ( ~n12491 & n12503 ) | ( ~n12491 & n12776 ) | ( n12503 & n12776 ) ;
  assign n12778 = ( n12766 & n12775 ) | ( n12766 & ~n12777 ) | ( n12775 & ~n12777 ) ;
  assign n12779 = ( n12503 & ~n12512 ) | ( n12503 & n12514 ) | ( ~n12512 & n12514 ) ;
  assign n12780 = ( ~n12503 & n12515 ) | ( ~n12503 & n12779 ) | ( n12515 & n12779 ) ;
  assign n12781 = n4202 & ~n12074 ;
  assign n12782 = n4201 & ~n9987 ;
  assign n12783 = n4200 & n9991 ;
  assign n12784 = n4345 & n9989 ;
  assign n12785 = n12783 | n12784 ;
  assign n12786 = ( ~n12781 & n12782 ) | ( ~n12781 & n12785 ) | ( n12782 & n12785 ) ;
  assign n12787 = ( ~x26 & n12781 ) | ( ~x26 & n12786 ) | ( n12781 & n12786 ) ;
  assign n12788 = ( n12781 & n12786 ) | ( n12781 & ~n12787 ) | ( n12786 & ~n12787 ) ;
  assign n12789 = ( x26 & n12787 ) | ( x26 & ~n12788 ) | ( n12787 & ~n12788 ) ;
  assign n12790 = ( n12778 & ~n12780 ) | ( n12778 & n12789 ) | ( ~n12780 & n12789 ) ;
  assign n12791 = ( ~n12515 & n12524 ) | ( ~n12515 & n12526 ) | ( n12524 & n12526 ) ;
  assign n12792 = ( n12515 & ~n12527 ) | ( n12515 & n12791 ) | ( ~n12527 & n12791 ) ;
  assign n12793 = n4202 & ~n12099 ;
  assign n12794 = n4201 & n9985 ;
  assign n12795 = n4200 & n9989 ;
  assign n12796 = n4345 & ~n9987 ;
  assign n12797 = n12795 | n12796 ;
  assign n12798 = ( ~n12793 & n12794 ) | ( ~n12793 & n12797 ) | ( n12794 & n12797 ) ;
  assign n12799 = ( ~x26 & n12793 ) | ( ~x26 & n12798 ) | ( n12793 & n12798 ) ;
  assign n12800 = ( n12793 & n12798 ) | ( n12793 & ~n12799 ) | ( n12798 & ~n12799 ) ;
  assign n12801 = ( x26 & n12799 ) | ( x26 & ~n12800 ) | ( n12799 & ~n12800 ) ;
  assign n12802 = ( n12790 & n12792 ) | ( n12790 & n12801 ) | ( n12792 & n12801 ) ;
  assign n12803 = ( n12527 & ~n12536 ) | ( n12527 & n12538 ) | ( ~n12536 & n12538 ) ;
  assign n12804 = ( ~n12527 & n12539 ) | ( ~n12527 & n12803 ) | ( n12539 & n12803 ) ;
  assign n12805 = n4202 & ~n12129 ;
  assign n12806 = n4201 & ~n9983 ;
  assign n12807 = n4200 & ~n9987 ;
  assign n12808 = n4345 & n9985 ;
  assign n12809 = n12807 | n12808 ;
  assign n12810 = ( ~n12805 & n12806 ) | ( ~n12805 & n12809 ) | ( n12806 & n12809 ) ;
  assign n12811 = ( ~x26 & n12805 ) | ( ~x26 & n12810 ) | ( n12805 & n12810 ) ;
  assign n12812 = ( n12805 & n12810 ) | ( n12805 & ~n12811 ) | ( n12810 & ~n12811 ) ;
  assign n12813 = ( x26 & n12811 ) | ( x26 & ~n12812 ) | ( n12811 & ~n12812 ) ;
  assign n12814 = ( n12802 & ~n12804 ) | ( n12802 & n12813 ) | ( ~n12804 & n12813 ) ;
  assign n12815 = ( n12539 & ~n12548 ) | ( n12539 & n12550 ) | ( ~n12548 & n12550 ) ;
  assign n12816 = ( ~n12539 & n12551 ) | ( ~n12539 & n12815 ) | ( n12551 & n12815 ) ;
  assign n12817 = n4202 & ~n11561 ;
  assign n12818 = n4201 & n9981 ;
  assign n12819 = n4200 & n9985 ;
  assign n12820 = n4345 & ~n9983 ;
  assign n12821 = n12819 | n12820 ;
  assign n12822 = ( ~n12817 & n12818 ) | ( ~n12817 & n12821 ) | ( n12818 & n12821 ) ;
  assign n12823 = ( ~x26 & n12817 ) | ( ~x26 & n12822 ) | ( n12817 & n12822 ) ;
  assign n12824 = ( n12817 & n12822 ) | ( n12817 & ~n12823 ) | ( n12822 & ~n12823 ) ;
  assign n12825 = ( x26 & n12823 ) | ( x26 & ~n12824 ) | ( n12823 & ~n12824 ) ;
  assign n12826 = ( n12814 & ~n12816 ) | ( n12814 & n12825 ) | ( ~n12816 & n12825 ) ;
  assign n12827 = ( ~n12551 & n12560 ) | ( ~n12551 & n12562 ) | ( n12560 & n12562 ) ;
  assign n12828 = ( n12551 & ~n12563 ) | ( n12551 & n12827 ) | ( ~n12563 & n12827 ) ;
  assign n12829 = n4202 & n12153 ;
  assign n12830 = n4201 & n9979 ;
  assign n12831 = n4200 & ~n9983 ;
  assign n12832 = n4345 & n9981 ;
  assign n12833 = n12831 | n12832 ;
  assign n12834 = ( ~n12829 & n12830 ) | ( ~n12829 & n12833 ) | ( n12830 & n12833 ) ;
  assign n12835 = ( ~x26 & n12829 ) | ( ~x26 & n12834 ) | ( n12829 & n12834 ) ;
  assign n12836 = ( n12829 & n12834 ) | ( n12829 & ~n12835 ) | ( n12834 & ~n12835 ) ;
  assign n12837 = ( x26 & n12835 ) | ( x26 & ~n12836 ) | ( n12835 & ~n12836 ) ;
  assign n12838 = ( n12826 & n12828 ) | ( n12826 & n12837 ) | ( n12828 & n12837 ) ;
  assign n12839 = ( ~n12563 & n12572 ) | ( ~n12563 & n12574 ) | ( n12572 & n12574 ) ;
  assign n12840 = ( n12563 & ~n12575 ) | ( n12563 & n12839 ) | ( ~n12575 & n12839 ) ;
  assign n12841 = n4202 & n12165 ;
  assign n12842 = n4201 & n9977 ;
  assign n12843 = n4200 & n9981 ;
  assign n12844 = n4345 & n9979 ;
  assign n12845 = n12843 | n12844 ;
  assign n12846 = ( ~n12841 & n12842 ) | ( ~n12841 & n12845 ) | ( n12842 & n12845 ) ;
  assign n12847 = ( ~x26 & n12841 ) | ( ~x26 & n12846 ) | ( n12841 & n12846 ) ;
  assign n12848 = ( n12841 & n12846 ) | ( n12841 & ~n12847 ) | ( n12846 & ~n12847 ) ;
  assign n12849 = ( x26 & n12847 ) | ( x26 & ~n12848 ) | ( n12847 & ~n12848 ) ;
  assign n12850 = ( n12838 & n12840 ) | ( n12838 & n12849 ) | ( n12840 & n12849 ) ;
  assign n12851 = ( ~n12575 & n12584 ) | ( ~n12575 & n12586 ) | ( n12584 & n12586 ) ;
  assign n12852 = ( n12575 & ~n12587 ) | ( n12575 & n12851 ) | ( ~n12587 & n12851 ) ;
  assign n12853 = n4202 & n11606 ;
  assign n12854 = n4201 & n9975 ;
  assign n12855 = n4200 & n9979 ;
  assign n12856 = n4345 & n9977 ;
  assign n12857 = n12855 | n12856 ;
  assign n12858 = ( ~n12853 & n12854 ) | ( ~n12853 & n12857 ) | ( n12854 & n12857 ) ;
  assign n12859 = ( ~x26 & n12853 ) | ( ~x26 & n12858 ) | ( n12853 & n12858 ) ;
  assign n12860 = ( n12853 & n12858 ) | ( n12853 & ~n12859 ) | ( n12858 & ~n12859 ) ;
  assign n12861 = ( x26 & n12859 ) | ( x26 & ~n12860 ) | ( n12859 & ~n12860 ) ;
  assign n12862 = ( n12850 & n12852 ) | ( n12850 & n12861 ) | ( n12852 & n12861 ) ;
  assign n12863 = ( ~n12587 & n12596 ) | ( ~n12587 & n12598 ) | ( n12596 & n12598 ) ;
  assign n12864 = ( n12587 & ~n12599 ) | ( n12587 & n12863 ) | ( ~n12599 & n12863 ) ;
  assign n12865 = n4202 & n11400 ;
  assign n12866 = n4201 & n9973 ;
  assign n12867 = n4200 & n9977 ;
  assign n12868 = n4345 & n9975 ;
  assign n12869 = n12867 | n12868 ;
  assign n12870 = ( ~n12865 & n12866 ) | ( ~n12865 & n12869 ) | ( n12866 & n12869 ) ;
  assign n12871 = ( ~x26 & n12865 ) | ( ~x26 & n12870 ) | ( n12865 & n12870 ) ;
  assign n12872 = ( n12865 & n12870 ) | ( n12865 & ~n12871 ) | ( n12870 & ~n12871 ) ;
  assign n12873 = ( x26 & n12871 ) | ( x26 & ~n12872 ) | ( n12871 & ~n12872 ) ;
  assign n12874 = ( n12862 & n12864 ) | ( n12862 & n12873 ) | ( n12864 & n12873 ) ;
  assign n12875 = ( ~n12599 & n12608 ) | ( ~n12599 & n12610 ) | ( n12608 & n12610 ) ;
  assign n12876 = ( n12599 & ~n12611 ) | ( n12599 & n12875 ) | ( ~n12611 & n12875 ) ;
  assign n12877 = n4202 & n11630 ;
  assign n12878 = n4201 & n9971 ;
  assign n12879 = n4200 & n9975 ;
  assign n12880 = n4345 & n9973 ;
  assign n12881 = n12879 | n12880 ;
  assign n12882 = ( ~n12877 & n12878 ) | ( ~n12877 & n12881 ) | ( n12878 & n12881 ) ;
  assign n12883 = ( ~x26 & n12877 ) | ( ~x26 & n12882 ) | ( n12877 & n12882 ) ;
  assign n12884 = ( n12877 & n12882 ) | ( n12877 & ~n12883 ) | ( n12882 & ~n12883 ) ;
  assign n12885 = ( x26 & n12883 ) | ( x26 & ~n12884 ) | ( n12883 & ~n12884 ) ;
  assign n12886 = ( n12874 & n12876 ) | ( n12874 & n12885 ) | ( n12876 & n12885 ) ;
  assign n12887 = ( ~n12611 & n12613 ) | ( ~n12611 & n12622 ) | ( n12613 & n12622 ) ;
  assign n12888 = ( ~n12622 & n12623 ) | ( ~n12622 & n12887 ) | ( n12623 & n12887 ) ;
  assign n12889 = n4713 & ~n11121 ;
  assign n12890 = n4712 & ~n9963 ;
  assign n12891 = n4709 & ~n9967 ;
  assign n12892 = n4792 & n9965 ;
  assign n12893 = n12891 | n12892 ;
  assign n12894 = ( ~n12889 & n12890 ) | ( ~n12889 & n12893 ) | ( n12890 & n12893 ) ;
  assign n12895 = ( ~x23 & n12889 ) | ( ~x23 & n12894 ) | ( n12889 & n12894 ) ;
  assign n12896 = ( n12889 & n12894 ) | ( n12889 & ~n12895 ) | ( n12894 & ~n12895 ) ;
  assign n12897 = ( x23 & n12895 ) | ( x23 & ~n12896 ) | ( n12895 & ~n12896 ) ;
  assign n12898 = ( n12886 & ~n12888 ) | ( n12886 & n12897 ) | ( ~n12888 & n12897 ) ;
  assign n12899 = ( ~n12623 & n12625 ) | ( ~n12623 & n12634 ) | ( n12625 & n12634 ) ;
  assign n12900 = ( n12623 & ~n12635 ) | ( n12623 & n12899 ) | ( ~n12635 & n12899 ) ;
  assign n12901 = n4974 & ~n10567 ;
  assign n12902 = n5398 & n9955 ;
  assign n12903 = n4973 & n9959 ;
  assign n12904 = n4972 & ~n9957 ;
  assign n12905 = n12903 | n12904 ;
  assign n12906 = ( ~n12901 & n12902 ) | ( ~n12901 & n12905 ) | ( n12902 & n12905 ) ;
  assign n12907 = ( ~x20 & n12901 ) | ( ~x20 & n12906 ) | ( n12901 & n12906 ) ;
  assign n12908 = ( n12901 & n12906 ) | ( n12901 & ~n12907 ) | ( n12906 & ~n12907 ) ;
  assign n12909 = ( x20 & n12907 ) | ( x20 & ~n12908 ) | ( n12907 & ~n12908 ) ;
  assign n12910 = ( n12898 & n12900 ) | ( n12898 & n12909 ) | ( n12900 & n12909 ) ;
  assign n12911 = ( ~n12635 & n12637 ) | ( ~n12635 & n12646 ) | ( n12637 & n12646 ) ;
  assign n12912 = ( ~n12646 & n12647 ) | ( ~n12646 & n12911 ) | ( n12647 & n12911 ) ;
  assign n12913 = n5508 & n10454 ;
  assign n12914 = n5507 & n9947 ;
  assign n12915 = n5504 & n9951 ;
  assign n12916 = n5666 & n9949 ;
  assign n12917 = n12915 | n12916 ;
  assign n12918 = ( ~n12913 & n12914 ) | ( ~n12913 & n12917 ) | ( n12914 & n12917 ) ;
  assign n12919 = ( ~x17 & n12913 ) | ( ~x17 & n12918 ) | ( n12913 & n12918 ) ;
  assign n12920 = ( n12913 & n12918 ) | ( n12913 & ~n12919 ) | ( n12918 & ~n12919 ) ;
  assign n12921 = ( x17 & n12919 ) | ( x17 & ~n12920 ) | ( n12919 & ~n12920 ) ;
  assign n12922 = ( n12910 & ~n12912 ) | ( n12910 & n12921 ) | ( ~n12912 & n12921 ) ;
  assign n12923 = ( ~n12647 & n12649 ) | ( ~n12647 & n12658 ) | ( n12649 & n12658 ) ;
  assign n12924 = ( ~n12658 & n12659 ) | ( ~n12658 & n12923 ) | ( n12659 & n12923 ) ;
  assign n12925 = n5508 & n10466 ;
  assign n12926 = n5507 & n9945 ;
  assign n12927 = n5504 & n9949 ;
  assign n12928 = n5666 & n9947 ;
  assign n12929 = n12927 | n12928 ;
  assign n12930 = ( ~n12925 & n12926 ) | ( ~n12925 & n12929 ) | ( n12926 & n12929 ) ;
  assign n12931 = ( ~x17 & n12925 ) | ( ~x17 & n12930 ) | ( n12925 & n12930 ) ;
  assign n12932 = ( n12925 & n12930 ) | ( n12925 & ~n12931 ) | ( n12930 & ~n12931 ) ;
  assign n12933 = ( x17 & n12931 ) | ( x17 & ~n12932 ) | ( n12931 & ~n12932 ) ;
  assign n12934 = ( n12922 & ~n12924 ) | ( n12922 & n12933 ) | ( ~n12924 & n12933 ) ;
  assign n12935 = ( n12659 & ~n12661 ) | ( n12659 & n12670 ) | ( ~n12661 & n12670 ) ;
  assign n12936 = ( n12661 & ~n12671 ) | ( n12661 & n12935 ) | ( ~n12671 & n12935 ) ;
  assign n12937 = n5966 & n10174 ;
  assign n12938 = n6464 & n9916 ;
  assign n12939 = n5969 | n9883 ;
  assign n12940 = n5970 & ~n9941 ;
  assign n12941 = ( ~n9883 & n12939 ) | ( ~n9883 & n12940 ) | ( n12939 & n12940 ) ;
  assign n12942 = ( ~n12937 & n12938 ) | ( ~n12937 & n12941 ) | ( n12938 & n12941 ) ;
  assign n12943 = ( ~x14 & n12937 ) | ( ~x14 & n12942 ) | ( n12937 & n12942 ) ;
  assign n12944 = ( n12937 & n12942 ) | ( n12937 & ~n12943 ) | ( n12942 & ~n12943 ) ;
  assign n12945 = ( x14 & n12943 ) | ( x14 & ~n12944 ) | ( n12943 & ~n12944 ) ;
  assign n12946 = ( n12934 & n12936 ) | ( n12934 & n12945 ) | ( n12936 & n12945 ) ;
  assign n12947 = ( ~n12671 & n12673 ) | ( ~n12671 & n12682 ) | ( n12673 & n12682 ) ;
  assign n12948 = ( ~n12682 & n12683 ) | ( ~n12682 & n12947 ) | ( n12683 & n12947 ) ;
  assign n12949 = n6584 & n10362 ;
  assign n12950 = n7022 & n10346 ;
  assign n12951 = n6588 & ~n10057 ;
  assign n12952 = n6587 & ~n10302 ;
  assign n12953 = n12951 | n12952 ;
  assign n12954 = ( ~n12949 & n12950 ) | ( ~n12949 & n12953 ) | ( n12950 & n12953 ) ;
  assign n12955 = ( ~x11 & n12949 ) | ( ~x11 & n12954 ) | ( n12949 & n12954 ) ;
  assign n12956 = ( n12949 & n12954 ) | ( n12949 & ~n12955 ) | ( n12954 & ~n12955 ) ;
  assign n12957 = ( x11 & n12955 ) | ( x11 & ~n12956 ) | ( n12955 & ~n12956 ) ;
  assign n12958 = ( n12946 & ~n12948 ) | ( n12946 & n12957 ) | ( ~n12948 & n12957 ) ;
  assign n12959 = n6584 & n10348 ;
  assign n12960 = n6587 & n10346 ;
  assign n12961 = n6588 & ~n10302 ;
  assign n12962 = n7022 | n12961 ;
  assign n12963 = ( ~n12959 & n12960 ) | ( ~n12959 & n12962 ) | ( n12960 & n12962 ) ;
  assign n12964 = ( ~x11 & n12959 ) | ( ~x11 & n12963 ) | ( n12959 & n12963 ) ;
  assign n12965 = ( n12959 & n12963 ) | ( n12959 & ~n12964 ) | ( n12963 & ~n12964 ) ;
  assign n12966 = ( x11 & n12964 ) | ( x11 & ~n12965 ) | ( n12964 & ~n12965 ) ;
  assign n12967 = ( ~n12683 & n12685 ) | ( ~n12683 & n12694 ) | ( n12685 & n12694 ) ;
  assign n12968 = ( ~n12694 & n12695 ) | ( ~n12694 & n12967 ) | ( n12695 & n12967 ) ;
  assign n12969 = ( n12958 & n12966 ) | ( n12958 & ~n12968 ) | ( n12966 & ~n12968 ) ;
  assign n12970 = n4713 & n11892 ;
  assign n12971 = n4712 & ~n9997 ;
  assign n12972 = n4709 & ~n10001 ;
  assign n12973 = n4792 & n9999 ;
  assign n12974 = n12972 | n12973 ;
  assign n12975 = ( ~n12970 & n12971 ) | ( ~n12970 & n12974 ) | ( n12971 & n12974 ) ;
  assign n12976 = ( ~x23 & n12970 ) | ( ~x23 & n12975 ) | ( n12970 & n12975 ) ;
  assign n12977 = ( n12970 & n12975 ) | ( n12970 & ~n12976 ) | ( n12975 & ~n12976 ) ;
  assign n12978 = ( x23 & n12976 ) | ( x23 & ~n12977 ) | ( n12976 & ~n12977 ) ;
  assign n12979 = n4709 & ~n10003 ;
  assign n12980 = n4792 & ~n10001 ;
  assign n12981 = n12979 | n12980 ;
  assign n12982 = n4712 & ~n9999 ;
  assign n12983 = ( n4712 & n12981 ) | ( n4712 & ~n12982 ) | ( n12981 & ~n12982 ) ;
  assign n12984 = n4713 & n11868 ;
  assign n12985 = n12983 | n12984 ;
  assign n12986 = n4711 & ~n10003 ;
  assign n12987 = x23 & n12986 ;
  assign n12988 = ( n4713 & n11804 ) | ( n4713 & n11805 ) | ( n11804 & n11805 ) ;
  assign n12989 = n4792 | n10003 ;
  assign n12990 = n4712 & ~n10001 ;
  assign n12991 = ( ~n10003 & n12989 ) | ( ~n10003 & n12990 ) | ( n12989 & n12990 ) ;
  assign n12992 = n12988 | n12991 ;
  assign n12993 = ( x23 & n12987 ) | ( x23 & n12992 ) | ( n12987 & n12992 ) ;
  assign n12994 = n12985 | n12993 ;
  assign n12995 = x23 & ~n12994 ;
  assign n12996 = ( n12720 & n12978 ) | ( n12720 & n12995 ) | ( n12978 & n12995 ) ;
  assign n12997 = n4713 & n11934 ;
  assign n12998 = n4712 & n9995 ;
  assign n12999 = n4709 & n9999 ;
  assign n13000 = n4792 & ~n9997 ;
  assign n13001 = n12999 | n13000 ;
  assign n13002 = ( ~n12997 & n12998 ) | ( ~n12997 & n13001 ) | ( n12998 & n13001 ) ;
  assign n13003 = ( ~x23 & n12997 ) | ( ~x23 & n13002 ) | ( n12997 & n13002 ) ;
  assign n13004 = ( n12997 & n13002 ) | ( n12997 & ~n13003 ) | ( n13002 & ~n13003 ) ;
  assign n13005 = ( x23 & n13003 ) | ( x23 & ~n13004 ) | ( n13003 & ~n13004 ) ;
  assign n13006 = ( n12722 & n12725 ) | ( n12722 & ~n12726 ) | ( n12725 & ~n12726 ) ;
  assign n13007 = ( n12721 & n12726 ) | ( n12721 & ~n13006 ) | ( n12726 & ~n13006 ) ;
  assign n13008 = ( n12996 & n13005 ) | ( n12996 & n13007 ) | ( n13005 & n13007 ) ;
  assign n13009 = n4713 & ~n11971 ;
  assign n13010 = n4712 & n9993 ;
  assign n13011 = n4709 & ~n9997 ;
  assign n13012 = n4792 & n9995 ;
  assign n13013 = n13011 | n13012 ;
  assign n13014 = ( ~n13009 & n13010 ) | ( ~n13009 & n13013 ) | ( n13010 & n13013 ) ;
  assign n13015 = ( ~x23 & n13009 ) | ( ~x23 & n13014 ) | ( n13009 & n13014 ) ;
  assign n13016 = ( n13009 & n13014 ) | ( n13009 & ~n13015 ) | ( n13014 & ~n13015 ) ;
  assign n13017 = ( x23 & n13015 ) | ( x23 & ~n13016 ) | ( n13015 & ~n13016 ) ;
  assign n13018 = ( n12719 & n12727 ) | ( n12719 & ~n12728 ) | ( n12727 & ~n12728 ) ;
  assign n13019 = n12728 & ~n13018 ;
  assign n13020 = ( n13008 & n13017 ) | ( n13008 & n13019 ) | ( n13017 & n13019 ) ;
  assign n13021 = n4713 & n12026 ;
  assign n13022 = n4712 & n9991 ;
  assign n13023 = n4709 & n9995 ;
  assign n13024 = n4792 & n9993 ;
  assign n13025 = n13023 | n13024 ;
  assign n13026 = ( ~n13021 & n13022 ) | ( ~n13021 & n13025 ) | ( n13022 & n13025 ) ;
  assign n13027 = ( ~x23 & n13021 ) | ( ~x23 & n13026 ) | ( n13021 & n13026 ) ;
  assign n13028 = ( n13021 & n13026 ) | ( n13021 & ~n13027 ) | ( n13026 & ~n13027 ) ;
  assign n13029 = ( x23 & n13027 ) | ( x23 & ~n13028 ) | ( n13027 & ~n13028 ) ;
  assign n13030 = ( n12481 & n12712 ) | ( n12481 & ~n12729 ) | ( n12712 & ~n12729 ) ;
  assign n13031 = ( n12729 & ~n12730 ) | ( n12729 & n13030 ) | ( ~n12730 & n13030 ) ;
  assign n13032 = ( n13020 & n13029 ) | ( n13020 & n13031 ) | ( n13029 & n13031 ) ;
  assign n13033 = n4713 & n12050 ;
  assign n13034 = n4712 & n9989 ;
  assign n13035 = n4709 & n9993 ;
  assign n13036 = n4792 & n9991 ;
  assign n13037 = n13035 | n13036 ;
  assign n13038 = ( ~n13033 & n13034 ) | ( ~n13033 & n13037 ) | ( n13034 & n13037 ) ;
  assign n13039 = ( ~x23 & n13033 ) | ( ~x23 & n13038 ) | ( n13033 & n13038 ) ;
  assign n13040 = ( n13033 & n13038 ) | ( n13033 & ~n13039 ) | ( n13038 & ~n13039 ) ;
  assign n13041 = ( x23 & n13039 ) | ( x23 & ~n13040 ) | ( n13039 & ~n13040 ) ;
  assign n13042 = ( ~n12730 & n12739 ) | ( ~n12730 & n12741 ) | ( n12739 & n12741 ) ;
  assign n13043 = ( n12730 & ~n12742 ) | ( n12730 & n13042 ) | ( ~n12742 & n13042 ) ;
  assign n13044 = ( n13032 & n13041 ) | ( n13032 & n13043 ) | ( n13041 & n13043 ) ;
  assign n13045 = ( ~n12742 & n12751 ) | ( ~n12742 & n12753 ) | ( n12751 & n12753 ) ;
  assign n13046 = ( n12742 & ~n12754 ) | ( n12742 & n13045 ) | ( ~n12754 & n13045 ) ;
  assign n13047 = n4713 & ~n12074 ;
  assign n13048 = n4712 & ~n9987 ;
  assign n13049 = n4709 & n9991 ;
  assign n13050 = n4792 & n9989 ;
  assign n13051 = n13049 | n13050 ;
  assign n13052 = ( ~n13047 & n13048 ) | ( ~n13047 & n13051 ) | ( n13048 & n13051 ) ;
  assign n13053 = ( ~x23 & n13047 ) | ( ~x23 & n13052 ) | ( n13047 & n13052 ) ;
  assign n13054 = ( n13047 & n13052 ) | ( n13047 & ~n13053 ) | ( n13052 & ~n13053 ) ;
  assign n13055 = ( x23 & n13053 ) | ( x23 & ~n13054 ) | ( n13053 & ~n13054 ) ;
  assign n13056 = ( n13044 & n13046 ) | ( n13044 & n13055 ) | ( n13046 & n13055 ) ;
  assign n13057 = ( ~n12754 & n12763 ) | ( ~n12754 & n12765 ) | ( n12763 & n12765 ) ;
  assign n13058 = ( n12754 & ~n12766 ) | ( n12754 & n13057 ) | ( ~n12766 & n13057 ) ;
  assign n13059 = n4713 & ~n12099 ;
  assign n13060 = n4712 & n9985 ;
  assign n13061 = n4709 & n9989 ;
  assign n13062 = n4792 & ~n9987 ;
  assign n13063 = n13061 | n13062 ;
  assign n13064 = ( ~n13059 & n13060 ) | ( ~n13059 & n13063 ) | ( n13060 & n13063 ) ;
  assign n13065 = ( ~x23 & n13059 ) | ( ~x23 & n13064 ) | ( n13059 & n13064 ) ;
  assign n13066 = ( n13059 & n13064 ) | ( n13059 & ~n13065 ) | ( n13064 & ~n13065 ) ;
  assign n13067 = ( x23 & n13065 ) | ( x23 & ~n13066 ) | ( n13065 & ~n13066 ) ;
  assign n13068 = ( n13056 & n13058 ) | ( n13056 & n13067 ) | ( n13058 & n13067 ) ;
  assign n13069 = n4713 & ~n12129 ;
  assign n13070 = n4712 & ~n9983 ;
  assign n13071 = n4709 & ~n9987 ;
  assign n13072 = n4792 & n9985 ;
  assign n13073 = n13071 | n13072 ;
  assign n13074 = ( ~n13069 & n13070 ) | ( ~n13069 & n13073 ) | ( n13070 & n13073 ) ;
  assign n13075 = ( ~x23 & n13069 ) | ( ~x23 & n13074 ) | ( n13069 & n13074 ) ;
  assign n13076 = ( n13069 & n13074 ) | ( n13069 & ~n13075 ) | ( n13074 & ~n13075 ) ;
  assign n13077 = ( x23 & n13075 ) | ( x23 & ~n13076 ) | ( n13075 & ~n13076 ) ;
  assign n13078 = ( n12766 & ~n12775 ) | ( n12766 & n12777 ) | ( ~n12775 & n12777 ) ;
  assign n13079 = ( ~n12766 & n12778 ) | ( ~n12766 & n13078 ) | ( n12778 & n13078 ) ;
  assign n13080 = ( n13068 & n13077 ) | ( n13068 & ~n13079 ) | ( n13077 & ~n13079 ) ;
  assign n13081 = n4713 & ~n11561 ;
  assign n13082 = n4712 & n9981 ;
  assign n13083 = n4709 & n9985 ;
  assign n13084 = n4792 & ~n9983 ;
  assign n13085 = n13083 | n13084 ;
  assign n13086 = ( ~n13081 & n13082 ) | ( ~n13081 & n13085 ) | ( n13082 & n13085 ) ;
  assign n13087 = ( ~x23 & n13081 ) | ( ~x23 & n13086 ) | ( n13081 & n13086 ) ;
  assign n13088 = ( n13081 & n13086 ) | ( n13081 & ~n13087 ) | ( n13086 & ~n13087 ) ;
  assign n13089 = ( x23 & n13087 ) | ( x23 & ~n13088 ) | ( n13087 & ~n13088 ) ;
  assign n13090 = ( ~n12778 & n12780 ) | ( ~n12778 & n12789 ) | ( n12780 & n12789 ) ;
  assign n13091 = ( ~n12789 & n12790 ) | ( ~n12789 & n13090 ) | ( n12790 & n13090 ) ;
  assign n13092 = ( n13080 & n13089 ) | ( n13080 & ~n13091 ) | ( n13089 & ~n13091 ) ;
  assign n13093 = n4713 & n12153 ;
  assign n13094 = n4712 & n9979 ;
  assign n13095 = n4709 & ~n9983 ;
  assign n13096 = n4792 & n9981 ;
  assign n13097 = n13095 | n13096 ;
  assign n13098 = ( ~n13093 & n13094 ) | ( ~n13093 & n13097 ) | ( n13094 & n13097 ) ;
  assign n13099 = ( ~x23 & n13093 ) | ( ~x23 & n13098 ) | ( n13093 & n13098 ) ;
  assign n13100 = ( n13093 & n13098 ) | ( n13093 & ~n13099 ) | ( n13098 & ~n13099 ) ;
  assign n13101 = ( x23 & n13099 ) | ( x23 & ~n13100 ) | ( n13099 & ~n13100 ) ;
  assign n13102 = ( ~n12790 & n12792 ) | ( ~n12790 & n12801 ) | ( n12792 & n12801 ) ;
  assign n13103 = ( n12790 & ~n12802 ) | ( n12790 & n13102 ) | ( ~n12802 & n13102 ) ;
  assign n13104 = ( n13092 & n13101 ) | ( n13092 & n13103 ) | ( n13101 & n13103 ) ;
  assign n13105 = n4713 & n12165 ;
  assign n13106 = n4712 & n9977 ;
  assign n13107 = n4709 & n9981 ;
  assign n13108 = n4792 & n9979 ;
  assign n13109 = n13107 | n13108 ;
  assign n13110 = ( ~n13105 & n13106 ) | ( ~n13105 & n13109 ) | ( n13106 & n13109 ) ;
  assign n13111 = ( ~x23 & n13105 ) | ( ~x23 & n13110 ) | ( n13105 & n13110 ) ;
  assign n13112 = ( n13105 & n13110 ) | ( n13105 & ~n13111 ) | ( n13110 & ~n13111 ) ;
  assign n13113 = ( x23 & n13111 ) | ( x23 & ~n13112 ) | ( n13111 & ~n13112 ) ;
  assign n13114 = ( ~n12802 & n12804 ) | ( ~n12802 & n12813 ) | ( n12804 & n12813 ) ;
  assign n13115 = ( ~n12813 & n12814 ) | ( ~n12813 & n13114 ) | ( n12814 & n13114 ) ;
  assign n13116 = ( n13104 & n13113 ) | ( n13104 & ~n13115 ) | ( n13113 & ~n13115 ) ;
  assign n13117 = n4713 & n11606 ;
  assign n13118 = n4712 & n9975 ;
  assign n13119 = n4709 & n9979 ;
  assign n13120 = n4792 & n9977 ;
  assign n13121 = n13119 | n13120 ;
  assign n13122 = ( ~n13117 & n13118 ) | ( ~n13117 & n13121 ) | ( n13118 & n13121 ) ;
  assign n13123 = ( ~x23 & n13117 ) | ( ~x23 & n13122 ) | ( n13117 & n13122 ) ;
  assign n13124 = ( n13117 & n13122 ) | ( n13117 & ~n13123 ) | ( n13122 & ~n13123 ) ;
  assign n13125 = ( x23 & n13123 ) | ( x23 & ~n13124 ) | ( n13123 & ~n13124 ) ;
  assign n13126 = ( ~n12814 & n12816 ) | ( ~n12814 & n12825 ) | ( n12816 & n12825 ) ;
  assign n13127 = ( ~n12825 & n12826 ) | ( ~n12825 & n13126 ) | ( n12826 & n13126 ) ;
  assign n13128 = ( n13116 & n13125 ) | ( n13116 & ~n13127 ) | ( n13125 & ~n13127 ) ;
  assign n13129 = n4713 & n11400 ;
  assign n13130 = n4712 & n9973 ;
  assign n13131 = n4709 & n9977 ;
  assign n13132 = n4792 & n9975 ;
  assign n13133 = n13131 | n13132 ;
  assign n13134 = ( ~n13129 & n13130 ) | ( ~n13129 & n13133 ) | ( n13130 & n13133 ) ;
  assign n13135 = ( ~x23 & n13129 ) | ( ~x23 & n13134 ) | ( n13129 & n13134 ) ;
  assign n13136 = ( n13129 & n13134 ) | ( n13129 & ~n13135 ) | ( n13134 & ~n13135 ) ;
  assign n13137 = ( x23 & n13135 ) | ( x23 & ~n13136 ) | ( n13135 & ~n13136 ) ;
  assign n13138 = ( ~n12826 & n12828 ) | ( ~n12826 & n12837 ) | ( n12828 & n12837 ) ;
  assign n13139 = ( n12826 & ~n12838 ) | ( n12826 & n13138 ) | ( ~n12838 & n13138 ) ;
  assign n13140 = ( n13128 & n13137 ) | ( n13128 & n13139 ) | ( n13137 & n13139 ) ;
  assign n13141 = n4713 & n11630 ;
  assign n13142 = n4712 & n9971 ;
  assign n13143 = n4709 & n9975 ;
  assign n13144 = n4792 & n9973 ;
  assign n13145 = n13143 | n13144 ;
  assign n13146 = ( ~n13141 & n13142 ) | ( ~n13141 & n13145 ) | ( n13142 & n13145 ) ;
  assign n13147 = ( ~x23 & n13141 ) | ( ~x23 & n13146 ) | ( n13141 & n13146 ) ;
  assign n13148 = ( n13141 & n13146 ) | ( n13141 & ~n13147 ) | ( n13146 & ~n13147 ) ;
  assign n13149 = ( x23 & n13147 ) | ( x23 & ~n13148 ) | ( n13147 & ~n13148 ) ;
  assign n13150 = ( ~n12838 & n12840 ) | ( ~n12838 & n12849 ) | ( n12840 & n12849 ) ;
  assign n13151 = ( n12838 & ~n12850 ) | ( n12838 & n13150 ) | ( ~n12850 & n13150 ) ;
  assign n13152 = ( n13140 & n13149 ) | ( n13140 & n13151 ) | ( n13149 & n13151 ) ;
  assign n13153 = n4713 & n11428 ;
  assign n13154 = n4712 & n9969 ;
  assign n13155 = n4709 & n9973 ;
  assign n13156 = n4792 & n9971 ;
  assign n13157 = n13155 | n13156 ;
  assign n13158 = ( ~n13153 & n13154 ) | ( ~n13153 & n13157 ) | ( n13154 & n13157 ) ;
  assign n13159 = ( ~x23 & n13153 ) | ( ~x23 & n13158 ) | ( n13153 & n13158 ) ;
  assign n13160 = ( n13153 & n13158 ) | ( n13153 & ~n13159 ) | ( n13158 & ~n13159 ) ;
  assign n13161 = ( x23 & n13159 ) | ( x23 & ~n13160 ) | ( n13159 & ~n13160 ) ;
  assign n13162 = ( ~n12850 & n12852 ) | ( ~n12850 & n12861 ) | ( n12852 & n12861 ) ;
  assign n13163 = ( n12850 & ~n12862 ) | ( n12850 & n13162 ) | ( ~n12862 & n13162 ) ;
  assign n13164 = ( n13152 & n13161 ) | ( n13152 & n13163 ) | ( n13161 & n13163 ) ;
  assign n13165 = n4713 & ~n10998 ;
  assign n13166 = n4712 & ~n9967 ;
  assign n13167 = n4709 & n9971 ;
  assign n13168 = n4792 & n9969 ;
  assign n13169 = n13167 | n13168 ;
  assign n13170 = ( ~n13165 & n13166 ) | ( ~n13165 & n13169 ) | ( n13166 & n13169 ) ;
  assign n13171 = ( ~x23 & n13165 ) | ( ~x23 & n13170 ) | ( n13165 & n13170 ) ;
  assign n13172 = ( n13165 & n13170 ) | ( n13165 & ~n13171 ) | ( n13170 & ~n13171 ) ;
  assign n13173 = ( x23 & n13171 ) | ( x23 & ~n13172 ) | ( n13171 & ~n13172 ) ;
  assign n13174 = ( ~n12862 & n12864 ) | ( ~n12862 & n12873 ) | ( n12864 & n12873 ) ;
  assign n13175 = ( n12862 & ~n12874 ) | ( n12862 & n13174 ) | ( ~n12874 & n13174 ) ;
  assign n13176 = ( n13164 & n13173 ) | ( n13164 & n13175 ) | ( n13173 & n13175 ) ;
  assign n13177 = n4713 & ~n11273 ;
  assign n13178 = n4712 & n9965 ;
  assign n13179 = n4709 & n9969 ;
  assign n13180 = n4792 & ~n9967 ;
  assign n13181 = n13179 | n13180 ;
  assign n13182 = ( ~n13177 & n13178 ) | ( ~n13177 & n13181 ) | ( n13178 & n13181 ) ;
  assign n13183 = ( ~x23 & n13177 ) | ( ~x23 & n13182 ) | ( n13177 & n13182 ) ;
  assign n13184 = ( n13177 & n13182 ) | ( n13177 & ~n13183 ) | ( n13182 & ~n13183 ) ;
  assign n13185 = ( x23 & n13183 ) | ( x23 & ~n13184 ) | ( n13183 & ~n13184 ) ;
  assign n13186 = ( ~n12874 & n12876 ) | ( ~n12874 & n12885 ) | ( n12876 & n12885 ) ;
  assign n13187 = ( n12874 & ~n12886 ) | ( n12874 & n13186 ) | ( ~n12886 & n13186 ) ;
  assign n13188 = ( n13176 & n13185 ) | ( n13176 & n13187 ) | ( n13185 & n13187 ) ;
  assign n13189 = ( ~n12886 & n12888 ) | ( ~n12886 & n12897 ) | ( n12888 & n12897 ) ;
  assign n13190 = ( ~n12897 & n12898 ) | ( ~n12897 & n13189 ) | ( n12898 & n13189 ) ;
  assign n13191 = n4974 & ~n10869 ;
  assign n13192 = n5398 & ~n9957 ;
  assign n13193 = n4973 & n9961 ;
  assign n13194 = n4972 & n9959 ;
  assign n13195 = n13193 | n13194 ;
  assign n13196 = ( ~n13191 & n13192 ) | ( ~n13191 & n13195 ) | ( n13192 & n13195 ) ;
  assign n13197 = ( ~x20 & n13191 ) | ( ~x20 & n13196 ) | ( n13191 & n13196 ) ;
  assign n13198 = ( n13191 & n13196 ) | ( n13191 & ~n13197 ) | ( n13196 & ~n13197 ) ;
  assign n13199 = ( x20 & n13197 ) | ( x20 & ~n13198 ) | ( n13197 & ~n13198 ) ;
  assign n13200 = ( n13188 & ~n13190 ) | ( n13188 & n13199 ) | ( ~n13190 & n13199 ) ;
  assign n13201 = ( n12898 & ~n12900 ) | ( n12898 & n12909 ) | ( ~n12900 & n12909 ) ;
  assign n13202 = ( n12900 & ~n12910 ) | ( n12900 & n13201 ) | ( ~n12910 & n13201 ) ;
  assign n13203 = n5508 & n10557 ;
  assign n13204 = n5507 & n9949 ;
  assign n13205 = n5504 & ~n9953 ;
  assign n13206 = n5666 & n9951 ;
  assign n13207 = n13205 | n13206 ;
  assign n13208 = ( ~n13203 & n13204 ) | ( ~n13203 & n13207 ) | ( n13204 & n13207 ) ;
  assign n13209 = ( ~x17 & n13203 ) | ( ~x17 & n13208 ) | ( n13203 & n13208 ) ;
  assign n13210 = ( n13203 & n13208 ) | ( n13203 & ~n13209 ) | ( n13208 & ~n13209 ) ;
  assign n13211 = ( x17 & n13209 ) | ( x17 & ~n13210 ) | ( n13209 & ~n13210 ) ;
  assign n13212 = ( n13200 & n13202 ) | ( n13200 & n13211 ) | ( n13202 & n13211 ) ;
  assign n13213 = ( ~n12910 & n12912 ) | ( ~n12910 & n12921 ) | ( n12912 & n12921 ) ;
  assign n13214 = ( ~n12921 & n12922 ) | ( ~n12921 & n13213 ) | ( n12922 & n13213 ) ;
  assign n13215 = n5966 & ~n10390 ;
  assign n13216 = n6464 & ~n9941 ;
  assign n13217 = n5970 & n9945 ;
  assign n13218 = n5969 & n9943 ;
  assign n13219 = n13217 | n13218 ;
  assign n13220 = ( ~n13215 & n13216 ) | ( ~n13215 & n13219 ) | ( n13216 & n13219 ) ;
  assign n13221 = ( ~x14 & n13215 ) | ( ~x14 & n13220 ) | ( n13215 & n13220 ) ;
  assign n13222 = ( n13215 & n13220 ) | ( n13215 & ~n13221 ) | ( n13220 & ~n13221 ) ;
  assign n13223 = ( x14 & n13221 ) | ( x14 & ~n13222 ) | ( n13221 & ~n13222 ) ;
  assign n13224 = ( n13212 & ~n13214 ) | ( n13212 & n13223 ) | ( ~n13214 & n13223 ) ;
  assign n13225 = ( ~n12922 & n12924 ) | ( ~n12922 & n12933 ) | ( n12924 & n12933 ) ;
  assign n13226 = ( ~n12933 & n12934 ) | ( ~n12933 & n13225 ) | ( n12934 & n13225 ) ;
  assign n13227 = n5966 & n10284 ;
  assign n13228 = n6464 & ~n9883 ;
  assign n13229 = n5970 & n9943 ;
  assign n13230 = n5969 & ~n9941 ;
  assign n13231 = n13229 | n13230 ;
  assign n13232 = ( ~n13227 & n13228 ) | ( ~n13227 & n13231 ) | ( n13228 & n13231 ) ;
  assign n13233 = ( ~x14 & n13227 ) | ( ~x14 & n13232 ) | ( n13227 & n13232 ) ;
  assign n13234 = ( n13227 & n13232 ) | ( n13227 & ~n13233 ) | ( n13232 & ~n13233 ) ;
  assign n13235 = ( x14 & n13233 ) | ( x14 & ~n13234 ) | ( n13233 & ~n13234 ) ;
  assign n13236 = ( n13224 & ~n13226 ) | ( n13224 & n13235 ) | ( ~n13226 & n13235 ) ;
  assign n13237 = ( n12934 & ~n12936 ) | ( n12934 & n12945 ) | ( ~n12936 & n12945 ) ;
  assign n13238 = ( n12936 & ~n12946 ) | ( n12936 & n13237 ) | ( ~n12946 & n13237 ) ;
  assign n13239 = n6584 & ~n10305 ;
  assign n13240 = n7022 & ~n10302 ;
  assign n13241 = n6588 & ~n9937 ;
  assign n13242 = n6587 & ~n10057 ;
  assign n13243 = n13241 | n13242 ;
  assign n13244 = ( ~n13239 & n13240 ) | ( ~n13239 & n13243 ) | ( n13240 & n13243 ) ;
  assign n13245 = ( ~x11 & n13239 ) | ( ~x11 & n13244 ) | ( n13239 & n13244 ) ;
  assign n13246 = ( n13239 & n13244 ) | ( n13239 & ~n13245 ) | ( n13244 & ~n13245 ) ;
  assign n13247 = ( x11 & n13245 ) | ( x11 & ~n13246 ) | ( n13245 & ~n13246 ) ;
  assign n13248 = ( n13236 & n13238 ) | ( n13236 & n13247 ) | ( n13238 & n13247 ) ;
  assign n13249 = x8 | n11067 ;
  assign n13250 = ( x8 & n11067 ) | ( x8 & ~n13249 ) | ( n11067 & ~n13249 ) ;
  assign n13251 = n13249 & ~n13250 ;
  assign n13252 = ( ~n12946 & n12948 ) | ( ~n12946 & n12957 ) | ( n12948 & n12957 ) ;
  assign n13253 = ( ~n12957 & n12958 ) | ( ~n12957 & n13252 ) | ( n12958 & n13252 ) ;
  assign n13254 = ( n13248 & n13251 ) | ( n13248 & ~n13253 ) | ( n13251 & ~n13253 ) ;
  assign n13255 = n4974 & n11892 ;
  assign n13256 = n5398 & ~n9997 ;
  assign n13257 = n4973 & ~n10001 ;
  assign n13258 = n4972 & n9999 ;
  assign n13259 = n13257 | n13258 ;
  assign n13260 = ( ~n13255 & n13256 ) | ( ~n13255 & n13259 ) | ( n13256 & n13259 ) ;
  assign n13261 = ( ~x20 & n13255 ) | ( ~x20 & n13260 ) | ( n13255 & n13260 ) ;
  assign n13262 = ( n13255 & n13260 ) | ( n13255 & ~n13261 ) | ( n13260 & ~n13261 ) ;
  assign n13263 = ( x20 & n13261 ) | ( x20 & ~n13262 ) | ( n13261 & ~n13262 ) ;
  assign n13264 = n4973 & ~n10003 ;
  assign n13265 = n4972 & ~n10001 ;
  assign n13266 = n13264 | n13265 ;
  assign n13267 = n5398 & ~n9999 ;
  assign n13268 = ( n5398 & n13266 ) | ( n5398 & ~n13267 ) | ( n13266 & ~n13267 ) ;
  assign n13269 = n4974 & n11868 ;
  assign n13270 = n13268 | n13269 ;
  assign n13271 = n5397 & ~n10003 ;
  assign n13272 = x20 & n13271 ;
  assign n13273 = ( n4974 & n11804 ) | ( n4974 & n11805 ) | ( n11804 & n11805 ) ;
  assign n13274 = n4972 | n10003 ;
  assign n13275 = n5398 & ~n10001 ;
  assign n13276 = ( ~n10003 & n13274 ) | ( ~n10003 & n13275 ) | ( n13274 & n13275 ) ;
  assign n13277 = n13273 | n13276 ;
  assign n13278 = ( x20 & n13272 ) | ( x20 & n13277 ) | ( n13272 & n13277 ) ;
  assign n13279 = n13270 | n13278 ;
  assign n13280 = x20 & ~n13279 ;
  assign n13281 = ( n12986 & n13263 ) | ( n12986 & n13280 ) | ( n13263 & n13280 ) ;
  assign n13282 = n4974 & n11934 ;
  assign n13283 = n5398 & n9995 ;
  assign n13284 = n4973 & n9999 ;
  assign n13285 = n4972 & ~n9997 ;
  assign n13286 = n13284 | n13285 ;
  assign n13287 = ( ~n13282 & n13283 ) | ( ~n13282 & n13286 ) | ( n13283 & n13286 ) ;
  assign n13288 = ( ~x20 & n13282 ) | ( ~x20 & n13287 ) | ( n13282 & n13287 ) ;
  assign n13289 = ( n13282 & n13287 ) | ( n13282 & ~n13288 ) | ( n13287 & ~n13288 ) ;
  assign n13290 = ( x20 & n13288 ) | ( x20 & ~n13289 ) | ( n13288 & ~n13289 ) ;
  assign n13291 = ( n12987 & n12988 ) | ( n12987 & n12991 ) | ( n12988 & n12991 ) ;
  assign n13292 = ~n12987 & n12992 ;
  assign n13293 = ( n12987 & ~n13291 ) | ( n12987 & n13292 ) | ( ~n13291 & n13292 ) ;
  assign n13294 = ( n13281 & n13290 ) | ( n13281 & n13293 ) | ( n13290 & n13293 ) ;
  assign n13295 = n4974 & ~n11971 ;
  assign n13296 = n5398 & n9993 ;
  assign n13297 = n4973 & ~n9997 ;
  assign n13298 = n4972 & n9995 ;
  assign n13299 = n13297 | n13298 ;
  assign n13300 = ( ~n13295 & n13296 ) | ( ~n13295 & n13299 ) | ( n13296 & n13299 ) ;
  assign n13301 = ( ~x20 & n13295 ) | ( ~x20 & n13300 ) | ( n13295 & n13300 ) ;
  assign n13302 = ( n13295 & n13300 ) | ( n13295 & ~n13301 ) | ( n13300 & ~n13301 ) ;
  assign n13303 = ( x20 & n13301 ) | ( x20 & ~n13302 ) | ( n13301 & ~n13302 ) ;
  assign n13304 = ( n12985 & n12993 ) | ( n12985 & ~n12994 ) | ( n12993 & ~n12994 ) ;
  assign n13305 = n12994 & ~n13304 ;
  assign n13306 = ( n13294 & n13303 ) | ( n13294 & n13305 ) | ( n13303 & n13305 ) ;
  assign n13307 = n4974 & n12026 ;
  assign n13308 = n5398 & n9991 ;
  assign n13309 = n4973 & n9995 ;
  assign n13310 = n4972 & n9993 ;
  assign n13311 = n13309 | n13310 ;
  assign n13312 = ( ~n13307 & n13308 ) | ( ~n13307 & n13311 ) | ( n13308 & n13311 ) ;
  assign n13313 = ( ~x20 & n13307 ) | ( ~x20 & n13312 ) | ( n13307 & n13312 ) ;
  assign n13314 = ( n13307 & n13312 ) | ( n13307 & ~n13313 ) | ( n13312 & ~n13313 ) ;
  assign n13315 = ( x20 & n13313 ) | ( x20 & ~n13314 ) | ( n13313 & ~n13314 ) ;
  assign n13316 = ( n12720 & n12978 ) | ( n12720 & ~n12995 ) | ( n12978 & ~n12995 ) ;
  assign n13317 = ( n12995 & ~n12996 ) | ( n12995 & n13316 ) | ( ~n12996 & n13316 ) ;
  assign n13318 = ( n13306 & n13315 ) | ( n13306 & n13317 ) | ( n13315 & n13317 ) ;
  assign n13319 = n4974 & n12050 ;
  assign n13320 = n5398 & n9989 ;
  assign n13321 = n4973 & n9993 ;
  assign n13322 = n4972 & n9991 ;
  assign n13323 = n13321 | n13322 ;
  assign n13324 = ( ~n13319 & n13320 ) | ( ~n13319 & n13323 ) | ( n13320 & n13323 ) ;
  assign n13325 = ( ~x20 & n13319 ) | ( ~x20 & n13324 ) | ( n13319 & n13324 ) ;
  assign n13326 = ( n13319 & n13324 ) | ( n13319 & ~n13325 ) | ( n13324 & ~n13325 ) ;
  assign n13327 = ( x20 & n13325 ) | ( x20 & ~n13326 ) | ( n13325 & ~n13326 ) ;
  assign n13328 = ( ~n12996 & n13005 ) | ( ~n12996 & n13007 ) | ( n13005 & n13007 ) ;
  assign n13329 = ( n12996 & ~n13008 ) | ( n12996 & n13328 ) | ( ~n13008 & n13328 ) ;
  assign n13330 = ( n13318 & n13327 ) | ( n13318 & n13329 ) | ( n13327 & n13329 ) ;
  assign n13331 = ( ~n13008 & n13017 ) | ( ~n13008 & n13019 ) | ( n13017 & n13019 ) ;
  assign n13332 = ( n13008 & ~n13020 ) | ( n13008 & n13331 ) | ( ~n13020 & n13331 ) ;
  assign n13333 = n4974 & ~n12074 ;
  assign n13334 = n5398 & ~n9987 ;
  assign n13335 = n4973 & n9991 ;
  assign n13336 = n4972 & n9989 ;
  assign n13337 = n13335 | n13336 ;
  assign n13338 = ( ~n13333 & n13334 ) | ( ~n13333 & n13337 ) | ( n13334 & n13337 ) ;
  assign n13339 = ( ~x20 & n13333 ) | ( ~x20 & n13338 ) | ( n13333 & n13338 ) ;
  assign n13340 = ( n13333 & n13338 ) | ( n13333 & ~n13339 ) | ( n13338 & ~n13339 ) ;
  assign n13341 = ( x20 & n13339 ) | ( x20 & ~n13340 ) | ( n13339 & ~n13340 ) ;
  assign n13342 = ( n13330 & n13332 ) | ( n13330 & n13341 ) | ( n13332 & n13341 ) ;
  assign n13343 = ( ~n13020 & n13029 ) | ( ~n13020 & n13031 ) | ( n13029 & n13031 ) ;
  assign n13344 = ( n13020 & ~n13032 ) | ( n13020 & n13343 ) | ( ~n13032 & n13343 ) ;
  assign n13345 = n4974 & ~n12099 ;
  assign n13346 = n5398 & n9985 ;
  assign n13347 = n4973 & n9989 ;
  assign n13348 = n4972 & ~n9987 ;
  assign n13349 = n13347 | n13348 ;
  assign n13350 = ( ~n13345 & n13346 ) | ( ~n13345 & n13349 ) | ( n13346 & n13349 ) ;
  assign n13351 = ( ~x20 & n13345 ) | ( ~x20 & n13350 ) | ( n13345 & n13350 ) ;
  assign n13352 = ( n13345 & n13350 ) | ( n13345 & ~n13351 ) | ( n13350 & ~n13351 ) ;
  assign n13353 = ( x20 & n13351 ) | ( x20 & ~n13352 ) | ( n13351 & ~n13352 ) ;
  assign n13354 = ( n13342 & n13344 ) | ( n13342 & n13353 ) | ( n13344 & n13353 ) ;
  assign n13355 = ( ~n13032 & n13041 ) | ( ~n13032 & n13043 ) | ( n13041 & n13043 ) ;
  assign n13356 = ( n13032 & ~n13044 ) | ( n13032 & n13355 ) | ( ~n13044 & n13355 ) ;
  assign n13357 = n4974 & ~n12129 ;
  assign n13358 = n5398 & ~n9983 ;
  assign n13359 = n4973 & ~n9987 ;
  assign n13360 = n4972 & n9985 ;
  assign n13361 = n13359 | n13360 ;
  assign n13362 = ( ~n13357 & n13358 ) | ( ~n13357 & n13361 ) | ( n13358 & n13361 ) ;
  assign n13363 = ( ~x20 & n13357 ) | ( ~x20 & n13362 ) | ( n13357 & n13362 ) ;
  assign n13364 = ( n13357 & n13362 ) | ( n13357 & ~n13363 ) | ( n13362 & ~n13363 ) ;
  assign n13365 = ( x20 & n13363 ) | ( x20 & ~n13364 ) | ( n13363 & ~n13364 ) ;
  assign n13366 = ( n13354 & n13356 ) | ( n13354 & n13365 ) | ( n13356 & n13365 ) ;
  assign n13367 = n4974 & ~n11561 ;
  assign n13368 = n5398 & n9981 ;
  assign n13369 = n4973 & n9985 ;
  assign n13370 = n4972 & ~n9983 ;
  assign n13371 = n13369 | n13370 ;
  assign n13372 = ( ~n13367 & n13368 ) | ( ~n13367 & n13371 ) | ( n13368 & n13371 ) ;
  assign n13373 = ( ~x20 & n13367 ) | ( ~x20 & n13372 ) | ( n13367 & n13372 ) ;
  assign n13374 = ( n13367 & n13372 ) | ( n13367 & ~n13373 ) | ( n13372 & ~n13373 ) ;
  assign n13375 = ( x20 & n13373 ) | ( x20 & ~n13374 ) | ( n13373 & ~n13374 ) ;
  assign n13376 = ( ~n13044 & n13046 ) | ( ~n13044 & n13055 ) | ( n13046 & n13055 ) ;
  assign n13377 = ( n13044 & ~n13056 ) | ( n13044 & n13376 ) | ( ~n13056 & n13376 ) ;
  assign n13378 = ( n13366 & n13375 ) | ( n13366 & n13377 ) | ( n13375 & n13377 ) ;
  assign n13379 = n4974 & n12153 ;
  assign n13380 = n5398 & n9979 ;
  assign n13381 = n4973 & ~n9983 ;
  assign n13382 = n4972 & n9981 ;
  assign n13383 = n13381 | n13382 ;
  assign n13384 = ( ~n13379 & n13380 ) | ( ~n13379 & n13383 ) | ( n13380 & n13383 ) ;
  assign n13385 = ( ~x20 & n13379 ) | ( ~x20 & n13384 ) | ( n13379 & n13384 ) ;
  assign n13386 = ( n13379 & n13384 ) | ( n13379 & ~n13385 ) | ( n13384 & ~n13385 ) ;
  assign n13387 = ( x20 & n13385 ) | ( x20 & ~n13386 ) | ( n13385 & ~n13386 ) ;
  assign n13388 = ( ~n13056 & n13058 ) | ( ~n13056 & n13067 ) | ( n13058 & n13067 ) ;
  assign n13389 = ( n13056 & ~n13068 ) | ( n13056 & n13388 ) | ( ~n13068 & n13388 ) ;
  assign n13390 = ( n13378 & n13387 ) | ( n13378 & n13389 ) | ( n13387 & n13389 ) ;
  assign n13391 = ( n13068 & ~n13077 ) | ( n13068 & n13079 ) | ( ~n13077 & n13079 ) ;
  assign n13392 = ( ~n13068 & n13080 ) | ( ~n13068 & n13391 ) | ( n13080 & n13391 ) ;
  assign n13393 = n4974 & n12165 ;
  assign n13394 = n5398 & n9977 ;
  assign n13395 = n4973 & n9981 ;
  assign n13396 = n4972 & n9979 ;
  assign n13397 = n13395 | n13396 ;
  assign n13398 = ( ~n13393 & n13394 ) | ( ~n13393 & n13397 ) | ( n13394 & n13397 ) ;
  assign n13399 = ( ~x20 & n13393 ) | ( ~x20 & n13398 ) | ( n13393 & n13398 ) ;
  assign n13400 = ( n13393 & n13398 ) | ( n13393 & ~n13399 ) | ( n13398 & ~n13399 ) ;
  assign n13401 = ( x20 & n13399 ) | ( x20 & ~n13400 ) | ( n13399 & ~n13400 ) ;
  assign n13402 = ( n13390 & ~n13392 ) | ( n13390 & n13401 ) | ( ~n13392 & n13401 ) ;
  assign n13403 = ( n13080 & ~n13089 ) | ( n13080 & n13091 ) | ( ~n13089 & n13091 ) ;
  assign n13404 = ( ~n13080 & n13092 ) | ( ~n13080 & n13403 ) | ( n13092 & n13403 ) ;
  assign n13405 = n4974 & n11606 ;
  assign n13406 = n5398 & n9975 ;
  assign n13407 = n4973 & n9979 ;
  assign n13408 = n4972 & n9977 ;
  assign n13409 = n13407 | n13408 ;
  assign n13410 = ( ~n13405 & n13406 ) | ( ~n13405 & n13409 ) | ( n13406 & n13409 ) ;
  assign n13411 = ( ~x20 & n13405 ) | ( ~x20 & n13410 ) | ( n13405 & n13410 ) ;
  assign n13412 = ( n13405 & n13410 ) | ( n13405 & ~n13411 ) | ( n13410 & ~n13411 ) ;
  assign n13413 = ( x20 & n13411 ) | ( x20 & ~n13412 ) | ( n13411 & ~n13412 ) ;
  assign n13414 = ( n13402 & ~n13404 ) | ( n13402 & n13413 ) | ( ~n13404 & n13413 ) ;
  assign n13415 = ( ~n13092 & n13101 ) | ( ~n13092 & n13103 ) | ( n13101 & n13103 ) ;
  assign n13416 = ( n13092 & ~n13104 ) | ( n13092 & n13415 ) | ( ~n13104 & n13415 ) ;
  assign n13417 = n4974 & n11400 ;
  assign n13418 = n5398 & n9973 ;
  assign n13419 = n4973 & n9977 ;
  assign n13420 = n4972 & n9975 ;
  assign n13421 = n13419 | n13420 ;
  assign n13422 = ( ~n13417 & n13418 ) | ( ~n13417 & n13421 ) | ( n13418 & n13421 ) ;
  assign n13423 = ( ~x20 & n13417 ) | ( ~x20 & n13422 ) | ( n13417 & n13422 ) ;
  assign n13424 = ( n13417 & n13422 ) | ( n13417 & ~n13423 ) | ( n13422 & ~n13423 ) ;
  assign n13425 = ( x20 & n13423 ) | ( x20 & ~n13424 ) | ( n13423 & ~n13424 ) ;
  assign n13426 = ( n13414 & n13416 ) | ( n13414 & n13425 ) | ( n13416 & n13425 ) ;
  assign n13427 = ( n13104 & ~n13113 ) | ( n13104 & n13115 ) | ( ~n13113 & n13115 ) ;
  assign n13428 = ( ~n13104 & n13116 ) | ( ~n13104 & n13427 ) | ( n13116 & n13427 ) ;
  assign n13429 = n4974 & n11630 ;
  assign n13430 = n5398 & n9971 ;
  assign n13431 = n4973 & n9975 ;
  assign n13432 = n4972 & n9973 ;
  assign n13433 = n13431 | n13432 ;
  assign n13434 = ( ~n13429 & n13430 ) | ( ~n13429 & n13433 ) | ( n13430 & n13433 ) ;
  assign n13435 = ( ~x20 & n13429 ) | ( ~x20 & n13434 ) | ( n13429 & n13434 ) ;
  assign n13436 = ( n13429 & n13434 ) | ( n13429 & ~n13435 ) | ( n13434 & ~n13435 ) ;
  assign n13437 = ( x20 & n13435 ) | ( x20 & ~n13436 ) | ( n13435 & ~n13436 ) ;
  assign n13438 = ( n13426 & ~n13428 ) | ( n13426 & n13437 ) | ( ~n13428 & n13437 ) ;
  assign n13439 = ( n13116 & ~n13125 ) | ( n13116 & n13127 ) | ( ~n13125 & n13127 ) ;
  assign n13440 = ( ~n13116 & n13128 ) | ( ~n13116 & n13439 ) | ( n13128 & n13439 ) ;
  assign n13441 = n4974 & n11428 ;
  assign n13442 = n5398 & n9969 ;
  assign n13443 = n4973 & n9973 ;
  assign n13444 = n4972 & n9971 ;
  assign n13445 = n13443 | n13444 ;
  assign n13446 = ( ~n13441 & n13442 ) | ( ~n13441 & n13445 ) | ( n13442 & n13445 ) ;
  assign n13447 = ( ~x20 & n13441 ) | ( ~x20 & n13446 ) | ( n13441 & n13446 ) ;
  assign n13448 = ( n13441 & n13446 ) | ( n13441 & ~n13447 ) | ( n13446 & ~n13447 ) ;
  assign n13449 = ( x20 & n13447 ) | ( x20 & ~n13448 ) | ( n13447 & ~n13448 ) ;
  assign n13450 = ( n13438 & ~n13440 ) | ( n13438 & n13449 ) | ( ~n13440 & n13449 ) ;
  assign n13451 = ( ~n13128 & n13137 ) | ( ~n13128 & n13139 ) | ( n13137 & n13139 ) ;
  assign n13452 = ( n13128 & ~n13140 ) | ( n13128 & n13451 ) | ( ~n13140 & n13451 ) ;
  assign n13453 = n4974 & ~n10998 ;
  assign n13454 = n5398 & ~n9967 ;
  assign n13455 = n4973 & n9971 ;
  assign n13456 = n4972 & n9969 ;
  assign n13457 = n13455 | n13456 ;
  assign n13458 = ( ~n13453 & n13454 ) | ( ~n13453 & n13457 ) | ( n13454 & n13457 ) ;
  assign n13459 = ( ~x20 & n13453 ) | ( ~x20 & n13458 ) | ( n13453 & n13458 ) ;
  assign n13460 = ( n13453 & n13458 ) | ( n13453 & ~n13459 ) | ( n13458 & ~n13459 ) ;
  assign n13461 = ( x20 & n13459 ) | ( x20 & ~n13460 ) | ( n13459 & ~n13460 ) ;
  assign n13462 = ( n13450 & n13452 ) | ( n13450 & n13461 ) | ( n13452 & n13461 ) ;
  assign n13463 = ( ~n13140 & n13149 ) | ( ~n13140 & n13151 ) | ( n13149 & n13151 ) ;
  assign n13464 = ( n13140 & ~n13152 ) | ( n13140 & n13463 ) | ( ~n13152 & n13463 ) ;
  assign n13465 = n4974 & ~n11273 ;
  assign n13466 = n5398 & n9965 ;
  assign n13467 = n4973 & n9969 ;
  assign n13468 = n4972 & ~n9967 ;
  assign n13469 = n13467 | n13468 ;
  assign n13470 = ( ~n13465 & n13466 ) | ( ~n13465 & n13469 ) | ( n13466 & n13469 ) ;
  assign n13471 = ( ~x20 & n13465 ) | ( ~x20 & n13470 ) | ( n13465 & n13470 ) ;
  assign n13472 = ( n13465 & n13470 ) | ( n13465 & ~n13471 ) | ( n13470 & ~n13471 ) ;
  assign n13473 = ( x20 & n13471 ) | ( x20 & ~n13472 ) | ( n13471 & ~n13472 ) ;
  assign n13474 = ( n13462 & n13464 ) | ( n13462 & n13473 ) | ( n13464 & n13473 ) ;
  assign n13475 = ( ~n13152 & n13161 ) | ( ~n13152 & n13163 ) | ( n13161 & n13163 ) ;
  assign n13476 = ( n13152 & ~n13164 ) | ( n13152 & n13475 ) | ( ~n13164 & n13475 ) ;
  assign n13477 = n4974 & ~n11121 ;
  assign n13478 = n5398 & ~n9963 ;
  assign n13479 = n4973 & ~n9967 ;
  assign n13480 = n4972 & n9965 ;
  assign n13481 = n13479 | n13480 ;
  assign n13482 = ( ~n13477 & n13478 ) | ( ~n13477 & n13481 ) | ( n13478 & n13481 ) ;
  assign n13483 = ( ~x20 & n13477 ) | ( ~x20 & n13482 ) | ( n13477 & n13482 ) ;
  assign n13484 = ( n13477 & n13482 ) | ( n13477 & ~n13483 ) | ( n13482 & ~n13483 ) ;
  assign n13485 = ( x20 & n13483 ) | ( x20 & ~n13484 ) | ( n13483 & ~n13484 ) ;
  assign n13486 = ( n13474 & n13476 ) | ( n13474 & n13485 ) | ( n13476 & n13485 ) ;
  assign n13487 = ( ~n13164 & n13173 ) | ( ~n13164 & n13175 ) | ( n13173 & n13175 ) ;
  assign n13488 = ( n13164 & ~n13176 ) | ( n13164 & n13487 ) | ( ~n13176 & n13487 ) ;
  assign n13489 = n4974 & ~n10929 ;
  assign n13490 = n5398 & n9961 ;
  assign n13491 = n4973 & n9965 ;
  assign n13492 = n4972 & ~n9963 ;
  assign n13493 = n13491 | n13492 ;
  assign n13494 = ( ~n13489 & n13490 ) | ( ~n13489 & n13493 ) | ( n13490 & n13493 ) ;
  assign n13495 = ( ~x20 & n13489 ) | ( ~x20 & n13494 ) | ( n13489 & n13494 ) ;
  assign n13496 = ( n13489 & n13494 ) | ( n13489 & ~n13495 ) | ( n13494 & ~n13495 ) ;
  assign n13497 = ( x20 & n13495 ) | ( x20 & ~n13496 ) | ( n13495 & ~n13496 ) ;
  assign n13498 = ( n13486 & n13488 ) | ( n13486 & n13497 ) | ( n13488 & n13497 ) ;
  assign n13499 = ( ~n13176 & n13185 ) | ( ~n13176 & n13187 ) | ( n13185 & n13187 ) ;
  assign n13500 = ( n13176 & ~n13188 ) | ( n13176 & n13499 ) | ( ~n13188 & n13499 ) ;
  assign n13501 = n4974 & n10859 ;
  assign n13502 = n5398 & n9959 ;
  assign n13503 = n4973 & ~n9963 ;
  assign n13504 = n4972 & n9961 ;
  assign n13505 = n13503 | n13504 ;
  assign n13506 = ( ~n13501 & n13502 ) | ( ~n13501 & n13505 ) | ( n13502 & n13505 ) ;
  assign n13507 = ( ~x20 & n13501 ) | ( ~x20 & n13506 ) | ( n13501 & n13506 ) ;
  assign n13508 = ( n13501 & n13506 ) | ( n13501 & ~n13507 ) | ( n13506 & ~n13507 ) ;
  assign n13509 = ( x20 & n13507 ) | ( x20 & ~n13508 ) | ( n13507 & ~n13508 ) ;
  assign n13510 = ( n13498 & n13500 ) | ( n13498 & n13509 ) | ( n13500 & n13509 ) ;
  assign n13511 = ( ~n13188 & n13190 ) | ( ~n13188 & n13199 ) | ( n13190 & n13199 ) ;
  assign n13512 = ( ~n13199 & n13200 ) | ( ~n13199 & n13511 ) | ( n13200 & n13511 ) ;
  assign n13513 = n5508 & ~n10652 ;
  assign n13514 = n5507 & n9951 ;
  assign n13515 = n5504 & n9955 ;
  assign n13516 = n5666 & ~n9953 ;
  assign n13517 = n13515 | n13516 ;
  assign n13518 = ( ~n13513 & n13514 ) | ( ~n13513 & n13517 ) | ( n13514 & n13517 ) ;
  assign n13519 = ( ~x17 & n13513 ) | ( ~x17 & n13518 ) | ( n13513 & n13518 ) ;
  assign n13520 = ( n13513 & n13518 ) | ( n13513 & ~n13519 ) | ( n13518 & ~n13519 ) ;
  assign n13521 = ( x17 & n13519 ) | ( x17 & ~n13520 ) | ( n13519 & ~n13520 ) ;
  assign n13522 = ( n13510 & ~n13512 ) | ( n13510 & n13521 ) | ( ~n13512 & n13521 ) ;
  assign n13523 = ( n13200 & ~n13202 ) | ( n13200 & n13211 ) | ( ~n13202 & n13211 ) ;
  assign n13524 = ( n13202 & ~n13212 ) | ( n13202 & n13523 ) | ( ~n13212 & n13523 ) ;
  assign n13525 = n5966 & n10271 ;
  assign n13526 = n6464 & n9943 ;
  assign n13527 = n5970 & n9947 ;
  assign n13528 = n5969 & n9945 ;
  assign n13529 = n13527 | n13528 ;
  assign n13530 = ( ~n13525 & n13526 ) | ( ~n13525 & n13529 ) | ( n13526 & n13529 ) ;
  assign n13531 = ( ~x14 & n13525 ) | ( ~x14 & n13530 ) | ( n13525 & n13530 ) ;
  assign n13532 = ( n13525 & n13530 ) | ( n13525 & ~n13531 ) | ( n13530 & ~n13531 ) ;
  assign n13533 = ( x14 & n13531 ) | ( x14 & ~n13532 ) | ( n13531 & ~n13532 ) ;
  assign n13534 = ( n13522 & n13524 ) | ( n13522 & n13533 ) | ( n13524 & n13533 ) ;
  assign n13535 = ( ~n13212 & n13214 ) | ( ~n13212 & n13223 ) | ( n13214 & n13223 ) ;
  assign n13536 = ( ~n13223 & n13224 ) | ( ~n13223 & n13535 ) | ( n13224 & n13535 ) ;
  assign n13537 = n6584 & n10040 ;
  assign n13538 = n7022 & ~n9937 ;
  assign n13539 = n6588 & ~n9883 ;
  assign n13540 = n6587 & n9916 ;
  assign n13541 = n13539 | n13540 ;
  assign n13542 = ( ~n13537 & n13538 ) | ( ~n13537 & n13541 ) | ( n13538 & n13541 ) ;
  assign n13543 = ( ~x11 & n13537 ) | ( ~x11 & n13542 ) | ( n13537 & n13542 ) ;
  assign n13544 = ( n13537 & n13542 ) | ( n13537 & ~n13543 ) | ( n13542 & ~n13543 ) ;
  assign n13545 = ( x11 & n13543 ) | ( x11 & ~n13544 ) | ( n13543 & ~n13544 ) ;
  assign n13546 = ( n13534 & ~n13536 ) | ( n13534 & n13545 ) | ( ~n13536 & n13545 ) ;
  assign n13547 = ( ~n13224 & n13226 ) | ( ~n13224 & n13235 ) | ( n13226 & n13235 ) ;
  assign n13548 = ( ~n13235 & n13236 ) | ( ~n13235 & n13547 ) | ( n13236 & n13547 ) ;
  assign n13549 = n6584 & ~n10064 ;
  assign n13550 = n7022 & ~n10057 ;
  assign n13551 = n6588 & n9916 ;
  assign n13552 = n6587 & ~n9937 ;
  assign n13553 = n13551 | n13552 ;
  assign n13554 = ( ~n13549 & n13550 ) | ( ~n13549 & n13553 ) | ( n13550 & n13553 ) ;
  assign n13555 = ( ~x11 & n13549 ) | ( ~x11 & n13554 ) | ( n13549 & n13554 ) ;
  assign n13556 = ( n13549 & n13554 ) | ( n13549 & ~n13555 ) | ( n13554 & ~n13555 ) ;
  assign n13557 = ( x11 & n13555 ) | ( x11 & ~n13556 ) | ( n13555 & ~n13556 ) ;
  assign n13558 = ( n13546 & ~n13548 ) | ( n13546 & n13557 ) | ( ~n13548 & n13557 ) ;
  assign n13559 = ( n13236 & ~n13238 ) | ( n13236 & n13247 ) | ( ~n13238 & n13247 ) ;
  assign n13560 = ( n13238 & ~n13248 ) | ( n13238 & n13559 ) | ( ~n13248 & n13559 ) ;
  assign n13561 = ~n7300 & n10346 ;
  assign n13562 = ( n10346 & n11065 ) | ( n10346 & ~n13561 ) | ( n11065 & ~n13561 ) ;
  assign n13563 = ( ~x8 & n7296 ) | ( ~x8 & n13562 ) | ( n7296 & n13562 ) ;
  assign n13564 = ( n7296 & n13562 ) | ( n7296 & ~n13563 ) | ( n13562 & ~n13563 ) ;
  assign n13565 = ( x8 & n13563 ) | ( x8 & ~n13564 ) | ( n13563 & ~n13564 ) ;
  assign n13566 = ( n13558 & n13560 ) | ( n13558 & n13565 ) | ( n13560 & n13565 ) ;
  assign n13567 = n5508 & n11892 ;
  assign n13568 = n5507 & ~n9997 ;
  assign n13569 = n5504 & ~n10001 ;
  assign n13570 = n5666 & n9999 ;
  assign n13571 = n13569 | n13570 ;
  assign n13572 = ( ~n13567 & n13568 ) | ( ~n13567 & n13571 ) | ( n13568 & n13571 ) ;
  assign n13573 = ( ~x17 & n13567 ) | ( ~x17 & n13572 ) | ( n13567 & n13572 ) ;
  assign n13574 = ( n13567 & n13572 ) | ( n13567 & ~n13573 ) | ( n13572 & ~n13573 ) ;
  assign n13575 = ( x17 & n13573 ) | ( x17 & ~n13574 ) | ( n13573 & ~n13574 ) ;
  assign n13576 = n5504 & ~n10003 ;
  assign n13577 = n5666 & ~n10001 ;
  assign n13578 = n13576 | n13577 ;
  assign n13579 = n5507 & ~n9999 ;
  assign n13580 = ( n5507 & n13578 ) | ( n5507 & ~n13579 ) | ( n13578 & ~n13579 ) ;
  assign n13581 = n5508 & n11868 ;
  assign n13582 = n13580 | n13581 ;
  assign n13583 = n5506 & ~n10003 ;
  assign n13584 = x17 & n13583 ;
  assign n13585 = ( n5508 & n11804 ) | ( n5508 & n11805 ) | ( n11804 & n11805 ) ;
  assign n13586 = n5666 | n10003 ;
  assign n13587 = n5507 & ~n10001 ;
  assign n13588 = ( ~n10003 & n13586 ) | ( ~n10003 & n13587 ) | ( n13586 & n13587 ) ;
  assign n13589 = n13585 | n13588 ;
  assign n13590 = ( x17 & n13584 ) | ( x17 & n13589 ) | ( n13584 & n13589 ) ;
  assign n13591 = n13582 | n13590 ;
  assign n13592 = x17 & ~n13591 ;
  assign n13593 = ( n13271 & n13575 ) | ( n13271 & n13592 ) | ( n13575 & n13592 ) ;
  assign n13594 = n5508 & n11934 ;
  assign n13595 = n5507 & n9995 ;
  assign n13596 = n5504 & n9999 ;
  assign n13597 = n5666 & ~n9997 ;
  assign n13598 = n13596 | n13597 ;
  assign n13599 = ( ~n13594 & n13595 ) | ( ~n13594 & n13598 ) | ( n13595 & n13598 ) ;
  assign n13600 = ( ~x17 & n13594 ) | ( ~x17 & n13599 ) | ( n13594 & n13599 ) ;
  assign n13601 = ( n13594 & n13599 ) | ( n13594 & ~n13600 ) | ( n13599 & ~n13600 ) ;
  assign n13602 = ( x17 & n13600 ) | ( x17 & ~n13601 ) | ( n13600 & ~n13601 ) ;
  assign n13603 = ( n13272 & n13273 ) | ( n13272 & n13276 ) | ( n13273 & n13276 ) ;
  assign n13604 = ~n13272 & n13277 ;
  assign n13605 = ( n13272 & ~n13603 ) | ( n13272 & n13604 ) | ( ~n13603 & n13604 ) ;
  assign n13606 = ( n13593 & n13602 ) | ( n13593 & n13605 ) | ( n13602 & n13605 ) ;
  assign n13607 = n5508 & ~n11971 ;
  assign n13608 = n5507 & n9993 ;
  assign n13609 = n5504 & ~n9997 ;
  assign n13610 = n5666 & n9995 ;
  assign n13611 = n13609 | n13610 ;
  assign n13612 = ( ~n13607 & n13608 ) | ( ~n13607 & n13611 ) | ( n13608 & n13611 ) ;
  assign n13613 = ( ~x17 & n13607 ) | ( ~x17 & n13612 ) | ( n13607 & n13612 ) ;
  assign n13614 = ( n13607 & n13612 ) | ( n13607 & ~n13613 ) | ( n13612 & ~n13613 ) ;
  assign n13615 = ( x17 & n13613 ) | ( x17 & ~n13614 ) | ( n13613 & ~n13614 ) ;
  assign n13616 = ( n13270 & n13278 ) | ( n13270 & ~n13279 ) | ( n13278 & ~n13279 ) ;
  assign n13617 = n13279 & ~n13616 ;
  assign n13618 = ( n13606 & n13615 ) | ( n13606 & n13617 ) | ( n13615 & n13617 ) ;
  assign n13619 = n5508 & n12026 ;
  assign n13620 = n5507 & n9991 ;
  assign n13621 = n5504 & n9995 ;
  assign n13622 = n5666 & n9993 ;
  assign n13623 = n13621 | n13622 ;
  assign n13624 = ( ~n13619 & n13620 ) | ( ~n13619 & n13623 ) | ( n13620 & n13623 ) ;
  assign n13625 = ( ~x17 & n13619 ) | ( ~x17 & n13624 ) | ( n13619 & n13624 ) ;
  assign n13626 = ( n13619 & n13624 ) | ( n13619 & ~n13625 ) | ( n13624 & ~n13625 ) ;
  assign n13627 = ( x17 & n13625 ) | ( x17 & ~n13626 ) | ( n13625 & ~n13626 ) ;
  assign n13628 = ( n12986 & n13263 ) | ( n12986 & ~n13280 ) | ( n13263 & ~n13280 ) ;
  assign n13629 = ( n13280 & ~n13281 ) | ( n13280 & n13628 ) | ( ~n13281 & n13628 ) ;
  assign n13630 = ( n13618 & n13627 ) | ( n13618 & n13629 ) | ( n13627 & n13629 ) ;
  assign n13631 = n5508 & n12050 ;
  assign n13632 = n5507 & n9989 ;
  assign n13633 = n5504 & n9993 ;
  assign n13634 = n5666 & n9991 ;
  assign n13635 = n13633 | n13634 ;
  assign n13636 = ( ~n13631 & n13632 ) | ( ~n13631 & n13635 ) | ( n13632 & n13635 ) ;
  assign n13637 = ( ~x17 & n13631 ) | ( ~x17 & n13636 ) | ( n13631 & n13636 ) ;
  assign n13638 = ( n13631 & n13636 ) | ( n13631 & ~n13637 ) | ( n13636 & ~n13637 ) ;
  assign n13639 = ( x17 & n13637 ) | ( x17 & ~n13638 ) | ( n13637 & ~n13638 ) ;
  assign n13640 = ( ~n13281 & n13290 ) | ( ~n13281 & n13293 ) | ( n13290 & n13293 ) ;
  assign n13641 = ( n13281 & ~n13294 ) | ( n13281 & n13640 ) | ( ~n13294 & n13640 ) ;
  assign n13642 = ( n13630 & n13639 ) | ( n13630 & n13641 ) | ( n13639 & n13641 ) ;
  assign n13643 = ( ~n13294 & n13303 ) | ( ~n13294 & n13305 ) | ( n13303 & n13305 ) ;
  assign n13644 = ( n13294 & ~n13306 ) | ( n13294 & n13643 ) | ( ~n13306 & n13643 ) ;
  assign n13645 = n5508 & ~n12074 ;
  assign n13646 = n5507 & ~n9987 ;
  assign n13647 = n5504 & n9991 ;
  assign n13648 = n5666 & n9989 ;
  assign n13649 = n13647 | n13648 ;
  assign n13650 = ( ~n13645 & n13646 ) | ( ~n13645 & n13649 ) | ( n13646 & n13649 ) ;
  assign n13651 = ( ~x17 & n13645 ) | ( ~x17 & n13650 ) | ( n13645 & n13650 ) ;
  assign n13652 = ( n13645 & n13650 ) | ( n13645 & ~n13651 ) | ( n13650 & ~n13651 ) ;
  assign n13653 = ( x17 & n13651 ) | ( x17 & ~n13652 ) | ( n13651 & ~n13652 ) ;
  assign n13654 = ( n13642 & n13644 ) | ( n13642 & n13653 ) | ( n13644 & n13653 ) ;
  assign n13655 = ( ~n13306 & n13315 ) | ( ~n13306 & n13317 ) | ( n13315 & n13317 ) ;
  assign n13656 = ( n13306 & ~n13318 ) | ( n13306 & n13655 ) | ( ~n13318 & n13655 ) ;
  assign n13657 = n5508 & ~n12099 ;
  assign n13658 = n5507 & n9985 ;
  assign n13659 = n5504 & n9989 ;
  assign n13660 = n5666 & ~n9987 ;
  assign n13661 = n13659 | n13660 ;
  assign n13662 = ( ~n13657 & n13658 ) | ( ~n13657 & n13661 ) | ( n13658 & n13661 ) ;
  assign n13663 = ( ~x17 & n13657 ) | ( ~x17 & n13662 ) | ( n13657 & n13662 ) ;
  assign n13664 = ( n13657 & n13662 ) | ( n13657 & ~n13663 ) | ( n13662 & ~n13663 ) ;
  assign n13665 = ( x17 & n13663 ) | ( x17 & ~n13664 ) | ( n13663 & ~n13664 ) ;
  assign n13666 = ( n13654 & n13656 ) | ( n13654 & n13665 ) | ( n13656 & n13665 ) ;
  assign n13667 = ( ~n13318 & n13327 ) | ( ~n13318 & n13329 ) | ( n13327 & n13329 ) ;
  assign n13668 = ( n13318 & ~n13330 ) | ( n13318 & n13667 ) | ( ~n13330 & n13667 ) ;
  assign n13669 = n5508 & ~n12129 ;
  assign n13670 = n5507 & ~n9983 ;
  assign n13671 = n5504 & ~n9987 ;
  assign n13672 = n5666 & n9985 ;
  assign n13673 = n13671 | n13672 ;
  assign n13674 = ( ~n13669 & n13670 ) | ( ~n13669 & n13673 ) | ( n13670 & n13673 ) ;
  assign n13675 = ( ~x17 & n13669 ) | ( ~x17 & n13674 ) | ( n13669 & n13674 ) ;
  assign n13676 = ( n13669 & n13674 ) | ( n13669 & ~n13675 ) | ( n13674 & ~n13675 ) ;
  assign n13677 = ( x17 & n13675 ) | ( x17 & ~n13676 ) | ( n13675 & ~n13676 ) ;
  assign n13678 = ( n13666 & n13668 ) | ( n13666 & n13677 ) | ( n13668 & n13677 ) ;
  assign n13679 = n5508 & ~n11561 ;
  assign n13680 = n5507 & n9981 ;
  assign n13681 = n5504 & n9985 ;
  assign n13682 = n5666 & ~n9983 ;
  assign n13683 = n13681 | n13682 ;
  assign n13684 = ( ~n13679 & n13680 ) | ( ~n13679 & n13683 ) | ( n13680 & n13683 ) ;
  assign n13685 = ( ~x17 & n13679 ) | ( ~x17 & n13684 ) | ( n13679 & n13684 ) ;
  assign n13686 = ( n13679 & n13684 ) | ( n13679 & ~n13685 ) | ( n13684 & ~n13685 ) ;
  assign n13687 = ( x17 & n13685 ) | ( x17 & ~n13686 ) | ( n13685 & ~n13686 ) ;
  assign n13688 = ( ~n13330 & n13332 ) | ( ~n13330 & n13341 ) | ( n13332 & n13341 ) ;
  assign n13689 = ( n13330 & ~n13342 ) | ( n13330 & n13688 ) | ( ~n13342 & n13688 ) ;
  assign n13690 = ( n13678 & n13687 ) | ( n13678 & n13689 ) | ( n13687 & n13689 ) ;
  assign n13691 = n5508 & n12153 ;
  assign n13692 = n5507 & n9979 ;
  assign n13693 = n5504 & ~n9983 ;
  assign n13694 = n5666 & n9981 ;
  assign n13695 = n13693 | n13694 ;
  assign n13696 = ( ~n13691 & n13692 ) | ( ~n13691 & n13695 ) | ( n13692 & n13695 ) ;
  assign n13697 = ( ~x17 & n13691 ) | ( ~x17 & n13696 ) | ( n13691 & n13696 ) ;
  assign n13698 = ( n13691 & n13696 ) | ( n13691 & ~n13697 ) | ( n13696 & ~n13697 ) ;
  assign n13699 = ( x17 & n13697 ) | ( x17 & ~n13698 ) | ( n13697 & ~n13698 ) ;
  assign n13700 = ( ~n13342 & n13344 ) | ( ~n13342 & n13353 ) | ( n13344 & n13353 ) ;
  assign n13701 = ( n13342 & ~n13354 ) | ( n13342 & n13700 ) | ( ~n13354 & n13700 ) ;
  assign n13702 = ( n13690 & n13699 ) | ( n13690 & n13701 ) | ( n13699 & n13701 ) ;
  assign n13703 = n5508 & n12165 ;
  assign n13704 = n5507 & n9977 ;
  assign n13705 = n5504 & n9981 ;
  assign n13706 = n5666 & n9979 ;
  assign n13707 = n13705 | n13706 ;
  assign n13708 = ( ~n13703 & n13704 ) | ( ~n13703 & n13707 ) | ( n13704 & n13707 ) ;
  assign n13709 = ( ~x17 & n13703 ) | ( ~x17 & n13708 ) | ( n13703 & n13708 ) ;
  assign n13710 = ( n13703 & n13708 ) | ( n13703 & ~n13709 ) | ( n13708 & ~n13709 ) ;
  assign n13711 = ( x17 & n13709 ) | ( x17 & ~n13710 ) | ( n13709 & ~n13710 ) ;
  assign n13712 = ( ~n13354 & n13356 ) | ( ~n13354 & n13365 ) | ( n13356 & n13365 ) ;
  assign n13713 = ( n13354 & ~n13366 ) | ( n13354 & n13712 ) | ( ~n13366 & n13712 ) ;
  assign n13714 = ( n13702 & n13711 ) | ( n13702 & n13713 ) | ( n13711 & n13713 ) ;
  assign n13715 = ( ~n13366 & n13375 ) | ( ~n13366 & n13377 ) | ( n13375 & n13377 ) ;
  assign n13716 = ( n13366 & ~n13378 ) | ( n13366 & n13715 ) | ( ~n13378 & n13715 ) ;
  assign n13717 = n5508 & n11606 ;
  assign n13718 = n5507 & n9975 ;
  assign n13719 = n5504 & n9979 ;
  assign n13720 = n5666 & n9977 ;
  assign n13721 = n13719 | n13720 ;
  assign n13722 = ( ~n13717 & n13718 ) | ( ~n13717 & n13721 ) | ( n13718 & n13721 ) ;
  assign n13723 = ( ~x17 & n13717 ) | ( ~x17 & n13722 ) | ( n13717 & n13722 ) ;
  assign n13724 = ( n13717 & n13722 ) | ( n13717 & ~n13723 ) | ( n13722 & ~n13723 ) ;
  assign n13725 = ( x17 & n13723 ) | ( x17 & ~n13724 ) | ( n13723 & ~n13724 ) ;
  assign n13726 = ( n13714 & n13716 ) | ( n13714 & n13725 ) | ( n13716 & n13725 ) ;
  assign n13727 = ( ~n13378 & n13387 ) | ( ~n13378 & n13389 ) | ( n13387 & n13389 ) ;
  assign n13728 = ( n13378 & ~n13390 ) | ( n13378 & n13727 ) | ( ~n13390 & n13727 ) ;
  assign n13729 = n5508 & n11400 ;
  assign n13730 = n5507 & n9973 ;
  assign n13731 = n5504 & n9977 ;
  assign n13732 = n5666 & n9975 ;
  assign n13733 = n13731 | n13732 ;
  assign n13734 = ( ~n13729 & n13730 ) | ( ~n13729 & n13733 ) | ( n13730 & n13733 ) ;
  assign n13735 = ( ~x17 & n13729 ) | ( ~x17 & n13734 ) | ( n13729 & n13734 ) ;
  assign n13736 = ( n13729 & n13734 ) | ( n13729 & ~n13735 ) | ( n13734 & ~n13735 ) ;
  assign n13737 = ( x17 & n13735 ) | ( x17 & ~n13736 ) | ( n13735 & ~n13736 ) ;
  assign n13738 = ( n13726 & n13728 ) | ( n13726 & n13737 ) | ( n13728 & n13737 ) ;
  assign n13739 = n5508 & n11630 ;
  assign n13740 = n5507 & n9971 ;
  assign n13741 = n5504 & n9975 ;
  assign n13742 = n5666 & n9973 ;
  assign n13743 = n13741 | n13742 ;
  assign n13744 = ( ~n13739 & n13740 ) | ( ~n13739 & n13743 ) | ( n13740 & n13743 ) ;
  assign n13745 = ( ~x17 & n13739 ) | ( ~x17 & n13744 ) | ( n13739 & n13744 ) ;
  assign n13746 = ( n13739 & n13744 ) | ( n13739 & ~n13745 ) | ( n13744 & ~n13745 ) ;
  assign n13747 = ( x17 & n13745 ) | ( x17 & ~n13746 ) | ( n13745 & ~n13746 ) ;
  assign n13748 = ( ~n13390 & n13392 ) | ( ~n13390 & n13401 ) | ( n13392 & n13401 ) ;
  assign n13749 = ( ~n13401 & n13402 ) | ( ~n13401 & n13748 ) | ( n13402 & n13748 ) ;
  assign n13750 = ( n13738 & n13747 ) | ( n13738 & ~n13749 ) | ( n13747 & ~n13749 ) ;
  assign n13751 = n5508 & n11428 ;
  assign n13752 = n5507 & n9969 ;
  assign n13753 = n5504 & n9973 ;
  assign n13754 = n5666 & n9971 ;
  assign n13755 = n13753 | n13754 ;
  assign n13756 = ( ~n13751 & n13752 ) | ( ~n13751 & n13755 ) | ( n13752 & n13755 ) ;
  assign n13757 = ( ~x17 & n13751 ) | ( ~x17 & n13756 ) | ( n13751 & n13756 ) ;
  assign n13758 = ( n13751 & n13756 ) | ( n13751 & ~n13757 ) | ( n13756 & ~n13757 ) ;
  assign n13759 = ( x17 & n13757 ) | ( x17 & ~n13758 ) | ( n13757 & ~n13758 ) ;
  assign n13760 = ( ~n13402 & n13404 ) | ( ~n13402 & n13413 ) | ( n13404 & n13413 ) ;
  assign n13761 = ( ~n13413 & n13414 ) | ( ~n13413 & n13760 ) | ( n13414 & n13760 ) ;
  assign n13762 = ( n13750 & n13759 ) | ( n13750 & ~n13761 ) | ( n13759 & ~n13761 ) ;
  assign n13763 = n5508 & ~n10998 ;
  assign n13764 = n5507 & ~n9967 ;
  assign n13765 = n5504 & n9971 ;
  assign n13766 = n5666 & n9969 ;
  assign n13767 = n13765 | n13766 ;
  assign n13768 = ( ~n13763 & n13764 ) | ( ~n13763 & n13767 ) | ( n13764 & n13767 ) ;
  assign n13769 = ( ~x17 & n13763 ) | ( ~x17 & n13768 ) | ( n13763 & n13768 ) ;
  assign n13770 = ( n13763 & n13768 ) | ( n13763 & ~n13769 ) | ( n13768 & ~n13769 ) ;
  assign n13771 = ( x17 & n13769 ) | ( x17 & ~n13770 ) | ( n13769 & ~n13770 ) ;
  assign n13772 = ( ~n13414 & n13416 ) | ( ~n13414 & n13425 ) | ( n13416 & n13425 ) ;
  assign n13773 = ( n13414 & ~n13426 ) | ( n13414 & n13772 ) | ( ~n13426 & n13772 ) ;
  assign n13774 = ( n13762 & n13771 ) | ( n13762 & n13773 ) | ( n13771 & n13773 ) ;
  assign n13775 = n5508 & ~n11273 ;
  assign n13776 = n5507 & n9965 ;
  assign n13777 = n5504 & n9969 ;
  assign n13778 = n5666 & ~n9967 ;
  assign n13779 = n13777 | n13778 ;
  assign n13780 = ( ~n13775 & n13776 ) | ( ~n13775 & n13779 ) | ( n13776 & n13779 ) ;
  assign n13781 = ( ~x17 & n13775 ) | ( ~x17 & n13780 ) | ( n13775 & n13780 ) ;
  assign n13782 = ( n13775 & n13780 ) | ( n13775 & ~n13781 ) | ( n13780 & ~n13781 ) ;
  assign n13783 = ( x17 & n13781 ) | ( x17 & ~n13782 ) | ( n13781 & ~n13782 ) ;
  assign n13784 = ( ~n13426 & n13428 ) | ( ~n13426 & n13437 ) | ( n13428 & n13437 ) ;
  assign n13785 = ( ~n13437 & n13438 ) | ( ~n13437 & n13784 ) | ( n13438 & n13784 ) ;
  assign n13786 = ( n13774 & n13783 ) | ( n13774 & ~n13785 ) | ( n13783 & ~n13785 ) ;
  assign n13787 = n5508 & ~n11121 ;
  assign n13788 = n5507 & ~n9963 ;
  assign n13789 = n5504 & ~n9967 ;
  assign n13790 = n5666 & n9965 ;
  assign n13791 = n13789 | n13790 ;
  assign n13792 = ( ~n13787 & n13788 ) | ( ~n13787 & n13791 ) | ( n13788 & n13791 ) ;
  assign n13793 = ( ~x17 & n13787 ) | ( ~x17 & n13792 ) | ( n13787 & n13792 ) ;
  assign n13794 = ( n13787 & n13792 ) | ( n13787 & ~n13793 ) | ( n13792 & ~n13793 ) ;
  assign n13795 = ( x17 & n13793 ) | ( x17 & ~n13794 ) | ( n13793 & ~n13794 ) ;
  assign n13796 = ( ~n13438 & n13440 ) | ( ~n13438 & n13449 ) | ( n13440 & n13449 ) ;
  assign n13797 = ( ~n13449 & n13450 ) | ( ~n13449 & n13796 ) | ( n13450 & n13796 ) ;
  assign n13798 = ( n13786 & n13795 ) | ( n13786 & ~n13797 ) | ( n13795 & ~n13797 ) ;
  assign n13799 = n5508 & ~n10929 ;
  assign n13800 = n5507 & n9961 ;
  assign n13801 = n5504 & n9965 ;
  assign n13802 = n5666 & ~n9963 ;
  assign n13803 = n13801 | n13802 ;
  assign n13804 = ( ~n13799 & n13800 ) | ( ~n13799 & n13803 ) | ( n13800 & n13803 ) ;
  assign n13805 = ( ~x17 & n13799 ) | ( ~x17 & n13804 ) | ( n13799 & n13804 ) ;
  assign n13806 = ( n13799 & n13804 ) | ( n13799 & ~n13805 ) | ( n13804 & ~n13805 ) ;
  assign n13807 = ( x17 & n13805 ) | ( x17 & ~n13806 ) | ( n13805 & ~n13806 ) ;
  assign n13808 = ( ~n13450 & n13452 ) | ( ~n13450 & n13461 ) | ( n13452 & n13461 ) ;
  assign n13809 = ( n13450 & ~n13462 ) | ( n13450 & n13808 ) | ( ~n13462 & n13808 ) ;
  assign n13810 = ( n13798 & n13807 ) | ( n13798 & n13809 ) | ( n13807 & n13809 ) ;
  assign n13811 = n5508 & n10859 ;
  assign n13812 = n5507 & n9959 ;
  assign n13813 = n5504 & ~n9963 ;
  assign n13814 = n5666 & n9961 ;
  assign n13815 = n13813 | n13814 ;
  assign n13816 = ( ~n13811 & n13812 ) | ( ~n13811 & n13815 ) | ( n13812 & n13815 ) ;
  assign n13817 = ( ~x17 & n13811 ) | ( ~x17 & n13816 ) | ( n13811 & n13816 ) ;
  assign n13818 = ( n13811 & n13816 ) | ( n13811 & ~n13817 ) | ( n13816 & ~n13817 ) ;
  assign n13819 = ( x17 & n13817 ) | ( x17 & ~n13818 ) | ( n13817 & ~n13818 ) ;
  assign n13820 = ( ~n13462 & n13464 ) | ( ~n13462 & n13473 ) | ( n13464 & n13473 ) ;
  assign n13821 = ( n13462 & ~n13474 ) | ( n13462 & n13820 ) | ( ~n13474 & n13820 ) ;
  assign n13822 = ( n13810 & n13819 ) | ( n13810 & n13821 ) | ( n13819 & n13821 ) ;
  assign n13823 = n5508 & ~n10869 ;
  assign n13824 = n5507 & ~n9957 ;
  assign n13825 = n5504 & n9961 ;
  assign n13826 = n5666 & n9959 ;
  assign n13827 = n13825 | n13826 ;
  assign n13828 = ( ~n13823 & n13824 ) | ( ~n13823 & n13827 ) | ( n13824 & n13827 ) ;
  assign n13829 = ( ~x17 & n13823 ) | ( ~x17 & n13828 ) | ( n13823 & n13828 ) ;
  assign n13830 = ( n13823 & n13828 ) | ( n13823 & ~n13829 ) | ( n13828 & ~n13829 ) ;
  assign n13831 = ( x17 & n13829 ) | ( x17 & ~n13830 ) | ( n13829 & ~n13830 ) ;
  assign n13832 = ( ~n13474 & n13476 ) | ( ~n13474 & n13485 ) | ( n13476 & n13485 ) ;
  assign n13833 = ( n13474 & ~n13486 ) | ( n13474 & n13832 ) | ( ~n13486 & n13832 ) ;
  assign n13834 = ( n13822 & n13831 ) | ( n13822 & n13833 ) | ( n13831 & n13833 ) ;
  assign n13835 = n5508 & ~n10567 ;
  assign n13836 = n5507 & n9955 ;
  assign n13837 = n5504 & n9959 ;
  assign n13838 = n5666 & ~n9957 ;
  assign n13839 = n13837 | n13838 ;
  assign n13840 = ( ~n13835 & n13836 ) | ( ~n13835 & n13839 ) | ( n13836 & n13839 ) ;
  assign n13841 = ( ~x17 & n13835 ) | ( ~x17 & n13840 ) | ( n13835 & n13840 ) ;
  assign n13842 = ( n13835 & n13840 ) | ( n13835 & ~n13841 ) | ( n13840 & ~n13841 ) ;
  assign n13843 = ( x17 & n13841 ) | ( x17 & ~n13842 ) | ( n13841 & ~n13842 ) ;
  assign n13844 = ( ~n13486 & n13488 ) | ( ~n13486 & n13497 ) | ( n13488 & n13497 ) ;
  assign n13845 = ( n13486 & ~n13498 ) | ( n13486 & n13844 ) | ( ~n13498 & n13844 ) ;
  assign n13846 = ( n13834 & n13843 ) | ( n13834 & n13845 ) | ( n13843 & n13845 ) ;
  assign n13847 = n5508 & ~n10750 ;
  assign n13848 = n5507 & ~n9953 ;
  assign n13849 = n5504 & ~n9957 ;
  assign n13850 = n5666 & n9955 ;
  assign n13851 = n13849 | n13850 ;
  assign n13852 = ( ~n13847 & n13848 ) | ( ~n13847 & n13851 ) | ( n13848 & n13851 ) ;
  assign n13853 = ( ~x17 & n13847 ) | ( ~x17 & n13852 ) | ( n13847 & n13852 ) ;
  assign n13854 = ( n13847 & n13852 ) | ( n13847 & ~n13853 ) | ( n13852 & ~n13853 ) ;
  assign n13855 = ( x17 & n13853 ) | ( x17 & ~n13854 ) | ( n13853 & ~n13854 ) ;
  assign n13856 = ( ~n13498 & n13500 ) | ( ~n13498 & n13509 ) | ( n13500 & n13509 ) ;
  assign n13857 = ( n13498 & ~n13510 ) | ( n13498 & n13856 ) | ( ~n13510 & n13856 ) ;
  assign n13858 = ( n13846 & n13855 ) | ( n13846 & n13857 ) | ( n13855 & n13857 ) ;
  assign n13859 = ( ~n13510 & n13512 ) | ( ~n13510 & n13521 ) | ( n13512 & n13521 ) ;
  assign n13860 = ( ~n13521 & n13522 ) | ( ~n13521 & n13859 ) | ( n13522 & n13859 ) ;
  assign n13861 = n5966 & n10466 ;
  assign n13862 = n6464 & n9945 ;
  assign n13863 = n5970 & n9949 ;
  assign n13864 = n5969 & n9947 ;
  assign n13865 = n13863 | n13864 ;
  assign n13866 = ( ~n13861 & n13862 ) | ( ~n13861 & n13865 ) | ( n13862 & n13865 ) ;
  assign n13867 = ( ~x14 & n13861 ) | ( ~x14 & n13866 ) | ( n13861 & n13866 ) ;
  assign n13868 = ( n13861 & n13866 ) | ( n13861 & ~n13867 ) | ( n13866 & ~n13867 ) ;
  assign n13869 = ( x14 & n13867 ) | ( x14 & ~n13868 ) | ( n13867 & ~n13868 ) ;
  assign n13870 = ( n13858 & ~n13860 ) | ( n13858 & n13869 ) | ( ~n13860 & n13869 ) ;
  assign n13871 = ( n13522 & ~n13524 ) | ( n13522 & n13533 ) | ( ~n13524 & n13533 ) ;
  assign n13872 = ( n13524 & ~n13534 ) | ( n13524 & n13871 ) | ( ~n13534 & n13871 ) ;
  assign n13873 = n6584 & n10174 ;
  assign n13874 = n7022 & n9916 ;
  assign n13875 = n6587 | n9883 ;
  assign n13876 = n6588 & ~n9941 ;
  assign n13877 = ( ~n9883 & n13875 ) | ( ~n9883 & n13876 ) | ( n13875 & n13876 ) ;
  assign n13878 = ( ~n13873 & n13874 ) | ( ~n13873 & n13877 ) | ( n13874 & n13877 ) ;
  assign n13879 = ( ~x11 & n13873 ) | ( ~x11 & n13878 ) | ( n13873 & n13878 ) ;
  assign n13880 = ( n13873 & n13878 ) | ( n13873 & ~n13879 ) | ( n13878 & ~n13879 ) ;
  assign n13881 = ( x11 & n13879 ) | ( x11 & ~n13880 ) | ( n13879 & ~n13880 ) ;
  assign n13882 = ( n13870 & n13872 ) | ( n13870 & n13881 ) | ( n13872 & n13881 ) ;
  assign n13883 = ( ~n13534 & n13536 ) | ( ~n13534 & n13545 ) | ( n13536 & n13545 ) ;
  assign n13884 = ( ~n13545 & n13546 ) | ( ~n13545 & n13883 ) | ( n13546 & n13883 ) ;
  assign n13885 = n7296 & n10362 ;
  assign n13886 = n7879 & n10346 ;
  assign n13887 = n7300 & ~n10057 ;
  assign n13888 = n7299 & ~n10302 ;
  assign n13889 = n13887 | n13888 ;
  assign n13890 = ( ~n13885 & n13886 ) | ( ~n13885 & n13889 ) | ( n13886 & n13889 ) ;
  assign n13891 = ( ~x8 & n13885 ) | ( ~x8 & n13890 ) | ( n13885 & n13890 ) ;
  assign n13892 = ( n13885 & n13890 ) | ( n13885 & ~n13891 ) | ( n13890 & ~n13891 ) ;
  assign n13893 = ( x8 & n13891 ) | ( x8 & ~n13892 ) | ( n13891 & ~n13892 ) ;
  assign n13894 = ( n13882 & ~n13884 ) | ( n13882 & n13893 ) | ( ~n13884 & n13893 ) ;
  assign n13895 = n7296 & n10348 ;
  assign n13896 = n7299 & n10346 ;
  assign n13897 = n7300 & ~n10302 ;
  assign n13898 = n7879 | n13897 ;
  assign n13899 = ( ~n13895 & n13896 ) | ( ~n13895 & n13898 ) | ( n13896 & n13898 ) ;
  assign n13900 = ( ~x8 & n13895 ) | ( ~x8 & n13899 ) | ( n13895 & n13899 ) ;
  assign n13901 = ( n13895 & n13899 ) | ( n13895 & ~n13900 ) | ( n13899 & ~n13900 ) ;
  assign n13902 = ( x8 & n13900 ) | ( x8 & ~n13901 ) | ( n13900 & ~n13901 ) ;
  assign n13903 = ( ~n13546 & n13548 ) | ( ~n13546 & n13557 ) | ( n13548 & n13557 ) ;
  assign n13904 = ( ~n13557 & n13558 ) | ( ~n13557 & n13903 ) | ( n13558 & n13903 ) ;
  assign n13905 = ( n13894 & n13902 ) | ( n13894 & ~n13904 ) | ( n13902 & ~n13904 ) ;
  assign n13906 = n5966 & n11892 ;
  assign n13907 = n6464 & ~n9997 ;
  assign n13908 = n5970 & ~n10001 ;
  assign n13909 = n5969 & n9999 ;
  assign n13910 = n13908 | n13909 ;
  assign n13911 = ( ~n13906 & n13907 ) | ( ~n13906 & n13910 ) | ( n13907 & n13910 ) ;
  assign n13912 = ( ~x14 & n13906 ) | ( ~x14 & n13911 ) | ( n13906 & n13911 ) ;
  assign n13913 = ( n13906 & n13911 ) | ( n13906 & ~n13912 ) | ( n13911 & ~n13912 ) ;
  assign n13914 = ( x14 & n13912 ) | ( x14 & ~n13913 ) | ( n13912 & ~n13913 ) ;
  assign n13915 = n5970 & ~n10003 ;
  assign n13916 = n5969 & ~n10001 ;
  assign n13917 = n13915 | n13916 ;
  assign n13918 = n6464 & ~n9999 ;
  assign n13919 = ( n6464 & n13917 ) | ( n6464 & ~n13918 ) | ( n13917 & ~n13918 ) ;
  assign n13920 = n5966 & n11868 ;
  assign n13921 = n13919 | n13920 ;
  assign n13922 = n6463 & ~n10003 ;
  assign n13923 = x14 & n13922 ;
  assign n13924 = ( n5966 & n11804 ) | ( n5966 & n11805 ) | ( n11804 & n11805 ) ;
  assign n13925 = n5969 | n10003 ;
  assign n13926 = n6464 & ~n10001 ;
  assign n13927 = ( ~n10003 & n13925 ) | ( ~n10003 & n13926 ) | ( n13925 & n13926 ) ;
  assign n13928 = n13924 | n13927 ;
  assign n13929 = ( x14 & n13923 ) | ( x14 & n13928 ) | ( n13923 & n13928 ) ;
  assign n13930 = n13921 | n13929 ;
  assign n13931 = x14 & ~n13930 ;
  assign n13932 = ( n13583 & n13914 ) | ( n13583 & n13931 ) | ( n13914 & n13931 ) ;
  assign n13933 = n5966 & n11934 ;
  assign n13934 = n6464 & n9995 ;
  assign n13935 = n5970 & n9999 ;
  assign n13936 = n5969 & ~n9997 ;
  assign n13937 = n13935 | n13936 ;
  assign n13938 = ( ~n13933 & n13934 ) | ( ~n13933 & n13937 ) | ( n13934 & n13937 ) ;
  assign n13939 = ( ~x14 & n13933 ) | ( ~x14 & n13938 ) | ( n13933 & n13938 ) ;
  assign n13940 = ( n13933 & n13938 ) | ( n13933 & ~n13939 ) | ( n13938 & ~n13939 ) ;
  assign n13941 = ( x14 & n13939 ) | ( x14 & ~n13940 ) | ( n13939 & ~n13940 ) ;
  assign n13942 = ( n13584 & n13585 ) | ( n13584 & n13588 ) | ( n13585 & n13588 ) ;
  assign n13943 = ~n13584 & n13589 ;
  assign n13944 = ( n13584 & ~n13942 ) | ( n13584 & n13943 ) | ( ~n13942 & n13943 ) ;
  assign n13945 = ( n13932 & n13941 ) | ( n13932 & n13944 ) | ( n13941 & n13944 ) ;
  assign n13946 = n5966 & ~n11971 ;
  assign n13947 = n6464 & n9993 ;
  assign n13948 = n5970 & ~n9997 ;
  assign n13949 = n5969 & n9995 ;
  assign n13950 = n13948 | n13949 ;
  assign n13951 = ( ~n13946 & n13947 ) | ( ~n13946 & n13950 ) | ( n13947 & n13950 ) ;
  assign n13952 = ( ~x14 & n13946 ) | ( ~x14 & n13951 ) | ( n13946 & n13951 ) ;
  assign n13953 = ( n13946 & n13951 ) | ( n13946 & ~n13952 ) | ( n13951 & ~n13952 ) ;
  assign n13954 = ( x14 & n13952 ) | ( x14 & ~n13953 ) | ( n13952 & ~n13953 ) ;
  assign n13955 = ( n13582 & n13590 ) | ( n13582 & ~n13591 ) | ( n13590 & ~n13591 ) ;
  assign n13956 = n13591 & ~n13955 ;
  assign n13957 = ( n13945 & n13954 ) | ( n13945 & n13956 ) | ( n13954 & n13956 ) ;
  assign n13958 = n5966 & n12026 ;
  assign n13959 = n6464 & n9991 ;
  assign n13960 = n5970 & n9995 ;
  assign n13961 = n5969 & n9993 ;
  assign n13962 = n13960 | n13961 ;
  assign n13963 = ( ~n13958 & n13959 ) | ( ~n13958 & n13962 ) | ( n13959 & n13962 ) ;
  assign n13964 = ( ~x14 & n13958 ) | ( ~x14 & n13963 ) | ( n13958 & n13963 ) ;
  assign n13965 = ( n13958 & n13963 ) | ( n13958 & ~n13964 ) | ( n13963 & ~n13964 ) ;
  assign n13966 = ( x14 & n13964 ) | ( x14 & ~n13965 ) | ( n13964 & ~n13965 ) ;
  assign n13967 = ( n13271 & n13575 ) | ( n13271 & ~n13592 ) | ( n13575 & ~n13592 ) ;
  assign n13968 = ( n13592 & ~n13593 ) | ( n13592 & n13967 ) | ( ~n13593 & n13967 ) ;
  assign n13969 = ( n13957 & n13966 ) | ( n13957 & n13968 ) | ( n13966 & n13968 ) ;
  assign n13970 = n5966 & n12050 ;
  assign n13971 = n6464 & n9989 ;
  assign n13972 = n5970 & n9993 ;
  assign n13973 = n5969 & n9991 ;
  assign n13974 = n13972 | n13973 ;
  assign n13975 = ( ~n13970 & n13971 ) | ( ~n13970 & n13974 ) | ( n13971 & n13974 ) ;
  assign n13976 = ( ~x14 & n13970 ) | ( ~x14 & n13975 ) | ( n13970 & n13975 ) ;
  assign n13977 = ( n13970 & n13975 ) | ( n13970 & ~n13976 ) | ( n13975 & ~n13976 ) ;
  assign n13978 = ( x14 & n13976 ) | ( x14 & ~n13977 ) | ( n13976 & ~n13977 ) ;
  assign n13979 = ( ~n13593 & n13602 ) | ( ~n13593 & n13605 ) | ( n13602 & n13605 ) ;
  assign n13980 = ( n13593 & ~n13606 ) | ( n13593 & n13979 ) | ( ~n13606 & n13979 ) ;
  assign n13981 = ( n13969 & n13978 ) | ( n13969 & n13980 ) | ( n13978 & n13980 ) ;
  assign n13982 = ( ~n13606 & n13615 ) | ( ~n13606 & n13617 ) | ( n13615 & n13617 ) ;
  assign n13983 = ( n13606 & ~n13618 ) | ( n13606 & n13982 ) | ( ~n13618 & n13982 ) ;
  assign n13984 = n5966 & ~n12074 ;
  assign n13985 = n6464 & ~n9987 ;
  assign n13986 = n5970 & n9991 ;
  assign n13987 = n5969 & n9989 ;
  assign n13988 = n13986 | n13987 ;
  assign n13989 = ( ~n13984 & n13985 ) | ( ~n13984 & n13988 ) | ( n13985 & n13988 ) ;
  assign n13990 = ( ~x14 & n13984 ) | ( ~x14 & n13989 ) | ( n13984 & n13989 ) ;
  assign n13991 = ( n13984 & n13989 ) | ( n13984 & ~n13990 ) | ( n13989 & ~n13990 ) ;
  assign n13992 = ( x14 & n13990 ) | ( x14 & ~n13991 ) | ( n13990 & ~n13991 ) ;
  assign n13993 = ( n13981 & n13983 ) | ( n13981 & n13992 ) | ( n13983 & n13992 ) ;
  assign n13994 = ( ~n13618 & n13627 ) | ( ~n13618 & n13629 ) | ( n13627 & n13629 ) ;
  assign n13995 = ( n13618 & ~n13630 ) | ( n13618 & n13994 ) | ( ~n13630 & n13994 ) ;
  assign n13996 = n5966 & ~n12099 ;
  assign n13997 = n6464 & n9985 ;
  assign n13998 = n5970 & n9989 ;
  assign n13999 = n5969 & ~n9987 ;
  assign n14000 = n13998 | n13999 ;
  assign n14001 = ( ~n13996 & n13997 ) | ( ~n13996 & n14000 ) | ( n13997 & n14000 ) ;
  assign n14002 = ( ~x14 & n13996 ) | ( ~x14 & n14001 ) | ( n13996 & n14001 ) ;
  assign n14003 = ( n13996 & n14001 ) | ( n13996 & ~n14002 ) | ( n14001 & ~n14002 ) ;
  assign n14004 = ( x14 & n14002 ) | ( x14 & ~n14003 ) | ( n14002 & ~n14003 ) ;
  assign n14005 = ( n13993 & n13995 ) | ( n13993 & n14004 ) | ( n13995 & n14004 ) ;
  assign n14006 = ( ~n13630 & n13639 ) | ( ~n13630 & n13641 ) | ( n13639 & n13641 ) ;
  assign n14007 = ( n13630 & ~n13642 ) | ( n13630 & n14006 ) | ( ~n13642 & n14006 ) ;
  assign n14008 = n5966 & ~n12129 ;
  assign n14009 = n6464 & ~n9983 ;
  assign n14010 = n5970 & ~n9987 ;
  assign n14011 = n5969 & n9985 ;
  assign n14012 = n14010 | n14011 ;
  assign n14013 = ( ~n14008 & n14009 ) | ( ~n14008 & n14012 ) | ( n14009 & n14012 ) ;
  assign n14014 = ( ~x14 & n14008 ) | ( ~x14 & n14013 ) | ( n14008 & n14013 ) ;
  assign n14015 = ( n14008 & n14013 ) | ( n14008 & ~n14014 ) | ( n14013 & ~n14014 ) ;
  assign n14016 = ( x14 & n14014 ) | ( x14 & ~n14015 ) | ( n14014 & ~n14015 ) ;
  assign n14017 = ( n14005 & n14007 ) | ( n14005 & n14016 ) | ( n14007 & n14016 ) ;
  assign n14018 = n5966 & ~n11561 ;
  assign n14019 = n6464 & n9981 ;
  assign n14020 = n5970 & n9985 ;
  assign n14021 = n5969 & ~n9983 ;
  assign n14022 = n14020 | n14021 ;
  assign n14023 = ( ~n14018 & n14019 ) | ( ~n14018 & n14022 ) | ( n14019 & n14022 ) ;
  assign n14024 = ( ~x14 & n14018 ) | ( ~x14 & n14023 ) | ( n14018 & n14023 ) ;
  assign n14025 = ( n14018 & n14023 ) | ( n14018 & ~n14024 ) | ( n14023 & ~n14024 ) ;
  assign n14026 = ( x14 & n14024 ) | ( x14 & ~n14025 ) | ( n14024 & ~n14025 ) ;
  assign n14027 = ( ~n13642 & n13644 ) | ( ~n13642 & n13653 ) | ( n13644 & n13653 ) ;
  assign n14028 = ( n13642 & ~n13654 ) | ( n13642 & n14027 ) | ( ~n13654 & n14027 ) ;
  assign n14029 = ( n14017 & n14026 ) | ( n14017 & n14028 ) | ( n14026 & n14028 ) ;
  assign n14030 = n5966 & n12153 ;
  assign n14031 = n6464 & n9979 ;
  assign n14032 = n5970 & ~n9983 ;
  assign n14033 = n5969 & n9981 ;
  assign n14034 = n14032 | n14033 ;
  assign n14035 = ( ~n14030 & n14031 ) | ( ~n14030 & n14034 ) | ( n14031 & n14034 ) ;
  assign n14036 = ( ~x14 & n14030 ) | ( ~x14 & n14035 ) | ( n14030 & n14035 ) ;
  assign n14037 = ( n14030 & n14035 ) | ( n14030 & ~n14036 ) | ( n14035 & ~n14036 ) ;
  assign n14038 = ( x14 & n14036 ) | ( x14 & ~n14037 ) | ( n14036 & ~n14037 ) ;
  assign n14039 = ( ~n13654 & n13656 ) | ( ~n13654 & n13665 ) | ( n13656 & n13665 ) ;
  assign n14040 = ( n13654 & ~n13666 ) | ( n13654 & n14039 ) | ( ~n13666 & n14039 ) ;
  assign n14041 = ( n14029 & n14038 ) | ( n14029 & n14040 ) | ( n14038 & n14040 ) ;
  assign n14042 = n5966 & n12165 ;
  assign n14043 = n6464 & n9977 ;
  assign n14044 = n5970 & n9981 ;
  assign n14045 = n5969 & n9979 ;
  assign n14046 = n14044 | n14045 ;
  assign n14047 = ( ~n14042 & n14043 ) | ( ~n14042 & n14046 ) | ( n14043 & n14046 ) ;
  assign n14048 = ( ~x14 & n14042 ) | ( ~x14 & n14047 ) | ( n14042 & n14047 ) ;
  assign n14049 = ( n14042 & n14047 ) | ( n14042 & ~n14048 ) | ( n14047 & ~n14048 ) ;
  assign n14050 = ( x14 & n14048 ) | ( x14 & ~n14049 ) | ( n14048 & ~n14049 ) ;
  assign n14051 = ( ~n13666 & n13668 ) | ( ~n13666 & n13677 ) | ( n13668 & n13677 ) ;
  assign n14052 = ( n13666 & ~n13678 ) | ( n13666 & n14051 ) | ( ~n13678 & n14051 ) ;
  assign n14053 = ( n14041 & n14050 ) | ( n14041 & n14052 ) | ( n14050 & n14052 ) ;
  assign n14054 = ( ~n13678 & n13687 ) | ( ~n13678 & n13689 ) | ( n13687 & n13689 ) ;
  assign n14055 = ( n13678 & ~n13690 ) | ( n13678 & n14054 ) | ( ~n13690 & n14054 ) ;
  assign n14056 = n5966 & n11606 ;
  assign n14057 = n6464 & n9975 ;
  assign n14058 = n5970 & n9979 ;
  assign n14059 = n5969 & n9977 ;
  assign n14060 = n14058 | n14059 ;
  assign n14061 = ( ~n14056 & n14057 ) | ( ~n14056 & n14060 ) | ( n14057 & n14060 ) ;
  assign n14062 = ( ~x14 & n14056 ) | ( ~x14 & n14061 ) | ( n14056 & n14061 ) ;
  assign n14063 = ( n14056 & n14061 ) | ( n14056 & ~n14062 ) | ( n14061 & ~n14062 ) ;
  assign n14064 = ( x14 & n14062 ) | ( x14 & ~n14063 ) | ( n14062 & ~n14063 ) ;
  assign n14065 = ( n14053 & n14055 ) | ( n14053 & n14064 ) | ( n14055 & n14064 ) ;
  assign n14066 = ( ~n13690 & n13699 ) | ( ~n13690 & n13701 ) | ( n13699 & n13701 ) ;
  assign n14067 = ( n13690 & ~n13702 ) | ( n13690 & n14066 ) | ( ~n13702 & n14066 ) ;
  assign n14068 = n5966 & n11400 ;
  assign n14069 = n6464 & n9973 ;
  assign n14070 = n5970 & n9977 ;
  assign n14071 = n5969 & n9975 ;
  assign n14072 = n14070 | n14071 ;
  assign n14073 = ( ~n14068 & n14069 ) | ( ~n14068 & n14072 ) | ( n14069 & n14072 ) ;
  assign n14074 = ( ~x14 & n14068 ) | ( ~x14 & n14073 ) | ( n14068 & n14073 ) ;
  assign n14075 = ( n14068 & n14073 ) | ( n14068 & ~n14074 ) | ( n14073 & ~n14074 ) ;
  assign n14076 = ( x14 & n14074 ) | ( x14 & ~n14075 ) | ( n14074 & ~n14075 ) ;
  assign n14077 = ( n14065 & n14067 ) | ( n14065 & n14076 ) | ( n14067 & n14076 ) ;
  assign n14078 = ( ~n13702 & n13711 ) | ( ~n13702 & n13713 ) | ( n13711 & n13713 ) ;
  assign n14079 = ( n13702 & ~n13714 ) | ( n13702 & n14078 ) | ( ~n13714 & n14078 ) ;
  assign n14080 = n5966 & n11630 ;
  assign n14081 = n6464 & n9971 ;
  assign n14082 = n5970 & n9975 ;
  assign n14083 = n5969 & n9973 ;
  assign n14084 = n14082 | n14083 ;
  assign n14085 = ( ~n14080 & n14081 ) | ( ~n14080 & n14084 ) | ( n14081 & n14084 ) ;
  assign n14086 = ( ~x14 & n14080 ) | ( ~x14 & n14085 ) | ( n14080 & n14085 ) ;
  assign n14087 = ( n14080 & n14085 ) | ( n14080 & ~n14086 ) | ( n14085 & ~n14086 ) ;
  assign n14088 = ( x14 & n14086 ) | ( x14 & ~n14087 ) | ( n14086 & ~n14087 ) ;
  assign n14089 = ( n14077 & n14079 ) | ( n14077 & n14088 ) | ( n14079 & n14088 ) ;
  assign n14090 = n5966 & n11428 ;
  assign n14091 = n6464 & n9969 ;
  assign n14092 = n5970 & n9973 ;
  assign n14093 = n5969 & n9971 ;
  assign n14094 = n14092 | n14093 ;
  assign n14095 = ( ~n14090 & n14091 ) | ( ~n14090 & n14094 ) | ( n14091 & n14094 ) ;
  assign n14096 = ( ~x14 & n14090 ) | ( ~x14 & n14095 ) | ( n14090 & n14095 ) ;
  assign n14097 = ( n14090 & n14095 ) | ( n14090 & ~n14096 ) | ( n14095 & ~n14096 ) ;
  assign n14098 = ( x14 & n14096 ) | ( x14 & ~n14097 ) | ( n14096 & ~n14097 ) ;
  assign n14099 = ( ~n13714 & n13716 ) | ( ~n13714 & n13725 ) | ( n13716 & n13725 ) ;
  assign n14100 = ( n13714 & ~n13726 ) | ( n13714 & n14099 ) | ( ~n13726 & n14099 ) ;
  assign n14101 = ( n14089 & n14098 ) | ( n14089 & n14100 ) | ( n14098 & n14100 ) ;
  assign n14102 = n5966 & ~n10998 ;
  assign n14103 = n6464 & ~n9967 ;
  assign n14104 = n5970 & n9971 ;
  assign n14105 = n5969 & n9969 ;
  assign n14106 = n14104 | n14105 ;
  assign n14107 = ( ~n14102 & n14103 ) | ( ~n14102 & n14106 ) | ( n14103 & n14106 ) ;
  assign n14108 = ( ~x14 & n14102 ) | ( ~x14 & n14107 ) | ( n14102 & n14107 ) ;
  assign n14109 = ( n14102 & n14107 ) | ( n14102 & ~n14108 ) | ( n14107 & ~n14108 ) ;
  assign n14110 = ( x14 & n14108 ) | ( x14 & ~n14109 ) | ( n14108 & ~n14109 ) ;
  assign n14111 = ( ~n13726 & n13728 ) | ( ~n13726 & n13737 ) | ( n13728 & n13737 ) ;
  assign n14112 = ( n13726 & ~n13738 ) | ( n13726 & n14111 ) | ( ~n13738 & n14111 ) ;
  assign n14113 = ( n14101 & n14110 ) | ( n14101 & n14112 ) | ( n14110 & n14112 ) ;
  assign n14114 = ( n13738 & ~n13747 ) | ( n13738 & n13749 ) | ( ~n13747 & n13749 ) ;
  assign n14115 = ( ~n13738 & n13750 ) | ( ~n13738 & n14114 ) | ( n13750 & n14114 ) ;
  assign n14116 = n5966 & ~n11273 ;
  assign n14117 = n6464 & n9965 ;
  assign n14118 = n5970 & n9969 ;
  assign n14119 = n5969 & ~n9967 ;
  assign n14120 = n14118 | n14119 ;
  assign n14121 = ( ~n14116 & n14117 ) | ( ~n14116 & n14120 ) | ( n14117 & n14120 ) ;
  assign n14122 = ( ~x14 & n14116 ) | ( ~x14 & n14121 ) | ( n14116 & n14121 ) ;
  assign n14123 = ( n14116 & n14121 ) | ( n14116 & ~n14122 ) | ( n14121 & ~n14122 ) ;
  assign n14124 = ( x14 & n14122 ) | ( x14 & ~n14123 ) | ( n14122 & ~n14123 ) ;
  assign n14125 = ( n14113 & ~n14115 ) | ( n14113 & n14124 ) | ( ~n14115 & n14124 ) ;
  assign n14126 = ( n13750 & ~n13759 ) | ( n13750 & n13761 ) | ( ~n13759 & n13761 ) ;
  assign n14127 = ( ~n13750 & n13762 ) | ( ~n13750 & n14126 ) | ( n13762 & n14126 ) ;
  assign n14128 = n5966 & ~n11121 ;
  assign n14129 = n6464 & ~n9963 ;
  assign n14130 = n5970 & ~n9967 ;
  assign n14131 = n5969 & n9965 ;
  assign n14132 = n14130 | n14131 ;
  assign n14133 = ( ~n14128 & n14129 ) | ( ~n14128 & n14132 ) | ( n14129 & n14132 ) ;
  assign n14134 = ( ~x14 & n14128 ) | ( ~x14 & n14133 ) | ( n14128 & n14133 ) ;
  assign n14135 = ( n14128 & n14133 ) | ( n14128 & ~n14134 ) | ( n14133 & ~n14134 ) ;
  assign n14136 = ( x14 & n14134 ) | ( x14 & ~n14135 ) | ( n14134 & ~n14135 ) ;
  assign n14137 = ( n14125 & ~n14127 ) | ( n14125 & n14136 ) | ( ~n14127 & n14136 ) ;
  assign n14138 = ( ~n13762 & n13771 ) | ( ~n13762 & n13773 ) | ( n13771 & n13773 ) ;
  assign n14139 = ( n13762 & ~n13774 ) | ( n13762 & n14138 ) | ( ~n13774 & n14138 ) ;
  assign n14140 = n5966 & ~n10929 ;
  assign n14141 = n6464 & n9961 ;
  assign n14142 = n5970 & n9965 ;
  assign n14143 = n5969 & ~n9963 ;
  assign n14144 = n14142 | n14143 ;
  assign n14145 = ( ~n14140 & n14141 ) | ( ~n14140 & n14144 ) | ( n14141 & n14144 ) ;
  assign n14146 = ( ~x14 & n14140 ) | ( ~x14 & n14145 ) | ( n14140 & n14145 ) ;
  assign n14147 = ( n14140 & n14145 ) | ( n14140 & ~n14146 ) | ( n14145 & ~n14146 ) ;
  assign n14148 = ( x14 & n14146 ) | ( x14 & ~n14147 ) | ( n14146 & ~n14147 ) ;
  assign n14149 = ( n14137 & n14139 ) | ( n14137 & n14148 ) | ( n14139 & n14148 ) ;
  assign n14150 = ( n13774 & ~n13783 ) | ( n13774 & n13785 ) | ( ~n13783 & n13785 ) ;
  assign n14151 = ( ~n13774 & n13786 ) | ( ~n13774 & n14150 ) | ( n13786 & n14150 ) ;
  assign n14152 = n5966 & n10859 ;
  assign n14153 = n6464 & n9959 ;
  assign n14154 = n5970 & ~n9963 ;
  assign n14155 = n5969 & n9961 ;
  assign n14156 = n14154 | n14155 ;
  assign n14157 = ( ~n14152 & n14153 ) | ( ~n14152 & n14156 ) | ( n14153 & n14156 ) ;
  assign n14158 = ( ~x14 & n14152 ) | ( ~x14 & n14157 ) | ( n14152 & n14157 ) ;
  assign n14159 = ( n14152 & n14157 ) | ( n14152 & ~n14158 ) | ( n14157 & ~n14158 ) ;
  assign n14160 = ( x14 & n14158 ) | ( x14 & ~n14159 ) | ( n14158 & ~n14159 ) ;
  assign n14161 = ( n14149 & ~n14151 ) | ( n14149 & n14160 ) | ( ~n14151 & n14160 ) ;
  assign n14162 = ( n13786 & ~n13795 ) | ( n13786 & n13797 ) | ( ~n13795 & n13797 ) ;
  assign n14163 = ( ~n13786 & n13798 ) | ( ~n13786 & n14162 ) | ( n13798 & n14162 ) ;
  assign n14164 = n5966 & ~n10869 ;
  assign n14165 = n6464 & ~n9957 ;
  assign n14166 = n5970 & n9961 ;
  assign n14167 = n5969 & n9959 ;
  assign n14168 = n14166 | n14167 ;
  assign n14169 = ( ~n14164 & n14165 ) | ( ~n14164 & n14168 ) | ( n14165 & n14168 ) ;
  assign n14170 = ( ~x14 & n14164 ) | ( ~x14 & n14169 ) | ( n14164 & n14169 ) ;
  assign n14171 = ( n14164 & n14169 ) | ( n14164 & ~n14170 ) | ( n14169 & ~n14170 ) ;
  assign n14172 = ( x14 & n14170 ) | ( x14 & ~n14171 ) | ( n14170 & ~n14171 ) ;
  assign n14173 = ( n14161 & ~n14163 ) | ( n14161 & n14172 ) | ( ~n14163 & n14172 ) ;
  assign n14174 = ( ~n13798 & n13807 ) | ( ~n13798 & n13809 ) | ( n13807 & n13809 ) ;
  assign n14175 = ( n13798 & ~n13810 ) | ( n13798 & n14174 ) | ( ~n13810 & n14174 ) ;
  assign n14176 = n5966 & ~n10567 ;
  assign n14177 = n6464 & n9955 ;
  assign n14178 = n5970 & n9959 ;
  assign n14179 = n5969 & ~n9957 ;
  assign n14180 = n14178 | n14179 ;
  assign n14181 = ( ~n14176 & n14177 ) | ( ~n14176 & n14180 ) | ( n14177 & n14180 ) ;
  assign n14182 = ( ~x14 & n14176 ) | ( ~x14 & n14181 ) | ( n14176 & n14181 ) ;
  assign n14183 = ( n14176 & n14181 ) | ( n14176 & ~n14182 ) | ( n14181 & ~n14182 ) ;
  assign n14184 = ( x14 & n14182 ) | ( x14 & ~n14183 ) | ( n14182 & ~n14183 ) ;
  assign n14185 = ( n14173 & n14175 ) | ( n14173 & n14184 ) | ( n14175 & n14184 ) ;
  assign n14186 = ( ~n13810 & n13819 ) | ( ~n13810 & n13821 ) | ( n13819 & n13821 ) ;
  assign n14187 = ( n13810 & ~n13822 ) | ( n13810 & n14186 ) | ( ~n13822 & n14186 ) ;
  assign n14188 = n5966 & ~n10750 ;
  assign n14189 = n6464 & ~n9953 ;
  assign n14190 = n5970 & ~n9957 ;
  assign n14191 = n5969 & n9955 ;
  assign n14192 = n14190 | n14191 ;
  assign n14193 = ( ~n14188 & n14189 ) | ( ~n14188 & n14192 ) | ( n14189 & n14192 ) ;
  assign n14194 = ( ~x14 & n14188 ) | ( ~x14 & n14193 ) | ( n14188 & n14193 ) ;
  assign n14195 = ( n14188 & n14193 ) | ( n14188 & ~n14194 ) | ( n14193 & ~n14194 ) ;
  assign n14196 = ( x14 & n14194 ) | ( x14 & ~n14195 ) | ( n14194 & ~n14195 ) ;
  assign n14197 = ( n14185 & n14187 ) | ( n14185 & n14196 ) | ( n14187 & n14196 ) ;
  assign n14198 = ( ~n13822 & n13831 ) | ( ~n13822 & n13833 ) | ( n13831 & n13833 ) ;
  assign n14199 = ( n13822 & ~n13834 ) | ( n13822 & n14198 ) | ( ~n13834 & n14198 ) ;
  assign n14200 = n5966 & ~n10652 ;
  assign n14201 = n6464 & n9951 ;
  assign n14202 = n5970 & n9955 ;
  assign n14203 = n5969 & ~n9953 ;
  assign n14204 = n14202 | n14203 ;
  assign n14205 = ( ~n14200 & n14201 ) | ( ~n14200 & n14204 ) | ( n14201 & n14204 ) ;
  assign n14206 = ( ~x14 & n14200 ) | ( ~x14 & n14205 ) | ( n14200 & n14205 ) ;
  assign n14207 = ( n14200 & n14205 ) | ( n14200 & ~n14206 ) | ( n14205 & ~n14206 ) ;
  assign n14208 = ( x14 & n14206 ) | ( x14 & ~n14207 ) | ( n14206 & ~n14207 ) ;
  assign n14209 = ( n14197 & n14199 ) | ( n14197 & n14208 ) | ( n14199 & n14208 ) ;
  assign n14210 = ( ~n13834 & n13843 ) | ( ~n13834 & n13845 ) | ( n13843 & n13845 ) ;
  assign n14211 = ( n13834 & ~n13846 ) | ( n13834 & n14210 ) | ( ~n13846 & n14210 ) ;
  assign n14212 = n5966 & n10557 ;
  assign n14213 = n6464 & n9949 ;
  assign n14214 = n5970 & ~n9953 ;
  assign n14215 = n5969 & n9951 ;
  assign n14216 = n14214 | n14215 ;
  assign n14217 = ( ~n14212 & n14213 ) | ( ~n14212 & n14216 ) | ( n14213 & n14216 ) ;
  assign n14218 = ( ~x14 & n14212 ) | ( ~x14 & n14217 ) | ( n14212 & n14217 ) ;
  assign n14219 = ( n14212 & n14217 ) | ( n14212 & ~n14218 ) | ( n14217 & ~n14218 ) ;
  assign n14220 = ( x14 & n14218 ) | ( x14 & ~n14219 ) | ( n14218 & ~n14219 ) ;
  assign n14221 = ( n14209 & n14211 ) | ( n14209 & n14220 ) | ( n14211 & n14220 ) ;
  assign n14222 = ( ~n13846 & n13855 ) | ( ~n13846 & n13857 ) | ( n13855 & n13857 ) ;
  assign n14223 = ( n13846 & ~n13858 ) | ( n13846 & n14222 ) | ( ~n13858 & n14222 ) ;
  assign n14224 = n5966 & n10454 ;
  assign n14225 = n6464 & n9947 ;
  assign n14226 = n5970 & n9951 ;
  assign n14227 = n5969 & n9949 ;
  assign n14228 = n14226 | n14227 ;
  assign n14229 = ( ~n14224 & n14225 ) | ( ~n14224 & n14228 ) | ( n14225 & n14228 ) ;
  assign n14230 = ( ~x14 & n14224 ) | ( ~x14 & n14229 ) | ( n14224 & n14229 ) ;
  assign n14231 = ( n14224 & n14229 ) | ( n14224 & ~n14230 ) | ( n14229 & ~n14230 ) ;
  assign n14232 = ( x14 & n14230 ) | ( x14 & ~n14231 ) | ( n14230 & ~n14231 ) ;
  assign n14233 = ( n14221 & n14223 ) | ( n14221 & n14232 ) | ( n14223 & n14232 ) ;
  assign n14234 = ( ~n13858 & n13860 ) | ( ~n13858 & n13869 ) | ( n13860 & n13869 ) ;
  assign n14235 = ( ~n13869 & n13870 ) | ( ~n13869 & n14234 ) | ( n13870 & n14234 ) ;
  assign n14236 = n6584 & n10284 ;
  assign n14237 = n7022 & ~n9883 ;
  assign n14238 = n6588 & n9943 ;
  assign n14239 = n6587 & ~n9941 ;
  assign n14240 = n14238 | n14239 ;
  assign n14241 = ( ~n14236 & n14237 ) | ( ~n14236 & n14240 ) | ( n14237 & n14240 ) ;
  assign n14242 = ( ~x11 & n14236 ) | ( ~x11 & n14241 ) | ( n14236 & n14241 ) ;
  assign n14243 = ( n14236 & n14241 ) | ( n14236 & ~n14242 ) | ( n14241 & ~n14242 ) ;
  assign n14244 = ( x11 & n14242 ) | ( x11 & ~n14243 ) | ( n14242 & ~n14243 ) ;
  assign n14245 = ( n14233 & ~n14235 ) | ( n14233 & n14244 ) | ( ~n14235 & n14244 ) ;
  assign n14246 = ( n13870 & ~n13872 ) | ( n13870 & n13881 ) | ( ~n13872 & n13881 ) ;
  assign n14247 = ( n13872 & ~n13882 ) | ( n13872 & n14246 ) | ( ~n13882 & n14246 ) ;
  assign n14248 = n7296 & ~n10305 ;
  assign n14249 = n7879 & ~n10302 ;
  assign n14250 = n7300 & ~n9937 ;
  assign n14251 = n7299 & ~n10057 ;
  assign n14252 = n14250 | n14251 ;
  assign n14253 = ( ~n14248 & n14249 ) | ( ~n14248 & n14252 ) | ( n14249 & n14252 ) ;
  assign n14254 = ( ~x8 & n14248 ) | ( ~x8 & n14253 ) | ( n14248 & n14253 ) ;
  assign n14255 = ( n14248 & n14253 ) | ( n14248 & ~n14254 ) | ( n14253 & ~n14254 ) ;
  assign n14256 = ( x8 & n14254 ) | ( x8 & ~n14255 ) | ( n14254 & ~n14255 ) ;
  assign n14257 = ( n14245 & n14247 ) | ( n14245 & n14256 ) | ( n14247 & n14256 ) ;
  assign n14258 = ( ~n13882 & n13884 ) | ( ~n13882 & n13893 ) | ( n13884 & n13893 ) ;
  assign n14259 = ( ~n13893 & n13894 ) | ( ~n13893 & n14258 ) | ( n13894 & n14258 ) ;
  assign n14260 = ( n11392 & n14257 ) | ( n11392 & ~n14259 ) | ( n14257 & ~n14259 ) ;
  assign n14261 = n6584 & n11892 ;
  assign n14262 = n7022 & ~n9997 ;
  assign n14263 = n6588 & ~n10001 ;
  assign n14264 = n6587 & n9999 ;
  assign n14265 = n14263 | n14264 ;
  assign n14266 = ( ~n14261 & n14262 ) | ( ~n14261 & n14265 ) | ( n14262 & n14265 ) ;
  assign n14267 = ( ~x11 & n14261 ) | ( ~x11 & n14266 ) | ( n14261 & n14266 ) ;
  assign n14268 = ( n14261 & n14266 ) | ( n14261 & ~n14267 ) | ( n14266 & ~n14267 ) ;
  assign n14269 = ( x11 & n14267 ) | ( x11 & ~n14268 ) | ( n14267 & ~n14268 ) ;
  assign n14270 = n6588 & ~n10003 ;
  assign n14271 = n6587 & ~n10001 ;
  assign n14272 = n14270 | n14271 ;
  assign n14273 = n7022 & ~n9999 ;
  assign n14274 = ( n7022 & n14272 ) | ( n7022 & ~n14273 ) | ( n14272 & ~n14273 ) ;
  assign n14275 = n6584 & n11868 ;
  assign n14276 = n14274 | n14275 ;
  assign n14277 = n7021 & ~n10003 ;
  assign n14278 = x11 & n14277 ;
  assign n14279 = ( n6584 & n11804 ) | ( n6584 & n11805 ) | ( n11804 & n11805 ) ;
  assign n14280 = n6587 | n10003 ;
  assign n14281 = n7022 & ~n10001 ;
  assign n14282 = ( ~n10003 & n14280 ) | ( ~n10003 & n14281 ) | ( n14280 & n14281 ) ;
  assign n14283 = n14279 | n14282 ;
  assign n14284 = ( x11 & n14278 ) | ( x11 & n14283 ) | ( n14278 & n14283 ) ;
  assign n14285 = n14276 | n14284 ;
  assign n14286 = x11 & ~n14285 ;
  assign n14287 = ( n13922 & n14269 ) | ( n13922 & n14286 ) | ( n14269 & n14286 ) ;
  assign n14288 = n6584 & n11934 ;
  assign n14289 = n7022 & n9995 ;
  assign n14290 = n6588 & n9999 ;
  assign n14291 = n6587 & ~n9997 ;
  assign n14292 = n14290 | n14291 ;
  assign n14293 = ( ~n14288 & n14289 ) | ( ~n14288 & n14292 ) | ( n14289 & n14292 ) ;
  assign n14294 = ( ~x11 & n14288 ) | ( ~x11 & n14293 ) | ( n14288 & n14293 ) ;
  assign n14295 = ( n14288 & n14293 ) | ( n14288 & ~n14294 ) | ( n14293 & ~n14294 ) ;
  assign n14296 = ( x11 & n14294 ) | ( x11 & ~n14295 ) | ( n14294 & ~n14295 ) ;
  assign n14297 = ( n13923 & n13924 ) | ( n13923 & n13927 ) | ( n13924 & n13927 ) ;
  assign n14298 = ~n13923 & n13928 ;
  assign n14299 = ( n13923 & ~n14297 ) | ( n13923 & n14298 ) | ( ~n14297 & n14298 ) ;
  assign n14300 = ( n14287 & n14296 ) | ( n14287 & n14299 ) | ( n14296 & n14299 ) ;
  assign n14301 = n6584 & ~n11971 ;
  assign n14302 = n7022 & n9993 ;
  assign n14303 = n6588 & ~n9997 ;
  assign n14304 = n6587 & n9995 ;
  assign n14305 = n14303 | n14304 ;
  assign n14306 = ( ~n14301 & n14302 ) | ( ~n14301 & n14305 ) | ( n14302 & n14305 ) ;
  assign n14307 = ( ~x11 & n14301 ) | ( ~x11 & n14306 ) | ( n14301 & n14306 ) ;
  assign n14308 = ( n14301 & n14306 ) | ( n14301 & ~n14307 ) | ( n14306 & ~n14307 ) ;
  assign n14309 = ( x11 & n14307 ) | ( x11 & ~n14308 ) | ( n14307 & ~n14308 ) ;
  assign n14310 = ( n13921 & n13929 ) | ( n13921 & ~n13930 ) | ( n13929 & ~n13930 ) ;
  assign n14311 = n13930 & ~n14310 ;
  assign n14312 = ( n14300 & n14309 ) | ( n14300 & n14311 ) | ( n14309 & n14311 ) ;
  assign n14313 = n6584 & n12026 ;
  assign n14314 = n7022 & n9991 ;
  assign n14315 = n6588 & n9995 ;
  assign n14316 = n6587 & n9993 ;
  assign n14317 = n14315 | n14316 ;
  assign n14318 = ( ~n14313 & n14314 ) | ( ~n14313 & n14317 ) | ( n14314 & n14317 ) ;
  assign n14319 = ( ~x11 & n14313 ) | ( ~x11 & n14318 ) | ( n14313 & n14318 ) ;
  assign n14320 = ( n14313 & n14318 ) | ( n14313 & ~n14319 ) | ( n14318 & ~n14319 ) ;
  assign n14321 = ( x11 & n14319 ) | ( x11 & ~n14320 ) | ( n14319 & ~n14320 ) ;
  assign n14322 = ( n13583 & n13914 ) | ( n13583 & ~n13931 ) | ( n13914 & ~n13931 ) ;
  assign n14323 = ( n13931 & ~n13932 ) | ( n13931 & n14322 ) | ( ~n13932 & n14322 ) ;
  assign n14324 = ( n14312 & n14321 ) | ( n14312 & n14323 ) | ( n14321 & n14323 ) ;
  assign n14325 = n6584 & n12050 ;
  assign n14326 = n7022 & n9989 ;
  assign n14327 = n6588 & n9993 ;
  assign n14328 = n6587 & n9991 ;
  assign n14329 = n14327 | n14328 ;
  assign n14330 = ( ~n14325 & n14326 ) | ( ~n14325 & n14329 ) | ( n14326 & n14329 ) ;
  assign n14331 = ( ~x11 & n14325 ) | ( ~x11 & n14330 ) | ( n14325 & n14330 ) ;
  assign n14332 = ( n14325 & n14330 ) | ( n14325 & ~n14331 ) | ( n14330 & ~n14331 ) ;
  assign n14333 = ( x11 & n14331 ) | ( x11 & ~n14332 ) | ( n14331 & ~n14332 ) ;
  assign n14334 = ( ~n13932 & n13941 ) | ( ~n13932 & n13944 ) | ( n13941 & n13944 ) ;
  assign n14335 = ( n13932 & ~n13945 ) | ( n13932 & n14334 ) | ( ~n13945 & n14334 ) ;
  assign n14336 = ( n14324 & n14333 ) | ( n14324 & n14335 ) | ( n14333 & n14335 ) ;
  assign n14337 = ( ~n13945 & n13954 ) | ( ~n13945 & n13956 ) | ( n13954 & n13956 ) ;
  assign n14338 = ( n13945 & ~n13957 ) | ( n13945 & n14337 ) | ( ~n13957 & n14337 ) ;
  assign n14339 = n6584 & ~n12074 ;
  assign n14340 = n7022 & ~n9987 ;
  assign n14341 = n6588 & n9991 ;
  assign n14342 = n6587 & n9989 ;
  assign n14343 = n14341 | n14342 ;
  assign n14344 = ( ~n14339 & n14340 ) | ( ~n14339 & n14343 ) | ( n14340 & n14343 ) ;
  assign n14345 = ( ~x11 & n14339 ) | ( ~x11 & n14344 ) | ( n14339 & n14344 ) ;
  assign n14346 = ( n14339 & n14344 ) | ( n14339 & ~n14345 ) | ( n14344 & ~n14345 ) ;
  assign n14347 = ( x11 & n14345 ) | ( x11 & ~n14346 ) | ( n14345 & ~n14346 ) ;
  assign n14348 = ( n14336 & n14338 ) | ( n14336 & n14347 ) | ( n14338 & n14347 ) ;
  assign n14349 = ( ~n13957 & n13966 ) | ( ~n13957 & n13968 ) | ( n13966 & n13968 ) ;
  assign n14350 = ( n13957 & ~n13969 ) | ( n13957 & n14349 ) | ( ~n13969 & n14349 ) ;
  assign n14351 = n6584 & ~n12099 ;
  assign n14352 = n7022 & n9985 ;
  assign n14353 = n6588 & n9989 ;
  assign n14354 = n6587 & ~n9987 ;
  assign n14355 = n14353 | n14354 ;
  assign n14356 = ( ~n14351 & n14352 ) | ( ~n14351 & n14355 ) | ( n14352 & n14355 ) ;
  assign n14357 = ( ~x11 & n14351 ) | ( ~x11 & n14356 ) | ( n14351 & n14356 ) ;
  assign n14358 = ( n14351 & n14356 ) | ( n14351 & ~n14357 ) | ( n14356 & ~n14357 ) ;
  assign n14359 = ( x11 & n14357 ) | ( x11 & ~n14358 ) | ( n14357 & ~n14358 ) ;
  assign n14360 = ( n14348 & n14350 ) | ( n14348 & n14359 ) | ( n14350 & n14359 ) ;
  assign n14361 = ( ~n13969 & n13978 ) | ( ~n13969 & n13980 ) | ( n13978 & n13980 ) ;
  assign n14362 = ( n13969 & ~n13981 ) | ( n13969 & n14361 ) | ( ~n13981 & n14361 ) ;
  assign n14363 = n6584 & ~n12129 ;
  assign n14364 = n7022 & ~n9983 ;
  assign n14365 = n6588 & ~n9987 ;
  assign n14366 = n6587 & n9985 ;
  assign n14367 = n14365 | n14366 ;
  assign n14368 = ( ~n14363 & n14364 ) | ( ~n14363 & n14367 ) | ( n14364 & n14367 ) ;
  assign n14369 = ( ~x11 & n14363 ) | ( ~x11 & n14368 ) | ( n14363 & n14368 ) ;
  assign n14370 = ( n14363 & n14368 ) | ( n14363 & ~n14369 ) | ( n14368 & ~n14369 ) ;
  assign n14371 = ( x11 & n14369 ) | ( x11 & ~n14370 ) | ( n14369 & ~n14370 ) ;
  assign n14372 = ( n14360 & n14362 ) | ( n14360 & n14371 ) | ( n14362 & n14371 ) ;
  assign n14373 = n6584 & ~n11561 ;
  assign n14374 = n7022 & n9981 ;
  assign n14375 = n6588 & n9985 ;
  assign n14376 = n6587 & ~n9983 ;
  assign n14377 = n14375 | n14376 ;
  assign n14378 = ( ~n14373 & n14374 ) | ( ~n14373 & n14377 ) | ( n14374 & n14377 ) ;
  assign n14379 = ( ~x11 & n14373 ) | ( ~x11 & n14378 ) | ( n14373 & n14378 ) ;
  assign n14380 = ( n14373 & n14378 ) | ( n14373 & ~n14379 ) | ( n14378 & ~n14379 ) ;
  assign n14381 = ( x11 & n14379 ) | ( x11 & ~n14380 ) | ( n14379 & ~n14380 ) ;
  assign n14382 = ( ~n13981 & n13983 ) | ( ~n13981 & n13992 ) | ( n13983 & n13992 ) ;
  assign n14383 = ( n13981 & ~n13993 ) | ( n13981 & n14382 ) | ( ~n13993 & n14382 ) ;
  assign n14384 = ( n14372 & n14381 ) | ( n14372 & n14383 ) | ( n14381 & n14383 ) ;
  assign n14385 = n6584 & n12153 ;
  assign n14386 = n7022 & n9979 ;
  assign n14387 = n6588 & ~n9983 ;
  assign n14388 = n6587 & n9981 ;
  assign n14389 = n14387 | n14388 ;
  assign n14390 = ( ~n14385 & n14386 ) | ( ~n14385 & n14389 ) | ( n14386 & n14389 ) ;
  assign n14391 = ( ~x11 & n14385 ) | ( ~x11 & n14390 ) | ( n14385 & n14390 ) ;
  assign n14392 = ( n14385 & n14390 ) | ( n14385 & ~n14391 ) | ( n14390 & ~n14391 ) ;
  assign n14393 = ( x11 & n14391 ) | ( x11 & ~n14392 ) | ( n14391 & ~n14392 ) ;
  assign n14394 = ( ~n13993 & n13995 ) | ( ~n13993 & n14004 ) | ( n13995 & n14004 ) ;
  assign n14395 = ( n13993 & ~n14005 ) | ( n13993 & n14394 ) | ( ~n14005 & n14394 ) ;
  assign n14396 = ( n14384 & n14393 ) | ( n14384 & n14395 ) | ( n14393 & n14395 ) ;
  assign n14397 = n6584 & n12165 ;
  assign n14398 = n7022 & n9977 ;
  assign n14399 = n6588 & n9981 ;
  assign n14400 = n6587 & n9979 ;
  assign n14401 = n14399 | n14400 ;
  assign n14402 = ( ~n14397 & n14398 ) | ( ~n14397 & n14401 ) | ( n14398 & n14401 ) ;
  assign n14403 = ( ~x11 & n14397 ) | ( ~x11 & n14402 ) | ( n14397 & n14402 ) ;
  assign n14404 = ( n14397 & n14402 ) | ( n14397 & ~n14403 ) | ( n14402 & ~n14403 ) ;
  assign n14405 = ( x11 & n14403 ) | ( x11 & ~n14404 ) | ( n14403 & ~n14404 ) ;
  assign n14406 = ( ~n14005 & n14007 ) | ( ~n14005 & n14016 ) | ( n14007 & n14016 ) ;
  assign n14407 = ( n14005 & ~n14017 ) | ( n14005 & n14406 ) | ( ~n14017 & n14406 ) ;
  assign n14408 = ( n14396 & n14405 ) | ( n14396 & n14407 ) | ( n14405 & n14407 ) ;
  assign n14409 = ( ~n14017 & n14026 ) | ( ~n14017 & n14028 ) | ( n14026 & n14028 ) ;
  assign n14410 = ( n14017 & ~n14029 ) | ( n14017 & n14409 ) | ( ~n14029 & n14409 ) ;
  assign n14411 = n6584 & n11606 ;
  assign n14412 = n7022 & n9975 ;
  assign n14413 = n6588 & n9979 ;
  assign n14414 = n6587 & n9977 ;
  assign n14415 = n14413 | n14414 ;
  assign n14416 = ( ~n14411 & n14412 ) | ( ~n14411 & n14415 ) | ( n14412 & n14415 ) ;
  assign n14417 = ( ~x11 & n14411 ) | ( ~x11 & n14416 ) | ( n14411 & n14416 ) ;
  assign n14418 = ( n14411 & n14416 ) | ( n14411 & ~n14417 ) | ( n14416 & ~n14417 ) ;
  assign n14419 = ( x11 & n14417 ) | ( x11 & ~n14418 ) | ( n14417 & ~n14418 ) ;
  assign n14420 = ( n14408 & n14410 ) | ( n14408 & n14419 ) | ( n14410 & n14419 ) ;
  assign n14421 = ( ~n14029 & n14038 ) | ( ~n14029 & n14040 ) | ( n14038 & n14040 ) ;
  assign n14422 = ( n14029 & ~n14041 ) | ( n14029 & n14421 ) | ( ~n14041 & n14421 ) ;
  assign n14423 = n6584 & n11400 ;
  assign n14424 = n7022 & n9973 ;
  assign n14425 = n6588 & n9977 ;
  assign n14426 = n6587 & n9975 ;
  assign n14427 = n14425 | n14426 ;
  assign n14428 = ( ~n14423 & n14424 ) | ( ~n14423 & n14427 ) | ( n14424 & n14427 ) ;
  assign n14429 = ( ~x11 & n14423 ) | ( ~x11 & n14428 ) | ( n14423 & n14428 ) ;
  assign n14430 = ( n14423 & n14428 ) | ( n14423 & ~n14429 ) | ( n14428 & ~n14429 ) ;
  assign n14431 = ( x11 & n14429 ) | ( x11 & ~n14430 ) | ( n14429 & ~n14430 ) ;
  assign n14432 = ( n14420 & n14422 ) | ( n14420 & n14431 ) | ( n14422 & n14431 ) ;
  assign n14433 = ( ~n14041 & n14050 ) | ( ~n14041 & n14052 ) | ( n14050 & n14052 ) ;
  assign n14434 = ( n14041 & ~n14053 ) | ( n14041 & n14433 ) | ( ~n14053 & n14433 ) ;
  assign n14435 = n6584 & n11630 ;
  assign n14436 = n7022 & n9971 ;
  assign n14437 = n6588 & n9975 ;
  assign n14438 = n6587 & n9973 ;
  assign n14439 = n14437 | n14438 ;
  assign n14440 = ( ~n14435 & n14436 ) | ( ~n14435 & n14439 ) | ( n14436 & n14439 ) ;
  assign n14441 = ( ~x11 & n14435 ) | ( ~x11 & n14440 ) | ( n14435 & n14440 ) ;
  assign n14442 = ( n14435 & n14440 ) | ( n14435 & ~n14441 ) | ( n14440 & ~n14441 ) ;
  assign n14443 = ( x11 & n14441 ) | ( x11 & ~n14442 ) | ( n14441 & ~n14442 ) ;
  assign n14444 = ( n14432 & n14434 ) | ( n14432 & n14443 ) | ( n14434 & n14443 ) ;
  assign n14445 = n6584 & n11428 ;
  assign n14446 = n7022 & n9969 ;
  assign n14447 = n6588 & n9973 ;
  assign n14448 = n6587 & n9971 ;
  assign n14449 = n14447 | n14448 ;
  assign n14450 = ( ~n14445 & n14446 ) | ( ~n14445 & n14449 ) | ( n14446 & n14449 ) ;
  assign n14451 = ( ~x11 & n14445 ) | ( ~x11 & n14450 ) | ( n14445 & n14450 ) ;
  assign n14452 = ( n14445 & n14450 ) | ( n14445 & ~n14451 ) | ( n14450 & ~n14451 ) ;
  assign n14453 = ( x11 & n14451 ) | ( x11 & ~n14452 ) | ( n14451 & ~n14452 ) ;
  assign n14454 = ( ~n14053 & n14055 ) | ( ~n14053 & n14064 ) | ( n14055 & n14064 ) ;
  assign n14455 = ( n14053 & ~n14065 ) | ( n14053 & n14454 ) | ( ~n14065 & n14454 ) ;
  assign n14456 = ( n14444 & n14453 ) | ( n14444 & n14455 ) | ( n14453 & n14455 ) ;
  assign n14457 = n6584 & ~n10998 ;
  assign n14458 = n7022 & ~n9967 ;
  assign n14459 = n6588 & n9971 ;
  assign n14460 = n6587 & n9969 ;
  assign n14461 = n14459 | n14460 ;
  assign n14462 = ( ~n14457 & n14458 ) | ( ~n14457 & n14461 ) | ( n14458 & n14461 ) ;
  assign n14463 = ( ~x11 & n14457 ) | ( ~x11 & n14462 ) | ( n14457 & n14462 ) ;
  assign n14464 = ( n14457 & n14462 ) | ( n14457 & ~n14463 ) | ( n14462 & ~n14463 ) ;
  assign n14465 = ( x11 & n14463 ) | ( x11 & ~n14464 ) | ( n14463 & ~n14464 ) ;
  assign n14466 = ( ~n14065 & n14067 ) | ( ~n14065 & n14076 ) | ( n14067 & n14076 ) ;
  assign n14467 = ( n14065 & ~n14077 ) | ( n14065 & n14466 ) | ( ~n14077 & n14466 ) ;
  assign n14468 = ( n14456 & n14465 ) | ( n14456 & n14467 ) | ( n14465 & n14467 ) ;
  assign n14469 = n6584 & ~n11273 ;
  assign n14470 = n7022 & n9965 ;
  assign n14471 = n6588 & n9969 ;
  assign n14472 = n6587 & ~n9967 ;
  assign n14473 = n14471 | n14472 ;
  assign n14474 = ( ~n14469 & n14470 ) | ( ~n14469 & n14473 ) | ( n14470 & n14473 ) ;
  assign n14475 = ( ~x11 & n14469 ) | ( ~x11 & n14474 ) | ( n14469 & n14474 ) ;
  assign n14476 = ( n14469 & n14474 ) | ( n14469 & ~n14475 ) | ( n14474 & ~n14475 ) ;
  assign n14477 = ( x11 & n14475 ) | ( x11 & ~n14476 ) | ( n14475 & ~n14476 ) ;
  assign n14478 = ( ~n14077 & n14079 ) | ( ~n14077 & n14088 ) | ( n14079 & n14088 ) ;
  assign n14479 = ( n14077 & ~n14089 ) | ( n14077 & n14478 ) | ( ~n14089 & n14478 ) ;
  assign n14480 = ( n14468 & n14477 ) | ( n14468 & n14479 ) | ( n14477 & n14479 ) ;
  assign n14481 = ( ~n14089 & n14098 ) | ( ~n14089 & n14100 ) | ( n14098 & n14100 ) ;
  assign n14482 = ( n14089 & ~n14101 ) | ( n14089 & n14481 ) | ( ~n14101 & n14481 ) ;
  assign n14483 = n6584 & ~n11121 ;
  assign n14484 = n7022 & ~n9963 ;
  assign n14485 = n6588 & ~n9967 ;
  assign n14486 = n6587 & n9965 ;
  assign n14487 = n14485 | n14486 ;
  assign n14488 = ( ~n14483 & n14484 ) | ( ~n14483 & n14487 ) | ( n14484 & n14487 ) ;
  assign n14489 = ( ~x11 & n14483 ) | ( ~x11 & n14488 ) | ( n14483 & n14488 ) ;
  assign n14490 = ( n14483 & n14488 ) | ( n14483 & ~n14489 ) | ( n14488 & ~n14489 ) ;
  assign n14491 = ( x11 & n14489 ) | ( x11 & ~n14490 ) | ( n14489 & ~n14490 ) ;
  assign n14492 = ( n14480 & n14482 ) | ( n14480 & n14491 ) | ( n14482 & n14491 ) ;
  assign n14493 = ( ~n14101 & n14110 ) | ( ~n14101 & n14112 ) | ( n14110 & n14112 ) ;
  assign n14494 = ( n14101 & ~n14113 ) | ( n14101 & n14493 ) | ( ~n14113 & n14493 ) ;
  assign n14495 = n6584 & ~n10929 ;
  assign n14496 = n7022 & n9961 ;
  assign n14497 = n6588 & n9965 ;
  assign n14498 = n6587 & ~n9963 ;
  assign n14499 = n14497 | n14498 ;
  assign n14500 = ( ~n14495 & n14496 ) | ( ~n14495 & n14499 ) | ( n14496 & n14499 ) ;
  assign n14501 = ( ~x11 & n14495 ) | ( ~x11 & n14500 ) | ( n14495 & n14500 ) ;
  assign n14502 = ( n14495 & n14500 ) | ( n14495 & ~n14501 ) | ( n14500 & ~n14501 ) ;
  assign n14503 = ( x11 & n14501 ) | ( x11 & ~n14502 ) | ( n14501 & ~n14502 ) ;
  assign n14504 = ( n14492 & n14494 ) | ( n14492 & n14503 ) | ( n14494 & n14503 ) ;
  assign n14505 = n6584 & n10859 ;
  assign n14506 = n7022 & n9959 ;
  assign n14507 = n6588 & ~n9963 ;
  assign n14508 = n6587 & n9961 ;
  assign n14509 = n14507 | n14508 ;
  assign n14510 = ( ~n14505 & n14506 ) | ( ~n14505 & n14509 ) | ( n14506 & n14509 ) ;
  assign n14511 = ( ~x11 & n14505 ) | ( ~x11 & n14510 ) | ( n14505 & n14510 ) ;
  assign n14512 = ( n14505 & n14510 ) | ( n14505 & ~n14511 ) | ( n14510 & ~n14511 ) ;
  assign n14513 = ( x11 & n14511 ) | ( x11 & ~n14512 ) | ( n14511 & ~n14512 ) ;
  assign n14514 = ( ~n14113 & n14115 ) | ( ~n14113 & n14124 ) | ( n14115 & n14124 ) ;
  assign n14515 = ( ~n14124 & n14125 ) | ( ~n14124 & n14514 ) | ( n14125 & n14514 ) ;
  assign n14516 = ( n14504 & n14513 ) | ( n14504 & ~n14515 ) | ( n14513 & ~n14515 ) ;
  assign n14517 = n6584 & ~n10869 ;
  assign n14518 = n7022 & ~n9957 ;
  assign n14519 = n6588 & n9961 ;
  assign n14520 = n6587 & n9959 ;
  assign n14521 = n14519 | n14520 ;
  assign n14522 = ( ~n14517 & n14518 ) | ( ~n14517 & n14521 ) | ( n14518 & n14521 ) ;
  assign n14523 = ( ~x11 & n14517 ) | ( ~x11 & n14522 ) | ( n14517 & n14522 ) ;
  assign n14524 = ( n14517 & n14522 ) | ( n14517 & ~n14523 ) | ( n14522 & ~n14523 ) ;
  assign n14525 = ( x11 & n14523 ) | ( x11 & ~n14524 ) | ( n14523 & ~n14524 ) ;
  assign n14526 = ( ~n14125 & n14127 ) | ( ~n14125 & n14136 ) | ( n14127 & n14136 ) ;
  assign n14527 = ( ~n14136 & n14137 ) | ( ~n14136 & n14526 ) | ( n14137 & n14526 ) ;
  assign n14528 = ( n14516 & n14525 ) | ( n14516 & ~n14527 ) | ( n14525 & ~n14527 ) ;
  assign n14529 = n6584 & ~n10567 ;
  assign n14530 = n7022 & n9955 ;
  assign n14531 = n6588 & n9959 ;
  assign n14532 = n6587 & ~n9957 ;
  assign n14533 = n14531 | n14532 ;
  assign n14534 = ( ~n14529 & n14530 ) | ( ~n14529 & n14533 ) | ( n14530 & n14533 ) ;
  assign n14535 = ( ~x11 & n14529 ) | ( ~x11 & n14534 ) | ( n14529 & n14534 ) ;
  assign n14536 = ( n14529 & n14534 ) | ( n14529 & ~n14535 ) | ( n14534 & ~n14535 ) ;
  assign n14537 = ( x11 & n14535 ) | ( x11 & ~n14536 ) | ( n14535 & ~n14536 ) ;
  assign n14538 = ( ~n14137 & n14139 ) | ( ~n14137 & n14148 ) | ( n14139 & n14148 ) ;
  assign n14539 = ( n14137 & ~n14149 ) | ( n14137 & n14538 ) | ( ~n14149 & n14538 ) ;
  assign n14540 = ( n14528 & n14537 ) | ( n14528 & n14539 ) | ( n14537 & n14539 ) ;
  assign n14541 = n6584 & ~n10750 ;
  assign n14542 = n7022 & ~n9953 ;
  assign n14543 = n6588 & ~n9957 ;
  assign n14544 = n6587 & n9955 ;
  assign n14545 = n14543 | n14544 ;
  assign n14546 = ( ~n14541 & n14542 ) | ( ~n14541 & n14545 ) | ( n14542 & n14545 ) ;
  assign n14547 = ( ~x11 & n14541 ) | ( ~x11 & n14546 ) | ( n14541 & n14546 ) ;
  assign n14548 = ( n14541 & n14546 ) | ( n14541 & ~n14547 ) | ( n14546 & ~n14547 ) ;
  assign n14549 = ( x11 & n14547 ) | ( x11 & ~n14548 ) | ( n14547 & ~n14548 ) ;
  assign n14550 = ( ~n14149 & n14151 ) | ( ~n14149 & n14160 ) | ( n14151 & n14160 ) ;
  assign n14551 = ( ~n14160 & n14161 ) | ( ~n14160 & n14550 ) | ( n14161 & n14550 ) ;
  assign n14552 = ( n14540 & n14549 ) | ( n14540 & ~n14551 ) | ( n14549 & ~n14551 ) ;
  assign n14553 = n6584 & ~n10652 ;
  assign n14554 = n7022 & n9951 ;
  assign n14555 = n6588 & n9955 ;
  assign n14556 = n6587 & ~n9953 ;
  assign n14557 = n14555 | n14556 ;
  assign n14558 = ( ~n14553 & n14554 ) | ( ~n14553 & n14557 ) | ( n14554 & n14557 ) ;
  assign n14559 = ( ~x11 & n14553 ) | ( ~x11 & n14558 ) | ( n14553 & n14558 ) ;
  assign n14560 = ( n14553 & n14558 ) | ( n14553 & ~n14559 ) | ( n14558 & ~n14559 ) ;
  assign n14561 = ( x11 & n14559 ) | ( x11 & ~n14560 ) | ( n14559 & ~n14560 ) ;
  assign n14562 = ( ~n14161 & n14163 ) | ( ~n14161 & n14172 ) | ( n14163 & n14172 ) ;
  assign n14563 = ( ~n14172 & n14173 ) | ( ~n14172 & n14562 ) | ( n14173 & n14562 ) ;
  assign n14564 = ( n14552 & n14561 ) | ( n14552 & ~n14563 ) | ( n14561 & ~n14563 ) ;
  assign n14565 = n6584 & n10557 ;
  assign n14566 = n7022 & n9949 ;
  assign n14567 = n6588 & ~n9953 ;
  assign n14568 = n6587 & n9951 ;
  assign n14569 = n14567 | n14568 ;
  assign n14570 = ( ~n14565 & n14566 ) | ( ~n14565 & n14569 ) | ( n14566 & n14569 ) ;
  assign n14571 = ( ~x11 & n14565 ) | ( ~x11 & n14570 ) | ( n14565 & n14570 ) ;
  assign n14572 = ( n14565 & n14570 ) | ( n14565 & ~n14571 ) | ( n14570 & ~n14571 ) ;
  assign n14573 = ( x11 & n14571 ) | ( x11 & ~n14572 ) | ( n14571 & ~n14572 ) ;
  assign n14574 = ( ~n14173 & n14175 ) | ( ~n14173 & n14184 ) | ( n14175 & n14184 ) ;
  assign n14575 = ( n14173 & ~n14185 ) | ( n14173 & n14574 ) | ( ~n14185 & n14574 ) ;
  assign n14576 = ( n14564 & n14573 ) | ( n14564 & n14575 ) | ( n14573 & n14575 ) ;
  assign n14577 = n6584 & n10454 ;
  assign n14578 = n7022 & n9947 ;
  assign n14579 = n6588 & n9951 ;
  assign n14580 = n6587 & n9949 ;
  assign n14581 = n14579 | n14580 ;
  assign n14582 = ( ~n14577 & n14578 ) | ( ~n14577 & n14581 ) | ( n14578 & n14581 ) ;
  assign n14583 = ( ~x11 & n14577 ) | ( ~x11 & n14582 ) | ( n14577 & n14582 ) ;
  assign n14584 = ( n14577 & n14582 ) | ( n14577 & ~n14583 ) | ( n14582 & ~n14583 ) ;
  assign n14585 = ( x11 & n14583 ) | ( x11 & ~n14584 ) | ( n14583 & ~n14584 ) ;
  assign n14586 = ( ~n14185 & n14187 ) | ( ~n14185 & n14196 ) | ( n14187 & n14196 ) ;
  assign n14587 = ( n14185 & ~n14197 ) | ( n14185 & n14586 ) | ( ~n14197 & n14586 ) ;
  assign n14588 = ( n14576 & n14585 ) | ( n14576 & n14587 ) | ( n14585 & n14587 ) ;
  assign n14589 = n6584 & n10466 ;
  assign n14590 = n7022 & n9945 ;
  assign n14591 = n6588 & n9949 ;
  assign n14592 = n6587 & n9947 ;
  assign n14593 = n14591 | n14592 ;
  assign n14594 = ( ~n14589 & n14590 ) | ( ~n14589 & n14593 ) | ( n14590 & n14593 ) ;
  assign n14595 = ( ~x11 & n14589 ) | ( ~x11 & n14594 ) | ( n14589 & n14594 ) ;
  assign n14596 = ( n14589 & n14594 ) | ( n14589 & ~n14595 ) | ( n14594 & ~n14595 ) ;
  assign n14597 = ( x11 & n14595 ) | ( x11 & ~n14596 ) | ( n14595 & ~n14596 ) ;
  assign n14598 = ( ~n14197 & n14199 ) | ( ~n14197 & n14208 ) | ( n14199 & n14208 ) ;
  assign n14599 = ( n14197 & ~n14209 ) | ( n14197 & n14598 ) | ( ~n14209 & n14598 ) ;
  assign n14600 = ( n14588 & n14597 ) | ( n14588 & n14599 ) | ( n14597 & n14599 ) ;
  assign n14601 = n6584 & n10271 ;
  assign n14602 = n7022 & n9943 ;
  assign n14603 = n6588 & n9947 ;
  assign n14604 = n6587 & n9945 ;
  assign n14605 = n14603 | n14604 ;
  assign n14606 = ( ~n14601 & n14602 ) | ( ~n14601 & n14605 ) | ( n14602 & n14605 ) ;
  assign n14607 = ( ~x11 & n14601 ) | ( ~x11 & n14606 ) | ( n14601 & n14606 ) ;
  assign n14608 = ( n14601 & n14606 ) | ( n14601 & ~n14607 ) | ( n14606 & ~n14607 ) ;
  assign n14609 = ( x11 & n14607 ) | ( x11 & ~n14608 ) | ( n14607 & ~n14608 ) ;
  assign n14610 = ( ~n14209 & n14211 ) | ( ~n14209 & n14220 ) | ( n14211 & n14220 ) ;
  assign n14611 = ( n14209 & ~n14221 ) | ( n14209 & n14610 ) | ( ~n14221 & n14610 ) ;
  assign n14612 = ( n14600 & n14609 ) | ( n14600 & n14611 ) | ( n14609 & n14611 ) ;
  assign n14613 = n6584 & ~n10390 ;
  assign n14614 = n7022 & ~n9941 ;
  assign n14615 = n6588 & n9945 ;
  assign n14616 = n6587 & n9943 ;
  assign n14617 = n14615 | n14616 ;
  assign n14618 = ( ~n14613 & n14614 ) | ( ~n14613 & n14617 ) | ( n14614 & n14617 ) ;
  assign n14619 = ( ~x11 & n14613 ) | ( ~x11 & n14618 ) | ( n14613 & n14618 ) ;
  assign n14620 = ( n14613 & n14618 ) | ( n14613 & ~n14619 ) | ( n14618 & ~n14619 ) ;
  assign n14621 = ( x11 & n14619 ) | ( x11 & ~n14620 ) | ( n14619 & ~n14620 ) ;
  assign n14622 = ( ~n14221 & n14223 ) | ( ~n14221 & n14232 ) | ( n14223 & n14232 ) ;
  assign n14623 = ( n14221 & ~n14233 ) | ( n14221 & n14622 ) | ( ~n14233 & n14622 ) ;
  assign n14624 = ( n14612 & n14621 ) | ( n14612 & n14623 ) | ( n14621 & n14623 ) ;
  assign n14625 = ( ~n14233 & n14235 ) | ( ~n14233 & n14244 ) | ( n14235 & n14244 ) ;
  assign n14626 = ( ~n14244 & n14245 ) | ( ~n14244 & n14625 ) | ( n14245 & n14625 ) ;
  assign n14627 = n7296 & ~n10064 ;
  assign n14628 = n7879 & ~n10057 ;
  assign n14629 = n7300 & n9916 ;
  assign n14630 = n7299 & ~n9937 ;
  assign n14631 = n14629 | n14630 ;
  assign n14632 = ( ~n14627 & n14628 ) | ( ~n14627 & n14631 ) | ( n14628 & n14631 ) ;
  assign n14633 = ( ~x8 & n14627 ) | ( ~x8 & n14632 ) | ( n14627 & n14632 ) ;
  assign n14634 = ( n14627 & n14632 ) | ( n14627 & ~n14633 ) | ( n14632 & ~n14633 ) ;
  assign n14635 = ( x8 & n14633 ) | ( x8 & ~n14634 ) | ( n14633 & ~n14634 ) ;
  assign n14636 = ( n14624 & ~n14626 ) | ( n14624 & n14635 ) | ( ~n14626 & n14635 ) ;
  assign n14637 = ( n14245 & ~n14247 ) | ( n14245 & n14256 ) | ( ~n14247 & n14256 ) ;
  assign n14638 = ( n14247 & ~n14257 ) | ( n14247 & n14637 ) | ( ~n14257 & n14637 ) ;
  assign n14639 = ~n8226 & n10346 ;
  assign n14640 = ( n10346 & n11389 ) | ( n10346 & ~n14639 ) | ( n11389 & ~n14639 ) ;
  assign n14641 = ( ~x5 & n8230 ) | ( ~x5 & n14640 ) | ( n8230 & n14640 ) ;
  assign n14642 = ( n8230 & n14640 ) | ( n8230 & ~n14641 ) | ( n14640 & ~n14641 ) ;
  assign n14643 = ( x5 & n14641 ) | ( x5 & ~n14642 ) | ( n14641 & ~n14642 ) ;
  assign n14644 = ( n14636 & n14638 ) | ( n14636 & n14643 ) | ( n14638 & n14643 ) ;
  assign n14645 = n7296 & n11892 ;
  assign n14646 = n7879 & ~n9997 ;
  assign n14647 = n7300 & ~n10001 ;
  assign n14648 = n7299 & n9999 ;
  assign n14649 = n14647 | n14648 ;
  assign n14650 = ( ~n14645 & n14646 ) | ( ~n14645 & n14649 ) | ( n14646 & n14649 ) ;
  assign n14651 = ( ~x8 & n14645 ) | ( ~x8 & n14650 ) | ( n14645 & n14650 ) ;
  assign n14652 = ( n14645 & n14650 ) | ( n14645 & ~n14651 ) | ( n14650 & ~n14651 ) ;
  assign n14653 = ( x8 & n14651 ) | ( x8 & ~n14652 ) | ( n14651 & ~n14652 ) ;
  assign n14654 = n7300 & ~n10003 ;
  assign n14655 = n7299 & ~n10001 ;
  assign n14656 = n14654 | n14655 ;
  assign n14657 = n7879 & ~n9999 ;
  assign n14658 = ( n7879 & n14656 ) | ( n7879 & ~n14657 ) | ( n14656 & ~n14657 ) ;
  assign n14659 = n7296 & n11868 ;
  assign n14660 = n14658 | n14659 ;
  assign n14661 = n7878 & ~n10003 ;
  assign n14662 = x8 & n14661 ;
  assign n14663 = ( n7296 & n11804 ) | ( n7296 & n11805 ) | ( n11804 & n11805 ) ;
  assign n14664 = n7299 | n10003 ;
  assign n14665 = n7879 & ~n10001 ;
  assign n14666 = ( ~n10003 & n14664 ) | ( ~n10003 & n14665 ) | ( n14664 & n14665 ) ;
  assign n14667 = n14663 | n14666 ;
  assign n14668 = ( x8 & n14662 ) | ( x8 & n14667 ) | ( n14662 & n14667 ) ;
  assign n14669 = n14660 | n14668 ;
  assign n14670 = x8 & ~n14669 ;
  assign n14671 = ( n14277 & n14653 ) | ( n14277 & n14670 ) | ( n14653 & n14670 ) ;
  assign n14672 = n7296 & n11934 ;
  assign n14673 = n7879 & n9995 ;
  assign n14674 = n7300 & n9999 ;
  assign n14675 = n7299 & ~n9997 ;
  assign n14676 = n14674 | n14675 ;
  assign n14677 = ( ~n14672 & n14673 ) | ( ~n14672 & n14676 ) | ( n14673 & n14676 ) ;
  assign n14678 = ( ~x8 & n14672 ) | ( ~x8 & n14677 ) | ( n14672 & n14677 ) ;
  assign n14679 = ( n14672 & n14677 ) | ( n14672 & ~n14678 ) | ( n14677 & ~n14678 ) ;
  assign n14680 = ( x8 & n14678 ) | ( x8 & ~n14679 ) | ( n14678 & ~n14679 ) ;
  assign n14681 = ( n14278 & n14279 ) | ( n14278 & n14282 ) | ( n14279 & n14282 ) ;
  assign n14682 = ~n14278 & n14283 ;
  assign n14683 = ( n14278 & ~n14681 ) | ( n14278 & n14682 ) | ( ~n14681 & n14682 ) ;
  assign n14684 = ( n14671 & n14680 ) | ( n14671 & n14683 ) | ( n14680 & n14683 ) ;
  assign n14685 = n7296 & ~n11971 ;
  assign n14686 = n7879 & n9993 ;
  assign n14687 = n7300 & ~n9997 ;
  assign n14688 = n7299 & n9995 ;
  assign n14689 = n14687 | n14688 ;
  assign n14690 = ( ~n14685 & n14686 ) | ( ~n14685 & n14689 ) | ( n14686 & n14689 ) ;
  assign n14691 = ( ~x8 & n14685 ) | ( ~x8 & n14690 ) | ( n14685 & n14690 ) ;
  assign n14692 = ( n14685 & n14690 ) | ( n14685 & ~n14691 ) | ( n14690 & ~n14691 ) ;
  assign n14693 = ( x8 & n14691 ) | ( x8 & ~n14692 ) | ( n14691 & ~n14692 ) ;
  assign n14694 = ( n14276 & n14284 ) | ( n14276 & ~n14285 ) | ( n14284 & ~n14285 ) ;
  assign n14695 = n14285 & ~n14694 ;
  assign n14696 = ( n14684 & n14693 ) | ( n14684 & n14695 ) | ( n14693 & n14695 ) ;
  assign n14697 = n7296 & n12026 ;
  assign n14698 = n7879 & n9991 ;
  assign n14699 = n7300 & n9995 ;
  assign n14700 = n7299 & n9993 ;
  assign n14701 = n14699 | n14700 ;
  assign n14702 = ( ~n14697 & n14698 ) | ( ~n14697 & n14701 ) | ( n14698 & n14701 ) ;
  assign n14703 = ( ~x8 & n14697 ) | ( ~x8 & n14702 ) | ( n14697 & n14702 ) ;
  assign n14704 = ( n14697 & n14702 ) | ( n14697 & ~n14703 ) | ( n14702 & ~n14703 ) ;
  assign n14705 = ( x8 & n14703 ) | ( x8 & ~n14704 ) | ( n14703 & ~n14704 ) ;
  assign n14706 = ( n13922 & n14269 ) | ( n13922 & ~n14286 ) | ( n14269 & ~n14286 ) ;
  assign n14707 = ( n14286 & ~n14287 ) | ( n14286 & n14706 ) | ( ~n14287 & n14706 ) ;
  assign n14708 = ( n14696 & n14705 ) | ( n14696 & n14707 ) | ( n14705 & n14707 ) ;
  assign n14709 = n7296 & n12050 ;
  assign n14710 = n7879 & n9989 ;
  assign n14711 = n7300 & n9993 ;
  assign n14712 = n7299 & n9991 ;
  assign n14713 = n14711 | n14712 ;
  assign n14714 = ( ~n14709 & n14710 ) | ( ~n14709 & n14713 ) | ( n14710 & n14713 ) ;
  assign n14715 = ( ~x8 & n14709 ) | ( ~x8 & n14714 ) | ( n14709 & n14714 ) ;
  assign n14716 = ( n14709 & n14714 ) | ( n14709 & ~n14715 ) | ( n14714 & ~n14715 ) ;
  assign n14717 = ( x8 & n14715 ) | ( x8 & ~n14716 ) | ( n14715 & ~n14716 ) ;
  assign n14718 = ( ~n14287 & n14296 ) | ( ~n14287 & n14299 ) | ( n14296 & n14299 ) ;
  assign n14719 = ( n14287 & ~n14300 ) | ( n14287 & n14718 ) | ( ~n14300 & n14718 ) ;
  assign n14720 = ( n14708 & n14717 ) | ( n14708 & n14719 ) | ( n14717 & n14719 ) ;
  assign n14721 = ( ~n14300 & n14309 ) | ( ~n14300 & n14311 ) | ( n14309 & n14311 ) ;
  assign n14722 = ( n14300 & ~n14312 ) | ( n14300 & n14721 ) | ( ~n14312 & n14721 ) ;
  assign n14723 = n7296 & ~n12074 ;
  assign n14724 = n7879 & ~n9987 ;
  assign n14725 = n7300 & n9991 ;
  assign n14726 = n7299 & n9989 ;
  assign n14727 = n14725 | n14726 ;
  assign n14728 = ( ~n14723 & n14724 ) | ( ~n14723 & n14727 ) | ( n14724 & n14727 ) ;
  assign n14729 = ( ~x8 & n14723 ) | ( ~x8 & n14728 ) | ( n14723 & n14728 ) ;
  assign n14730 = ( n14723 & n14728 ) | ( n14723 & ~n14729 ) | ( n14728 & ~n14729 ) ;
  assign n14731 = ( x8 & n14729 ) | ( x8 & ~n14730 ) | ( n14729 & ~n14730 ) ;
  assign n14732 = ( n14720 & n14722 ) | ( n14720 & n14731 ) | ( n14722 & n14731 ) ;
  assign n14733 = ( ~n14312 & n14321 ) | ( ~n14312 & n14323 ) | ( n14321 & n14323 ) ;
  assign n14734 = ( n14312 & ~n14324 ) | ( n14312 & n14733 ) | ( ~n14324 & n14733 ) ;
  assign n14735 = n7296 & ~n12099 ;
  assign n14736 = n7879 & n9985 ;
  assign n14737 = n7300 & n9989 ;
  assign n14738 = n7299 & ~n9987 ;
  assign n14739 = n14737 | n14738 ;
  assign n14740 = ( ~n14735 & n14736 ) | ( ~n14735 & n14739 ) | ( n14736 & n14739 ) ;
  assign n14741 = ( ~x8 & n14735 ) | ( ~x8 & n14740 ) | ( n14735 & n14740 ) ;
  assign n14742 = ( n14735 & n14740 ) | ( n14735 & ~n14741 ) | ( n14740 & ~n14741 ) ;
  assign n14743 = ( x8 & n14741 ) | ( x8 & ~n14742 ) | ( n14741 & ~n14742 ) ;
  assign n14744 = ( n14732 & n14734 ) | ( n14732 & n14743 ) | ( n14734 & n14743 ) ;
  assign n14745 = ( ~n14324 & n14333 ) | ( ~n14324 & n14335 ) | ( n14333 & n14335 ) ;
  assign n14746 = ( n14324 & ~n14336 ) | ( n14324 & n14745 ) | ( ~n14336 & n14745 ) ;
  assign n14747 = n7296 & ~n12129 ;
  assign n14748 = n7879 & ~n9983 ;
  assign n14749 = n7300 & ~n9987 ;
  assign n14750 = n7299 & n9985 ;
  assign n14751 = n14749 | n14750 ;
  assign n14752 = ( ~n14747 & n14748 ) | ( ~n14747 & n14751 ) | ( n14748 & n14751 ) ;
  assign n14753 = ( ~x8 & n14747 ) | ( ~x8 & n14752 ) | ( n14747 & n14752 ) ;
  assign n14754 = ( n14747 & n14752 ) | ( n14747 & ~n14753 ) | ( n14752 & ~n14753 ) ;
  assign n14755 = ( x8 & n14753 ) | ( x8 & ~n14754 ) | ( n14753 & ~n14754 ) ;
  assign n14756 = ( n14744 & n14746 ) | ( n14744 & n14755 ) | ( n14746 & n14755 ) ;
  assign n14757 = n7296 & ~n11561 ;
  assign n14758 = n7879 & n9981 ;
  assign n14759 = n7300 & n9985 ;
  assign n14760 = n7299 & ~n9983 ;
  assign n14761 = n14759 | n14760 ;
  assign n14762 = ( ~n14757 & n14758 ) | ( ~n14757 & n14761 ) | ( n14758 & n14761 ) ;
  assign n14763 = ( ~x8 & n14757 ) | ( ~x8 & n14762 ) | ( n14757 & n14762 ) ;
  assign n14764 = ( n14757 & n14762 ) | ( n14757 & ~n14763 ) | ( n14762 & ~n14763 ) ;
  assign n14765 = ( x8 & n14763 ) | ( x8 & ~n14764 ) | ( n14763 & ~n14764 ) ;
  assign n14766 = ( ~n14336 & n14338 ) | ( ~n14336 & n14347 ) | ( n14338 & n14347 ) ;
  assign n14767 = ( n14336 & ~n14348 ) | ( n14336 & n14766 ) | ( ~n14348 & n14766 ) ;
  assign n14768 = ( n14756 & n14765 ) | ( n14756 & n14767 ) | ( n14765 & n14767 ) ;
  assign n14769 = n7296 & n12153 ;
  assign n14770 = n7879 & n9979 ;
  assign n14771 = n7300 & ~n9983 ;
  assign n14772 = n7299 & n9981 ;
  assign n14773 = n14771 | n14772 ;
  assign n14774 = ( ~n14769 & n14770 ) | ( ~n14769 & n14773 ) | ( n14770 & n14773 ) ;
  assign n14775 = ( ~x8 & n14769 ) | ( ~x8 & n14774 ) | ( n14769 & n14774 ) ;
  assign n14776 = ( n14769 & n14774 ) | ( n14769 & ~n14775 ) | ( n14774 & ~n14775 ) ;
  assign n14777 = ( x8 & n14775 ) | ( x8 & ~n14776 ) | ( n14775 & ~n14776 ) ;
  assign n14778 = ( ~n14348 & n14350 ) | ( ~n14348 & n14359 ) | ( n14350 & n14359 ) ;
  assign n14779 = ( n14348 & ~n14360 ) | ( n14348 & n14778 ) | ( ~n14360 & n14778 ) ;
  assign n14780 = ( n14768 & n14777 ) | ( n14768 & n14779 ) | ( n14777 & n14779 ) ;
  assign n14781 = n7296 & n12165 ;
  assign n14782 = n7879 & n9977 ;
  assign n14783 = n7300 & n9981 ;
  assign n14784 = n7299 & n9979 ;
  assign n14785 = n14783 | n14784 ;
  assign n14786 = ( ~n14781 & n14782 ) | ( ~n14781 & n14785 ) | ( n14782 & n14785 ) ;
  assign n14787 = ( ~x8 & n14781 ) | ( ~x8 & n14786 ) | ( n14781 & n14786 ) ;
  assign n14788 = ( n14781 & n14786 ) | ( n14781 & ~n14787 ) | ( n14786 & ~n14787 ) ;
  assign n14789 = ( x8 & n14787 ) | ( x8 & ~n14788 ) | ( n14787 & ~n14788 ) ;
  assign n14790 = ( ~n14360 & n14362 ) | ( ~n14360 & n14371 ) | ( n14362 & n14371 ) ;
  assign n14791 = ( n14360 & ~n14372 ) | ( n14360 & n14790 ) | ( ~n14372 & n14790 ) ;
  assign n14792 = ( n14780 & n14789 ) | ( n14780 & n14791 ) | ( n14789 & n14791 ) ;
  assign n14793 = ( ~n14372 & n14381 ) | ( ~n14372 & n14383 ) | ( n14381 & n14383 ) ;
  assign n14794 = ( n14372 & ~n14384 ) | ( n14372 & n14793 ) | ( ~n14384 & n14793 ) ;
  assign n14795 = n7296 & n11606 ;
  assign n14796 = n7879 & n9975 ;
  assign n14797 = n7300 & n9979 ;
  assign n14798 = n7299 & n9977 ;
  assign n14799 = n14797 | n14798 ;
  assign n14800 = ( ~n14795 & n14796 ) | ( ~n14795 & n14799 ) | ( n14796 & n14799 ) ;
  assign n14801 = ( ~x8 & n14795 ) | ( ~x8 & n14800 ) | ( n14795 & n14800 ) ;
  assign n14802 = ( n14795 & n14800 ) | ( n14795 & ~n14801 ) | ( n14800 & ~n14801 ) ;
  assign n14803 = ( x8 & n14801 ) | ( x8 & ~n14802 ) | ( n14801 & ~n14802 ) ;
  assign n14804 = ( n14792 & n14794 ) | ( n14792 & n14803 ) | ( n14794 & n14803 ) ;
  assign n14805 = ( ~n14384 & n14393 ) | ( ~n14384 & n14395 ) | ( n14393 & n14395 ) ;
  assign n14806 = ( n14384 & ~n14396 ) | ( n14384 & n14805 ) | ( ~n14396 & n14805 ) ;
  assign n14807 = n7296 & n11400 ;
  assign n14808 = n7879 & n9973 ;
  assign n14809 = n7300 & n9977 ;
  assign n14810 = n7299 & n9975 ;
  assign n14811 = n14809 | n14810 ;
  assign n14812 = ( ~n14807 & n14808 ) | ( ~n14807 & n14811 ) | ( n14808 & n14811 ) ;
  assign n14813 = ( ~x8 & n14807 ) | ( ~x8 & n14812 ) | ( n14807 & n14812 ) ;
  assign n14814 = ( n14807 & n14812 ) | ( n14807 & ~n14813 ) | ( n14812 & ~n14813 ) ;
  assign n14815 = ( x8 & n14813 ) | ( x8 & ~n14814 ) | ( n14813 & ~n14814 ) ;
  assign n14816 = ( n14804 & n14806 ) | ( n14804 & n14815 ) | ( n14806 & n14815 ) ;
  assign n14817 = ( ~n14396 & n14405 ) | ( ~n14396 & n14407 ) | ( n14405 & n14407 ) ;
  assign n14818 = ( n14396 & ~n14408 ) | ( n14396 & n14817 ) | ( ~n14408 & n14817 ) ;
  assign n14819 = n7296 & n11630 ;
  assign n14820 = n7879 & n9971 ;
  assign n14821 = n7300 & n9975 ;
  assign n14822 = n7299 & n9973 ;
  assign n14823 = n14821 | n14822 ;
  assign n14824 = ( ~n14819 & n14820 ) | ( ~n14819 & n14823 ) | ( n14820 & n14823 ) ;
  assign n14825 = ( ~x8 & n14819 ) | ( ~x8 & n14824 ) | ( n14819 & n14824 ) ;
  assign n14826 = ( n14819 & n14824 ) | ( n14819 & ~n14825 ) | ( n14824 & ~n14825 ) ;
  assign n14827 = ( x8 & n14825 ) | ( x8 & ~n14826 ) | ( n14825 & ~n14826 ) ;
  assign n14828 = ( n14816 & n14818 ) | ( n14816 & n14827 ) | ( n14818 & n14827 ) ;
  assign n14829 = n7296 & n11428 ;
  assign n14830 = n7879 & n9969 ;
  assign n14831 = n7300 & n9973 ;
  assign n14832 = n7299 & n9971 ;
  assign n14833 = n14831 | n14832 ;
  assign n14834 = ( ~n14829 & n14830 ) | ( ~n14829 & n14833 ) | ( n14830 & n14833 ) ;
  assign n14835 = ( ~x8 & n14829 ) | ( ~x8 & n14834 ) | ( n14829 & n14834 ) ;
  assign n14836 = ( n14829 & n14834 ) | ( n14829 & ~n14835 ) | ( n14834 & ~n14835 ) ;
  assign n14837 = ( x8 & n14835 ) | ( x8 & ~n14836 ) | ( n14835 & ~n14836 ) ;
  assign n14838 = ( ~n14408 & n14410 ) | ( ~n14408 & n14419 ) | ( n14410 & n14419 ) ;
  assign n14839 = ( n14408 & ~n14420 ) | ( n14408 & n14838 ) | ( ~n14420 & n14838 ) ;
  assign n14840 = ( n14828 & n14837 ) | ( n14828 & n14839 ) | ( n14837 & n14839 ) ;
  assign n14841 = n7296 & ~n10998 ;
  assign n14842 = n7879 & ~n9967 ;
  assign n14843 = n7300 & n9971 ;
  assign n14844 = n7299 & n9969 ;
  assign n14845 = n14843 | n14844 ;
  assign n14846 = ( ~n14841 & n14842 ) | ( ~n14841 & n14845 ) | ( n14842 & n14845 ) ;
  assign n14847 = ( ~x8 & n14841 ) | ( ~x8 & n14846 ) | ( n14841 & n14846 ) ;
  assign n14848 = ( n14841 & n14846 ) | ( n14841 & ~n14847 ) | ( n14846 & ~n14847 ) ;
  assign n14849 = ( x8 & n14847 ) | ( x8 & ~n14848 ) | ( n14847 & ~n14848 ) ;
  assign n14850 = ( ~n14420 & n14422 ) | ( ~n14420 & n14431 ) | ( n14422 & n14431 ) ;
  assign n14851 = ( n14420 & ~n14432 ) | ( n14420 & n14850 ) | ( ~n14432 & n14850 ) ;
  assign n14852 = ( n14840 & n14849 ) | ( n14840 & n14851 ) | ( n14849 & n14851 ) ;
  assign n14853 = n7296 & ~n11273 ;
  assign n14854 = n7879 & n9965 ;
  assign n14855 = n7300 & n9969 ;
  assign n14856 = n7299 & ~n9967 ;
  assign n14857 = n14855 | n14856 ;
  assign n14858 = ( ~n14853 & n14854 ) | ( ~n14853 & n14857 ) | ( n14854 & n14857 ) ;
  assign n14859 = ( ~x8 & n14853 ) | ( ~x8 & n14858 ) | ( n14853 & n14858 ) ;
  assign n14860 = ( n14853 & n14858 ) | ( n14853 & ~n14859 ) | ( n14858 & ~n14859 ) ;
  assign n14861 = ( x8 & n14859 ) | ( x8 & ~n14860 ) | ( n14859 & ~n14860 ) ;
  assign n14862 = ( ~n14432 & n14434 ) | ( ~n14432 & n14443 ) | ( n14434 & n14443 ) ;
  assign n14863 = ( n14432 & ~n14444 ) | ( n14432 & n14862 ) | ( ~n14444 & n14862 ) ;
  assign n14864 = ( n14852 & n14861 ) | ( n14852 & n14863 ) | ( n14861 & n14863 ) ;
  assign n14865 = ( ~n14444 & n14453 ) | ( ~n14444 & n14455 ) | ( n14453 & n14455 ) ;
  assign n14866 = ( n14444 & ~n14456 ) | ( n14444 & n14865 ) | ( ~n14456 & n14865 ) ;
  assign n14867 = n7296 & ~n11121 ;
  assign n14868 = n7879 & ~n9963 ;
  assign n14869 = n7300 & ~n9967 ;
  assign n14870 = n7299 & n9965 ;
  assign n14871 = n14869 | n14870 ;
  assign n14872 = ( ~n14867 & n14868 ) | ( ~n14867 & n14871 ) | ( n14868 & n14871 ) ;
  assign n14873 = ( ~x8 & n14867 ) | ( ~x8 & n14872 ) | ( n14867 & n14872 ) ;
  assign n14874 = ( n14867 & n14872 ) | ( n14867 & ~n14873 ) | ( n14872 & ~n14873 ) ;
  assign n14875 = ( x8 & n14873 ) | ( x8 & ~n14874 ) | ( n14873 & ~n14874 ) ;
  assign n14876 = ( n14864 & n14866 ) | ( n14864 & n14875 ) | ( n14866 & n14875 ) ;
  assign n14877 = ( ~n14456 & n14465 ) | ( ~n14456 & n14467 ) | ( n14465 & n14467 ) ;
  assign n14878 = ( n14456 & ~n14468 ) | ( n14456 & n14877 ) | ( ~n14468 & n14877 ) ;
  assign n14879 = n7296 & ~n10929 ;
  assign n14880 = n7879 & n9961 ;
  assign n14881 = n7300 & n9965 ;
  assign n14882 = n7299 & ~n9963 ;
  assign n14883 = n14881 | n14882 ;
  assign n14884 = ( ~n14879 & n14880 ) | ( ~n14879 & n14883 ) | ( n14880 & n14883 ) ;
  assign n14885 = ( ~x8 & n14879 ) | ( ~x8 & n14884 ) | ( n14879 & n14884 ) ;
  assign n14886 = ( n14879 & n14884 ) | ( n14879 & ~n14885 ) | ( n14884 & ~n14885 ) ;
  assign n14887 = ( x8 & n14885 ) | ( x8 & ~n14886 ) | ( n14885 & ~n14886 ) ;
  assign n14888 = ( n14876 & n14878 ) | ( n14876 & n14887 ) | ( n14878 & n14887 ) ;
  assign n14889 = ( ~n14468 & n14477 ) | ( ~n14468 & n14479 ) | ( n14477 & n14479 ) ;
  assign n14890 = ( n14468 & ~n14480 ) | ( n14468 & n14889 ) | ( ~n14480 & n14889 ) ;
  assign n14891 = n7296 & n10859 ;
  assign n14892 = n7879 & n9959 ;
  assign n14893 = n7300 & ~n9963 ;
  assign n14894 = n7299 & n9961 ;
  assign n14895 = n14893 | n14894 ;
  assign n14896 = ( ~n14891 & n14892 ) | ( ~n14891 & n14895 ) | ( n14892 & n14895 ) ;
  assign n14897 = ( ~x8 & n14891 ) | ( ~x8 & n14896 ) | ( n14891 & n14896 ) ;
  assign n14898 = ( n14891 & n14896 ) | ( n14891 & ~n14897 ) | ( n14896 & ~n14897 ) ;
  assign n14899 = ( x8 & n14897 ) | ( x8 & ~n14898 ) | ( n14897 & ~n14898 ) ;
  assign n14900 = ( n14888 & n14890 ) | ( n14888 & n14899 ) | ( n14890 & n14899 ) ;
  assign n14901 = n7296 & ~n10869 ;
  assign n14902 = n7879 & ~n9957 ;
  assign n14903 = n7300 & n9961 ;
  assign n14904 = n7299 & n9959 ;
  assign n14905 = n14903 | n14904 ;
  assign n14906 = ( ~n14901 & n14902 ) | ( ~n14901 & n14905 ) | ( n14902 & n14905 ) ;
  assign n14907 = ( ~x8 & n14901 ) | ( ~x8 & n14906 ) | ( n14901 & n14906 ) ;
  assign n14908 = ( n14901 & n14906 ) | ( n14901 & ~n14907 ) | ( n14906 & ~n14907 ) ;
  assign n14909 = ( x8 & n14907 ) | ( x8 & ~n14908 ) | ( n14907 & ~n14908 ) ;
  assign n14910 = ( ~n14480 & n14482 ) | ( ~n14480 & n14491 ) | ( n14482 & n14491 ) ;
  assign n14911 = ( n14480 & ~n14492 ) | ( n14480 & n14910 ) | ( ~n14492 & n14910 ) ;
  assign n14912 = ( n14900 & n14909 ) | ( n14900 & n14911 ) | ( n14909 & n14911 ) ;
  assign n14913 = n7296 & ~n10567 ;
  assign n14914 = n7879 & n9955 ;
  assign n14915 = n7300 & n9959 ;
  assign n14916 = n7299 & ~n9957 ;
  assign n14917 = n14915 | n14916 ;
  assign n14918 = ( ~n14913 & n14914 ) | ( ~n14913 & n14917 ) | ( n14914 & n14917 ) ;
  assign n14919 = ( ~x8 & n14913 ) | ( ~x8 & n14918 ) | ( n14913 & n14918 ) ;
  assign n14920 = ( n14913 & n14918 ) | ( n14913 & ~n14919 ) | ( n14918 & ~n14919 ) ;
  assign n14921 = ( x8 & n14919 ) | ( x8 & ~n14920 ) | ( n14919 & ~n14920 ) ;
  assign n14922 = ( ~n14492 & n14494 ) | ( ~n14492 & n14503 ) | ( n14494 & n14503 ) ;
  assign n14923 = ( n14492 & ~n14504 ) | ( n14492 & n14922 ) | ( ~n14504 & n14922 ) ;
  assign n14924 = ( n14912 & n14921 ) | ( n14912 & n14923 ) | ( n14921 & n14923 ) ;
  assign n14925 = ( n14504 & ~n14513 ) | ( n14504 & n14515 ) | ( ~n14513 & n14515 ) ;
  assign n14926 = ( ~n14504 & n14516 ) | ( ~n14504 & n14925 ) | ( n14516 & n14925 ) ;
  assign n14927 = n7296 & ~n10750 ;
  assign n14928 = n7879 & ~n9953 ;
  assign n14929 = n7300 & ~n9957 ;
  assign n14930 = n7299 & n9955 ;
  assign n14931 = n14929 | n14930 ;
  assign n14932 = ( ~n14927 & n14928 ) | ( ~n14927 & n14931 ) | ( n14928 & n14931 ) ;
  assign n14933 = ( ~x8 & n14927 ) | ( ~x8 & n14932 ) | ( n14927 & n14932 ) ;
  assign n14934 = ( n14927 & n14932 ) | ( n14927 & ~n14933 ) | ( n14932 & ~n14933 ) ;
  assign n14935 = ( x8 & n14933 ) | ( x8 & ~n14934 ) | ( n14933 & ~n14934 ) ;
  assign n14936 = ( n14924 & ~n14926 ) | ( n14924 & n14935 ) | ( ~n14926 & n14935 ) ;
  assign n14937 = ( n14516 & ~n14525 ) | ( n14516 & n14527 ) | ( ~n14525 & n14527 ) ;
  assign n14938 = ( ~n14516 & n14528 ) | ( ~n14516 & n14937 ) | ( n14528 & n14937 ) ;
  assign n14939 = n7296 & ~n10652 ;
  assign n14940 = n7879 & n9951 ;
  assign n14941 = n7300 & n9955 ;
  assign n14942 = n7299 & ~n9953 ;
  assign n14943 = n14941 | n14942 ;
  assign n14944 = ( ~n14939 & n14940 ) | ( ~n14939 & n14943 ) | ( n14940 & n14943 ) ;
  assign n14945 = ( ~x8 & n14939 ) | ( ~x8 & n14944 ) | ( n14939 & n14944 ) ;
  assign n14946 = ( n14939 & n14944 ) | ( n14939 & ~n14945 ) | ( n14944 & ~n14945 ) ;
  assign n14947 = ( x8 & n14945 ) | ( x8 & ~n14946 ) | ( n14945 & ~n14946 ) ;
  assign n14948 = ( n14936 & ~n14938 ) | ( n14936 & n14947 ) | ( ~n14938 & n14947 ) ;
  assign n14949 = ( ~n14528 & n14537 ) | ( ~n14528 & n14539 ) | ( n14537 & n14539 ) ;
  assign n14950 = ( n14528 & ~n14540 ) | ( n14528 & n14949 ) | ( ~n14540 & n14949 ) ;
  assign n14951 = n7296 & n10557 ;
  assign n14952 = n7879 & n9949 ;
  assign n14953 = n7300 & ~n9953 ;
  assign n14954 = n7299 & n9951 ;
  assign n14955 = n14953 | n14954 ;
  assign n14956 = ( ~n14951 & n14952 ) | ( ~n14951 & n14955 ) | ( n14952 & n14955 ) ;
  assign n14957 = ( ~x8 & n14951 ) | ( ~x8 & n14956 ) | ( n14951 & n14956 ) ;
  assign n14958 = ( n14951 & n14956 ) | ( n14951 & ~n14957 ) | ( n14956 & ~n14957 ) ;
  assign n14959 = ( x8 & n14957 ) | ( x8 & ~n14958 ) | ( n14957 & ~n14958 ) ;
  assign n14960 = ( n14948 & n14950 ) | ( n14948 & n14959 ) | ( n14950 & n14959 ) ;
  assign n14961 = ( n14540 & ~n14549 ) | ( n14540 & n14551 ) | ( ~n14549 & n14551 ) ;
  assign n14962 = ( ~n14540 & n14552 ) | ( ~n14540 & n14961 ) | ( n14552 & n14961 ) ;
  assign n14963 = n7296 & n10454 ;
  assign n14964 = n7879 & n9947 ;
  assign n14965 = n7300 & n9951 ;
  assign n14966 = n7299 & n9949 ;
  assign n14967 = n14965 | n14966 ;
  assign n14968 = ( ~n14963 & n14964 ) | ( ~n14963 & n14967 ) | ( n14964 & n14967 ) ;
  assign n14969 = ( ~x8 & n14963 ) | ( ~x8 & n14968 ) | ( n14963 & n14968 ) ;
  assign n14970 = ( n14963 & n14968 ) | ( n14963 & ~n14969 ) | ( n14968 & ~n14969 ) ;
  assign n14971 = ( x8 & n14969 ) | ( x8 & ~n14970 ) | ( n14969 & ~n14970 ) ;
  assign n14972 = ( n14960 & ~n14962 ) | ( n14960 & n14971 ) | ( ~n14962 & n14971 ) ;
  assign n14973 = ( n14552 & ~n14561 ) | ( n14552 & n14563 ) | ( ~n14561 & n14563 ) ;
  assign n14974 = ( ~n14552 & n14564 ) | ( ~n14552 & n14973 ) | ( n14564 & n14973 ) ;
  assign n14975 = n7296 & n10466 ;
  assign n14976 = n7879 & n9945 ;
  assign n14977 = n7300 & n9949 ;
  assign n14978 = n7299 & n9947 ;
  assign n14979 = n14977 | n14978 ;
  assign n14980 = ( ~n14975 & n14976 ) | ( ~n14975 & n14979 ) | ( n14976 & n14979 ) ;
  assign n14981 = ( ~x8 & n14975 ) | ( ~x8 & n14980 ) | ( n14975 & n14980 ) ;
  assign n14982 = ( n14975 & n14980 ) | ( n14975 & ~n14981 ) | ( n14980 & ~n14981 ) ;
  assign n14983 = ( x8 & n14981 ) | ( x8 & ~n14982 ) | ( n14981 & ~n14982 ) ;
  assign n14984 = ( n14972 & ~n14974 ) | ( n14972 & n14983 ) | ( ~n14974 & n14983 ) ;
  assign n14985 = ( ~n14564 & n14573 ) | ( ~n14564 & n14575 ) | ( n14573 & n14575 ) ;
  assign n14986 = ( n14564 & ~n14576 ) | ( n14564 & n14985 ) | ( ~n14576 & n14985 ) ;
  assign n14987 = n7296 & n10271 ;
  assign n14988 = n7879 & n9943 ;
  assign n14989 = n7300 & n9947 ;
  assign n14990 = n7299 & n9945 ;
  assign n14991 = n14989 | n14990 ;
  assign n14992 = ( ~n14987 & n14988 ) | ( ~n14987 & n14991 ) | ( n14988 & n14991 ) ;
  assign n14993 = ( ~x8 & n14987 ) | ( ~x8 & n14992 ) | ( n14987 & n14992 ) ;
  assign n14994 = ( n14987 & n14992 ) | ( n14987 & ~n14993 ) | ( n14992 & ~n14993 ) ;
  assign n14995 = ( x8 & n14993 ) | ( x8 & ~n14994 ) | ( n14993 & ~n14994 ) ;
  assign n14996 = ( n14984 & n14986 ) | ( n14984 & n14995 ) | ( n14986 & n14995 ) ;
  assign n14997 = ( ~n14576 & n14585 ) | ( ~n14576 & n14587 ) | ( n14585 & n14587 ) ;
  assign n14998 = ( n14576 & ~n14588 ) | ( n14576 & n14997 ) | ( ~n14588 & n14997 ) ;
  assign n14999 = n7296 & ~n10390 ;
  assign n15000 = n7879 & ~n9941 ;
  assign n15001 = n7300 & n9945 ;
  assign n15002 = n7299 & n9943 ;
  assign n15003 = n15001 | n15002 ;
  assign n15004 = ( ~n14999 & n15000 ) | ( ~n14999 & n15003 ) | ( n15000 & n15003 ) ;
  assign n15005 = ( ~x8 & n14999 ) | ( ~x8 & n15004 ) | ( n14999 & n15004 ) ;
  assign n15006 = ( n14999 & n15004 ) | ( n14999 & ~n15005 ) | ( n15004 & ~n15005 ) ;
  assign n15007 = ( x8 & n15005 ) | ( x8 & ~n15006 ) | ( n15005 & ~n15006 ) ;
  assign n15008 = ( n14996 & n14998 ) | ( n14996 & n15007 ) | ( n14998 & n15007 ) ;
  assign n15009 = ( ~n14588 & n14597 ) | ( ~n14588 & n14599 ) | ( n14597 & n14599 ) ;
  assign n15010 = ( n14588 & ~n14600 ) | ( n14588 & n15009 ) | ( ~n14600 & n15009 ) ;
  assign n15011 = n7296 & n10284 ;
  assign n15012 = n7879 & ~n9883 ;
  assign n15013 = n7300 & n9943 ;
  assign n15014 = n7299 & ~n9941 ;
  assign n15015 = n15013 | n15014 ;
  assign n15016 = ( ~n15011 & n15012 ) | ( ~n15011 & n15015 ) | ( n15012 & n15015 ) ;
  assign n15017 = ( ~x8 & n15011 ) | ( ~x8 & n15016 ) | ( n15011 & n15016 ) ;
  assign n15018 = ( n15011 & n15016 ) | ( n15011 & ~n15017 ) | ( n15016 & ~n15017 ) ;
  assign n15019 = ( x8 & n15017 ) | ( x8 & ~n15018 ) | ( n15017 & ~n15018 ) ;
  assign n15020 = ( n15008 & n15010 ) | ( n15008 & n15019 ) | ( n15010 & n15019 ) ;
  assign n15021 = ( ~n14600 & n14609 ) | ( ~n14600 & n14611 ) | ( n14609 & n14611 ) ;
  assign n15022 = ( n14600 & ~n14612 ) | ( n14600 & n15021 ) | ( ~n14612 & n15021 ) ;
  assign n15023 = n7296 & n10174 ;
  assign n15024 = n7879 & n9916 ;
  assign n15025 = n7299 | n9883 ;
  assign n15026 = n7300 & ~n9941 ;
  assign n15027 = ( ~n9883 & n15025 ) | ( ~n9883 & n15026 ) | ( n15025 & n15026 ) ;
  assign n15028 = ( ~n15023 & n15024 ) | ( ~n15023 & n15027 ) | ( n15024 & n15027 ) ;
  assign n15029 = ( ~x8 & n15023 ) | ( ~x8 & n15028 ) | ( n15023 & n15028 ) ;
  assign n15030 = ( n15023 & n15028 ) | ( n15023 & ~n15029 ) | ( n15028 & ~n15029 ) ;
  assign n15031 = ( x8 & n15029 ) | ( x8 & ~n15030 ) | ( n15029 & ~n15030 ) ;
  assign n15032 = ( n15020 & n15022 ) | ( n15020 & n15031 ) | ( n15022 & n15031 ) ;
  assign n15033 = ( ~n14612 & n14621 ) | ( ~n14612 & n14623 ) | ( n14621 & n14623 ) ;
  assign n15034 = ( n14612 & ~n14624 ) | ( n14612 & n15033 ) | ( ~n14624 & n15033 ) ;
  assign n15035 = n7296 & n10040 ;
  assign n15036 = n7879 & ~n9937 ;
  assign n15037 = n7300 & ~n9883 ;
  assign n15038 = n7299 & n9916 ;
  assign n15039 = n15037 | n15038 ;
  assign n15040 = ( ~n15035 & n15036 ) | ( ~n15035 & n15039 ) | ( n15036 & n15039 ) ;
  assign n15041 = ( ~x8 & n15035 ) | ( ~x8 & n15040 ) | ( n15035 & n15040 ) ;
  assign n15042 = ( n15035 & n15040 ) | ( n15035 & ~n15041 ) | ( n15040 & ~n15041 ) ;
  assign n15043 = ( x8 & n15041 ) | ( x8 & ~n15042 ) | ( n15041 & ~n15042 ) ;
  assign n15044 = ( n15032 & n15034 ) | ( n15032 & n15043 ) | ( n15034 & n15043 ) ;
  assign n15045 = ( ~n14624 & n14626 ) | ( ~n14624 & n14635 ) | ( n14626 & n14635 ) ;
  assign n15046 = ( ~n14635 & n14636 ) | ( ~n14635 & n15045 ) | ( n14636 & n15045 ) ;
  assign n15047 = n8230 & n10348 ;
  assign n15048 = n8225 & n10346 ;
  assign n15049 = n8226 & ~n10302 ;
  assign n15050 = n8229 | n15049 ;
  assign n15051 = ( ~n15047 & n15048 ) | ( ~n15047 & n15050 ) | ( n15048 & n15050 ) ;
  assign n15052 = ( ~x5 & n15047 ) | ( ~x5 & n15051 ) | ( n15047 & n15051 ) ;
  assign n15053 = ( n15047 & n15051 ) | ( n15047 & ~n15052 ) | ( n15051 & ~n15052 ) ;
  assign n15054 = ( x5 & n15052 ) | ( x5 & ~n15053 ) | ( n15052 & ~n15053 ) ;
  assign n15055 = ( n15044 & ~n15046 ) | ( n15044 & n15054 ) | ( ~n15046 & n15054 ) ;
  assign n15056 = n8230 & n10362 ;
  assign n15057 = n8229 & n10346 ;
  assign n15058 = n8226 & ~n10057 ;
  assign n15059 = n8225 & ~n10302 ;
  assign n15060 = n15058 | n15059 ;
  assign n15061 = ( ~n15056 & n15057 ) | ( ~n15056 & n15060 ) | ( n15057 & n15060 ) ;
  assign n15062 = ( ~x5 & n15056 ) | ( ~x5 & n15061 ) | ( n15056 & n15061 ) ;
  assign n15063 = ( n15056 & n15061 ) | ( n15056 & ~n15062 ) | ( n15061 & ~n15062 ) ;
  assign n15064 = ( x5 & n15062 ) | ( x5 & ~n15063 ) | ( n15062 & ~n15063 ) ;
  assign n15065 = ( ~n15032 & n15034 ) | ( ~n15032 & n15043 ) | ( n15034 & n15043 ) ;
  assign n15066 = ( n15032 & ~n15044 ) | ( n15032 & n15065 ) | ( ~n15044 & n15065 ) ;
  assign n15067 = ( n11351 & n15064 ) | ( n11351 & n15066 ) | ( n15064 & n15066 ) ;
  assign n15068 = n8230 & n11892 ;
  assign n15069 = n8229 & ~n9997 ;
  assign n15070 = n8226 & ~n10001 ;
  assign n15071 = n8225 & n9999 ;
  assign n15072 = n15070 | n15071 ;
  assign n15073 = ( ~n15068 & n15069 ) | ( ~n15068 & n15072 ) | ( n15069 & n15072 ) ;
  assign n15074 = ( ~x5 & n15068 ) | ( ~x5 & n15073 ) | ( n15068 & n15073 ) ;
  assign n15075 = ( n15068 & n15073 ) | ( n15068 & ~n15074 ) | ( n15073 & ~n15074 ) ;
  assign n15076 = ( x5 & n15074 ) | ( x5 & ~n15075 ) | ( n15074 & ~n15075 ) ;
  assign n15077 = n8226 & ~n10003 ;
  assign n15078 = n8225 & ~n10001 ;
  assign n15079 = n15077 | n15078 ;
  assign n15080 = n8229 & ~n9999 ;
  assign n15081 = ( n8229 & n15079 ) | ( n8229 & ~n15080 ) | ( n15079 & ~n15080 ) ;
  assign n15082 = n8230 & n11868 ;
  assign n15083 = n15081 | n15082 ;
  assign n15084 = n8228 & ~n10003 ;
  assign n15085 = x5 & n15084 ;
  assign n15086 = ( n8230 & n11804 ) | ( n8230 & n11805 ) | ( n11804 & n11805 ) ;
  assign n15087 = n8225 | n10003 ;
  assign n15088 = n8229 & ~n10001 ;
  assign n15089 = ( ~n10003 & n15087 ) | ( ~n10003 & n15088 ) | ( n15087 & n15088 ) ;
  assign n15090 = n15086 | n15089 ;
  assign n15091 = ( x5 & n15085 ) | ( x5 & n15090 ) | ( n15085 & n15090 ) ;
  assign n15092 = n15083 | n15091 ;
  assign n15093 = x5 & ~n15092 ;
  assign n15094 = ( n14661 & n15076 ) | ( n14661 & n15093 ) | ( n15076 & n15093 ) ;
  assign n15095 = n8230 & n11934 ;
  assign n15096 = n8229 & n9995 ;
  assign n15097 = n8226 & n9999 ;
  assign n15098 = n8225 & ~n9997 ;
  assign n15099 = n15097 | n15098 ;
  assign n15100 = ( ~n15095 & n15096 ) | ( ~n15095 & n15099 ) | ( n15096 & n15099 ) ;
  assign n15101 = ( ~x5 & n15095 ) | ( ~x5 & n15100 ) | ( n15095 & n15100 ) ;
  assign n15102 = ( n15095 & n15100 ) | ( n15095 & ~n15101 ) | ( n15100 & ~n15101 ) ;
  assign n15103 = ( x5 & n15101 ) | ( x5 & ~n15102 ) | ( n15101 & ~n15102 ) ;
  assign n15104 = ( n14662 & n14663 ) | ( n14662 & n14666 ) | ( n14663 & n14666 ) ;
  assign n15105 = ~n14662 & n14667 ;
  assign n15106 = ( n14662 & ~n15104 ) | ( n14662 & n15105 ) | ( ~n15104 & n15105 ) ;
  assign n15107 = ( n15094 & n15103 ) | ( n15094 & n15106 ) | ( n15103 & n15106 ) ;
  assign n15108 = n8230 & ~n11971 ;
  assign n15109 = n8229 & n9993 ;
  assign n15110 = n8226 & ~n9997 ;
  assign n15111 = n8225 & n9995 ;
  assign n15112 = n15110 | n15111 ;
  assign n15113 = ( ~n15108 & n15109 ) | ( ~n15108 & n15112 ) | ( n15109 & n15112 ) ;
  assign n15114 = ( ~x5 & n15108 ) | ( ~x5 & n15113 ) | ( n15108 & n15113 ) ;
  assign n15115 = ( n15108 & n15113 ) | ( n15108 & ~n15114 ) | ( n15113 & ~n15114 ) ;
  assign n15116 = ( x5 & n15114 ) | ( x5 & ~n15115 ) | ( n15114 & ~n15115 ) ;
  assign n15117 = ( n14660 & n14668 ) | ( n14660 & ~n14669 ) | ( n14668 & ~n14669 ) ;
  assign n15118 = n14669 & ~n15117 ;
  assign n15119 = ( n15107 & n15116 ) | ( n15107 & n15118 ) | ( n15116 & n15118 ) ;
  assign n15120 = n8230 & n12026 ;
  assign n15121 = n8229 & n9991 ;
  assign n15122 = n8226 & n9995 ;
  assign n15123 = n8225 & n9993 ;
  assign n15124 = n15122 | n15123 ;
  assign n15125 = ( ~n15120 & n15121 ) | ( ~n15120 & n15124 ) | ( n15121 & n15124 ) ;
  assign n15126 = ( ~x5 & n15120 ) | ( ~x5 & n15125 ) | ( n15120 & n15125 ) ;
  assign n15127 = ( n15120 & n15125 ) | ( n15120 & ~n15126 ) | ( n15125 & ~n15126 ) ;
  assign n15128 = ( x5 & n15126 ) | ( x5 & ~n15127 ) | ( n15126 & ~n15127 ) ;
  assign n15129 = ( n14277 & n14653 ) | ( n14277 & ~n14670 ) | ( n14653 & ~n14670 ) ;
  assign n15130 = ( n14670 & ~n14671 ) | ( n14670 & n15129 ) | ( ~n14671 & n15129 ) ;
  assign n15131 = ( n15119 & n15128 ) | ( n15119 & n15130 ) | ( n15128 & n15130 ) ;
  assign n15132 = n8230 & n12050 ;
  assign n15133 = n8229 & n9989 ;
  assign n15134 = n8226 & n9993 ;
  assign n15135 = n8225 & n9991 ;
  assign n15136 = n15134 | n15135 ;
  assign n15137 = ( ~n15132 & n15133 ) | ( ~n15132 & n15136 ) | ( n15133 & n15136 ) ;
  assign n15138 = ( ~x5 & n15132 ) | ( ~x5 & n15137 ) | ( n15132 & n15137 ) ;
  assign n15139 = ( n15132 & n15137 ) | ( n15132 & ~n15138 ) | ( n15137 & ~n15138 ) ;
  assign n15140 = ( x5 & n15138 ) | ( x5 & ~n15139 ) | ( n15138 & ~n15139 ) ;
  assign n15141 = ( ~n14671 & n14680 ) | ( ~n14671 & n14683 ) | ( n14680 & n14683 ) ;
  assign n15142 = ( n14671 & ~n14684 ) | ( n14671 & n15141 ) | ( ~n14684 & n15141 ) ;
  assign n15143 = ( n15131 & n15140 ) | ( n15131 & n15142 ) | ( n15140 & n15142 ) ;
  assign n15144 = ( ~n14684 & n14693 ) | ( ~n14684 & n14695 ) | ( n14693 & n14695 ) ;
  assign n15145 = ( n14684 & ~n14696 ) | ( n14684 & n15144 ) | ( ~n14696 & n15144 ) ;
  assign n15146 = n8230 & ~n12074 ;
  assign n15147 = n8229 & ~n9987 ;
  assign n15148 = n8226 & n9991 ;
  assign n15149 = n8225 & n9989 ;
  assign n15150 = n15148 | n15149 ;
  assign n15151 = ( ~n15146 & n15147 ) | ( ~n15146 & n15150 ) | ( n15147 & n15150 ) ;
  assign n15152 = ( ~x5 & n15146 ) | ( ~x5 & n15151 ) | ( n15146 & n15151 ) ;
  assign n15153 = ( n15146 & n15151 ) | ( n15146 & ~n15152 ) | ( n15151 & ~n15152 ) ;
  assign n15154 = ( x5 & n15152 ) | ( x5 & ~n15153 ) | ( n15152 & ~n15153 ) ;
  assign n15155 = ( n15143 & n15145 ) | ( n15143 & n15154 ) | ( n15145 & n15154 ) ;
  assign n15156 = ( ~n14696 & n14705 ) | ( ~n14696 & n14707 ) | ( n14705 & n14707 ) ;
  assign n15157 = ( n14696 & ~n14708 ) | ( n14696 & n15156 ) | ( ~n14708 & n15156 ) ;
  assign n15158 = n8230 & ~n12099 ;
  assign n15159 = n8229 & n9985 ;
  assign n15160 = n8226 & n9989 ;
  assign n15161 = n8225 & ~n9987 ;
  assign n15162 = n15160 | n15161 ;
  assign n15163 = ( ~n15158 & n15159 ) | ( ~n15158 & n15162 ) | ( n15159 & n15162 ) ;
  assign n15164 = ( ~x5 & n15158 ) | ( ~x5 & n15163 ) | ( n15158 & n15163 ) ;
  assign n15165 = ( n15158 & n15163 ) | ( n15158 & ~n15164 ) | ( n15163 & ~n15164 ) ;
  assign n15166 = ( x5 & n15164 ) | ( x5 & ~n15165 ) | ( n15164 & ~n15165 ) ;
  assign n15167 = ( n15155 & n15157 ) | ( n15155 & n15166 ) | ( n15157 & n15166 ) ;
  assign n15168 = ( ~n14708 & n14717 ) | ( ~n14708 & n14719 ) | ( n14717 & n14719 ) ;
  assign n15169 = ( n14708 & ~n14720 ) | ( n14708 & n15168 ) | ( ~n14720 & n15168 ) ;
  assign n15170 = n8230 & ~n12129 ;
  assign n15171 = n8229 & ~n9983 ;
  assign n15172 = n8226 & ~n9987 ;
  assign n15173 = n8225 & n9985 ;
  assign n15174 = n15172 | n15173 ;
  assign n15175 = ( ~n15170 & n15171 ) | ( ~n15170 & n15174 ) | ( n15171 & n15174 ) ;
  assign n15176 = ( ~x5 & n15170 ) | ( ~x5 & n15175 ) | ( n15170 & n15175 ) ;
  assign n15177 = ( n15170 & n15175 ) | ( n15170 & ~n15176 ) | ( n15175 & ~n15176 ) ;
  assign n15178 = ( x5 & n15176 ) | ( x5 & ~n15177 ) | ( n15176 & ~n15177 ) ;
  assign n15179 = ( n15167 & n15169 ) | ( n15167 & n15178 ) | ( n15169 & n15178 ) ;
  assign n15180 = n8230 & ~n11561 ;
  assign n15181 = n8229 & n9981 ;
  assign n15182 = n8226 & n9985 ;
  assign n15183 = n8225 & ~n9983 ;
  assign n15184 = n15182 | n15183 ;
  assign n15185 = ( ~n15180 & n15181 ) | ( ~n15180 & n15184 ) | ( n15181 & n15184 ) ;
  assign n15186 = ( ~x5 & n15180 ) | ( ~x5 & n15185 ) | ( n15180 & n15185 ) ;
  assign n15187 = ( n15180 & n15185 ) | ( n15180 & ~n15186 ) | ( n15185 & ~n15186 ) ;
  assign n15188 = ( x5 & n15186 ) | ( x5 & ~n15187 ) | ( n15186 & ~n15187 ) ;
  assign n15189 = ( ~n14720 & n14722 ) | ( ~n14720 & n14731 ) | ( n14722 & n14731 ) ;
  assign n15190 = ( n14720 & ~n14732 ) | ( n14720 & n15189 ) | ( ~n14732 & n15189 ) ;
  assign n15191 = ( n15179 & n15188 ) | ( n15179 & n15190 ) | ( n15188 & n15190 ) ;
  assign n15192 = n8230 & n12153 ;
  assign n15193 = n8229 & n9979 ;
  assign n15194 = n8226 & ~n9983 ;
  assign n15195 = n8225 & n9981 ;
  assign n15196 = n15194 | n15195 ;
  assign n15197 = ( ~n15192 & n15193 ) | ( ~n15192 & n15196 ) | ( n15193 & n15196 ) ;
  assign n15198 = ( ~x5 & n15192 ) | ( ~x5 & n15197 ) | ( n15192 & n15197 ) ;
  assign n15199 = ( n15192 & n15197 ) | ( n15192 & ~n15198 ) | ( n15197 & ~n15198 ) ;
  assign n15200 = ( x5 & n15198 ) | ( x5 & ~n15199 ) | ( n15198 & ~n15199 ) ;
  assign n15201 = ( ~n14732 & n14734 ) | ( ~n14732 & n14743 ) | ( n14734 & n14743 ) ;
  assign n15202 = ( n14732 & ~n14744 ) | ( n14732 & n15201 ) | ( ~n14744 & n15201 ) ;
  assign n15203 = ( n15191 & n15200 ) | ( n15191 & n15202 ) | ( n15200 & n15202 ) ;
  assign n15204 = n8230 & n12165 ;
  assign n15205 = n8229 & n9977 ;
  assign n15206 = n8226 & n9981 ;
  assign n15207 = n8225 & n9979 ;
  assign n15208 = n15206 | n15207 ;
  assign n15209 = ( ~n15204 & n15205 ) | ( ~n15204 & n15208 ) | ( n15205 & n15208 ) ;
  assign n15210 = ( ~x5 & n15204 ) | ( ~x5 & n15209 ) | ( n15204 & n15209 ) ;
  assign n15211 = ( n15204 & n15209 ) | ( n15204 & ~n15210 ) | ( n15209 & ~n15210 ) ;
  assign n15212 = ( x5 & n15210 ) | ( x5 & ~n15211 ) | ( n15210 & ~n15211 ) ;
  assign n15213 = ( ~n14744 & n14746 ) | ( ~n14744 & n14755 ) | ( n14746 & n14755 ) ;
  assign n15214 = ( n14744 & ~n14756 ) | ( n14744 & n15213 ) | ( ~n14756 & n15213 ) ;
  assign n15215 = ( n15203 & n15212 ) | ( n15203 & n15214 ) | ( n15212 & n15214 ) ;
  assign n15216 = ( ~n14756 & n14765 ) | ( ~n14756 & n14767 ) | ( n14765 & n14767 ) ;
  assign n15217 = ( n14756 & ~n14768 ) | ( n14756 & n15216 ) | ( ~n14768 & n15216 ) ;
  assign n15218 = n8230 & n11606 ;
  assign n15219 = n8229 & n9975 ;
  assign n15220 = n8226 & n9979 ;
  assign n15221 = n8225 & n9977 ;
  assign n15222 = n15220 | n15221 ;
  assign n15223 = ( ~n15218 & n15219 ) | ( ~n15218 & n15222 ) | ( n15219 & n15222 ) ;
  assign n15224 = ( ~x5 & n15218 ) | ( ~x5 & n15223 ) | ( n15218 & n15223 ) ;
  assign n15225 = ( n15218 & n15223 ) | ( n15218 & ~n15224 ) | ( n15223 & ~n15224 ) ;
  assign n15226 = ( x5 & n15224 ) | ( x5 & ~n15225 ) | ( n15224 & ~n15225 ) ;
  assign n15227 = ( n15215 & n15217 ) | ( n15215 & n15226 ) | ( n15217 & n15226 ) ;
  assign n15228 = ( ~n14768 & n14777 ) | ( ~n14768 & n14779 ) | ( n14777 & n14779 ) ;
  assign n15229 = ( n14768 & ~n14780 ) | ( n14768 & n15228 ) | ( ~n14780 & n15228 ) ;
  assign n15230 = n8230 & n11400 ;
  assign n15231 = n8229 & n9973 ;
  assign n15232 = n8226 & n9977 ;
  assign n15233 = n8225 & n9975 ;
  assign n15234 = n15232 | n15233 ;
  assign n15235 = ( ~n15230 & n15231 ) | ( ~n15230 & n15234 ) | ( n15231 & n15234 ) ;
  assign n15236 = ( ~x5 & n15230 ) | ( ~x5 & n15235 ) | ( n15230 & n15235 ) ;
  assign n15237 = ( n15230 & n15235 ) | ( n15230 & ~n15236 ) | ( n15235 & ~n15236 ) ;
  assign n15238 = ( x5 & n15236 ) | ( x5 & ~n15237 ) | ( n15236 & ~n15237 ) ;
  assign n15239 = ( n15227 & n15229 ) | ( n15227 & n15238 ) | ( n15229 & n15238 ) ;
  assign n15240 = ( ~n14780 & n14789 ) | ( ~n14780 & n14791 ) | ( n14789 & n14791 ) ;
  assign n15241 = ( n14780 & ~n14792 ) | ( n14780 & n15240 ) | ( ~n14792 & n15240 ) ;
  assign n15242 = n8230 & n11630 ;
  assign n15243 = n8229 & n9971 ;
  assign n15244 = n8226 & n9975 ;
  assign n15245 = n8225 & n9973 ;
  assign n15246 = n15244 | n15245 ;
  assign n15247 = ( ~n15242 & n15243 ) | ( ~n15242 & n15246 ) | ( n15243 & n15246 ) ;
  assign n15248 = ( ~x5 & n15242 ) | ( ~x5 & n15247 ) | ( n15242 & n15247 ) ;
  assign n15249 = ( n15242 & n15247 ) | ( n15242 & ~n15248 ) | ( n15247 & ~n15248 ) ;
  assign n15250 = ( x5 & n15248 ) | ( x5 & ~n15249 ) | ( n15248 & ~n15249 ) ;
  assign n15251 = ( n15239 & n15241 ) | ( n15239 & n15250 ) | ( n15241 & n15250 ) ;
  assign n15252 = n8230 & n11428 ;
  assign n15253 = n8229 & n9969 ;
  assign n15254 = n8226 & n9973 ;
  assign n15255 = n8225 & n9971 ;
  assign n15256 = n15254 | n15255 ;
  assign n15257 = ( ~n15252 & n15253 ) | ( ~n15252 & n15256 ) | ( n15253 & n15256 ) ;
  assign n15258 = ( ~x5 & n15252 ) | ( ~x5 & n15257 ) | ( n15252 & n15257 ) ;
  assign n15259 = ( n15252 & n15257 ) | ( n15252 & ~n15258 ) | ( n15257 & ~n15258 ) ;
  assign n15260 = ( x5 & n15258 ) | ( x5 & ~n15259 ) | ( n15258 & ~n15259 ) ;
  assign n15261 = ( ~n14792 & n14794 ) | ( ~n14792 & n14803 ) | ( n14794 & n14803 ) ;
  assign n15262 = ( n14792 & ~n14804 ) | ( n14792 & n15261 ) | ( ~n14804 & n15261 ) ;
  assign n15263 = ( n15251 & n15260 ) | ( n15251 & n15262 ) | ( n15260 & n15262 ) ;
  assign n15264 = n8230 & ~n10998 ;
  assign n15265 = n8229 & ~n9967 ;
  assign n15266 = n8226 & n9971 ;
  assign n15267 = n8225 & n9969 ;
  assign n15268 = n15266 | n15267 ;
  assign n15269 = ( ~n15264 & n15265 ) | ( ~n15264 & n15268 ) | ( n15265 & n15268 ) ;
  assign n15270 = ( ~x5 & n15264 ) | ( ~x5 & n15269 ) | ( n15264 & n15269 ) ;
  assign n15271 = ( n15264 & n15269 ) | ( n15264 & ~n15270 ) | ( n15269 & ~n15270 ) ;
  assign n15272 = ( x5 & n15270 ) | ( x5 & ~n15271 ) | ( n15270 & ~n15271 ) ;
  assign n15273 = ( ~n14804 & n14806 ) | ( ~n14804 & n14815 ) | ( n14806 & n14815 ) ;
  assign n15274 = ( n14804 & ~n14816 ) | ( n14804 & n15273 ) | ( ~n14816 & n15273 ) ;
  assign n15275 = ( n15263 & n15272 ) | ( n15263 & n15274 ) | ( n15272 & n15274 ) ;
  assign n15276 = n8230 & ~n11273 ;
  assign n15277 = n8229 & n9965 ;
  assign n15278 = n8226 & n9969 ;
  assign n15279 = n8225 & ~n9967 ;
  assign n15280 = n15278 | n15279 ;
  assign n15281 = ( ~n15276 & n15277 ) | ( ~n15276 & n15280 ) | ( n15277 & n15280 ) ;
  assign n15282 = ( ~x5 & n15276 ) | ( ~x5 & n15281 ) | ( n15276 & n15281 ) ;
  assign n15283 = ( n15276 & n15281 ) | ( n15276 & ~n15282 ) | ( n15281 & ~n15282 ) ;
  assign n15284 = ( x5 & n15282 ) | ( x5 & ~n15283 ) | ( n15282 & ~n15283 ) ;
  assign n15285 = ( ~n14816 & n14818 ) | ( ~n14816 & n14827 ) | ( n14818 & n14827 ) ;
  assign n15286 = ( n14816 & ~n14828 ) | ( n14816 & n15285 ) | ( ~n14828 & n15285 ) ;
  assign n15287 = ( n15275 & n15284 ) | ( n15275 & n15286 ) | ( n15284 & n15286 ) ;
  assign n15288 = ( ~n14828 & n14837 ) | ( ~n14828 & n14839 ) | ( n14837 & n14839 ) ;
  assign n15289 = ( n14828 & ~n14840 ) | ( n14828 & n15288 ) | ( ~n14840 & n15288 ) ;
  assign n15290 = n8230 & ~n11121 ;
  assign n15291 = n8229 & ~n9963 ;
  assign n15292 = n8226 & ~n9967 ;
  assign n15293 = n8225 & n9965 ;
  assign n15294 = n15292 | n15293 ;
  assign n15295 = ( ~n15290 & n15291 ) | ( ~n15290 & n15294 ) | ( n15291 & n15294 ) ;
  assign n15296 = ( ~x5 & n15290 ) | ( ~x5 & n15295 ) | ( n15290 & n15295 ) ;
  assign n15297 = ( n15290 & n15295 ) | ( n15290 & ~n15296 ) | ( n15295 & ~n15296 ) ;
  assign n15298 = ( x5 & n15296 ) | ( x5 & ~n15297 ) | ( n15296 & ~n15297 ) ;
  assign n15299 = ( n15287 & n15289 ) | ( n15287 & n15298 ) | ( n15289 & n15298 ) ;
  assign n15300 = ( ~n14840 & n14849 ) | ( ~n14840 & n14851 ) | ( n14849 & n14851 ) ;
  assign n15301 = ( n14840 & ~n14852 ) | ( n14840 & n15300 ) | ( ~n14852 & n15300 ) ;
  assign n15302 = n8230 & ~n10929 ;
  assign n15303 = n8229 & n9961 ;
  assign n15304 = n8226 & n9965 ;
  assign n15305 = n8225 & ~n9963 ;
  assign n15306 = n15304 | n15305 ;
  assign n15307 = ( ~n15302 & n15303 ) | ( ~n15302 & n15306 ) | ( n15303 & n15306 ) ;
  assign n15308 = ( ~x5 & n15302 ) | ( ~x5 & n15307 ) | ( n15302 & n15307 ) ;
  assign n15309 = ( n15302 & n15307 ) | ( n15302 & ~n15308 ) | ( n15307 & ~n15308 ) ;
  assign n15310 = ( x5 & n15308 ) | ( x5 & ~n15309 ) | ( n15308 & ~n15309 ) ;
  assign n15311 = ( n15299 & n15301 ) | ( n15299 & n15310 ) | ( n15301 & n15310 ) ;
  assign n15312 = ( ~n14852 & n14861 ) | ( ~n14852 & n14863 ) | ( n14861 & n14863 ) ;
  assign n15313 = ( n14852 & ~n14864 ) | ( n14852 & n15312 ) | ( ~n14864 & n15312 ) ;
  assign n15314 = n8230 & n10859 ;
  assign n15315 = n8229 & n9959 ;
  assign n15316 = n8226 & ~n9963 ;
  assign n15317 = n8225 & n9961 ;
  assign n15318 = n15316 | n15317 ;
  assign n15319 = ( ~n15314 & n15315 ) | ( ~n15314 & n15318 ) | ( n15315 & n15318 ) ;
  assign n15320 = ( ~x5 & n15314 ) | ( ~x5 & n15319 ) | ( n15314 & n15319 ) ;
  assign n15321 = ( n15314 & n15319 ) | ( n15314 & ~n15320 ) | ( n15319 & ~n15320 ) ;
  assign n15322 = ( x5 & n15320 ) | ( x5 & ~n15321 ) | ( n15320 & ~n15321 ) ;
  assign n15323 = ( n15311 & n15313 ) | ( n15311 & n15322 ) | ( n15313 & n15322 ) ;
  assign n15324 = n8230 & ~n10869 ;
  assign n15325 = n8229 & ~n9957 ;
  assign n15326 = n8226 & n9961 ;
  assign n15327 = n8225 & n9959 ;
  assign n15328 = n15326 | n15327 ;
  assign n15329 = ( ~n15324 & n15325 ) | ( ~n15324 & n15328 ) | ( n15325 & n15328 ) ;
  assign n15330 = ( ~x5 & n15324 ) | ( ~x5 & n15329 ) | ( n15324 & n15329 ) ;
  assign n15331 = ( n15324 & n15329 ) | ( n15324 & ~n15330 ) | ( n15329 & ~n15330 ) ;
  assign n15332 = ( x5 & n15330 ) | ( x5 & ~n15331 ) | ( n15330 & ~n15331 ) ;
  assign n15333 = ( ~n14864 & n14866 ) | ( ~n14864 & n14875 ) | ( n14866 & n14875 ) ;
  assign n15334 = ( n14864 & ~n14876 ) | ( n14864 & n15333 ) | ( ~n14876 & n15333 ) ;
  assign n15335 = ( n15323 & n15332 ) | ( n15323 & n15334 ) | ( n15332 & n15334 ) ;
  assign n15336 = n8230 & ~n10567 ;
  assign n15337 = n8229 & n9955 ;
  assign n15338 = n8226 & n9959 ;
  assign n15339 = n8225 & ~n9957 ;
  assign n15340 = n15338 | n15339 ;
  assign n15341 = ( ~n15336 & n15337 ) | ( ~n15336 & n15340 ) | ( n15337 & n15340 ) ;
  assign n15342 = ( ~x5 & n15336 ) | ( ~x5 & n15341 ) | ( n15336 & n15341 ) ;
  assign n15343 = ( n15336 & n15341 ) | ( n15336 & ~n15342 ) | ( n15341 & ~n15342 ) ;
  assign n15344 = ( x5 & n15342 ) | ( x5 & ~n15343 ) | ( n15342 & ~n15343 ) ;
  assign n15345 = ( ~n14876 & n14878 ) | ( ~n14876 & n14887 ) | ( n14878 & n14887 ) ;
  assign n15346 = ( n14876 & ~n14888 ) | ( n14876 & n15345 ) | ( ~n14888 & n15345 ) ;
  assign n15347 = ( n15335 & n15344 ) | ( n15335 & n15346 ) | ( n15344 & n15346 ) ;
  assign n15348 = n8230 & ~n10750 ;
  assign n15349 = n8229 & ~n9953 ;
  assign n15350 = n8226 & ~n9957 ;
  assign n15351 = n8225 & n9955 ;
  assign n15352 = n15350 | n15351 ;
  assign n15353 = ( ~n15348 & n15349 ) | ( ~n15348 & n15352 ) | ( n15349 & n15352 ) ;
  assign n15354 = ( ~x5 & n15348 ) | ( ~x5 & n15353 ) | ( n15348 & n15353 ) ;
  assign n15355 = ( n15348 & n15353 ) | ( n15348 & ~n15354 ) | ( n15353 & ~n15354 ) ;
  assign n15356 = ( x5 & n15354 ) | ( x5 & ~n15355 ) | ( n15354 & ~n15355 ) ;
  assign n15357 = ( ~n14888 & n14890 ) | ( ~n14888 & n14899 ) | ( n14890 & n14899 ) ;
  assign n15358 = ( n14888 & ~n14900 ) | ( n14888 & n15357 ) | ( ~n14900 & n15357 ) ;
  assign n15359 = ( n15347 & n15356 ) | ( n15347 & n15358 ) | ( n15356 & n15358 ) ;
  assign n15360 = ( ~n14900 & n14909 ) | ( ~n14900 & n14911 ) | ( n14909 & n14911 ) ;
  assign n15361 = ( n14900 & ~n14912 ) | ( n14900 & n15360 ) | ( ~n14912 & n15360 ) ;
  assign n15362 = n8230 & ~n10652 ;
  assign n15363 = n8229 & n9951 ;
  assign n15364 = n8226 & n9955 ;
  assign n15365 = n8225 & ~n9953 ;
  assign n15366 = n15364 | n15365 ;
  assign n15367 = ( ~n15362 & n15363 ) | ( ~n15362 & n15366 ) | ( n15363 & n15366 ) ;
  assign n15368 = ( ~x5 & n15362 ) | ( ~x5 & n15367 ) | ( n15362 & n15367 ) ;
  assign n15369 = ( n15362 & n15367 ) | ( n15362 & ~n15368 ) | ( n15367 & ~n15368 ) ;
  assign n15370 = ( x5 & n15368 ) | ( x5 & ~n15369 ) | ( n15368 & ~n15369 ) ;
  assign n15371 = ( n15359 & n15361 ) | ( n15359 & n15370 ) | ( n15361 & n15370 ) ;
  assign n15372 = ( ~n14912 & n14921 ) | ( ~n14912 & n14923 ) | ( n14921 & n14923 ) ;
  assign n15373 = ( n14912 & ~n14924 ) | ( n14912 & n15372 ) | ( ~n14924 & n15372 ) ;
  assign n15374 = n8230 & n10557 ;
  assign n15375 = n8229 & n9949 ;
  assign n15376 = n8226 & ~n9953 ;
  assign n15377 = n8225 & n9951 ;
  assign n15378 = n15376 | n15377 ;
  assign n15379 = ( ~n15374 & n15375 ) | ( ~n15374 & n15378 ) | ( n15375 & n15378 ) ;
  assign n15380 = ( ~x5 & n15374 ) | ( ~x5 & n15379 ) | ( n15374 & n15379 ) ;
  assign n15381 = ( n15374 & n15379 ) | ( n15374 & ~n15380 ) | ( n15379 & ~n15380 ) ;
  assign n15382 = ( x5 & n15380 ) | ( x5 & ~n15381 ) | ( n15380 & ~n15381 ) ;
  assign n15383 = ( n15371 & n15373 ) | ( n15371 & n15382 ) | ( n15373 & n15382 ) ;
  assign n15384 = n8230 & n10454 ;
  assign n15385 = n8229 & n9947 ;
  assign n15386 = n8226 & n9951 ;
  assign n15387 = n8225 & n9949 ;
  assign n15388 = n15386 | n15387 ;
  assign n15389 = ( ~n15384 & n15385 ) | ( ~n15384 & n15388 ) | ( n15385 & n15388 ) ;
  assign n15390 = ( ~x5 & n15384 ) | ( ~x5 & n15389 ) | ( n15384 & n15389 ) ;
  assign n15391 = ( n15384 & n15389 ) | ( n15384 & ~n15390 ) | ( n15389 & ~n15390 ) ;
  assign n15392 = ( x5 & n15390 ) | ( x5 & ~n15391 ) | ( n15390 & ~n15391 ) ;
  assign n15393 = ( ~n14924 & n14926 ) | ( ~n14924 & n14935 ) | ( n14926 & n14935 ) ;
  assign n15394 = ( ~n14935 & n14936 ) | ( ~n14935 & n15393 ) | ( n14936 & n15393 ) ;
  assign n15395 = ( n15383 & n15392 ) | ( n15383 & ~n15394 ) | ( n15392 & ~n15394 ) ;
  assign n15396 = n8230 & n10466 ;
  assign n15397 = n8229 & n9945 ;
  assign n15398 = n8226 & n9949 ;
  assign n15399 = n8225 & n9947 ;
  assign n15400 = n15398 | n15399 ;
  assign n15401 = ( ~n15396 & n15397 ) | ( ~n15396 & n15400 ) | ( n15397 & n15400 ) ;
  assign n15402 = ( ~x5 & n15396 ) | ( ~x5 & n15401 ) | ( n15396 & n15401 ) ;
  assign n15403 = ( n15396 & n15401 ) | ( n15396 & ~n15402 ) | ( n15401 & ~n15402 ) ;
  assign n15404 = ( x5 & n15402 ) | ( x5 & ~n15403 ) | ( n15402 & ~n15403 ) ;
  assign n15405 = ( ~n14936 & n14938 ) | ( ~n14936 & n14947 ) | ( n14938 & n14947 ) ;
  assign n15406 = ( ~n14947 & n14948 ) | ( ~n14947 & n15405 ) | ( n14948 & n15405 ) ;
  assign n15407 = ( n15395 & n15404 ) | ( n15395 & ~n15406 ) | ( n15404 & ~n15406 ) ;
  assign n15408 = n8230 & n10271 ;
  assign n15409 = n8229 & n9943 ;
  assign n15410 = n8226 & n9947 ;
  assign n15411 = n8225 & n9945 ;
  assign n15412 = n15410 | n15411 ;
  assign n15413 = ( ~n15408 & n15409 ) | ( ~n15408 & n15412 ) | ( n15409 & n15412 ) ;
  assign n15414 = ( ~x5 & n15408 ) | ( ~x5 & n15413 ) | ( n15408 & n15413 ) ;
  assign n15415 = ( n15408 & n15413 ) | ( n15408 & ~n15414 ) | ( n15413 & ~n15414 ) ;
  assign n15416 = ( x5 & n15414 ) | ( x5 & ~n15415 ) | ( n15414 & ~n15415 ) ;
  assign n15417 = ( ~n14948 & n14950 ) | ( ~n14948 & n14959 ) | ( n14950 & n14959 ) ;
  assign n15418 = ( n14948 & ~n14960 ) | ( n14948 & n15417 ) | ( ~n14960 & n15417 ) ;
  assign n15419 = ( n15407 & n15416 ) | ( n15407 & n15418 ) | ( n15416 & n15418 ) ;
  assign n15420 = n8230 & ~n10390 ;
  assign n15421 = n8229 & ~n9941 ;
  assign n15422 = n8226 & n9945 ;
  assign n15423 = n8225 & n9943 ;
  assign n15424 = n15422 | n15423 ;
  assign n15425 = ( ~n15420 & n15421 ) | ( ~n15420 & n15424 ) | ( n15421 & n15424 ) ;
  assign n15426 = ( ~x5 & n15420 ) | ( ~x5 & n15425 ) | ( n15420 & n15425 ) ;
  assign n15427 = ( n15420 & n15425 ) | ( n15420 & ~n15426 ) | ( n15425 & ~n15426 ) ;
  assign n15428 = ( x5 & n15426 ) | ( x5 & ~n15427 ) | ( n15426 & ~n15427 ) ;
  assign n15429 = ( ~n14960 & n14962 ) | ( ~n14960 & n14971 ) | ( n14962 & n14971 ) ;
  assign n15430 = ( ~n14971 & n14972 ) | ( ~n14971 & n15429 ) | ( n14972 & n15429 ) ;
  assign n15431 = ( n15419 & n15428 ) | ( n15419 & ~n15430 ) | ( n15428 & ~n15430 ) ;
  assign n15432 = n8230 & n10284 ;
  assign n15433 = n8229 & ~n9883 ;
  assign n15434 = n8226 & n9943 ;
  assign n15435 = n8225 & ~n9941 ;
  assign n15436 = n15434 | n15435 ;
  assign n15437 = ( ~n15432 & n15433 ) | ( ~n15432 & n15436 ) | ( n15433 & n15436 ) ;
  assign n15438 = ( ~x5 & n15432 ) | ( ~x5 & n15437 ) | ( n15432 & n15437 ) ;
  assign n15439 = ( n15432 & n15437 ) | ( n15432 & ~n15438 ) | ( n15437 & ~n15438 ) ;
  assign n15440 = ( x5 & n15438 ) | ( x5 & ~n15439 ) | ( n15438 & ~n15439 ) ;
  assign n15441 = ( ~n14972 & n14974 ) | ( ~n14972 & n14983 ) | ( n14974 & n14983 ) ;
  assign n15442 = ( ~n14983 & n14984 ) | ( ~n14983 & n15441 ) | ( n14984 & n15441 ) ;
  assign n15443 = ( n15431 & n15440 ) | ( n15431 & ~n15442 ) | ( n15440 & ~n15442 ) ;
  assign n15444 = n8230 & n10174 ;
  assign n15445 = n8229 & n9916 ;
  assign n15446 = n8225 | n9883 ;
  assign n15447 = n8226 & ~n9941 ;
  assign n15448 = ( ~n9883 & n15446 ) | ( ~n9883 & n15447 ) | ( n15446 & n15447 ) ;
  assign n15449 = ( ~n15444 & n15445 ) | ( ~n15444 & n15448 ) | ( n15445 & n15448 ) ;
  assign n15450 = ( ~x5 & n15444 ) | ( ~x5 & n15449 ) | ( n15444 & n15449 ) ;
  assign n15451 = ( n15444 & n15449 ) | ( n15444 & ~n15450 ) | ( n15449 & ~n15450 ) ;
  assign n15452 = ( x5 & n15450 ) | ( x5 & ~n15451 ) | ( n15450 & ~n15451 ) ;
  assign n15453 = ( ~n14984 & n14986 ) | ( ~n14984 & n14995 ) | ( n14986 & n14995 ) ;
  assign n15454 = ( n14984 & ~n14996 ) | ( n14984 & n15453 ) | ( ~n14996 & n15453 ) ;
  assign n15455 = ( n15443 & n15452 ) | ( n15443 & n15454 ) | ( n15452 & n15454 ) ;
  assign n15456 = n8230 & n10040 ;
  assign n15457 = n8229 & ~n9937 ;
  assign n15458 = n8226 & ~n9883 ;
  assign n15459 = n8225 & n9916 ;
  assign n15460 = n15458 | n15459 ;
  assign n15461 = ( ~n15456 & n15457 ) | ( ~n15456 & n15460 ) | ( n15457 & n15460 ) ;
  assign n15462 = ( ~x5 & n15456 ) | ( ~x5 & n15461 ) | ( n15456 & n15461 ) ;
  assign n15463 = ( n15456 & n15461 ) | ( n15456 & ~n15462 ) | ( n15461 & ~n15462 ) ;
  assign n15464 = ( x5 & n15462 ) | ( x5 & ~n15463 ) | ( n15462 & ~n15463 ) ;
  assign n15465 = ( ~n14996 & n14998 ) | ( ~n14996 & n15007 ) | ( n14998 & n15007 ) ;
  assign n15466 = ( n14996 & ~n15008 ) | ( n14996 & n15465 ) | ( ~n15008 & n15465 ) ;
  assign n15467 = ( n15455 & n15464 ) | ( n15455 & n15466 ) | ( n15464 & n15466 ) ;
  assign n15468 = n8230 & ~n10064 ;
  assign n15469 = n8229 & ~n10057 ;
  assign n15470 = n8226 & n9916 ;
  assign n15471 = n8225 & ~n9937 ;
  assign n15472 = n15470 | n15471 ;
  assign n15473 = ( ~n15468 & n15469 ) | ( ~n15468 & n15472 ) | ( n15469 & n15472 ) ;
  assign n15474 = ( ~x5 & n15468 ) | ( ~x5 & n15473 ) | ( n15468 & n15473 ) ;
  assign n15475 = ( n15468 & n15473 ) | ( n15468 & ~n15474 ) | ( n15473 & ~n15474 ) ;
  assign n15476 = ( x5 & n15474 ) | ( x5 & ~n15475 ) | ( n15474 & ~n15475 ) ;
  assign n15477 = ( ~n15008 & n15010 ) | ( ~n15008 & n15019 ) | ( n15010 & n15019 ) ;
  assign n15478 = ( n15008 & ~n15020 ) | ( n15008 & n15477 ) | ( ~n15020 & n15477 ) ;
  assign n15479 = ( n15467 & n15476 ) | ( n15467 & n15478 ) | ( n15476 & n15478 ) ;
  assign n15480 = n8230 & ~n10305 ;
  assign n15481 = n8229 & ~n10302 ;
  assign n15482 = n8226 & ~n9937 ;
  assign n15483 = n8225 & ~n10057 ;
  assign n15484 = n15482 | n15483 ;
  assign n15485 = ( ~n15480 & n15481 ) | ( ~n15480 & n15484 ) | ( n15481 & n15484 ) ;
  assign n15486 = ( ~x5 & n15480 ) | ( ~x5 & n15485 ) | ( n15480 & n15485 ) ;
  assign n15487 = ( n15480 & n15485 ) | ( n15480 & ~n15486 ) | ( n15485 & ~n15486 ) ;
  assign n15488 = ( x5 & n15486 ) | ( x5 & ~n15487 ) | ( n15486 & ~n15487 ) ;
  assign n15489 = ( ~n15020 & n15022 ) | ( ~n15020 & n15031 ) | ( n15022 & n15031 ) ;
  assign n15490 = ( n15020 & ~n15032 ) | ( n15020 & n15489 ) | ( ~n15032 & n15489 ) ;
  assign n15491 = ( n15479 & n15488 ) | ( n15479 & n15490 ) | ( n15488 & n15490 ) ;
  assign n15492 = n36 & n12026 ;
  assign n15493 = ~n8967 & n9995 ;
  assign n15494 = n9378 & n9993 ;
  assign n15495 = ( n9995 & ~n15493 ) | ( n9995 & n15494 ) | ( ~n15493 & n15494 ) ;
  assign n15496 = n35 & ~n9991 ;
  assign n15497 = ( n35 & n15495 ) | ( n35 & ~n15496 ) | ( n15495 & ~n15496 ) ;
  assign n15498 = ( ~x2 & n15492 ) | ( ~x2 & n15497 ) | ( n15492 & n15497 ) ;
  assign n15499 = ( n15492 & n15497 ) | ( n15492 & ~n15498 ) | ( n15497 & ~n15498 ) ;
  assign n15500 = ( x2 & n15498 ) | ( x2 & ~n15499 ) | ( n15498 & ~n15499 ) ;
  assign n15501 = ( n36 & n10004 ) | ( n36 & n11804 ) | ( n10004 & n11804 ) ;
  assign n15502 = n35 & n9999 ;
  assign n15503 = x1 & ~n10001 ;
  assign n15504 = ( ~x2 & n10003 ) | ( ~x2 & n15503 ) | ( n10003 & n15503 ) ;
  assign n15505 = n10003 & ~n15504 ;
  assign n15506 = ( n15501 & ~n15502 ) | ( n15501 & n15505 ) | ( ~n15502 & n15505 ) ;
  assign n15507 = ( n15084 & ~n15501 ) | ( n15084 & n15506 ) | ( ~n15501 & n15506 ) ;
  assign n15508 = n8967 & ~n10001 ;
  assign n15509 = ( x0 & n8966 ) | ( x0 & ~n9999 ) | ( n8966 & ~n9999 ) ;
  assign n15510 = ( n8966 & n15508 ) | ( n8966 & ~n15509 ) | ( n15508 & ~n15509 ) ;
  assign n15511 = n35 & n9997 ;
  assign n15512 = ( n35 & n15510 ) | ( n35 & ~n15511 ) | ( n15510 & ~n15511 ) ;
  assign n15513 = n36 & n11892 ;
  assign n15514 = n15512 | n15513 ;
  assign n15515 = ( x2 & n15507 ) | ( x2 & n15514 ) | ( n15507 & n15514 ) ;
  assign n15516 = x2 & ~n15514 ;
  assign n15517 = ( ~x2 & n15515 ) | ( ~x2 & n15516 ) | ( n15515 & n15516 ) ;
  assign n15518 = n36 & n11934 ;
  assign n15519 = n8967 & n9999 ;
  assign n15520 = ( x0 & n8966 ) | ( x0 & n9997 ) | ( n8966 & n9997 ) ;
  assign n15521 = ( n8966 & n15519 ) | ( n8966 & ~n15520 ) | ( n15519 & ~n15520 ) ;
  assign n15522 = n35 & ~n9995 ;
  assign n15523 = ( n35 & n15521 ) | ( n35 & ~n15522 ) | ( n15521 & ~n15522 ) ;
  assign n15524 = ( ~x2 & n15518 ) | ( ~x2 & n15523 ) | ( n15518 & n15523 ) ;
  assign n15525 = ( n15518 & n15523 ) | ( n15518 & ~n15524 ) | ( n15523 & ~n15524 ) ;
  assign n15526 = ( x2 & n15524 ) | ( x2 & ~n15525 ) | ( n15524 & ~n15525 ) ;
  assign n15527 = ( n15085 & n15086 ) | ( n15085 & n15089 ) | ( n15086 & n15089 ) ;
  assign n15528 = ~n15085 & n15090 ;
  assign n15529 = ( n15085 & ~n15527 ) | ( n15085 & n15528 ) | ( ~n15527 & n15528 ) ;
  assign n15530 = ( n15517 & n15526 ) | ( n15517 & n15529 ) | ( n15526 & n15529 ) ;
  assign n15531 = n36 & ~n11971 ;
  assign n15532 = n8967 & ~n9997 ;
  assign n15533 = ( x0 & n8966 ) | ( x0 & ~n9995 ) | ( n8966 & ~n9995 ) ;
  assign n15534 = ( n8966 & n15532 ) | ( n8966 & ~n15533 ) | ( n15532 & ~n15533 ) ;
  assign n15535 = n35 & ~n9993 ;
  assign n15536 = ( n35 & n15534 ) | ( n35 & ~n15535 ) | ( n15534 & ~n15535 ) ;
  assign n15537 = ( ~x2 & n15531 ) | ( ~x2 & n15536 ) | ( n15531 & n15536 ) ;
  assign n15538 = ( n15531 & n15536 ) | ( n15531 & ~n15537 ) | ( n15536 & ~n15537 ) ;
  assign n15539 = ( x2 & n15537 ) | ( x2 & ~n15538 ) | ( n15537 & ~n15538 ) ;
  assign n15540 = ~n15083 & n15091 ;
  assign n15541 = ( ~n15091 & n15092 ) | ( ~n15091 & n15540 ) | ( n15092 & n15540 ) ;
  assign n15542 = ( n15530 & n15539 ) | ( n15530 & n15541 ) | ( n15539 & n15541 ) ;
  assign n15543 = ( n14661 & n15076 ) | ( n14661 & ~n15093 ) | ( n15076 & ~n15093 ) ;
  assign n15544 = ( n15093 & ~n15094 ) | ( n15093 & n15543 ) | ( ~n15094 & n15543 ) ;
  assign n15545 = ( n15500 & n15542 ) | ( n15500 & n15544 ) | ( n15542 & n15544 ) ;
  assign n15546 = ( ~n15094 & n15103 ) | ( ~n15094 & n15106 ) | ( n15103 & n15106 ) ;
  assign n15547 = ( n15094 & ~n15107 ) | ( n15094 & n15546 ) | ( ~n15107 & n15546 ) ;
  assign n15548 = n36 & n12050 ;
  assign n15549 = n8967 & n9993 ;
  assign n15550 = ( x0 & n8966 ) | ( x0 & ~n9991 ) | ( n8966 & ~n9991 ) ;
  assign n15551 = ( n8966 & n15549 ) | ( n8966 & ~n15550 ) | ( n15549 & ~n15550 ) ;
  assign n15552 = n35 & ~n9989 ;
  assign n15553 = ( n35 & n15551 ) | ( n35 & ~n15552 ) | ( n15551 & ~n15552 ) ;
  assign n15554 = ( ~x2 & n15548 ) | ( ~x2 & n15553 ) | ( n15548 & n15553 ) ;
  assign n15555 = ( n15548 & n15553 ) | ( n15548 & ~n15554 ) | ( n15553 & ~n15554 ) ;
  assign n15556 = ( x2 & n15554 ) | ( x2 & ~n15555 ) | ( n15554 & ~n15555 ) ;
  assign n15557 = ( n15545 & n15547 ) | ( n15545 & n15556 ) | ( n15547 & n15556 ) ;
  assign n15558 = n36 & ~n12074 ;
  assign n15559 = n8967 & n9991 ;
  assign n15560 = ( x0 & n8966 ) | ( x0 & ~n9989 ) | ( n8966 & ~n9989 ) ;
  assign n15561 = ( n8966 & n15559 ) | ( n8966 & ~n15560 ) | ( n15559 & ~n15560 ) ;
  assign n15562 = n35 & n9987 ;
  assign n15563 = ( n35 & n15561 ) | ( n35 & ~n15562 ) | ( n15561 & ~n15562 ) ;
  assign n15564 = ( ~x2 & n15558 ) | ( ~x2 & n15563 ) | ( n15558 & n15563 ) ;
  assign n15565 = ( n15558 & n15563 ) | ( n15558 & ~n15564 ) | ( n15563 & ~n15564 ) ;
  assign n15566 = ( x2 & n15564 ) | ( x2 & ~n15565 ) | ( n15564 & ~n15565 ) ;
  assign n15567 = ( ~n15107 & n15116 ) | ( ~n15107 & n15118 ) | ( n15116 & n15118 ) ;
  assign n15568 = ( n15107 & ~n15119 ) | ( n15107 & n15567 ) | ( ~n15119 & n15567 ) ;
  assign n15569 = ( n15557 & n15566 ) | ( n15557 & n15568 ) | ( n15566 & n15568 ) ;
  assign n15570 = n36 & ~n12099 ;
  assign n15571 = n8967 & n9989 ;
  assign n15572 = ( x0 & n8966 ) | ( x0 & n9987 ) | ( n8966 & n9987 ) ;
  assign n15573 = ( n8966 & n15571 ) | ( n8966 & ~n15572 ) | ( n15571 & ~n15572 ) ;
  assign n15574 = n35 & ~n9985 ;
  assign n15575 = ( n35 & n15573 ) | ( n35 & ~n15574 ) | ( n15573 & ~n15574 ) ;
  assign n15576 = ( ~x2 & n15570 ) | ( ~x2 & n15575 ) | ( n15570 & n15575 ) ;
  assign n15577 = ( n15570 & n15575 ) | ( n15570 & ~n15576 ) | ( n15575 & ~n15576 ) ;
  assign n15578 = ( x2 & n15576 ) | ( x2 & ~n15577 ) | ( n15576 & ~n15577 ) ;
  assign n15579 = ( ~n15119 & n15128 ) | ( ~n15119 & n15130 ) | ( n15128 & n15130 ) ;
  assign n15580 = ( n15119 & ~n15131 ) | ( n15119 & n15579 ) | ( ~n15131 & n15579 ) ;
  assign n15581 = ( n15569 & n15578 ) | ( n15569 & n15580 ) | ( n15578 & n15580 ) ;
  assign n15582 = n36 & ~n12129 ;
  assign n15583 = n8967 & ~n9987 ;
  assign n15584 = ( x0 & n8966 ) | ( x0 & ~n9985 ) | ( n8966 & ~n9985 ) ;
  assign n15585 = ( n8966 & n15583 ) | ( n8966 & ~n15584 ) | ( n15583 & ~n15584 ) ;
  assign n15586 = n35 & n9983 ;
  assign n15587 = ( n35 & n15585 ) | ( n35 & ~n15586 ) | ( n15585 & ~n15586 ) ;
  assign n15588 = ( ~x2 & n15582 ) | ( ~x2 & n15587 ) | ( n15582 & n15587 ) ;
  assign n15589 = ( n15582 & n15587 ) | ( n15582 & ~n15588 ) | ( n15587 & ~n15588 ) ;
  assign n15590 = ( x2 & n15588 ) | ( x2 & ~n15589 ) | ( n15588 & ~n15589 ) ;
  assign n15591 = ( ~n15131 & n15140 ) | ( ~n15131 & n15142 ) | ( n15140 & n15142 ) ;
  assign n15592 = ( n15131 & ~n15143 ) | ( n15131 & n15591 ) | ( ~n15143 & n15591 ) ;
  assign n15593 = ( n15581 & n15590 ) | ( n15581 & n15592 ) | ( n15590 & n15592 ) ;
  assign n15594 = ( ~n15143 & n15145 ) | ( ~n15143 & n15154 ) | ( n15145 & n15154 ) ;
  assign n15595 = ( n15143 & ~n15155 ) | ( n15143 & n15594 ) | ( ~n15155 & n15594 ) ;
  assign n15596 = n36 & ~n11561 ;
  assign n15597 = n8967 & n9985 ;
  assign n15598 = ( x0 & n8966 ) | ( x0 & n9983 ) | ( n8966 & n9983 ) ;
  assign n15599 = ( n8966 & n15597 ) | ( n8966 & ~n15598 ) | ( n15597 & ~n15598 ) ;
  assign n15600 = n35 & ~n9981 ;
  assign n15601 = ( n35 & n15599 ) | ( n35 & ~n15600 ) | ( n15599 & ~n15600 ) ;
  assign n15602 = ( ~x2 & n15596 ) | ( ~x2 & n15601 ) | ( n15596 & n15601 ) ;
  assign n15603 = ( n15596 & n15601 ) | ( n15596 & ~n15602 ) | ( n15601 & ~n15602 ) ;
  assign n15604 = ( x2 & n15602 ) | ( x2 & ~n15603 ) | ( n15602 & ~n15603 ) ;
  assign n15605 = ( n15593 & n15595 ) | ( n15593 & n15604 ) | ( n15595 & n15604 ) ;
  assign n15606 = ( ~n15155 & n15157 ) | ( ~n15155 & n15166 ) | ( n15157 & n15166 ) ;
  assign n15607 = ( n15155 & ~n15167 ) | ( n15155 & n15606 ) | ( ~n15167 & n15606 ) ;
  assign n15608 = n36 & n12153 ;
  assign n15609 = n8967 & ~n9983 ;
  assign n15610 = ( x0 & n8966 ) | ( x0 & ~n9981 ) | ( n8966 & ~n9981 ) ;
  assign n15611 = ( n8966 & n15609 ) | ( n8966 & ~n15610 ) | ( n15609 & ~n15610 ) ;
  assign n15612 = n35 & ~n9979 ;
  assign n15613 = ( n35 & n15611 ) | ( n35 & ~n15612 ) | ( n15611 & ~n15612 ) ;
  assign n15614 = ( ~x2 & n15608 ) | ( ~x2 & n15613 ) | ( n15608 & n15613 ) ;
  assign n15615 = ( n15608 & n15613 ) | ( n15608 & ~n15614 ) | ( n15613 & ~n15614 ) ;
  assign n15616 = ( x2 & n15614 ) | ( x2 & ~n15615 ) | ( n15614 & ~n15615 ) ;
  assign n15617 = ( n15605 & n15607 ) | ( n15605 & n15616 ) | ( n15607 & n15616 ) ;
  assign n15618 = ( ~n15167 & n15169 ) | ( ~n15167 & n15178 ) | ( n15169 & n15178 ) ;
  assign n15619 = ( n15167 & ~n15179 ) | ( n15167 & n15618 ) | ( ~n15179 & n15618 ) ;
  assign n15620 = n36 & n12165 ;
  assign n15621 = n8967 & n9981 ;
  assign n15622 = ( x0 & n8966 ) | ( x0 & ~n9979 ) | ( n8966 & ~n9979 ) ;
  assign n15623 = ( n8966 & n15621 ) | ( n8966 & ~n15622 ) | ( n15621 & ~n15622 ) ;
  assign n15624 = n35 & ~n9977 ;
  assign n15625 = ( n35 & n15623 ) | ( n35 & ~n15624 ) | ( n15623 & ~n15624 ) ;
  assign n15626 = ( ~x2 & n15620 ) | ( ~x2 & n15625 ) | ( n15620 & n15625 ) ;
  assign n15627 = ( n15620 & n15625 ) | ( n15620 & ~n15626 ) | ( n15625 & ~n15626 ) ;
  assign n15628 = ( x2 & n15626 ) | ( x2 & ~n15627 ) | ( n15626 & ~n15627 ) ;
  assign n15629 = ( n15617 & n15619 ) | ( n15617 & n15628 ) | ( n15619 & n15628 ) ;
  assign n15630 = n36 & n11606 ;
  assign n15631 = n8967 & n9979 ;
  assign n15632 = ( x0 & n8966 ) | ( x0 & ~n9977 ) | ( n8966 & ~n9977 ) ;
  assign n15633 = ( n8966 & n15631 ) | ( n8966 & ~n15632 ) | ( n15631 & ~n15632 ) ;
  assign n15634 = n35 & ~n9975 ;
  assign n15635 = ( n35 & n15633 ) | ( n35 & ~n15634 ) | ( n15633 & ~n15634 ) ;
  assign n15636 = ( ~x2 & n15630 ) | ( ~x2 & n15635 ) | ( n15630 & n15635 ) ;
  assign n15637 = ( n15630 & n15635 ) | ( n15630 & ~n15636 ) | ( n15635 & ~n15636 ) ;
  assign n15638 = ( x2 & n15636 ) | ( x2 & ~n15637 ) | ( n15636 & ~n15637 ) ;
  assign n15639 = ( ~n15179 & n15188 ) | ( ~n15179 & n15190 ) | ( n15188 & n15190 ) ;
  assign n15640 = ( n15179 & ~n15191 ) | ( n15179 & n15639 ) | ( ~n15191 & n15639 ) ;
  assign n15641 = ( n15629 & n15638 ) | ( n15629 & n15640 ) | ( n15638 & n15640 ) ;
  assign n15642 = n36 & n11400 ;
  assign n15643 = n8967 & n9977 ;
  assign n15644 = ( x0 & n8966 ) | ( x0 & ~n9975 ) | ( n8966 & ~n9975 ) ;
  assign n15645 = ( n8966 & n15643 ) | ( n8966 & ~n15644 ) | ( n15643 & ~n15644 ) ;
  assign n15646 = n35 & ~n9973 ;
  assign n15647 = ( n35 & n15645 ) | ( n35 & ~n15646 ) | ( n15645 & ~n15646 ) ;
  assign n15648 = ( ~x2 & n15642 ) | ( ~x2 & n15647 ) | ( n15642 & n15647 ) ;
  assign n15649 = ( n15642 & n15647 ) | ( n15642 & ~n15648 ) | ( n15647 & ~n15648 ) ;
  assign n15650 = ( x2 & n15648 ) | ( x2 & ~n15649 ) | ( n15648 & ~n15649 ) ;
  assign n15651 = ( ~n15191 & n15200 ) | ( ~n15191 & n15202 ) | ( n15200 & n15202 ) ;
  assign n15652 = ( n15191 & ~n15203 ) | ( n15191 & n15651 ) | ( ~n15203 & n15651 ) ;
  assign n15653 = ( n15641 & n15650 ) | ( n15641 & n15652 ) | ( n15650 & n15652 ) ;
  assign n15654 = n36 & n11630 ;
  assign n15655 = n8967 & n9975 ;
  assign n15656 = ( x0 & n8966 ) | ( x0 & ~n9973 ) | ( n8966 & ~n9973 ) ;
  assign n15657 = ( n8966 & n15655 ) | ( n8966 & ~n15656 ) | ( n15655 & ~n15656 ) ;
  assign n15658 = n35 & ~n9971 ;
  assign n15659 = ( n35 & n15657 ) | ( n35 & ~n15658 ) | ( n15657 & ~n15658 ) ;
  assign n15660 = ( ~x2 & n15654 ) | ( ~x2 & n15659 ) | ( n15654 & n15659 ) ;
  assign n15661 = ( n15654 & n15659 ) | ( n15654 & ~n15660 ) | ( n15659 & ~n15660 ) ;
  assign n15662 = ( x2 & n15660 ) | ( x2 & ~n15661 ) | ( n15660 & ~n15661 ) ;
  assign n15663 = ( ~n15203 & n15212 ) | ( ~n15203 & n15214 ) | ( n15212 & n15214 ) ;
  assign n15664 = ( n15203 & ~n15215 ) | ( n15203 & n15663 ) | ( ~n15215 & n15663 ) ;
  assign n15665 = ( n15653 & n15662 ) | ( n15653 & n15664 ) | ( n15662 & n15664 ) ;
  assign n15666 = ( ~n15215 & n15217 ) | ( ~n15215 & n15226 ) | ( n15217 & n15226 ) ;
  assign n15667 = ( n15215 & ~n15227 ) | ( n15215 & n15666 ) | ( ~n15227 & n15666 ) ;
  assign n15668 = n36 & n11428 ;
  assign n15669 = n8967 & n9973 ;
  assign n15670 = ( x0 & n8966 ) | ( x0 & ~n9971 ) | ( n8966 & ~n9971 ) ;
  assign n15671 = ( n8966 & n15669 ) | ( n8966 & ~n15670 ) | ( n15669 & ~n15670 ) ;
  assign n15672 = n35 & ~n9969 ;
  assign n15673 = ( n35 & n15671 ) | ( n35 & ~n15672 ) | ( n15671 & ~n15672 ) ;
  assign n15674 = ( ~x2 & n15668 ) | ( ~x2 & n15673 ) | ( n15668 & n15673 ) ;
  assign n15675 = ( n15668 & n15673 ) | ( n15668 & ~n15674 ) | ( n15673 & ~n15674 ) ;
  assign n15676 = ( x2 & n15674 ) | ( x2 & ~n15675 ) | ( n15674 & ~n15675 ) ;
  assign n15677 = ( n15665 & n15667 ) | ( n15665 & n15676 ) | ( n15667 & n15676 ) ;
  assign n15678 = ( ~n15227 & n15229 ) | ( ~n15227 & n15238 ) | ( n15229 & n15238 ) ;
  assign n15679 = ( n15227 & ~n15239 ) | ( n15227 & n15678 ) | ( ~n15239 & n15678 ) ;
  assign n15680 = n36 & ~n10998 ;
  assign n15681 = n8967 & n9971 ;
  assign n15682 = ( x0 & n8966 ) | ( x0 & ~n9969 ) | ( n8966 & ~n9969 ) ;
  assign n15683 = ( n8966 & n15681 ) | ( n8966 & ~n15682 ) | ( n15681 & ~n15682 ) ;
  assign n15684 = n35 & n9967 ;
  assign n15685 = ( n35 & n15683 ) | ( n35 & ~n15684 ) | ( n15683 & ~n15684 ) ;
  assign n15686 = ( ~x2 & n15680 ) | ( ~x2 & n15685 ) | ( n15680 & n15685 ) ;
  assign n15687 = ( n15680 & n15685 ) | ( n15680 & ~n15686 ) | ( n15685 & ~n15686 ) ;
  assign n15688 = ( x2 & n15686 ) | ( x2 & ~n15687 ) | ( n15686 & ~n15687 ) ;
  assign n15689 = ( n15677 & n15679 ) | ( n15677 & n15688 ) | ( n15679 & n15688 ) ;
  assign n15690 = ( ~n15239 & n15241 ) | ( ~n15239 & n15250 ) | ( n15241 & n15250 ) ;
  assign n15691 = ( n15239 & ~n15251 ) | ( n15239 & n15690 ) | ( ~n15251 & n15690 ) ;
  assign n15692 = n36 & ~n11273 ;
  assign n15693 = n8967 & n9969 ;
  assign n15694 = ( x0 & n8966 ) | ( x0 & n9967 ) | ( n8966 & n9967 ) ;
  assign n15695 = ( n8966 & n15693 ) | ( n8966 & ~n15694 ) | ( n15693 & ~n15694 ) ;
  assign n15696 = n35 & ~n9965 ;
  assign n15697 = ( n35 & n15695 ) | ( n35 & ~n15696 ) | ( n15695 & ~n15696 ) ;
  assign n15698 = ( ~x2 & n15692 ) | ( ~x2 & n15697 ) | ( n15692 & n15697 ) ;
  assign n15699 = ( n15692 & n15697 ) | ( n15692 & ~n15698 ) | ( n15697 & ~n15698 ) ;
  assign n15700 = ( x2 & n15698 ) | ( x2 & ~n15699 ) | ( n15698 & ~n15699 ) ;
  assign n15701 = ( n15689 & n15691 ) | ( n15689 & n15700 ) | ( n15691 & n15700 ) ;
  assign n15702 = n36 & ~n11121 ;
  assign n15703 = n8967 & ~n9967 ;
  assign n15704 = ( x0 & n8966 ) | ( x0 & ~n9965 ) | ( n8966 & ~n9965 ) ;
  assign n15705 = ( n8966 & n15703 ) | ( n8966 & ~n15704 ) | ( n15703 & ~n15704 ) ;
  assign n15706 = n35 & n9963 ;
  assign n15707 = ( n35 & n15705 ) | ( n35 & ~n15706 ) | ( n15705 & ~n15706 ) ;
  assign n15708 = ( ~x2 & n15702 ) | ( ~x2 & n15707 ) | ( n15702 & n15707 ) ;
  assign n15709 = ( n15702 & n15707 ) | ( n15702 & ~n15708 ) | ( n15707 & ~n15708 ) ;
  assign n15710 = ( x2 & n15708 ) | ( x2 & ~n15709 ) | ( n15708 & ~n15709 ) ;
  assign n15711 = ( ~n15251 & n15260 ) | ( ~n15251 & n15262 ) | ( n15260 & n15262 ) ;
  assign n15712 = ( n15251 & ~n15263 ) | ( n15251 & n15711 ) | ( ~n15263 & n15711 ) ;
  assign n15713 = ( n15701 & n15710 ) | ( n15701 & n15712 ) | ( n15710 & n15712 ) ;
  assign n15714 = n36 & ~n10929 ;
  assign n15715 = n8967 & n9965 ;
  assign n15716 = ( x0 & n8966 ) | ( x0 & n9963 ) | ( n8966 & n9963 ) ;
  assign n15717 = ( n8966 & n15715 ) | ( n8966 & ~n15716 ) | ( n15715 & ~n15716 ) ;
  assign n15718 = n35 & ~n9961 ;
  assign n15719 = ( n35 & n15717 ) | ( n35 & ~n15718 ) | ( n15717 & ~n15718 ) ;
  assign n15720 = ( ~x2 & n15714 ) | ( ~x2 & n15719 ) | ( n15714 & n15719 ) ;
  assign n15721 = ( n15714 & n15719 ) | ( n15714 & ~n15720 ) | ( n15719 & ~n15720 ) ;
  assign n15722 = ( x2 & n15720 ) | ( x2 & ~n15721 ) | ( n15720 & ~n15721 ) ;
  assign n15723 = ( ~n15263 & n15272 ) | ( ~n15263 & n15274 ) | ( n15272 & n15274 ) ;
  assign n15724 = ( n15263 & ~n15275 ) | ( n15263 & n15723 ) | ( ~n15275 & n15723 ) ;
  assign n15725 = ( n15713 & n15722 ) | ( n15713 & n15724 ) | ( n15722 & n15724 ) ;
  assign n15726 = n36 & n10859 ;
  assign n15727 = n8967 & ~n9963 ;
  assign n15728 = ( x0 & n8966 ) | ( x0 & ~n9961 ) | ( n8966 & ~n9961 ) ;
  assign n15729 = ( n8966 & n15727 ) | ( n8966 & ~n15728 ) | ( n15727 & ~n15728 ) ;
  assign n15730 = n35 & ~n9959 ;
  assign n15731 = ( n35 & n15729 ) | ( n35 & ~n15730 ) | ( n15729 & ~n15730 ) ;
  assign n15732 = ( ~x2 & n15726 ) | ( ~x2 & n15731 ) | ( n15726 & n15731 ) ;
  assign n15733 = ( n15726 & n15731 ) | ( n15726 & ~n15732 ) | ( n15731 & ~n15732 ) ;
  assign n15734 = ( x2 & n15732 ) | ( x2 & ~n15733 ) | ( n15732 & ~n15733 ) ;
  assign n15735 = ( ~n15275 & n15284 ) | ( ~n15275 & n15286 ) | ( n15284 & n15286 ) ;
  assign n15736 = ( n15275 & ~n15287 ) | ( n15275 & n15735 ) | ( ~n15287 & n15735 ) ;
  assign n15737 = ( n15725 & n15734 ) | ( n15725 & n15736 ) | ( n15734 & n15736 ) ;
  assign n15738 = ( ~n15287 & n15289 ) | ( ~n15287 & n15298 ) | ( n15289 & n15298 ) ;
  assign n15739 = ( n15287 & ~n15299 ) | ( n15287 & n15738 ) | ( ~n15299 & n15738 ) ;
  assign n15740 = n36 & ~n10869 ;
  assign n15741 = n8967 & n9961 ;
  assign n15742 = ( x0 & n8966 ) | ( x0 & ~n9959 ) | ( n8966 & ~n9959 ) ;
  assign n15743 = ( n8966 & n15741 ) | ( n8966 & ~n15742 ) | ( n15741 & ~n15742 ) ;
  assign n15744 = n35 & n9957 ;
  assign n15745 = ( n35 & n15743 ) | ( n35 & ~n15744 ) | ( n15743 & ~n15744 ) ;
  assign n15746 = ( ~x2 & n15740 ) | ( ~x2 & n15745 ) | ( n15740 & n15745 ) ;
  assign n15747 = ( n15740 & n15745 ) | ( n15740 & ~n15746 ) | ( n15745 & ~n15746 ) ;
  assign n15748 = ( x2 & n15746 ) | ( x2 & ~n15747 ) | ( n15746 & ~n15747 ) ;
  assign n15749 = ( n15737 & n15739 ) | ( n15737 & n15748 ) | ( n15739 & n15748 ) ;
  assign n15750 = ( ~n15299 & n15301 ) | ( ~n15299 & n15310 ) | ( n15301 & n15310 ) ;
  assign n15751 = ( n15299 & ~n15311 ) | ( n15299 & n15750 ) | ( ~n15311 & n15750 ) ;
  assign n15752 = n36 & ~n10567 ;
  assign n15753 = n8967 & n9959 ;
  assign n15754 = ( x0 & n8966 ) | ( x0 & n9957 ) | ( n8966 & n9957 ) ;
  assign n15755 = ( n8966 & n15753 ) | ( n8966 & ~n15754 ) | ( n15753 & ~n15754 ) ;
  assign n15756 = n35 & ~n9955 ;
  assign n15757 = ( n35 & n15755 ) | ( n35 & ~n15756 ) | ( n15755 & ~n15756 ) ;
  assign n15758 = ( ~x2 & n15752 ) | ( ~x2 & n15757 ) | ( n15752 & n15757 ) ;
  assign n15759 = ( n15752 & n15757 ) | ( n15752 & ~n15758 ) | ( n15757 & ~n15758 ) ;
  assign n15760 = ( x2 & n15758 ) | ( x2 & ~n15759 ) | ( n15758 & ~n15759 ) ;
  assign n15761 = ( n15749 & n15751 ) | ( n15749 & n15760 ) | ( n15751 & n15760 ) ;
  assign n15762 = ( ~n15311 & n15313 ) | ( ~n15311 & n15322 ) | ( n15313 & n15322 ) ;
  assign n15763 = ( n15311 & ~n15323 ) | ( n15311 & n15762 ) | ( ~n15323 & n15762 ) ;
  assign n15764 = n36 & ~n10750 ;
  assign n15765 = n8967 & ~n9957 ;
  assign n15766 = ( x0 & n8966 ) | ( x0 & ~n9955 ) | ( n8966 & ~n9955 ) ;
  assign n15767 = ( n8966 & n15765 ) | ( n8966 & ~n15766 ) | ( n15765 & ~n15766 ) ;
  assign n15768 = n35 & n9953 ;
  assign n15769 = ( n35 & n15767 ) | ( n35 & ~n15768 ) | ( n15767 & ~n15768 ) ;
  assign n15770 = ( ~x2 & n15764 ) | ( ~x2 & n15769 ) | ( n15764 & n15769 ) ;
  assign n15771 = ( n15764 & n15769 ) | ( n15764 & ~n15770 ) | ( n15769 & ~n15770 ) ;
  assign n15772 = ( x2 & n15770 ) | ( x2 & ~n15771 ) | ( n15770 & ~n15771 ) ;
  assign n15773 = ( n15761 & n15763 ) | ( n15761 & n15772 ) | ( n15763 & n15772 ) ;
  assign n15774 = n36 & ~n10652 ;
  assign n15775 = n8967 & n9955 ;
  assign n15776 = ( x0 & n8966 ) | ( x0 & n9953 ) | ( n8966 & n9953 ) ;
  assign n15777 = ( n8966 & n15775 ) | ( n8966 & ~n15776 ) | ( n15775 & ~n15776 ) ;
  assign n15778 = n35 & ~n9951 ;
  assign n15779 = ( n35 & n15777 ) | ( n35 & ~n15778 ) | ( n15777 & ~n15778 ) ;
  assign n15780 = ( ~x2 & n15774 ) | ( ~x2 & n15779 ) | ( n15774 & n15779 ) ;
  assign n15781 = ( n15774 & n15779 ) | ( n15774 & ~n15780 ) | ( n15779 & ~n15780 ) ;
  assign n15782 = ( x2 & n15780 ) | ( x2 & ~n15781 ) | ( n15780 & ~n15781 ) ;
  assign n15783 = ( ~n15323 & n15332 ) | ( ~n15323 & n15334 ) | ( n15332 & n15334 ) ;
  assign n15784 = ( n15323 & ~n15335 ) | ( n15323 & n15783 ) | ( ~n15335 & n15783 ) ;
  assign n15785 = ( n15773 & n15782 ) | ( n15773 & n15784 ) | ( n15782 & n15784 ) ;
  assign n15786 = n36 & n10557 ;
  assign n15787 = n8967 & ~n9953 ;
  assign n15788 = ( x0 & n8966 ) | ( x0 & ~n9951 ) | ( n8966 & ~n9951 ) ;
  assign n15789 = ( n8966 & n15787 ) | ( n8966 & ~n15788 ) | ( n15787 & ~n15788 ) ;
  assign n15790 = n35 & ~n9949 ;
  assign n15791 = ( n35 & n15789 ) | ( n35 & ~n15790 ) | ( n15789 & ~n15790 ) ;
  assign n15792 = ( ~x2 & n15786 ) | ( ~x2 & n15791 ) | ( n15786 & n15791 ) ;
  assign n15793 = ( n15786 & n15791 ) | ( n15786 & ~n15792 ) | ( n15791 & ~n15792 ) ;
  assign n15794 = ( x2 & n15792 ) | ( x2 & ~n15793 ) | ( n15792 & ~n15793 ) ;
  assign n15795 = ( ~n15335 & n15344 ) | ( ~n15335 & n15346 ) | ( n15344 & n15346 ) ;
  assign n15796 = ( n15335 & ~n15347 ) | ( n15335 & n15795 ) | ( ~n15347 & n15795 ) ;
  assign n15797 = ( n15785 & n15794 ) | ( n15785 & n15796 ) | ( n15794 & n15796 ) ;
  assign n15798 = n36 & n10454 ;
  assign n15799 = n8967 & n9951 ;
  assign n15800 = ( x0 & n8966 ) | ( x0 & ~n9949 ) | ( n8966 & ~n9949 ) ;
  assign n15801 = ( n8966 & n15799 ) | ( n8966 & ~n15800 ) | ( n15799 & ~n15800 ) ;
  assign n15802 = n35 & ~n9947 ;
  assign n15803 = ( n35 & n15801 ) | ( n35 & ~n15802 ) | ( n15801 & ~n15802 ) ;
  assign n15804 = ( ~x2 & n15798 ) | ( ~x2 & n15803 ) | ( n15798 & n15803 ) ;
  assign n15805 = ( n15798 & n15803 ) | ( n15798 & ~n15804 ) | ( n15803 & ~n15804 ) ;
  assign n15806 = ( x2 & n15804 ) | ( x2 & ~n15805 ) | ( n15804 & ~n15805 ) ;
  assign n15807 = ( ~n15347 & n15356 ) | ( ~n15347 & n15358 ) | ( n15356 & n15358 ) ;
  assign n15808 = ( n15347 & ~n15359 ) | ( n15347 & n15807 ) | ( ~n15359 & n15807 ) ;
  assign n15809 = ( n15797 & n15806 ) | ( n15797 & n15808 ) | ( n15806 & n15808 ) ;
  assign n15810 = ( ~n15359 & n15361 ) | ( ~n15359 & n15370 ) | ( n15361 & n15370 ) ;
  assign n15811 = ( n15359 & ~n15371 ) | ( n15359 & n15810 ) | ( ~n15371 & n15810 ) ;
  assign n15812 = n36 & n10466 ;
  assign n15813 = n8967 & n9949 ;
  assign n15814 = ( x0 & n8966 ) | ( x0 & ~n9947 ) | ( n8966 & ~n9947 ) ;
  assign n15815 = ( n8966 & n15813 ) | ( n8966 & ~n15814 ) | ( n15813 & ~n15814 ) ;
  assign n15816 = n35 & ~n9945 ;
  assign n15817 = ( n35 & n15815 ) | ( n35 & ~n15816 ) | ( n15815 & ~n15816 ) ;
  assign n15818 = ( ~x2 & n15812 ) | ( ~x2 & n15817 ) | ( n15812 & n15817 ) ;
  assign n15819 = ( n15812 & n15817 ) | ( n15812 & ~n15818 ) | ( n15817 & ~n15818 ) ;
  assign n15820 = ( x2 & n15818 ) | ( x2 & ~n15819 ) | ( n15818 & ~n15819 ) ;
  assign n15821 = ( n15809 & n15811 ) | ( n15809 & n15820 ) | ( n15811 & n15820 ) ;
  assign n15822 = ( ~n15371 & n15373 ) | ( ~n15371 & n15382 ) | ( n15373 & n15382 ) ;
  assign n15823 = ( n15371 & ~n15383 ) | ( n15371 & n15822 ) | ( ~n15383 & n15822 ) ;
  assign n15824 = n36 & n10271 ;
  assign n15825 = n8967 & n9947 ;
  assign n15826 = ( x0 & n8966 ) | ( x0 & ~n9945 ) | ( n8966 & ~n9945 ) ;
  assign n15827 = ( n8966 & n15825 ) | ( n8966 & ~n15826 ) | ( n15825 & ~n15826 ) ;
  assign n15828 = n35 & ~n9943 ;
  assign n15829 = ( n35 & n15827 ) | ( n35 & ~n15828 ) | ( n15827 & ~n15828 ) ;
  assign n15830 = ( ~x2 & n15824 ) | ( ~x2 & n15829 ) | ( n15824 & n15829 ) ;
  assign n15831 = ( n15824 & n15829 ) | ( n15824 & ~n15830 ) | ( n15829 & ~n15830 ) ;
  assign n15832 = ( x2 & n15830 ) | ( x2 & ~n15831 ) | ( n15830 & ~n15831 ) ;
  assign n15833 = ( n15821 & n15823 ) | ( n15821 & n15832 ) | ( n15823 & n15832 ) ;
  assign n15834 = ( n15383 & ~n15392 ) | ( n15383 & n15394 ) | ( ~n15392 & n15394 ) ;
  assign n15835 = ( ~n15383 & n15395 ) | ( ~n15383 & n15834 ) | ( n15395 & n15834 ) ;
  assign n15836 = n36 & ~n10390 ;
  assign n15837 = n8967 & n9945 ;
  assign n15838 = ( x0 & n8966 ) | ( x0 & ~n9943 ) | ( n8966 & ~n9943 ) ;
  assign n15839 = ( n8966 & n15837 ) | ( n8966 & ~n15838 ) | ( n15837 & ~n15838 ) ;
  assign n15840 = n35 & n9941 ;
  assign n15841 = ( n35 & n15839 ) | ( n35 & ~n15840 ) | ( n15839 & ~n15840 ) ;
  assign n15842 = ( ~x2 & n15836 ) | ( ~x2 & n15841 ) | ( n15836 & n15841 ) ;
  assign n15843 = ( n15836 & n15841 ) | ( n15836 & ~n15842 ) | ( n15841 & ~n15842 ) ;
  assign n15844 = ( x2 & n15842 ) | ( x2 & ~n15843 ) | ( n15842 & ~n15843 ) ;
  assign n15845 = ( n15833 & ~n15835 ) | ( n15833 & n15844 ) | ( ~n15835 & n15844 ) ;
  assign n15846 = ( n15395 & ~n15404 ) | ( n15395 & n15406 ) | ( ~n15404 & n15406 ) ;
  assign n15847 = ( ~n15395 & n15407 ) | ( ~n15395 & n15846 ) | ( n15407 & n15846 ) ;
  assign n15848 = n36 & n10284 ;
  assign n15849 = n8967 & n9943 ;
  assign n15850 = ( x0 & n8966 ) | ( x0 & n9941 ) | ( n8966 & n9941 ) ;
  assign n15851 = ( n8966 & n15849 ) | ( n8966 & ~n15850 ) | ( n15849 & ~n15850 ) ;
  assign n15852 = n35 & n9883 ;
  assign n15853 = ( n35 & n15851 ) | ( n35 & ~n15852 ) | ( n15851 & ~n15852 ) ;
  assign n15854 = ( ~x2 & n15848 ) | ( ~x2 & n15853 ) | ( n15848 & n15853 ) ;
  assign n15855 = ( n15848 & n15853 ) | ( n15848 & ~n15854 ) | ( n15853 & ~n15854 ) ;
  assign n15856 = ( x2 & n15854 ) | ( x2 & ~n15855 ) | ( n15854 & ~n15855 ) ;
  assign n15857 = ( n15845 & ~n15847 ) | ( n15845 & n15856 ) | ( ~n15847 & n15856 ) ;
  assign n15858 = ( ~n15407 & n15416 ) | ( ~n15407 & n15418 ) | ( n15416 & n15418 ) ;
  assign n15859 = ( n15407 & ~n15419 ) | ( n15407 & n15858 ) | ( ~n15419 & n15858 ) ;
  assign n15860 = n36 & n10174 ;
  assign n15861 = n8967 & ~n9941 ;
  assign n15862 = ( x0 & n8966 ) | ( x0 & n9883 ) | ( n8966 & n9883 ) ;
  assign n15863 = ( n8966 & n15861 ) | ( n8966 & ~n15862 ) | ( n15861 & ~n15862 ) ;
  assign n15864 = n35 & ~n9916 ;
  assign n15865 = ( n35 & n15863 ) | ( n35 & ~n15864 ) | ( n15863 & ~n15864 ) ;
  assign n15866 = ( ~x2 & n15860 ) | ( ~x2 & n15865 ) | ( n15860 & n15865 ) ;
  assign n15867 = ( n15860 & n15865 ) | ( n15860 & ~n15866 ) | ( n15865 & ~n15866 ) ;
  assign n15868 = ( x2 & n15866 ) | ( x2 & ~n15867 ) | ( n15866 & ~n15867 ) ;
  assign n15869 = ( n15857 & n15859 ) | ( n15857 & n15868 ) | ( n15859 & n15868 ) ;
  assign n15870 = ( n15419 & ~n15428 ) | ( n15419 & n15430 ) | ( ~n15428 & n15430 ) ;
  assign n15871 = ( ~n15419 & n15431 ) | ( ~n15419 & n15870 ) | ( n15431 & n15870 ) ;
  assign n15872 = n36 & n10040 ;
  assign n15873 = n8967 & ~n9883 ;
  assign n15874 = ( x0 & n8966 ) | ( x0 & ~n9916 ) | ( n8966 & ~n9916 ) ;
  assign n15875 = ( n8966 & n15873 ) | ( n8966 & ~n15874 ) | ( n15873 & ~n15874 ) ;
  assign n15876 = n35 & n9937 ;
  assign n15877 = ( n35 & n15875 ) | ( n35 & ~n15876 ) | ( n15875 & ~n15876 ) ;
  assign n15878 = ( ~x2 & n15872 ) | ( ~x2 & n15877 ) | ( n15872 & n15877 ) ;
  assign n15879 = ( n15872 & n15877 ) | ( n15872 & ~n15878 ) | ( n15877 & ~n15878 ) ;
  assign n15880 = ( x2 & n15878 ) | ( x2 & ~n15879 ) | ( n15878 & ~n15879 ) ;
  assign n15881 = ( n15869 & ~n15871 ) | ( n15869 & n15880 ) | ( ~n15871 & n15880 ) ;
  assign n15882 = ( n15431 & ~n15440 ) | ( n15431 & n15442 ) | ( ~n15440 & n15442 ) ;
  assign n15883 = ( ~n15431 & n15443 ) | ( ~n15431 & n15882 ) | ( n15443 & n15882 ) ;
  assign n15884 = n36 & ~n10064 ;
  assign n15885 = n8967 & n9916 ;
  assign n15886 = ( x0 & n8966 ) | ( x0 & n9937 ) | ( n8966 & n9937 ) ;
  assign n15887 = ( n8966 & n15885 ) | ( n8966 & ~n15886 ) | ( n15885 & ~n15886 ) ;
  assign n15888 = n35 & n10057 ;
  assign n15889 = ( n35 & n15887 ) | ( n35 & ~n15888 ) | ( n15887 & ~n15888 ) ;
  assign n15890 = ( ~x2 & n15884 ) | ( ~x2 & n15889 ) | ( n15884 & n15889 ) ;
  assign n15891 = ( n15884 & n15889 ) | ( n15884 & ~n15890 ) | ( n15889 & ~n15890 ) ;
  assign n15892 = ( x2 & n15890 ) | ( x2 & ~n15891 ) | ( n15890 & ~n15891 ) ;
  assign n15893 = ( n15881 & ~n15883 ) | ( n15881 & n15892 ) | ( ~n15883 & n15892 ) ;
  assign n15894 = ( ~n15443 & n15452 ) | ( ~n15443 & n15454 ) | ( n15452 & n15454 ) ;
  assign n15895 = ( n15443 & ~n15455 ) | ( n15443 & n15894 ) | ( ~n15455 & n15894 ) ;
  assign n15896 = n36 & ~n10305 ;
  assign n15897 = n8967 & ~n9937 ;
  assign n15898 = ( x0 & n8966 ) | ( x0 & n10057 ) | ( n8966 & n10057 ) ;
  assign n15899 = ( n8966 & n15897 ) | ( n8966 & ~n15898 ) | ( n15897 & ~n15898 ) ;
  assign n15900 = n35 & n10302 ;
  assign n15901 = ( n35 & n15899 ) | ( n35 & ~n15900 ) | ( n15899 & ~n15900 ) ;
  assign n15902 = ( ~x2 & n15896 ) | ( ~x2 & n15901 ) | ( n15896 & n15901 ) ;
  assign n15903 = ( n15896 & n15901 ) | ( n15896 & ~n15902 ) | ( n15901 & ~n15902 ) ;
  assign n15904 = ( x2 & n15902 ) | ( x2 & ~n15903 ) | ( n15902 & ~n15903 ) ;
  assign n15905 = ( n15893 & n15895 ) | ( n15893 & n15904 ) | ( n15895 & n15904 ) ;
  assign n15906 = ( ~n15455 & n15464 ) | ( ~n15455 & n15466 ) | ( n15464 & n15466 ) ;
  assign n15907 = ( n15455 & ~n15467 ) | ( n15455 & n15906 ) | ( ~n15467 & n15906 ) ;
  assign n15908 = n36 & n10362 ;
  assign n15909 = n8967 & ~n10057 ;
  assign n15910 = ( x0 & n8966 ) | ( x0 & n10302 ) | ( n8966 & n10302 ) ;
  assign n15911 = ( n8966 & n15909 ) | ( n8966 & ~n15910 ) | ( n15909 & ~n15910 ) ;
  assign n15912 = n35 & ~n10346 ;
  assign n15913 = ( n35 & n15911 ) | ( n35 & ~n15912 ) | ( n15911 & ~n15912 ) ;
  assign n15914 = ( ~x2 & n15908 ) | ( ~x2 & n15913 ) | ( n15908 & n15913 ) ;
  assign n15915 = ( n15908 & n15913 ) | ( n15908 & ~n15914 ) | ( n15913 & ~n15914 ) ;
  assign n15916 = ( x2 & n15914 ) | ( x2 & ~n15915 ) | ( n15914 & ~n15915 ) ;
  assign n15917 = ( n15905 & n15907 ) | ( n15905 & n15916 ) | ( n15907 & n15916 ) ;
  assign n15918 = ( ~n15467 & n15476 ) | ( ~n15467 & n15478 ) | ( n15476 & n15478 ) ;
  assign n15919 = ( n15467 & ~n15479 ) | ( n15467 & n15918 ) | ( ~n15479 & n15918 ) ;
  assign n15920 = n36 & n10348 ;
  assign n15921 = n8967 & ~n10302 ;
  assign n15922 = n35 | n15921 ;
  assign n15923 = n9378 & ~n10346 ;
  assign n15924 = ( n9378 & n15922 ) | ( n9378 & ~n15923 ) | ( n15922 & ~n15923 ) ;
  assign n15925 = ( ~x2 & n15920 ) | ( ~x2 & n15924 ) | ( n15920 & n15924 ) ;
  assign n15926 = ( n15920 & n15924 ) | ( n15920 & ~n15925 ) | ( n15924 & ~n15925 ) ;
  assign n15927 = ( x2 & n15925 ) | ( x2 & ~n15926 ) | ( n15925 & ~n15926 ) ;
  assign n15928 = ( n15917 & n15919 ) | ( n15917 & n15927 ) | ( n15919 & n15927 ) ;
  assign n15929 = ( ~n15479 & n15488 ) | ( ~n15479 & n15490 ) | ( n15488 & n15490 ) ;
  assign n15930 = ( n15479 & ~n15491 ) | ( n15479 & n15929 ) | ( ~n15491 & n15929 ) ;
  assign n15931 = ~n8967 & n10346 ;
  assign n15932 = ( n9406 & n10346 ) | ( n9406 & ~n15931 ) | ( n10346 & ~n15931 ) ;
  assign n15933 = ( n36 & ~n11351 ) | ( n36 & n15932 ) | ( ~n11351 & n15932 ) ;
  assign n15934 = ( x2 & n11351 ) | ( x2 & ~n15933 ) | ( n11351 & ~n15933 ) ;
  assign n15935 = ( n15928 & n15930 ) | ( n15928 & n15934 ) | ( n15930 & n15934 ) ;
  assign n15936 = ( n11351 & n15064 ) | ( n11351 & ~n15066 ) | ( n15064 & ~n15066 ) ;
  assign n15937 = ( n15066 & ~n15067 ) | ( n15066 & n15936 ) | ( ~n15067 & n15936 ) ;
  assign n15938 = ( n15491 & n15935 ) | ( n15491 & n15937 ) | ( n15935 & n15937 ) ;
  assign n15939 = ( n15044 & n15046 ) | ( n15044 & n15054 ) | ( n15046 & n15054 ) ;
  assign n15940 = ( n15046 & n15055 ) | ( n15046 & ~n15939 ) | ( n15055 & ~n15939 ) ;
  assign n15941 = ( n15067 & n15938 ) | ( n15067 & ~n15940 ) | ( n15938 & ~n15940 ) ;
  assign n15942 = ( n14636 & ~n14638 ) | ( n14636 & n14643 ) | ( ~n14638 & n14643 ) ;
  assign n15943 = ( n14638 & ~n14644 ) | ( n14638 & n15942 ) | ( ~n14644 & n15942 ) ;
  assign n15944 = ( n15055 & n15941 ) | ( n15055 & n15943 ) | ( n15941 & n15943 ) ;
  assign n15945 = ( n11392 & n14257 ) | ( n11392 & n14259 ) | ( n14257 & n14259 ) ;
  assign n15946 = ( n14259 & n14260 ) | ( n14259 & ~n15945 ) | ( n14260 & ~n15945 ) ;
  assign n15947 = ( n14644 & n15944 ) | ( n14644 & ~n15946 ) | ( n15944 & ~n15946 ) ;
  assign n15948 = ( n13894 & n13902 ) | ( n13894 & n13904 ) | ( n13902 & n13904 ) ;
  assign n15949 = ( n13904 & n13905 ) | ( n13904 & ~n15948 ) | ( n13905 & ~n15948 ) ;
  assign n15950 = ( n14260 & n15947 ) | ( n14260 & ~n15949 ) | ( n15947 & ~n15949 ) ;
  assign n15951 = ( n13558 & ~n13560 ) | ( n13558 & n13565 ) | ( ~n13560 & n13565 ) ;
  assign n15952 = ( n13560 & ~n13566 ) | ( n13560 & n15951 ) | ( ~n13566 & n15951 ) ;
  assign n15953 = ( n13905 & n15950 ) | ( n13905 & n15952 ) | ( n15950 & n15952 ) ;
  assign n15954 = ( n13248 & n13251 ) | ( n13248 & n13253 ) | ( n13251 & n13253 ) ;
  assign n15955 = ( n13253 & n13254 ) | ( n13253 & ~n15954 ) | ( n13254 & ~n15954 ) ;
  assign n15956 = ( n13566 & n15953 ) | ( n13566 & ~n15955 ) | ( n15953 & ~n15955 ) ;
  assign n15957 = ( n12958 & n12966 ) | ( n12958 & n12968 ) | ( n12966 & n12968 ) ;
  assign n15958 = ( n12968 & n12969 ) | ( n12968 & ~n15957 ) | ( n12969 & ~n15957 ) ;
  assign n15959 = ( n13254 & n15956 ) | ( n13254 & ~n15958 ) | ( n15956 & ~n15958 ) ;
  assign n15960 = ( n12695 & n12697 ) | ( n12695 & n12702 ) | ( n12697 & n12702 ) ;
  assign n15961 = ( n12697 & n12703 ) | ( n12697 & ~n15960 ) | ( n12703 & ~n15960 ) ;
  assign n15962 = ( n12969 & n15959 ) | ( n12969 & ~n15961 ) | ( n15959 & ~n15961 ) ;
  assign n15963 = ( n12457 & n12460 ) | ( n12457 & n12462 ) | ( n12460 & n12462 ) ;
  assign n15964 = ( n12462 & n12463 ) | ( n12462 & ~n15963 ) | ( n12463 & ~n15963 ) ;
  assign n15965 = ( n12703 & n15962 ) | ( n12703 & ~n15964 ) | ( n15962 & ~n15964 ) ;
  assign n15966 = ( n12353 & n12361 ) | ( n12353 & n12363 ) | ( n12361 & n12363 ) ;
  assign n15967 = ( n12363 & n12364 ) | ( n12363 & ~n15966 ) | ( n12364 & ~n15966 ) ;
  assign n15968 = ( n12463 & n15965 ) | ( n12463 & ~n15967 ) | ( n15965 & ~n15967 ) ;
  assign n15969 = ( n12252 & ~n12254 ) | ( n12252 & n12259 ) | ( ~n12254 & n12259 ) ;
  assign n15970 = ( n12254 & ~n12260 ) | ( n12254 & n15969 ) | ( ~n12260 & n15969 ) ;
  assign n15971 = ( n12364 & n15968 ) | ( n12364 & n15970 ) | ( n15968 & n15970 ) ;
  assign n15972 = ( n11797 & ~n11800 ) | ( n11797 & n11802 ) | ( ~n11800 & n11802 ) ;
  assign n15973 = ( n11800 & ~n11803 ) | ( n11800 & n15972 ) | ( ~n11803 & n15972 ) ;
  assign n15974 = ( n12260 & n15971 ) | ( n12260 & n15973 ) | ( n15971 & n15973 ) ;
  assign n15975 = ( n11705 & n11713 ) | ( n11705 & n11715 ) | ( n11713 & n11715 ) ;
  assign n15976 = ( n11715 & n11716 ) | ( n11715 & ~n15975 ) | ( n11716 & ~n15975 ) ;
  assign n15977 = ( n11803 & n15974 ) | ( n11803 & ~n15976 ) | ( n15974 & ~n15976 ) ;
  assign n15978 = ( n11503 & ~n11505 ) | ( n11503 & n11510 ) | ( ~n11505 & n11510 ) ;
  assign n15979 = ( n11505 & ~n11511 ) | ( n11505 & n15978 ) | ( ~n11511 & n15978 ) ;
  assign n15980 = ( n11716 & n15977 ) | ( n11716 & n15979 ) | ( n15977 & n15979 ) ;
  assign n15981 = ( n11345 & n11347 ) | ( n11345 & n11349 ) | ( n11347 & n11349 ) ;
  assign n15982 = ( n11347 & n11350 ) | ( n11347 & ~n15981 ) | ( n11350 & ~n15981 ) ;
  assign n15983 = ( n11511 & n15980 ) | ( n11511 & ~n15982 ) | ( n15980 & ~n15982 ) ;
  assign n15984 = ( n11253 & ~n11261 ) | ( n11253 & n11263 ) | ( ~n11261 & n11263 ) ;
  assign n15985 = ( n11261 & ~n11264 ) | ( n11261 & n15984 ) | ( ~n11264 & n15984 ) ;
  assign n15986 = ( n11350 & n15983 ) | ( n11350 & n15985 ) | ( n15983 & n15985 ) ;
  assign n15987 = ( n11187 & n11189 ) | ( n11187 & n11195 ) | ( n11189 & n11195 ) ;
  assign n15988 = ( n11189 & n11196 ) | ( n11189 & ~n15987 ) | ( n11196 & ~n15987 ) ;
  assign n15989 = ( n11264 & n15986 ) | ( n11264 & ~n15988 ) | ( n15986 & ~n15988 ) ;
  assign n15990 = ( n10242 & n10919 ) | ( n10242 & n10921 ) | ( n10919 & n10921 ) ;
  assign n15991 = ( n10921 & n10922 ) | ( n10921 & ~n15990 ) | ( n10922 & ~n15990 ) ;
  assign n15992 = ( n11196 & n15989 ) | ( n11196 & ~n15991 ) | ( n15989 & ~n15991 ) ;
  assign n15993 = ( ~n10798 & n10800 ) | ( ~n10798 & n10808 ) | ( n10800 & n10808 ) ;
  assign n15994 = ( ~n10808 & n10809 ) | ( ~n10808 & n15993 ) | ( n10809 & n15993 ) ;
  assign n15995 = ( n10922 & n15992 ) | ( n10922 & ~n15994 ) | ( n15992 & ~n15994 ) ;
  assign n15996 = ( ~n10732 & n10734 ) | ( ~n10732 & n10739 ) | ( n10734 & n10739 ) ;
  assign n15997 = ( n10732 & ~n10740 ) | ( n10732 & n15996 ) | ( ~n10740 & n15996 ) ;
  assign n15998 = ( n10809 & n15995 ) | ( n10809 & n15997 ) | ( n15995 & n15997 ) ;
  assign n15999 = ( ~n10694 & n10696 ) | ( ~n10694 & n10698 ) | ( n10696 & n10698 ) ;
  assign n16000 = ( n10694 & ~n10699 ) | ( n10694 & n15999 ) | ( ~n10699 & n15999 ) ;
  assign n16001 = ( n10740 & n15998 ) | ( n10740 & n16000 ) | ( n15998 & n16000 ) ;
  assign n16002 = ( ~n10493 & n10495 ) | ( ~n10493 & n10503 ) | ( n10495 & n10503 ) ;
  assign n16003 = ( n10493 & ~n10504 ) | ( n10493 & n16002 ) | ( ~n10504 & n16002 ) ;
  assign n16004 = ( n10699 & n16001 ) | ( n10699 & n16003 ) | ( n16001 & n16003 ) ;
  assign n16005 = ( n10405 & n10411 ) | ( n10405 & n10413 ) | ( n10411 & n10413 ) ;
  assign n16006 = ( n10413 & n10414 ) | ( n10413 & ~n16005 ) | ( n10414 & ~n16005 ) ;
  assign n16007 = ( n10504 & n16004 ) | ( n10504 & ~n16006 ) | ( n16004 & ~n16006 ) ;
  assign n16008 = ( n38 & n10360 ) | ( n38 & ~n10371 ) | ( n10360 & ~n10371 ) ;
  assign n16009 = ( n10371 & ~n10372 ) | ( n10371 & n16008 ) | ( ~n10372 & n16008 ) ;
  assign n16010 = ( n10414 & n16007 ) | ( n10414 & n16009 ) | ( n16007 & n16009 ) ;
  assign n16011 = ( ~n10358 & n10372 ) | ( ~n10358 & n16010 ) | ( n10372 & n16010 ) ;
  assign n16012 = ( n10358 & n10372 ) | ( n10358 & n16010 ) | ( n10372 & n16010 ) ;
  assign n16013 = ( n10358 & n16011 ) | ( n10358 & ~n16012 ) | ( n16011 & ~n16012 ) ;
  assign n16014 = ( ~n10414 & n16007 ) | ( ~n10414 & n16009 ) | ( n16007 & n16009 ) ;
  assign n16015 = ( n10414 & ~n16010 ) | ( n10414 & n16014 ) | ( ~n16010 & n16014 ) ;
  assign n16016 = ( n10504 & ~n16004 ) | ( n10504 & n16006 ) | ( ~n16004 & n16006 ) ;
  assign n16017 = ( ~n10504 & n16007 ) | ( ~n10504 & n16016 ) | ( n16007 & n16016 ) ;
  assign n16018 = ( ~n10699 & n16001 ) | ( ~n10699 & n16003 ) | ( n16001 & n16003 ) ;
  assign n16019 = ( n10699 & ~n16004 ) | ( n10699 & n16018 ) | ( ~n16004 & n16018 ) ;
  assign n16020 = ( ~n10740 & n15998 ) | ( ~n10740 & n16000 ) | ( n15998 & n16000 ) ;
  assign n16021 = ( n10740 & ~n16001 ) | ( n10740 & n16020 ) | ( ~n16001 & n16020 ) ;
  assign n16022 = ( ~n10809 & n15995 ) | ( ~n10809 & n15997 ) | ( n15995 & n15997 ) ;
  assign n16023 = ( n10809 & ~n15998 ) | ( n10809 & n16022 ) | ( ~n15998 & n16022 ) ;
  assign n16024 = ( n10922 & ~n15992 ) | ( n10922 & n15994 ) | ( ~n15992 & n15994 ) ;
  assign n16025 = ( ~n10922 & n15995 ) | ( ~n10922 & n16024 ) | ( n15995 & n16024 ) ;
  assign n16026 = ( n11196 & ~n15989 ) | ( n11196 & n15991 ) | ( ~n15989 & n15991 ) ;
  assign n16027 = ( ~n11196 & n15992 ) | ( ~n11196 & n16026 ) | ( n15992 & n16026 ) ;
  assign n16028 = ( n11264 & ~n15986 ) | ( n11264 & n15988 ) | ( ~n15986 & n15988 ) ;
  assign n16029 = ( ~n11264 & n15989 ) | ( ~n11264 & n16028 ) | ( n15989 & n16028 ) ;
  assign n16030 = ( n11350 & ~n15983 ) | ( n11350 & n15985 ) | ( ~n15983 & n15985 ) ;
  assign n16031 = ( n15983 & ~n15986 ) | ( n15983 & n16030 ) | ( ~n15986 & n16030 ) ;
  assign n16032 = ( n11511 & ~n15980 ) | ( n11511 & n15982 ) | ( ~n15980 & n15982 ) ;
  assign n16033 = ( ~n11511 & n15983 ) | ( ~n11511 & n16032 ) | ( n15983 & n16032 ) ;
  assign n16034 = ( n11716 & ~n15977 ) | ( n11716 & n15979 ) | ( ~n15977 & n15979 ) ;
  assign n16035 = ( n15977 & ~n15980 ) | ( n15977 & n16034 ) | ( ~n15980 & n16034 ) ;
  assign n16036 = ( n11803 & ~n15974 ) | ( n11803 & n15976 ) | ( ~n15974 & n15976 ) ;
  assign n16037 = ( ~n11803 & n15977 ) | ( ~n11803 & n16036 ) | ( n15977 & n16036 ) ;
  assign n16038 = ( n12260 & ~n15971 ) | ( n12260 & n15973 ) | ( ~n15971 & n15973 ) ;
  assign n16039 = ( n15971 & ~n15974 ) | ( n15971 & n16038 ) | ( ~n15974 & n16038 ) ;
  assign n16040 = ( n12364 & ~n15968 ) | ( n12364 & n15970 ) | ( ~n15968 & n15970 ) ;
  assign n16041 = ( n15968 & ~n15971 ) | ( n15968 & n16040 ) | ( ~n15971 & n16040 ) ;
  assign n16042 = ( n12463 & ~n15965 ) | ( n12463 & n15967 ) | ( ~n15965 & n15967 ) ;
  assign n16043 = ( ~n12463 & n15968 ) | ( ~n12463 & n16042 ) | ( n15968 & n16042 ) ;
  assign n16044 = ( n12703 & ~n15962 ) | ( n12703 & n15964 ) | ( ~n15962 & n15964 ) ;
  assign n16045 = ( ~n12703 & n15965 ) | ( ~n12703 & n16044 ) | ( n15965 & n16044 ) ;
  assign n16046 = ( n12969 & ~n15959 ) | ( n12969 & n15961 ) | ( ~n15959 & n15961 ) ;
  assign n16047 = ( ~n12969 & n15962 ) | ( ~n12969 & n16046 ) | ( n15962 & n16046 ) ;
  assign n16048 = ( n13254 & ~n15956 ) | ( n13254 & n15958 ) | ( ~n15956 & n15958 ) ;
  assign n16049 = ( ~n13254 & n15959 ) | ( ~n13254 & n16048 ) | ( n15959 & n16048 ) ;
  assign n16050 = ( n13566 & ~n15953 ) | ( n13566 & n15955 ) | ( ~n15953 & n15955 ) ;
  assign n16051 = ( ~n13566 & n15956 ) | ( ~n13566 & n16050 ) | ( n15956 & n16050 ) ;
  assign n16052 = ( n13905 & ~n15950 ) | ( n13905 & n15952 ) | ( ~n15950 & n15952 ) ;
  assign n16053 = ( n15950 & ~n15953 ) | ( n15950 & n16052 ) | ( ~n15953 & n16052 ) ;
  assign n16054 = ( n14260 & ~n15947 ) | ( n14260 & n15949 ) | ( ~n15947 & n15949 ) ;
  assign n16055 = ( ~n14260 & n15950 ) | ( ~n14260 & n16054 ) | ( n15950 & n16054 ) ;
  assign n16056 = ( n14644 & ~n15944 ) | ( n14644 & n15946 ) | ( ~n15944 & n15946 ) ;
  assign n16057 = ( ~n14644 & n15947 ) | ( ~n14644 & n16056 ) | ( n15947 & n16056 ) ;
  assign n16058 = ( n15055 & ~n15941 ) | ( n15055 & n15943 ) | ( ~n15941 & n15943 ) ;
  assign n16059 = ( n15941 & ~n15944 ) | ( n15941 & n16058 ) | ( ~n15944 & n16058 ) ;
  assign n16060 = ( n15067 & ~n15938 ) | ( n15067 & n15940 ) | ( ~n15938 & n15940 ) ;
  assign n16061 = ( ~n15067 & n15941 ) | ( ~n15067 & n16060 ) | ( n15941 & n16060 ) ;
  assign n16062 = ( n15491 & ~n15935 ) | ( n15491 & n15937 ) | ( ~n15935 & n15937 ) ;
  assign n16063 = ( n15935 & ~n15938 ) | ( n15935 & n16062 ) | ( ~n15938 & n16062 ) ;
  assign n16064 = ( ~n15928 & n15930 ) | ( ~n15928 & n15934 ) | ( n15930 & n15934 ) ;
  assign n16065 = ( n15928 & ~n15935 ) | ( n15928 & n16064 ) | ( ~n15935 & n16064 ) ;
  assign n16066 = ( ~n15917 & n15919 ) | ( ~n15917 & n15927 ) | ( n15919 & n15927 ) ;
  assign n16067 = ( n15917 & ~n15928 ) | ( n15917 & n16066 ) | ( ~n15928 & n16066 ) ;
  assign n16068 = ( ~n15905 & n15907 ) | ( ~n15905 & n15916 ) | ( n15907 & n15916 ) ;
  assign n16069 = ( n15905 & ~n15917 ) | ( n15905 & n16068 ) | ( ~n15917 & n16068 ) ;
  assign n16070 = ( ~n15893 & n15895 ) | ( ~n15893 & n15904 ) | ( n15895 & n15904 ) ;
  assign n16071 = ( n15893 & ~n15905 ) | ( n15893 & n16070 ) | ( ~n15905 & n16070 ) ;
  assign n16072 = ( ~n15881 & n15883 ) | ( ~n15881 & n15892 ) | ( n15883 & n15892 ) ;
  assign n16073 = ( ~n15892 & n15893 ) | ( ~n15892 & n16072 ) | ( n15893 & n16072 ) ;
  assign n16074 = ( ~n15869 & n15871 ) | ( ~n15869 & n15880 ) | ( n15871 & n15880 ) ;
  assign n16075 = ( ~n15880 & n15881 ) | ( ~n15880 & n16074 ) | ( n15881 & n16074 ) ;
  assign n16076 = ( ~n15857 & n15859 ) | ( ~n15857 & n15868 ) | ( n15859 & n15868 ) ;
  assign n16077 = ( n15857 & ~n15869 ) | ( n15857 & n16076 ) | ( ~n15869 & n16076 ) ;
  assign n16078 = ( ~n15845 & n15847 ) | ( ~n15845 & n15856 ) | ( n15847 & n15856 ) ;
  assign n16079 = ( ~n15856 & n15857 ) | ( ~n15856 & n16078 ) | ( n15857 & n16078 ) ;
  assign n16080 = ( ~n15833 & n15835 ) | ( ~n15833 & n15844 ) | ( n15835 & n15844 ) ;
  assign n16081 = ( ~n15844 & n15845 ) | ( ~n15844 & n16080 ) | ( n15845 & n16080 ) ;
  assign n16082 = ( n16077 & ~n16079 ) | ( n16077 & n16081 ) | ( ~n16079 & n16081 ) ;
  assign n16083 = ~n16077 & n16082 ;
  assign n16084 = n16079 | n16083 ;
  assign n16085 = ( n16075 & ~n16077 ) | ( n16075 & n16084 ) | ( ~n16077 & n16084 ) ;
  assign n16086 = ( n16073 & n16075 ) | ( n16073 & n16085 ) | ( n16075 & n16085 ) ;
  assign n16087 = ( ~n16071 & n16073 ) | ( ~n16071 & n16086 ) | ( n16073 & n16086 ) ;
  assign n16088 = ( n16069 & n16071 ) | ( n16069 & ~n16087 ) | ( n16071 & ~n16087 ) ;
  assign n16089 = ( n16067 & n16069 ) | ( n16067 & n16088 ) | ( n16069 & n16088 ) ;
  assign n16090 = ( n16065 & n16067 ) | ( n16065 & n16089 ) | ( n16067 & n16089 ) ;
  assign n16091 = ( n16063 & n16065 ) | ( n16063 & n16090 ) | ( n16065 & n16090 ) ;
  assign n16092 = ( ~n16061 & n16063 ) | ( ~n16061 & n16091 ) | ( n16063 & n16091 ) ;
  assign n16093 = ( n16059 & ~n16061 ) | ( n16059 & n16092 ) | ( ~n16061 & n16092 ) ;
  assign n16094 = ( ~n16057 & n16059 ) | ( ~n16057 & n16093 ) | ( n16059 & n16093 ) ;
  assign n16095 = ( n16055 & n16057 ) | ( n16055 & ~n16094 ) | ( n16057 & ~n16094 ) ;
  assign n16096 = ( ~n16053 & n16055 ) | ( ~n16053 & n16095 ) | ( n16055 & n16095 ) ;
  assign n16097 = ( n16051 & ~n16053 ) | ( n16051 & n16096 ) | ( ~n16053 & n16096 ) ;
  assign n16098 = ( n16049 & n16051 ) | ( n16049 & n16097 ) | ( n16051 & n16097 ) ;
  assign n16099 = ( n16047 & n16049 ) | ( n16047 & n16098 ) | ( n16049 & n16098 ) ;
  assign n16100 = ( n16045 & n16047 ) | ( n16045 & n16099 ) | ( n16047 & n16099 ) ;
  assign n16101 = ( n16043 & n16045 ) | ( n16043 & n16100 ) | ( n16045 & n16100 ) ;
  assign n16102 = ( ~n16041 & n16043 ) | ( ~n16041 & n16101 ) | ( n16043 & n16101 ) ;
  assign n16103 = ( n16039 & n16041 ) | ( n16039 & ~n16102 ) | ( n16041 & ~n16102 ) ;
  assign n16104 = ( ~n16037 & n16039 ) | ( ~n16037 & n16103 ) | ( n16039 & n16103 ) ;
  assign n16105 = ( n16035 & ~n16037 ) | ( n16035 & n16104 ) | ( ~n16037 & n16104 ) ;
  assign n16106 = ( ~n16033 & n16035 ) | ( ~n16033 & n16105 ) | ( n16035 & n16105 ) ;
  assign n16107 = ( n16031 & ~n16033 ) | ( n16031 & n16106 ) | ( ~n16033 & n16106 ) ;
  assign n16108 = ( ~n16029 & n16031 ) | ( ~n16029 & n16107 ) | ( n16031 & n16107 ) ;
  assign n16109 = ( n16027 & n16029 ) | ( n16027 & ~n16108 ) | ( n16029 & ~n16108 ) ;
  assign n16110 = ( n16025 & n16027 ) | ( n16025 & n16109 ) | ( n16027 & n16109 ) ;
  assign n16111 = ( ~n16023 & n16025 ) | ( ~n16023 & n16110 ) | ( n16025 & n16110 ) ;
  assign n16112 = ( n16021 & n16023 ) | ( n16021 & ~n16111 ) | ( n16023 & ~n16111 ) ;
  assign n16113 = ( n16019 & n16021 ) | ( n16019 & n16112 ) | ( n16021 & n16112 ) ;
  assign n16114 = ( ~n16017 & n16019 ) | ( ~n16017 & n16113 ) | ( n16019 & n16113 ) ;
  assign n16115 = ( n16015 & ~n16017 ) | ( n16015 & n16114 ) | ( ~n16017 & n16114 ) ;
  assign n16116 = ( ~n16013 & n16015 ) | ( ~n16013 & n16115 ) | ( n16015 & n16115 ) ;
  assign n16117 = n607 & ~n9937 ;
  assign n16118 = n1250 & ~n10057 ;
  assign n16119 = n16117 | n16118 ;
  assign n16120 = n606 & n10302 ;
  assign n16121 = ( n606 & n16119 ) | ( n606 & ~n16120 ) | ( n16119 & ~n16120 ) ;
  assign n16122 = n1248 & ~n10305 ;
  assign n16123 = n16121 | n16122 ;
  assign n16124 = ( n414 & ~n455 ) | ( n414 & n1286 ) | ( ~n455 & n1286 ) ;
  assign n16125 = ( n455 & ~n3687 ) | ( n455 & n16124 ) | ( ~n3687 & n16124 ) ;
  assign n16126 = n3687 | n16125 ;
  assign n16127 = ( n460 & n16123 ) | ( n460 & n16126 ) | ( n16123 & n16126 ) ;
  assign n16128 = ( n460 & ~n16123 ) | ( n460 & n16126 ) | ( ~n16123 & n16126 ) ;
  assign n16129 = ( n16123 & ~n16127 ) | ( n16123 & n16128 ) | ( ~n16127 & n16128 ) ;
  assign n16130 = x29 & n3698 ;
  assign n16131 = n53 | n3698 ;
  assign n16132 = ~n16130 & n16131 ;
  assign n16133 = ( n10067 & n16129 ) | ( n10067 & n16132 ) | ( n16129 & n16132 ) ;
  assign n16134 = ( n10067 & ~n16129 ) | ( n10067 & n16132 ) | ( ~n16129 & n16132 ) ;
  assign n16135 = ( n16129 & ~n16133 ) | ( n16129 & n16134 ) | ( ~n16133 & n16134 ) ;
  assign n16136 = ( n10356 & n16011 ) | ( n10356 & n16135 ) | ( n16011 & n16135 ) ;
  assign n16137 = ( ~n10356 & n16011 ) | ( ~n10356 & n16135 ) | ( n16011 & n16135 ) ;
  assign n16138 = ( n10356 & ~n16136 ) | ( n10356 & n16137 ) | ( ~n16136 & n16137 ) ;
  assign n16139 = ( ~n16013 & n16116 ) | ( ~n16013 & n16138 ) | ( n16116 & n16138 ) ;
  assign n16140 = ( n16017 & n16019 ) | ( n16017 & ~n16113 ) | ( n16019 & ~n16113 ) ;
  assign n16141 = ( ~n16015 & n16113 ) | ( ~n16015 & n16140 ) | ( n16113 & n16140 ) ;
  assign n16142 = ( n16013 & ~n16017 ) | ( n16013 & n16141 ) | ( ~n16017 & n16141 ) ;
  assign n16143 = ( n16015 & n16138 ) | ( n16015 & n16142 ) | ( n16138 & n16142 ) ;
  assign n16144 = ( n16013 & n16139 ) | ( n16013 & ~n16143 ) | ( n16139 & ~n16143 ) ;
  assign n16145 = n36 & ~n16144 ;
  assign n16146 = n8967 & n16015 ;
  assign n16147 = ( x0 & n8966 ) | ( x0 & n16013 ) | ( n8966 & n16013 ) ;
  assign n16148 = ( n8966 & n16146 ) | ( n8966 & ~n16147 ) | ( n16146 & ~n16147 ) ;
  assign n16149 = n35 & ~n16138 ;
  assign n16150 = ( n35 & n16148 ) | ( n35 & ~n16149 ) | ( n16148 & ~n16149 ) ;
  assign n16151 = ( ~x2 & n16145 ) | ( ~x2 & n16150 ) | ( n16145 & n16150 ) ;
  assign n16152 = ( n16145 & n16150 ) | ( n16145 & ~n16151 ) | ( n16150 & ~n16151 ) ;
  assign n16153 = ( x2 & n16151 ) | ( x2 & ~n16152 ) | ( n16151 & ~n16152 ) ;
  assign n16154 = n8228 & ~n16081 ;
  assign n16155 = n16079 & ~n16081 ;
  assign n16156 = ( n36 & n16082 ) | ( n36 & n16155 ) | ( n16082 & n16155 ) ;
  assign n16157 = n35 & n16077 ;
  assign n16158 = x1 & ~n16079 ;
  assign n16159 = ( ~x2 & n16081 ) | ( ~x2 & n16158 ) | ( n16081 & n16158 ) ;
  assign n16160 = n16081 & ~n16159 ;
  assign n16161 = ( n16156 & ~n16157 ) | ( n16156 & n16160 ) | ( ~n16157 & n16160 ) ;
  assign n16162 = ( n16154 & ~n16156 ) | ( n16154 & n16161 ) | ( ~n16156 & n16161 ) ;
  assign n16163 = n8967 & ~n16079 ;
  assign n16164 = ( x0 & n8966 ) | ( x0 & ~n16077 ) | ( n8966 & ~n16077 ) ;
  assign n16165 = ( n8966 & n16163 ) | ( n8966 & ~n16164 ) | ( n16163 & ~n16164 ) ;
  assign n16166 = n35 & n16075 ;
  assign n16167 = ( n35 & n16165 ) | ( n35 & ~n16166 ) | ( n16165 & ~n16166 ) ;
  assign n16168 = ( n16075 & n16077 ) | ( n16075 & n16084 ) | ( n16077 & n16084 ) ;
  assign n16169 = ( n16077 & n16085 ) | ( n16077 & ~n16168 ) | ( n16085 & ~n16168 ) ;
  assign n16170 = n36 & n16169 ;
  assign n16171 = n16167 | n16170 ;
  assign n16172 = ( x2 & n16162 ) | ( x2 & n16171 ) | ( n16162 & n16171 ) ;
  assign n16173 = x2 & ~n16171 ;
  assign n16174 = ( ~x2 & n16172 ) | ( ~x2 & n16173 ) | ( n16172 & n16173 ) ;
  assign n16175 = ( n16073 & n16075 ) | ( n16073 & ~n16085 ) | ( n16075 & ~n16085 ) ;
  assign n16176 = ( n16085 & ~n16086 ) | ( n16085 & n16175 ) | ( ~n16086 & n16175 ) ;
  assign n16177 = n36 & ~n16176 ;
  assign n16178 = n8967 & n16077 ;
  assign n16179 = ( x0 & n8966 ) | ( x0 & n16075 ) | ( n8966 & n16075 ) ;
  assign n16180 = ( n8966 & n16178 ) | ( n8966 & ~n16179 ) | ( n16178 & ~n16179 ) ;
  assign n16181 = n35 & n16073 ;
  assign n16182 = ( n35 & n16180 ) | ( n35 & ~n16181 ) | ( n16180 & ~n16181 ) ;
  assign n16183 = ( ~x2 & n16177 ) | ( ~x2 & n16182 ) | ( n16177 & n16182 ) ;
  assign n16184 = ( n16177 & n16182 ) | ( n16177 & ~n16183 ) | ( n16182 & ~n16183 ) ;
  assign n16185 = ( x2 & n16183 ) | ( x2 & ~n16184 ) | ( n16183 & ~n16184 ) ;
  assign n16186 = x5 & n16154 ;
  assign n16187 = ~n16079 & n16081 ;
  assign n16188 = ( n8230 & n16155 ) | ( n8230 & n16187 ) | ( n16155 & n16187 ) ;
  assign n16189 = n8225 | n16081 ;
  assign n16190 = n8229 & ~n16079 ;
  assign n16191 = ( ~n16081 & n16189 ) | ( ~n16081 & n16190 ) | ( n16189 & n16190 ) ;
  assign n16192 = ( n16186 & n16188 ) | ( n16186 & n16191 ) | ( n16188 & n16191 ) ;
  assign n16193 = n16188 | n16191 ;
  assign n16194 = ~n16186 & n16193 ;
  assign n16195 = ( n16186 & ~n16192 ) | ( n16186 & n16194 ) | ( ~n16192 & n16194 ) ;
  assign n16196 = ( n16174 & n16185 ) | ( n16174 & n16195 ) | ( n16185 & n16195 ) ;
  assign n16197 = ( x5 & n16186 ) | ( x5 & n16193 ) | ( n16186 & n16193 ) ;
  assign n16198 = n16077 & ~n16187 ;
  assign n16199 = ( n8230 & n16083 ) | ( n8230 & n16198 ) | ( n16083 & n16198 ) ;
  assign n16200 = n8226 & ~n16081 ;
  assign n16201 = n8225 & ~n16079 ;
  assign n16202 = n16200 | n16201 ;
  assign n16203 = n8229 & ~n16077 ;
  assign n16204 = ( n8229 & n16202 ) | ( n8229 & ~n16203 ) | ( n16202 & ~n16203 ) ;
  assign n16205 = ( ~n16197 & n16199 ) | ( ~n16197 & n16204 ) | ( n16199 & n16204 ) ;
  assign n16206 = ( n16199 & n16204 ) | ( n16199 & ~n16205 ) | ( n16204 & ~n16205 ) ;
  assign n16207 = ( n16197 & n16205 ) | ( n16197 & ~n16206 ) | ( n16205 & ~n16206 ) ;
  assign n16208 = ( n16071 & n16073 ) | ( n16071 & ~n16086 ) | ( n16073 & ~n16086 ) ;
  assign n16209 = ( ~n16073 & n16087 ) | ( ~n16073 & n16208 ) | ( n16087 & n16208 ) ;
  assign n16210 = n36 & n16209 ;
  assign n16211 = n8967 & ~n16075 ;
  assign n16212 = ( x0 & n8966 ) | ( x0 & n16073 ) | ( n8966 & n16073 ) ;
  assign n16213 = ( n8966 & n16211 ) | ( n8966 & ~n16212 ) | ( n16211 & ~n16212 ) ;
  assign n16214 = n35 & ~n16071 ;
  assign n16215 = ( n35 & n16213 ) | ( n35 & ~n16214 ) | ( n16213 & ~n16214 ) ;
  assign n16216 = ( ~x2 & n16210 ) | ( ~x2 & n16215 ) | ( n16210 & n16215 ) ;
  assign n16217 = ( n16210 & n16215 ) | ( n16210 & ~n16216 ) | ( n16215 & ~n16216 ) ;
  assign n16218 = ( x2 & n16216 ) | ( x2 & ~n16217 ) | ( n16216 & ~n16217 ) ;
  assign n16219 = ( n16196 & n16207 ) | ( n16196 & n16218 ) | ( n16207 & n16218 ) ;
  assign n16220 = ( n16069 & n16071 ) | ( n16069 & ~n16088 ) | ( n16071 & ~n16088 ) ;
  assign n16221 = ( n16087 & n16088 ) | ( n16087 & ~n16220 ) | ( n16088 & ~n16220 ) ;
  assign n16222 = n36 & ~n16221 ;
  assign n16223 = n8967 & ~n16073 ;
  assign n16224 = ( x0 & n8966 ) | ( x0 & ~n16071 ) | ( n8966 & ~n16071 ) ;
  assign n16225 = ( n8966 & n16223 ) | ( n8966 & ~n16224 ) | ( n16223 & ~n16224 ) ;
  assign n16226 = n35 & ~n16069 ;
  assign n16227 = ( n35 & n16225 ) | ( n35 & ~n16226 ) | ( n16225 & ~n16226 ) ;
  assign n16228 = ( ~x2 & n16222 ) | ( ~x2 & n16227 ) | ( n16222 & n16227 ) ;
  assign n16229 = ( n16222 & n16227 ) | ( n16222 & ~n16228 ) | ( n16227 & ~n16228 ) ;
  assign n16230 = ( x2 & n16228 ) | ( x2 & ~n16229 ) | ( n16228 & ~n16229 ) ;
  assign n16231 = x5 & ~n16205 ;
  assign n16232 = ~n16197 & n16231 ;
  assign n16233 = n7878 & ~n16081 ;
  assign n16234 = n8230 & n16169 ;
  assign n16235 = n8229 & ~n16075 ;
  assign n16236 = n8226 & ~n16079 ;
  assign n16237 = n8225 & n16077 ;
  assign n16238 = n16236 | n16237 ;
  assign n16239 = ( ~n16234 & n16235 ) | ( ~n16234 & n16238 ) | ( n16235 & n16238 ) ;
  assign n16240 = ( ~x5 & n16234 ) | ( ~x5 & n16239 ) | ( n16234 & n16239 ) ;
  assign n16241 = ( n16234 & n16239 ) | ( n16234 & ~n16240 ) | ( n16239 & ~n16240 ) ;
  assign n16242 = ( x5 & n16240 ) | ( x5 & ~n16241 ) | ( n16240 & ~n16241 ) ;
  assign n16243 = ( n16232 & n16233 ) | ( n16232 & n16242 ) | ( n16233 & n16242 ) ;
  assign n16244 = ( ~n16232 & n16233 ) | ( ~n16232 & n16242 ) | ( n16233 & n16242 ) ;
  assign n16245 = ( n16232 & ~n16243 ) | ( n16232 & n16244 ) | ( ~n16243 & n16244 ) ;
  assign n16246 = ( n16219 & n16230 ) | ( n16219 & n16245 ) | ( n16230 & n16245 ) ;
  assign n16247 = n8230 & ~n16176 ;
  assign n16248 = n8229 & ~n16073 ;
  assign n16249 = n8226 & n16077 ;
  assign n16250 = n8225 & ~n16075 ;
  assign n16251 = n16249 | n16250 ;
  assign n16252 = ( ~n16247 & n16248 ) | ( ~n16247 & n16251 ) | ( n16248 & n16251 ) ;
  assign n16253 = ( ~x5 & n16247 ) | ( ~x5 & n16252 ) | ( n16247 & n16252 ) ;
  assign n16254 = ( n16247 & n16252 ) | ( n16247 & ~n16253 ) | ( n16252 & ~n16253 ) ;
  assign n16255 = ( x5 & n16253 ) | ( x5 & ~n16254 ) | ( n16253 & ~n16254 ) ;
  assign n16256 = x8 & n16233 ;
  assign n16257 = ( n7296 & n16155 ) | ( n7296 & n16187 ) | ( n16155 & n16187 ) ;
  assign n16258 = n7299 | n16081 ;
  assign n16259 = n7879 & ~n16079 ;
  assign n16260 = ( ~n16081 & n16258 ) | ( ~n16081 & n16259 ) | ( n16258 & n16259 ) ;
  assign n16261 = ( n16256 & n16257 ) | ( n16256 & n16260 ) | ( n16257 & n16260 ) ;
  assign n16262 = n16257 | n16260 ;
  assign n16263 = ~n16256 & n16262 ;
  assign n16264 = ( n16256 & ~n16261 ) | ( n16256 & n16263 ) | ( ~n16261 & n16263 ) ;
  assign n16265 = ( n16243 & n16255 ) | ( n16243 & n16264 ) | ( n16255 & n16264 ) ;
  assign n16266 = ( ~n16243 & n16255 ) | ( ~n16243 & n16264 ) | ( n16255 & n16264 ) ;
  assign n16267 = ( n16243 & ~n16265 ) | ( n16243 & n16266 ) | ( ~n16265 & n16266 ) ;
  assign n16268 = ( n16067 & n16069 ) | ( n16067 & ~n16088 ) | ( n16069 & ~n16088 ) ;
  assign n16269 = ( n16088 & ~n16089 ) | ( n16088 & n16268 ) | ( ~n16089 & n16268 ) ;
  assign n16270 = n36 & n16269 ;
  assign n16271 = n8967 & n16071 ;
  assign n16272 = ( x0 & n8966 ) | ( x0 & ~n16069 ) | ( n8966 & ~n16069 ) ;
  assign n16273 = ( n8966 & n16271 ) | ( n8966 & ~n16272 ) | ( n16271 & ~n16272 ) ;
  assign n16274 = n35 & ~n16067 ;
  assign n16275 = ( n35 & n16273 ) | ( n35 & ~n16274 ) | ( n16273 & ~n16274 ) ;
  assign n16276 = ( ~x2 & n16270 ) | ( ~x2 & n16275 ) | ( n16270 & n16275 ) ;
  assign n16277 = ( n16270 & n16275 ) | ( n16270 & ~n16276 ) | ( n16275 & ~n16276 ) ;
  assign n16278 = ( x2 & n16276 ) | ( x2 & ~n16277 ) | ( n16276 & ~n16277 ) ;
  assign n16279 = ( n16246 & n16267 ) | ( n16246 & n16278 ) | ( n16267 & n16278 ) ;
  assign n16280 = ( n16065 & n16067 ) | ( n16065 & ~n16089 ) | ( n16067 & ~n16089 ) ;
  assign n16281 = ( n16089 & ~n16090 ) | ( n16089 & n16280 ) | ( ~n16090 & n16280 ) ;
  assign n16282 = n36 & n16281 ;
  assign n16283 = n8967 & n16069 ;
  assign n16284 = ( x0 & n8966 ) | ( x0 & ~n16067 ) | ( n8966 & ~n16067 ) ;
  assign n16285 = ( n8966 & n16283 ) | ( n8966 & ~n16284 ) | ( n16283 & ~n16284 ) ;
  assign n16286 = n35 & ~n16065 ;
  assign n16287 = ( n35 & n16285 ) | ( n35 & ~n16286 ) | ( n16285 & ~n16286 ) ;
  assign n16288 = ( ~x2 & n16282 ) | ( ~x2 & n16287 ) | ( n16282 & n16287 ) ;
  assign n16289 = ( n16282 & n16287 ) | ( n16282 & ~n16288 ) | ( n16287 & ~n16288 ) ;
  assign n16290 = ( x2 & n16288 ) | ( x2 & ~n16289 ) | ( n16288 & ~n16289 ) ;
  assign n16291 = n8230 & n16209 ;
  assign n16292 = n8229 & n16071 ;
  assign n16293 = n8226 & ~n16075 ;
  assign n16294 = n8225 & ~n16073 ;
  assign n16295 = n16293 | n16294 ;
  assign n16296 = ( ~n16291 & n16292 ) | ( ~n16291 & n16295 ) | ( n16292 & n16295 ) ;
  assign n16297 = ( ~x5 & n16291 ) | ( ~x5 & n16296 ) | ( n16291 & n16296 ) ;
  assign n16298 = ( n16291 & n16296 ) | ( n16291 & ~n16297 ) | ( n16296 & ~n16297 ) ;
  assign n16299 = ( x5 & n16297 ) | ( x5 & ~n16298 ) | ( n16297 & ~n16298 ) ;
  assign n16300 = ( x8 & n16256 ) | ( x8 & n16262 ) | ( n16256 & n16262 ) ;
  assign n16301 = ( n7296 & n16083 ) | ( n7296 & n16198 ) | ( n16083 & n16198 ) ;
  assign n16302 = n7300 & ~n16081 ;
  assign n16303 = n7299 & ~n16079 ;
  assign n16304 = n16302 | n16303 ;
  assign n16305 = n7879 & ~n16077 ;
  assign n16306 = ( n7879 & n16304 ) | ( n7879 & ~n16305 ) | ( n16304 & ~n16305 ) ;
  assign n16307 = ( ~n16300 & n16301 ) | ( ~n16300 & n16306 ) | ( n16301 & n16306 ) ;
  assign n16308 = ( n16301 & n16306 ) | ( n16301 & ~n16307 ) | ( n16306 & ~n16307 ) ;
  assign n16309 = ( n16300 & n16307 ) | ( n16300 & ~n16308 ) | ( n16307 & ~n16308 ) ;
  assign n16310 = ( n16265 & n16299 ) | ( n16265 & n16309 ) | ( n16299 & n16309 ) ;
  assign n16311 = ( ~n16265 & n16299 ) | ( ~n16265 & n16309 ) | ( n16299 & n16309 ) ;
  assign n16312 = ( n16265 & ~n16310 ) | ( n16265 & n16311 ) | ( ~n16310 & n16311 ) ;
  assign n16313 = ( n16279 & n16290 ) | ( n16279 & n16312 ) | ( n16290 & n16312 ) ;
  assign n16314 = ( n16063 & n16065 ) | ( n16063 & ~n16090 ) | ( n16065 & ~n16090 ) ;
  assign n16315 = ( n16090 & ~n16091 ) | ( n16090 & n16314 ) | ( ~n16091 & n16314 ) ;
  assign n16316 = n36 & n16315 ;
  assign n16317 = n8967 & n16067 ;
  assign n16318 = ( x0 & n8966 ) | ( x0 & ~n16065 ) | ( n8966 & ~n16065 ) ;
  assign n16319 = ( n8966 & n16317 ) | ( n8966 & ~n16318 ) | ( n16317 & ~n16318 ) ;
  assign n16320 = n35 & ~n16063 ;
  assign n16321 = ( n35 & n16319 ) | ( n35 & ~n16320 ) | ( n16319 & ~n16320 ) ;
  assign n16322 = ( ~x2 & n16316 ) | ( ~x2 & n16321 ) | ( n16316 & n16321 ) ;
  assign n16323 = ( n16316 & n16321 ) | ( n16316 & ~n16322 ) | ( n16321 & ~n16322 ) ;
  assign n16324 = ( x2 & n16322 ) | ( x2 & ~n16323 ) | ( n16322 & ~n16323 ) ;
  assign n16325 = n8230 & ~n16221 ;
  assign n16326 = n8229 & n16069 ;
  assign n16327 = n8226 & ~n16073 ;
  assign n16328 = n8225 & n16071 ;
  assign n16329 = n16327 | n16328 ;
  assign n16330 = ( ~n16325 & n16326 ) | ( ~n16325 & n16329 ) | ( n16326 & n16329 ) ;
  assign n16331 = ( ~x5 & n16325 ) | ( ~x5 & n16330 ) | ( n16325 & n16330 ) ;
  assign n16332 = ( n16325 & n16330 ) | ( n16325 & ~n16331 ) | ( n16330 & ~n16331 ) ;
  assign n16333 = ( x5 & n16331 ) | ( x5 & ~n16332 ) | ( n16331 & ~n16332 ) ;
  assign n16334 = x8 & ~n16307 ;
  assign n16335 = ~n16300 & n16334 ;
  assign n16336 = n7021 & ~n16081 ;
  assign n16337 = n7296 & n16169 ;
  assign n16338 = n7879 & ~n16075 ;
  assign n16339 = n7300 & ~n16079 ;
  assign n16340 = n7299 & n16077 ;
  assign n16341 = n16339 | n16340 ;
  assign n16342 = ( ~n16337 & n16338 ) | ( ~n16337 & n16341 ) | ( n16338 & n16341 ) ;
  assign n16343 = ( ~x8 & n16337 ) | ( ~x8 & n16342 ) | ( n16337 & n16342 ) ;
  assign n16344 = ( n16337 & n16342 ) | ( n16337 & ~n16343 ) | ( n16342 & ~n16343 ) ;
  assign n16345 = ( x8 & n16343 ) | ( x8 & ~n16344 ) | ( n16343 & ~n16344 ) ;
  assign n16346 = ( n16335 & n16336 ) | ( n16335 & n16345 ) | ( n16336 & n16345 ) ;
  assign n16347 = ( ~n16335 & n16336 ) | ( ~n16335 & n16345 ) | ( n16336 & n16345 ) ;
  assign n16348 = ( n16335 & ~n16346 ) | ( n16335 & n16347 ) | ( ~n16346 & n16347 ) ;
  assign n16349 = ( n16310 & n16333 ) | ( n16310 & n16348 ) | ( n16333 & n16348 ) ;
  assign n16350 = ( ~n16310 & n16333 ) | ( ~n16310 & n16348 ) | ( n16333 & n16348 ) ;
  assign n16351 = ( n16310 & ~n16349 ) | ( n16310 & n16350 ) | ( ~n16349 & n16350 ) ;
  assign n16352 = ( n16313 & n16324 ) | ( n16313 & n16351 ) | ( n16324 & n16351 ) ;
  assign n16353 = ( n16061 & n16063 ) | ( n16061 & ~n16091 ) | ( n16063 & ~n16091 ) ;
  assign n16354 = ( ~n16063 & n16092 ) | ( ~n16063 & n16353 ) | ( n16092 & n16353 ) ;
  assign n16355 = n36 & ~n16354 ;
  assign n16356 = n8967 & n16065 ;
  assign n16357 = ( x0 & n8966 ) | ( x0 & ~n16063 ) | ( n8966 & ~n16063 ) ;
  assign n16358 = ( n8966 & n16356 ) | ( n8966 & ~n16357 ) | ( n16356 & ~n16357 ) ;
  assign n16359 = n35 & ~n16061 ;
  assign n16360 = n16358 | n16359 ;
  assign n16361 = ( ~x2 & n16355 ) | ( ~x2 & n16360 ) | ( n16355 & n16360 ) ;
  assign n16362 = ( n16355 & n16360 ) | ( n16355 & ~n16361 ) | ( n16360 & ~n16361 ) ;
  assign n16363 = ( x2 & n16361 ) | ( x2 & ~n16362 ) | ( n16361 & ~n16362 ) ;
  assign n16364 = n8230 & n16269 ;
  assign n16365 = n8229 & n16067 ;
  assign n16366 = n8226 & n16071 ;
  assign n16367 = n8225 & n16069 ;
  assign n16368 = n16366 | n16367 ;
  assign n16369 = ( ~n16364 & n16365 ) | ( ~n16364 & n16368 ) | ( n16365 & n16368 ) ;
  assign n16370 = ( ~x5 & n16364 ) | ( ~x5 & n16369 ) | ( n16364 & n16369 ) ;
  assign n16371 = ( n16364 & n16369 ) | ( n16364 & ~n16370 ) | ( n16369 & ~n16370 ) ;
  assign n16372 = ( x5 & n16370 ) | ( x5 & ~n16371 ) | ( n16370 & ~n16371 ) ;
  assign n16373 = n7296 & ~n16176 ;
  assign n16374 = n7879 & ~n16073 ;
  assign n16375 = n7300 & n16077 ;
  assign n16376 = n7299 & ~n16075 ;
  assign n16377 = n16375 | n16376 ;
  assign n16378 = ( ~n16373 & n16374 ) | ( ~n16373 & n16377 ) | ( n16374 & n16377 ) ;
  assign n16379 = ( ~x8 & n16373 ) | ( ~x8 & n16378 ) | ( n16373 & n16378 ) ;
  assign n16380 = ( n16373 & n16378 ) | ( n16373 & ~n16379 ) | ( n16378 & ~n16379 ) ;
  assign n16381 = ( x8 & n16379 ) | ( x8 & ~n16380 ) | ( n16379 & ~n16380 ) ;
  assign n16382 = x11 & n16336 ;
  assign n16383 = ( n6584 & n16155 ) | ( n6584 & n16187 ) | ( n16155 & n16187 ) ;
  assign n16384 = n6587 | n16081 ;
  assign n16385 = n7022 & ~n16079 ;
  assign n16386 = ( ~n16081 & n16384 ) | ( ~n16081 & n16385 ) | ( n16384 & n16385 ) ;
  assign n16387 = ( n16382 & n16383 ) | ( n16382 & n16386 ) | ( n16383 & n16386 ) ;
  assign n16388 = n16383 | n16386 ;
  assign n16389 = ~n16382 & n16388 ;
  assign n16390 = ( n16382 & ~n16387 ) | ( n16382 & n16389 ) | ( ~n16387 & n16389 ) ;
  assign n16391 = ( n16346 & n16381 ) | ( n16346 & n16390 ) | ( n16381 & n16390 ) ;
  assign n16392 = ( ~n16346 & n16381 ) | ( ~n16346 & n16390 ) | ( n16381 & n16390 ) ;
  assign n16393 = ( n16346 & ~n16391 ) | ( n16346 & n16392 ) | ( ~n16391 & n16392 ) ;
  assign n16394 = ( n16349 & n16372 ) | ( n16349 & n16393 ) | ( n16372 & n16393 ) ;
  assign n16395 = ( ~n16349 & n16372 ) | ( ~n16349 & n16393 ) | ( n16372 & n16393 ) ;
  assign n16396 = ( n16349 & ~n16394 ) | ( n16349 & n16395 ) | ( ~n16394 & n16395 ) ;
  assign n16397 = ( n16352 & n16363 ) | ( n16352 & n16396 ) | ( n16363 & n16396 ) ;
  assign n16398 = n7296 & n16209 ;
  assign n16399 = n7879 & n16071 ;
  assign n16400 = n7300 & ~n16075 ;
  assign n16401 = n7299 & ~n16073 ;
  assign n16402 = n16400 | n16401 ;
  assign n16403 = ( ~n16398 & n16399 ) | ( ~n16398 & n16402 ) | ( n16399 & n16402 ) ;
  assign n16404 = ( ~x8 & n16398 ) | ( ~x8 & n16403 ) | ( n16398 & n16403 ) ;
  assign n16405 = ( n16398 & n16403 ) | ( n16398 & ~n16404 ) | ( n16403 & ~n16404 ) ;
  assign n16406 = ( x8 & n16404 ) | ( x8 & ~n16405 ) | ( n16404 & ~n16405 ) ;
  assign n16407 = ( x11 & n16382 ) | ( x11 & n16388 ) | ( n16382 & n16388 ) ;
  assign n16408 = ( n6584 & n16083 ) | ( n6584 & n16198 ) | ( n16083 & n16198 ) ;
  assign n16409 = n6588 & ~n16081 ;
  assign n16410 = n6587 & ~n16079 ;
  assign n16411 = n16409 | n16410 ;
  assign n16412 = n7022 & ~n16077 ;
  assign n16413 = ( n7022 & n16411 ) | ( n7022 & ~n16412 ) | ( n16411 & ~n16412 ) ;
  assign n16414 = ( ~n16407 & n16408 ) | ( ~n16407 & n16413 ) | ( n16408 & n16413 ) ;
  assign n16415 = ( n16408 & n16413 ) | ( n16408 & ~n16414 ) | ( n16413 & ~n16414 ) ;
  assign n16416 = ( n16407 & n16414 ) | ( n16407 & ~n16415 ) | ( n16414 & ~n16415 ) ;
  assign n16417 = ( n16391 & n16406 ) | ( n16391 & n16416 ) | ( n16406 & n16416 ) ;
  assign n16418 = ( ~n16391 & n16406 ) | ( ~n16391 & n16416 ) | ( n16406 & n16416 ) ;
  assign n16419 = ( n16391 & ~n16417 ) | ( n16391 & n16418 ) | ( ~n16417 & n16418 ) ;
  assign n16420 = n8230 & n16281 ;
  assign n16421 = n8229 & n16065 ;
  assign n16422 = n8226 & n16069 ;
  assign n16423 = n8225 & n16067 ;
  assign n16424 = n16422 | n16423 ;
  assign n16425 = ( ~n16420 & n16421 ) | ( ~n16420 & n16424 ) | ( n16421 & n16424 ) ;
  assign n16426 = ( ~x5 & n16420 ) | ( ~x5 & n16425 ) | ( n16420 & n16425 ) ;
  assign n16427 = ( n16420 & n16425 ) | ( n16420 & ~n16426 ) | ( n16425 & ~n16426 ) ;
  assign n16428 = ( x5 & n16426 ) | ( x5 & ~n16427 ) | ( n16426 & ~n16427 ) ;
  assign n16429 = ( n16394 & n16419 ) | ( n16394 & n16428 ) | ( n16419 & n16428 ) ;
  assign n16430 = ( ~n16394 & n16419 ) | ( ~n16394 & n16428 ) | ( n16419 & n16428 ) ;
  assign n16431 = ( n16394 & ~n16429 ) | ( n16394 & n16430 ) | ( ~n16429 & n16430 ) ;
  assign n16432 = ( ~n16059 & n16061 ) | ( ~n16059 & n16092 ) | ( n16061 & n16092 ) ;
  assign n16433 = ( ~n16092 & n16093 ) | ( ~n16092 & n16432 ) | ( n16093 & n16432 ) ;
  assign n16434 = n36 & ~n16433 ;
  assign n16435 = n8967 & n16063 ;
  assign n16436 = n9378 & ~n16061 ;
  assign n16437 = n16435 | n16436 ;
  assign n16438 = n35 & ~n16059 ;
  assign n16439 = ( n35 & n16437 ) | ( n35 & ~n16438 ) | ( n16437 & ~n16438 ) ;
  assign n16440 = ( ~x2 & n16434 ) | ( ~x2 & n16439 ) | ( n16434 & n16439 ) ;
  assign n16441 = ( n16434 & n16439 ) | ( n16434 & ~n16440 ) | ( n16439 & ~n16440 ) ;
  assign n16442 = ( x2 & n16440 ) | ( x2 & ~n16441 ) | ( n16440 & ~n16441 ) ;
  assign n16443 = ( n16397 & n16431 ) | ( n16397 & n16442 ) | ( n16431 & n16442 ) ;
  assign n16444 = n7296 & ~n16221 ;
  assign n16445 = n7879 & n16069 ;
  assign n16446 = n7300 & ~n16073 ;
  assign n16447 = n7299 & n16071 ;
  assign n16448 = n16446 | n16447 ;
  assign n16449 = ( ~n16444 & n16445 ) | ( ~n16444 & n16448 ) | ( n16445 & n16448 ) ;
  assign n16450 = ( ~x8 & n16444 ) | ( ~x8 & n16449 ) | ( n16444 & n16449 ) ;
  assign n16451 = ( n16444 & n16449 ) | ( n16444 & ~n16450 ) | ( n16449 & ~n16450 ) ;
  assign n16452 = ( x8 & n16450 ) | ( x8 & ~n16451 ) | ( n16450 & ~n16451 ) ;
  assign n16453 = x11 & ~n16414 ;
  assign n16454 = ~n16407 & n16453 ;
  assign n16455 = n6463 & ~n16081 ;
  assign n16456 = n6584 & n16169 ;
  assign n16457 = n7022 & ~n16075 ;
  assign n16458 = n6588 & ~n16079 ;
  assign n16459 = n6587 & n16077 ;
  assign n16460 = n16458 | n16459 ;
  assign n16461 = ( ~n16456 & n16457 ) | ( ~n16456 & n16460 ) | ( n16457 & n16460 ) ;
  assign n16462 = ( ~x11 & n16456 ) | ( ~x11 & n16461 ) | ( n16456 & n16461 ) ;
  assign n16463 = ( n16456 & n16461 ) | ( n16456 & ~n16462 ) | ( n16461 & ~n16462 ) ;
  assign n16464 = ( x11 & n16462 ) | ( x11 & ~n16463 ) | ( n16462 & ~n16463 ) ;
  assign n16465 = ( n16454 & n16455 ) | ( n16454 & n16464 ) | ( n16455 & n16464 ) ;
  assign n16466 = ( ~n16454 & n16455 ) | ( ~n16454 & n16464 ) | ( n16455 & n16464 ) ;
  assign n16467 = ( n16454 & ~n16465 ) | ( n16454 & n16466 ) | ( ~n16465 & n16466 ) ;
  assign n16468 = ( n16417 & n16452 ) | ( n16417 & n16467 ) | ( n16452 & n16467 ) ;
  assign n16469 = ( ~n16417 & n16452 ) | ( ~n16417 & n16467 ) | ( n16452 & n16467 ) ;
  assign n16470 = ( n16417 & ~n16468 ) | ( n16417 & n16469 ) | ( ~n16468 & n16469 ) ;
  assign n16471 = n8230 & n16315 ;
  assign n16472 = n8229 & n16063 ;
  assign n16473 = n8226 & n16067 ;
  assign n16474 = n8225 & n16065 ;
  assign n16475 = n16473 | n16474 ;
  assign n16476 = ( ~n16471 & n16472 ) | ( ~n16471 & n16475 ) | ( n16472 & n16475 ) ;
  assign n16477 = ( ~x5 & n16471 ) | ( ~x5 & n16476 ) | ( n16471 & n16476 ) ;
  assign n16478 = ( n16471 & n16476 ) | ( n16471 & ~n16477 ) | ( n16476 & ~n16477 ) ;
  assign n16479 = ( x5 & n16477 ) | ( x5 & ~n16478 ) | ( n16477 & ~n16478 ) ;
  assign n16480 = ( n16429 & n16470 ) | ( n16429 & n16479 ) | ( n16470 & n16479 ) ;
  assign n16481 = ( ~n16429 & n16470 ) | ( ~n16429 & n16479 ) | ( n16470 & n16479 ) ;
  assign n16482 = ( n16429 & ~n16480 ) | ( n16429 & n16481 ) | ( ~n16480 & n16481 ) ;
  assign n16483 = ( n16057 & ~n16059 ) | ( n16057 & n16093 ) | ( ~n16059 & n16093 ) ;
  assign n16484 = ( ~n16093 & n16094 ) | ( ~n16093 & n16483 ) | ( n16094 & n16483 ) ;
  assign n16485 = n36 & ~n16484 ;
  assign n16486 = n8967 & ~n16061 ;
  assign n16487 = ( x0 & n8966 ) | ( x0 & ~n16059 ) | ( n8966 & ~n16059 ) ;
  assign n16488 = ( n8966 & n16486 ) | ( n8966 & ~n16487 ) | ( n16486 & ~n16487 ) ;
  assign n16489 = n35 & n16057 ;
  assign n16490 = ( n35 & n16488 ) | ( n35 & ~n16489 ) | ( n16488 & ~n16489 ) ;
  assign n16491 = ( ~x2 & n16485 ) | ( ~x2 & n16490 ) | ( n16485 & n16490 ) ;
  assign n16492 = ( n16485 & n16490 ) | ( n16485 & ~n16491 ) | ( n16490 & ~n16491 ) ;
  assign n16493 = ( x2 & n16491 ) | ( x2 & ~n16492 ) | ( n16491 & ~n16492 ) ;
  assign n16494 = ( n16443 & n16482 ) | ( n16443 & n16493 ) | ( n16482 & n16493 ) ;
  assign n16495 = n7296 & n16269 ;
  assign n16496 = n7879 & n16067 ;
  assign n16497 = n7300 & n16071 ;
  assign n16498 = n7299 & n16069 ;
  assign n16499 = n16497 | n16498 ;
  assign n16500 = ( ~n16495 & n16496 ) | ( ~n16495 & n16499 ) | ( n16496 & n16499 ) ;
  assign n16501 = ( ~x8 & n16495 ) | ( ~x8 & n16500 ) | ( n16495 & n16500 ) ;
  assign n16502 = ( n16495 & n16500 ) | ( n16495 & ~n16501 ) | ( n16500 & ~n16501 ) ;
  assign n16503 = ( x8 & n16501 ) | ( x8 & ~n16502 ) | ( n16501 & ~n16502 ) ;
  assign n16504 = n6584 & ~n16176 ;
  assign n16505 = n7022 & ~n16073 ;
  assign n16506 = n6588 & n16077 ;
  assign n16507 = n6587 & ~n16075 ;
  assign n16508 = n16506 | n16507 ;
  assign n16509 = ( ~n16504 & n16505 ) | ( ~n16504 & n16508 ) | ( n16505 & n16508 ) ;
  assign n16510 = ( ~x11 & n16504 ) | ( ~x11 & n16509 ) | ( n16504 & n16509 ) ;
  assign n16511 = ( n16504 & n16509 ) | ( n16504 & ~n16510 ) | ( n16509 & ~n16510 ) ;
  assign n16512 = ( x11 & n16510 ) | ( x11 & ~n16511 ) | ( n16510 & ~n16511 ) ;
  assign n16513 = x14 & n16455 ;
  assign n16514 = ( n5966 & n16155 ) | ( n5966 & n16187 ) | ( n16155 & n16187 ) ;
  assign n16515 = n5969 | n16081 ;
  assign n16516 = n6464 & ~n16079 ;
  assign n16517 = ( ~n16081 & n16515 ) | ( ~n16081 & n16516 ) | ( n16515 & n16516 ) ;
  assign n16518 = ( n16513 & n16514 ) | ( n16513 & n16517 ) | ( n16514 & n16517 ) ;
  assign n16519 = n16514 | n16517 ;
  assign n16520 = ~n16513 & n16519 ;
  assign n16521 = ( n16513 & ~n16518 ) | ( n16513 & n16520 ) | ( ~n16518 & n16520 ) ;
  assign n16522 = ( n16465 & n16512 ) | ( n16465 & n16521 ) | ( n16512 & n16521 ) ;
  assign n16523 = ( ~n16465 & n16512 ) | ( ~n16465 & n16521 ) | ( n16512 & n16521 ) ;
  assign n16524 = ( n16465 & ~n16522 ) | ( n16465 & n16523 ) | ( ~n16522 & n16523 ) ;
  assign n16525 = ( n16468 & n16503 ) | ( n16468 & n16524 ) | ( n16503 & n16524 ) ;
  assign n16526 = ( ~n16468 & n16503 ) | ( ~n16468 & n16524 ) | ( n16503 & n16524 ) ;
  assign n16527 = ( n16468 & ~n16525 ) | ( n16468 & n16526 ) | ( ~n16525 & n16526 ) ;
  assign n16528 = n8230 & ~n16354 ;
  assign n16529 = n8229 & ~n16061 ;
  assign n16530 = n8226 & n16065 ;
  assign n16531 = n8225 & n16063 ;
  assign n16532 = n16530 | n16531 ;
  assign n16533 = ( ~n16528 & n16529 ) | ( ~n16528 & n16532 ) | ( n16529 & n16532 ) ;
  assign n16534 = ( ~x5 & n16528 ) | ( ~x5 & n16533 ) | ( n16528 & n16533 ) ;
  assign n16535 = ( n16528 & n16533 ) | ( n16528 & ~n16534 ) | ( n16533 & ~n16534 ) ;
  assign n16536 = ( x5 & n16534 ) | ( x5 & ~n16535 ) | ( n16534 & ~n16535 ) ;
  assign n16537 = ( n16480 & n16527 ) | ( n16480 & n16536 ) | ( n16527 & n16536 ) ;
  assign n16538 = ( ~n16480 & n16527 ) | ( ~n16480 & n16536 ) | ( n16527 & n16536 ) ;
  assign n16539 = ( n16480 & ~n16537 ) | ( n16480 & n16538 ) | ( ~n16537 & n16538 ) ;
  assign n16540 = ( n16055 & n16057 ) | ( n16055 & ~n16095 ) | ( n16057 & ~n16095 ) ;
  assign n16541 = ( n16094 & n16095 ) | ( n16094 & ~n16540 ) | ( n16095 & ~n16540 ) ;
  assign n16542 = n36 & n16541 ;
  assign n16543 = n8967 & n16059 ;
  assign n16544 = ( x0 & n8966 ) | ( x0 & n16057 ) | ( n8966 & n16057 ) ;
  assign n16545 = ( n8966 & n16543 ) | ( n8966 & ~n16544 ) | ( n16543 & ~n16544 ) ;
  assign n16546 = n35 & n16055 ;
  assign n16547 = ( n35 & n16545 ) | ( n35 & ~n16546 ) | ( n16545 & ~n16546 ) ;
  assign n16548 = ( ~x2 & n16542 ) | ( ~x2 & n16547 ) | ( n16542 & n16547 ) ;
  assign n16549 = ( n16542 & n16547 ) | ( n16542 & ~n16548 ) | ( n16547 & ~n16548 ) ;
  assign n16550 = ( x2 & n16548 ) | ( x2 & ~n16549 ) | ( n16548 & ~n16549 ) ;
  assign n16551 = ( n16494 & n16539 ) | ( n16494 & n16550 ) | ( n16539 & n16550 ) ;
  assign n16552 = ( n16053 & n16055 ) | ( n16053 & ~n16095 ) | ( n16055 & ~n16095 ) ;
  assign n16553 = ( ~n16055 & n16096 ) | ( ~n16055 & n16552 ) | ( n16096 & n16552 ) ;
  assign n16554 = n36 & n16553 ;
  assign n16555 = n8967 & ~n16057 ;
  assign n16556 = ( x0 & n8966 ) | ( x0 & n16055 ) | ( n8966 & n16055 ) ;
  assign n16557 = ( n8966 & n16555 ) | ( n8966 & ~n16556 ) | ( n16555 & ~n16556 ) ;
  assign n16558 = n35 & ~n16053 ;
  assign n16559 = ( n35 & n16557 ) | ( n35 & ~n16558 ) | ( n16557 & ~n16558 ) ;
  assign n16560 = ( ~x2 & n16554 ) | ( ~x2 & n16559 ) | ( n16554 & n16559 ) ;
  assign n16561 = ( n16554 & n16559 ) | ( n16554 & ~n16560 ) | ( n16559 & ~n16560 ) ;
  assign n16562 = ( x2 & n16560 ) | ( x2 & ~n16561 ) | ( n16560 & ~n16561 ) ;
  assign n16563 = n8230 & ~n16433 ;
  assign n16564 = n8229 & n16059 ;
  assign n16565 = n8226 & n16063 ;
  assign n16566 = n8225 & ~n16061 ;
  assign n16567 = n16565 | n16566 ;
  assign n16568 = ( ~n16563 & n16564 ) | ( ~n16563 & n16567 ) | ( n16564 & n16567 ) ;
  assign n16569 = ( ~x5 & n16563 ) | ( ~x5 & n16568 ) | ( n16563 & n16568 ) ;
  assign n16570 = ( n16563 & n16568 ) | ( n16563 & ~n16569 ) | ( n16568 & ~n16569 ) ;
  assign n16571 = ( x5 & n16569 ) | ( x5 & ~n16570 ) | ( n16569 & ~n16570 ) ;
  assign n16572 = n6584 & n16209 ;
  assign n16573 = n7022 & n16071 ;
  assign n16574 = n6588 & ~n16075 ;
  assign n16575 = n6587 & ~n16073 ;
  assign n16576 = n16574 | n16575 ;
  assign n16577 = ( ~n16572 & n16573 ) | ( ~n16572 & n16576 ) | ( n16573 & n16576 ) ;
  assign n16578 = ( ~x11 & n16572 ) | ( ~x11 & n16577 ) | ( n16572 & n16577 ) ;
  assign n16579 = ( n16572 & n16577 ) | ( n16572 & ~n16578 ) | ( n16577 & ~n16578 ) ;
  assign n16580 = ( x11 & n16578 ) | ( x11 & ~n16579 ) | ( n16578 & ~n16579 ) ;
  assign n16581 = ( x14 & n16513 ) | ( x14 & n16519 ) | ( n16513 & n16519 ) ;
  assign n16582 = ( n5966 & n16083 ) | ( n5966 & n16198 ) | ( n16083 & n16198 ) ;
  assign n16583 = n5970 & ~n16081 ;
  assign n16584 = n5969 & ~n16079 ;
  assign n16585 = n16583 | n16584 ;
  assign n16586 = n6464 & ~n16077 ;
  assign n16587 = ( n6464 & n16585 ) | ( n6464 & ~n16586 ) | ( n16585 & ~n16586 ) ;
  assign n16588 = ( ~n16581 & n16582 ) | ( ~n16581 & n16587 ) | ( n16582 & n16587 ) ;
  assign n16589 = ( n16582 & n16587 ) | ( n16582 & ~n16588 ) | ( n16587 & ~n16588 ) ;
  assign n16590 = ( n16581 & n16588 ) | ( n16581 & ~n16589 ) | ( n16588 & ~n16589 ) ;
  assign n16591 = ( n16522 & n16580 ) | ( n16522 & n16590 ) | ( n16580 & n16590 ) ;
  assign n16592 = ( ~n16522 & n16580 ) | ( ~n16522 & n16590 ) | ( n16580 & n16590 ) ;
  assign n16593 = ( n16522 & ~n16591 ) | ( n16522 & n16592 ) | ( ~n16591 & n16592 ) ;
  assign n16594 = n7296 & n16281 ;
  assign n16595 = n7879 & n16065 ;
  assign n16596 = n7300 & n16069 ;
  assign n16597 = n7299 & n16067 ;
  assign n16598 = n16596 | n16597 ;
  assign n16599 = ( ~n16594 & n16595 ) | ( ~n16594 & n16598 ) | ( n16595 & n16598 ) ;
  assign n16600 = ( ~x8 & n16594 ) | ( ~x8 & n16599 ) | ( n16594 & n16599 ) ;
  assign n16601 = ( n16594 & n16599 ) | ( n16594 & ~n16600 ) | ( n16599 & ~n16600 ) ;
  assign n16602 = ( x8 & n16600 ) | ( x8 & ~n16601 ) | ( n16600 & ~n16601 ) ;
  assign n16603 = ( n16525 & n16593 ) | ( n16525 & n16602 ) | ( n16593 & n16602 ) ;
  assign n16604 = ( ~n16525 & n16593 ) | ( ~n16525 & n16602 ) | ( n16593 & n16602 ) ;
  assign n16605 = ( n16525 & ~n16603 ) | ( n16525 & n16604 ) | ( ~n16603 & n16604 ) ;
  assign n16606 = ( n16537 & n16571 ) | ( n16537 & n16605 ) | ( n16571 & n16605 ) ;
  assign n16607 = ( ~n16537 & n16571 ) | ( ~n16537 & n16605 ) | ( n16571 & n16605 ) ;
  assign n16608 = ( n16537 & ~n16606 ) | ( n16537 & n16607 ) | ( ~n16606 & n16607 ) ;
  assign n16609 = ( n16551 & n16562 ) | ( n16551 & n16608 ) | ( n16562 & n16608 ) ;
  assign n16610 = ( ~n16051 & n16053 ) | ( ~n16051 & n16096 ) | ( n16053 & n16096 ) ;
  assign n16611 = ( ~n16096 & n16097 ) | ( ~n16096 & n16610 ) | ( n16097 & n16610 ) ;
  assign n16612 = n36 & n16611 ;
  assign n16613 = n8967 & ~n16055 ;
  assign n16614 = ( x0 & n8966 ) | ( x0 & ~n16053 ) | ( n8966 & ~n16053 ) ;
  assign n16615 = ( n8966 & n16613 ) | ( n8966 & ~n16614 ) | ( n16613 & ~n16614 ) ;
  assign n16616 = n35 & n16051 ;
  assign n16617 = ( n35 & n16615 ) | ( n35 & ~n16616 ) | ( n16615 & ~n16616 ) ;
  assign n16618 = ( ~x2 & n16612 ) | ( ~x2 & n16617 ) | ( n16612 & n16617 ) ;
  assign n16619 = ( n16612 & n16617 ) | ( n16612 & ~n16618 ) | ( n16617 & ~n16618 ) ;
  assign n16620 = ( x2 & n16618 ) | ( x2 & ~n16619 ) | ( n16618 & ~n16619 ) ;
  assign n16621 = n8230 & ~n16484 ;
  assign n16622 = n8229 & ~n16057 ;
  assign n16623 = n8226 & ~n16061 ;
  assign n16624 = n8225 & n16059 ;
  assign n16625 = n16623 | n16624 ;
  assign n16626 = ( ~n16621 & n16622 ) | ( ~n16621 & n16625 ) | ( n16622 & n16625 ) ;
  assign n16627 = ( ~x5 & n16621 ) | ( ~x5 & n16626 ) | ( n16621 & n16626 ) ;
  assign n16628 = ( n16621 & n16626 ) | ( n16621 & ~n16627 ) | ( n16626 & ~n16627 ) ;
  assign n16629 = ( x5 & n16627 ) | ( x5 & ~n16628 ) | ( n16627 & ~n16628 ) ;
  assign n16630 = n6584 & ~n16221 ;
  assign n16631 = n7022 & n16069 ;
  assign n16632 = n6588 & ~n16073 ;
  assign n16633 = n6587 & n16071 ;
  assign n16634 = n16632 | n16633 ;
  assign n16635 = ( ~n16630 & n16631 ) | ( ~n16630 & n16634 ) | ( n16631 & n16634 ) ;
  assign n16636 = ( ~x11 & n16630 ) | ( ~x11 & n16635 ) | ( n16630 & n16635 ) ;
  assign n16637 = ( n16630 & n16635 ) | ( n16630 & ~n16636 ) | ( n16635 & ~n16636 ) ;
  assign n16638 = ( x11 & n16636 ) | ( x11 & ~n16637 ) | ( n16636 & ~n16637 ) ;
  assign n16639 = x14 & ~n16588 ;
  assign n16640 = ~n16581 & n16639 ;
  assign n16641 = n5506 & ~n16081 ;
  assign n16642 = n5966 & n16169 ;
  assign n16643 = n6464 & ~n16075 ;
  assign n16644 = n5970 & ~n16079 ;
  assign n16645 = n5969 & n16077 ;
  assign n16646 = n16644 | n16645 ;
  assign n16647 = ( ~n16642 & n16643 ) | ( ~n16642 & n16646 ) | ( n16643 & n16646 ) ;
  assign n16648 = ( ~x14 & n16642 ) | ( ~x14 & n16647 ) | ( n16642 & n16647 ) ;
  assign n16649 = ( n16642 & n16647 ) | ( n16642 & ~n16648 ) | ( n16647 & ~n16648 ) ;
  assign n16650 = ( x14 & n16648 ) | ( x14 & ~n16649 ) | ( n16648 & ~n16649 ) ;
  assign n16651 = ( n16640 & n16641 ) | ( n16640 & n16650 ) | ( n16641 & n16650 ) ;
  assign n16652 = ( ~n16640 & n16641 ) | ( ~n16640 & n16650 ) | ( n16641 & n16650 ) ;
  assign n16653 = ( n16640 & ~n16651 ) | ( n16640 & n16652 ) | ( ~n16651 & n16652 ) ;
  assign n16654 = ( n16591 & n16638 ) | ( n16591 & n16653 ) | ( n16638 & n16653 ) ;
  assign n16655 = ( ~n16591 & n16638 ) | ( ~n16591 & n16653 ) | ( n16638 & n16653 ) ;
  assign n16656 = ( n16591 & ~n16654 ) | ( n16591 & n16655 ) | ( ~n16654 & n16655 ) ;
  assign n16657 = n7296 & n16315 ;
  assign n16658 = n7879 & n16063 ;
  assign n16659 = n7300 & n16067 ;
  assign n16660 = n7299 & n16065 ;
  assign n16661 = n16659 | n16660 ;
  assign n16662 = ( ~n16657 & n16658 ) | ( ~n16657 & n16661 ) | ( n16658 & n16661 ) ;
  assign n16663 = ( ~x8 & n16657 ) | ( ~x8 & n16662 ) | ( n16657 & n16662 ) ;
  assign n16664 = ( n16657 & n16662 ) | ( n16657 & ~n16663 ) | ( n16662 & ~n16663 ) ;
  assign n16665 = ( x8 & n16663 ) | ( x8 & ~n16664 ) | ( n16663 & ~n16664 ) ;
  assign n16666 = ( n16603 & n16656 ) | ( n16603 & n16665 ) | ( n16656 & n16665 ) ;
  assign n16667 = ( ~n16603 & n16656 ) | ( ~n16603 & n16665 ) | ( n16656 & n16665 ) ;
  assign n16668 = ( n16603 & ~n16666 ) | ( n16603 & n16667 ) | ( ~n16666 & n16667 ) ;
  assign n16669 = ( n16606 & n16629 ) | ( n16606 & n16668 ) | ( n16629 & n16668 ) ;
  assign n16670 = ( ~n16606 & n16629 ) | ( ~n16606 & n16668 ) | ( n16629 & n16668 ) ;
  assign n16671 = ( n16606 & ~n16669 ) | ( n16606 & n16670 ) | ( ~n16669 & n16670 ) ;
  assign n16672 = ( n16609 & n16620 ) | ( n16609 & n16671 ) | ( n16620 & n16671 ) ;
  assign n16673 = ( n16049 & ~n16051 ) | ( n16049 & n16097 ) | ( ~n16051 & n16097 ) ;
  assign n16674 = ( n16051 & ~n16098 ) | ( n16051 & n16673 ) | ( ~n16098 & n16673 ) ;
  assign n16675 = n36 & ~n16674 ;
  assign n16676 = n8967 & n16053 ;
  assign n16677 = ( x0 & n8966 ) | ( x0 & n16051 ) | ( n8966 & n16051 ) ;
  assign n16678 = ( n8966 & n16676 ) | ( n8966 & ~n16677 ) | ( n16676 & ~n16677 ) ;
  assign n16679 = n35 & n16049 ;
  assign n16680 = ( n35 & n16678 ) | ( n35 & ~n16679 ) | ( n16678 & ~n16679 ) ;
  assign n16681 = ( ~x2 & n16675 ) | ( ~x2 & n16680 ) | ( n16675 & n16680 ) ;
  assign n16682 = ( n16675 & n16680 ) | ( n16675 & ~n16681 ) | ( n16680 & ~n16681 ) ;
  assign n16683 = ( x2 & n16681 ) | ( x2 & ~n16682 ) | ( n16681 & ~n16682 ) ;
  assign n16684 = n8230 & n16541 ;
  assign n16685 = n8229 & ~n16055 ;
  assign n16686 = n8226 & n16059 ;
  assign n16687 = n8225 & ~n16057 ;
  assign n16688 = n16686 | n16687 ;
  assign n16689 = ( ~n16684 & n16685 ) | ( ~n16684 & n16688 ) | ( n16685 & n16688 ) ;
  assign n16690 = ( ~x5 & n16684 ) | ( ~x5 & n16689 ) | ( n16684 & n16689 ) ;
  assign n16691 = ( n16684 & n16689 ) | ( n16684 & ~n16690 ) | ( n16689 & ~n16690 ) ;
  assign n16692 = ( x5 & n16690 ) | ( x5 & ~n16691 ) | ( n16690 & ~n16691 ) ;
  assign n16693 = n6584 & n16269 ;
  assign n16694 = n7022 & n16067 ;
  assign n16695 = n6588 & n16071 ;
  assign n16696 = n6587 & n16069 ;
  assign n16697 = n16695 | n16696 ;
  assign n16698 = ( ~n16693 & n16694 ) | ( ~n16693 & n16697 ) | ( n16694 & n16697 ) ;
  assign n16699 = ( ~x11 & n16693 ) | ( ~x11 & n16698 ) | ( n16693 & n16698 ) ;
  assign n16700 = ( n16693 & n16698 ) | ( n16693 & ~n16699 ) | ( n16698 & ~n16699 ) ;
  assign n16701 = ( x11 & n16699 ) | ( x11 & ~n16700 ) | ( n16699 & ~n16700 ) ;
  assign n16702 = n5966 & ~n16176 ;
  assign n16703 = n6464 & ~n16073 ;
  assign n16704 = n5970 & n16077 ;
  assign n16705 = n5969 & ~n16075 ;
  assign n16706 = n16704 | n16705 ;
  assign n16707 = ( ~n16702 & n16703 ) | ( ~n16702 & n16706 ) | ( n16703 & n16706 ) ;
  assign n16708 = ( ~x14 & n16702 ) | ( ~x14 & n16707 ) | ( n16702 & n16707 ) ;
  assign n16709 = ( n16702 & n16707 ) | ( n16702 & ~n16708 ) | ( n16707 & ~n16708 ) ;
  assign n16710 = ( x14 & n16708 ) | ( x14 & ~n16709 ) | ( n16708 & ~n16709 ) ;
  assign n16711 = x17 & n16641 ;
  assign n16712 = ( n5508 & n16155 ) | ( n5508 & n16187 ) | ( n16155 & n16187 ) ;
  assign n16713 = n5666 | n16081 ;
  assign n16714 = n5507 & ~n16079 ;
  assign n16715 = ( ~n16081 & n16713 ) | ( ~n16081 & n16714 ) | ( n16713 & n16714 ) ;
  assign n16716 = ( n16711 & n16712 ) | ( n16711 & n16715 ) | ( n16712 & n16715 ) ;
  assign n16717 = n16712 | n16715 ;
  assign n16718 = ~n16711 & n16717 ;
  assign n16719 = ( n16711 & ~n16716 ) | ( n16711 & n16718 ) | ( ~n16716 & n16718 ) ;
  assign n16720 = ( n16651 & n16710 ) | ( n16651 & n16719 ) | ( n16710 & n16719 ) ;
  assign n16721 = ( ~n16651 & n16710 ) | ( ~n16651 & n16719 ) | ( n16710 & n16719 ) ;
  assign n16722 = ( n16651 & ~n16720 ) | ( n16651 & n16721 ) | ( ~n16720 & n16721 ) ;
  assign n16723 = ( n16654 & n16701 ) | ( n16654 & n16722 ) | ( n16701 & n16722 ) ;
  assign n16724 = ( ~n16654 & n16701 ) | ( ~n16654 & n16722 ) | ( n16701 & n16722 ) ;
  assign n16725 = ( n16654 & ~n16723 ) | ( n16654 & n16724 ) | ( ~n16723 & n16724 ) ;
  assign n16726 = n7296 & ~n16354 ;
  assign n16727 = n7879 & ~n16061 ;
  assign n16728 = n7300 & n16065 ;
  assign n16729 = n7299 & n16063 ;
  assign n16730 = n16728 | n16729 ;
  assign n16731 = ( ~n16726 & n16727 ) | ( ~n16726 & n16730 ) | ( n16727 & n16730 ) ;
  assign n16732 = ( ~x8 & n16726 ) | ( ~x8 & n16731 ) | ( n16726 & n16731 ) ;
  assign n16733 = ( n16726 & n16731 ) | ( n16726 & ~n16732 ) | ( n16731 & ~n16732 ) ;
  assign n16734 = ( x8 & n16732 ) | ( x8 & ~n16733 ) | ( n16732 & ~n16733 ) ;
  assign n16735 = ( n16666 & n16725 ) | ( n16666 & n16734 ) | ( n16725 & n16734 ) ;
  assign n16736 = ( ~n16666 & n16725 ) | ( ~n16666 & n16734 ) | ( n16725 & n16734 ) ;
  assign n16737 = ( n16666 & ~n16735 ) | ( n16666 & n16736 ) | ( ~n16735 & n16736 ) ;
  assign n16738 = ( n16669 & n16692 ) | ( n16669 & n16737 ) | ( n16692 & n16737 ) ;
  assign n16739 = ( ~n16669 & n16692 ) | ( ~n16669 & n16737 ) | ( n16692 & n16737 ) ;
  assign n16740 = ( n16669 & ~n16738 ) | ( n16669 & n16739 ) | ( ~n16738 & n16739 ) ;
  assign n16741 = ( n16672 & n16683 ) | ( n16672 & n16740 ) | ( n16683 & n16740 ) ;
  assign n16742 = n7296 & ~n16433 ;
  assign n16743 = n7879 & n16059 ;
  assign n16744 = n7300 & n16063 ;
  assign n16745 = n7299 & ~n16061 ;
  assign n16746 = n16744 | n16745 ;
  assign n16747 = ( ~n16742 & n16743 ) | ( ~n16742 & n16746 ) | ( n16743 & n16746 ) ;
  assign n16748 = ( ~x8 & n16742 ) | ( ~x8 & n16747 ) | ( n16742 & n16747 ) ;
  assign n16749 = ( n16742 & n16747 ) | ( n16742 & ~n16748 ) | ( n16747 & ~n16748 ) ;
  assign n16750 = ( x8 & n16748 ) | ( x8 & ~n16749 ) | ( n16748 & ~n16749 ) ;
  assign n16751 = n5966 & n16209 ;
  assign n16752 = n6464 & n16071 ;
  assign n16753 = n5970 & ~n16075 ;
  assign n16754 = n5969 & ~n16073 ;
  assign n16755 = n16753 | n16754 ;
  assign n16756 = ( ~n16751 & n16752 ) | ( ~n16751 & n16755 ) | ( n16752 & n16755 ) ;
  assign n16757 = ( ~x14 & n16751 ) | ( ~x14 & n16756 ) | ( n16751 & n16756 ) ;
  assign n16758 = ( n16751 & n16756 ) | ( n16751 & ~n16757 ) | ( n16756 & ~n16757 ) ;
  assign n16759 = ( x14 & n16757 ) | ( x14 & ~n16758 ) | ( n16757 & ~n16758 ) ;
  assign n16760 = ( x17 & n16711 ) | ( x17 & n16717 ) | ( n16711 & n16717 ) ;
  assign n16761 = ( n5508 & n16083 ) | ( n5508 & n16198 ) | ( n16083 & n16198 ) ;
  assign n16762 = n5504 & ~n16081 ;
  assign n16763 = n5666 & ~n16079 ;
  assign n16764 = n16762 | n16763 ;
  assign n16765 = n5507 & ~n16077 ;
  assign n16766 = ( n5507 & n16764 ) | ( n5507 & ~n16765 ) | ( n16764 & ~n16765 ) ;
  assign n16767 = ( ~n16760 & n16761 ) | ( ~n16760 & n16766 ) | ( n16761 & n16766 ) ;
  assign n16768 = ( n16761 & n16766 ) | ( n16761 & ~n16767 ) | ( n16766 & ~n16767 ) ;
  assign n16769 = ( n16760 & n16767 ) | ( n16760 & ~n16768 ) | ( n16767 & ~n16768 ) ;
  assign n16770 = ( n16720 & n16759 ) | ( n16720 & n16769 ) | ( n16759 & n16769 ) ;
  assign n16771 = ( ~n16720 & n16759 ) | ( ~n16720 & n16769 ) | ( n16759 & n16769 ) ;
  assign n16772 = ( n16720 & ~n16770 ) | ( n16720 & n16771 ) | ( ~n16770 & n16771 ) ;
  assign n16773 = n6584 & n16281 ;
  assign n16774 = n7022 & n16065 ;
  assign n16775 = n6588 & n16069 ;
  assign n16776 = n6587 & n16067 ;
  assign n16777 = n16775 | n16776 ;
  assign n16778 = ( ~n16773 & n16774 ) | ( ~n16773 & n16777 ) | ( n16774 & n16777 ) ;
  assign n16779 = ( ~x11 & n16773 ) | ( ~x11 & n16778 ) | ( n16773 & n16778 ) ;
  assign n16780 = ( n16773 & n16778 ) | ( n16773 & ~n16779 ) | ( n16778 & ~n16779 ) ;
  assign n16781 = ( x11 & n16779 ) | ( x11 & ~n16780 ) | ( n16779 & ~n16780 ) ;
  assign n16782 = ( n16723 & n16772 ) | ( n16723 & n16781 ) | ( n16772 & n16781 ) ;
  assign n16783 = ( ~n16723 & n16772 ) | ( ~n16723 & n16781 ) | ( n16772 & n16781 ) ;
  assign n16784 = ( n16723 & ~n16782 ) | ( n16723 & n16783 ) | ( ~n16782 & n16783 ) ;
  assign n16785 = ( n16735 & n16750 ) | ( n16735 & n16784 ) | ( n16750 & n16784 ) ;
  assign n16786 = ( ~n16735 & n16750 ) | ( ~n16735 & n16784 ) | ( n16750 & n16784 ) ;
  assign n16787 = ( n16735 & ~n16785 ) | ( n16735 & n16786 ) | ( ~n16785 & n16786 ) ;
  assign n16788 = n8230 & n16553 ;
  assign n16789 = n8229 & n16053 ;
  assign n16790 = n8226 & ~n16057 ;
  assign n16791 = n8225 & ~n16055 ;
  assign n16792 = n16790 | n16791 ;
  assign n16793 = ( ~n16788 & n16789 ) | ( ~n16788 & n16792 ) | ( n16789 & n16792 ) ;
  assign n16794 = ( ~x5 & n16788 ) | ( ~x5 & n16793 ) | ( n16788 & n16793 ) ;
  assign n16795 = ( n16788 & n16793 ) | ( n16788 & ~n16794 ) | ( n16793 & ~n16794 ) ;
  assign n16796 = ( x5 & n16794 ) | ( x5 & ~n16795 ) | ( n16794 & ~n16795 ) ;
  assign n16797 = ( n16738 & n16787 ) | ( n16738 & n16796 ) | ( n16787 & n16796 ) ;
  assign n16798 = ( ~n16738 & n16787 ) | ( ~n16738 & n16796 ) | ( n16787 & n16796 ) ;
  assign n16799 = ( n16738 & ~n16797 ) | ( n16738 & n16798 ) | ( ~n16797 & n16798 ) ;
  assign n16800 = ( n16047 & ~n16049 ) | ( n16047 & n16098 ) | ( ~n16049 & n16098 ) ;
  assign n16801 = ( n16049 & ~n16099 ) | ( n16049 & n16800 ) | ( ~n16099 & n16800 ) ;
  assign n16802 = n36 & ~n16801 ;
  assign n16803 = n8967 & ~n16051 ;
  assign n16804 = ( x0 & n8966 ) | ( x0 & n16049 ) | ( n8966 & n16049 ) ;
  assign n16805 = ( n8966 & n16803 ) | ( n8966 & ~n16804 ) | ( n16803 & ~n16804 ) ;
  assign n16806 = n35 & n16047 ;
  assign n16807 = ( n35 & n16805 ) | ( n35 & ~n16806 ) | ( n16805 & ~n16806 ) ;
  assign n16808 = ( ~x2 & n16802 ) | ( ~x2 & n16807 ) | ( n16802 & n16807 ) ;
  assign n16809 = ( n16802 & n16807 ) | ( n16802 & ~n16808 ) | ( n16807 & ~n16808 ) ;
  assign n16810 = ( x2 & n16808 ) | ( x2 & ~n16809 ) | ( n16808 & ~n16809 ) ;
  assign n16811 = ( n16741 & n16799 ) | ( n16741 & n16810 ) | ( n16799 & n16810 ) ;
  assign n16812 = n7296 & ~n16484 ;
  assign n16813 = n7879 & ~n16057 ;
  assign n16814 = n7300 & ~n16061 ;
  assign n16815 = n7299 & n16059 ;
  assign n16816 = n16814 | n16815 ;
  assign n16817 = ( ~n16812 & n16813 ) | ( ~n16812 & n16816 ) | ( n16813 & n16816 ) ;
  assign n16818 = ( ~x8 & n16812 ) | ( ~x8 & n16817 ) | ( n16812 & n16817 ) ;
  assign n16819 = ( n16812 & n16817 ) | ( n16812 & ~n16818 ) | ( n16817 & ~n16818 ) ;
  assign n16820 = ( x8 & n16818 ) | ( x8 & ~n16819 ) | ( n16818 & ~n16819 ) ;
  assign n16821 = n5966 & ~n16221 ;
  assign n16822 = n6464 & n16069 ;
  assign n16823 = n5970 & ~n16073 ;
  assign n16824 = n5969 & n16071 ;
  assign n16825 = n16823 | n16824 ;
  assign n16826 = ( ~n16821 & n16822 ) | ( ~n16821 & n16825 ) | ( n16822 & n16825 ) ;
  assign n16827 = ( ~x14 & n16821 ) | ( ~x14 & n16826 ) | ( n16821 & n16826 ) ;
  assign n16828 = ( n16821 & n16826 ) | ( n16821 & ~n16827 ) | ( n16826 & ~n16827 ) ;
  assign n16829 = ( x14 & n16827 ) | ( x14 & ~n16828 ) | ( n16827 & ~n16828 ) ;
  assign n16830 = x17 & ~n16767 ;
  assign n16831 = ~n16760 & n16830 ;
  assign n16832 = n5397 & ~n16081 ;
  assign n16833 = n5508 & n16169 ;
  assign n16834 = n5507 & ~n16075 ;
  assign n16835 = n5504 & ~n16079 ;
  assign n16836 = n5666 & n16077 ;
  assign n16837 = n16835 | n16836 ;
  assign n16838 = ( ~n16833 & n16834 ) | ( ~n16833 & n16837 ) | ( n16834 & n16837 ) ;
  assign n16839 = ( ~x17 & n16833 ) | ( ~x17 & n16838 ) | ( n16833 & n16838 ) ;
  assign n16840 = ( n16833 & n16838 ) | ( n16833 & ~n16839 ) | ( n16838 & ~n16839 ) ;
  assign n16841 = ( x17 & n16839 ) | ( x17 & ~n16840 ) | ( n16839 & ~n16840 ) ;
  assign n16842 = ( n16831 & n16832 ) | ( n16831 & n16841 ) | ( n16832 & n16841 ) ;
  assign n16843 = ( ~n16831 & n16832 ) | ( ~n16831 & n16841 ) | ( n16832 & n16841 ) ;
  assign n16844 = ( n16831 & ~n16842 ) | ( n16831 & n16843 ) | ( ~n16842 & n16843 ) ;
  assign n16845 = ( n16770 & n16829 ) | ( n16770 & n16844 ) | ( n16829 & n16844 ) ;
  assign n16846 = ( ~n16770 & n16829 ) | ( ~n16770 & n16844 ) | ( n16829 & n16844 ) ;
  assign n16847 = ( n16770 & ~n16845 ) | ( n16770 & n16846 ) | ( ~n16845 & n16846 ) ;
  assign n16848 = n6584 & n16315 ;
  assign n16849 = n7022 & n16063 ;
  assign n16850 = n6588 & n16067 ;
  assign n16851 = n6587 & n16065 ;
  assign n16852 = n16850 | n16851 ;
  assign n16853 = ( ~n16848 & n16849 ) | ( ~n16848 & n16852 ) | ( n16849 & n16852 ) ;
  assign n16854 = ( ~x11 & n16848 ) | ( ~x11 & n16853 ) | ( n16848 & n16853 ) ;
  assign n16855 = ( n16848 & n16853 ) | ( n16848 & ~n16854 ) | ( n16853 & ~n16854 ) ;
  assign n16856 = ( x11 & n16854 ) | ( x11 & ~n16855 ) | ( n16854 & ~n16855 ) ;
  assign n16857 = ( n16782 & n16847 ) | ( n16782 & n16856 ) | ( n16847 & n16856 ) ;
  assign n16858 = ( ~n16782 & n16847 ) | ( ~n16782 & n16856 ) | ( n16847 & n16856 ) ;
  assign n16859 = ( n16782 & ~n16857 ) | ( n16782 & n16858 ) | ( ~n16857 & n16858 ) ;
  assign n16860 = ( n16785 & n16820 ) | ( n16785 & n16859 ) | ( n16820 & n16859 ) ;
  assign n16861 = ( ~n16785 & n16820 ) | ( ~n16785 & n16859 ) | ( n16820 & n16859 ) ;
  assign n16862 = ( n16785 & ~n16860 ) | ( n16785 & n16861 ) | ( ~n16860 & n16861 ) ;
  assign n16863 = n8230 & n16611 ;
  assign n16864 = n8229 & ~n16051 ;
  assign n16865 = n8226 & ~n16055 ;
  assign n16866 = n8225 & n16053 ;
  assign n16867 = n16865 | n16866 ;
  assign n16868 = ( ~n16863 & n16864 ) | ( ~n16863 & n16867 ) | ( n16864 & n16867 ) ;
  assign n16869 = ( ~x5 & n16863 ) | ( ~x5 & n16868 ) | ( n16863 & n16868 ) ;
  assign n16870 = ( n16863 & n16868 ) | ( n16863 & ~n16869 ) | ( n16868 & ~n16869 ) ;
  assign n16871 = ( x5 & n16869 ) | ( x5 & ~n16870 ) | ( n16869 & ~n16870 ) ;
  assign n16872 = ( n16797 & n16862 ) | ( n16797 & n16871 ) | ( n16862 & n16871 ) ;
  assign n16873 = ( ~n16797 & n16862 ) | ( ~n16797 & n16871 ) | ( n16862 & n16871 ) ;
  assign n16874 = ( n16797 & ~n16872 ) | ( n16797 & n16873 ) | ( ~n16872 & n16873 ) ;
  assign n16875 = ( n16045 & ~n16047 ) | ( n16045 & n16099 ) | ( ~n16047 & n16099 ) ;
  assign n16876 = ( n16047 & ~n16100 ) | ( n16047 & n16875 ) | ( ~n16100 & n16875 ) ;
  assign n16877 = n36 & ~n16876 ;
  assign n16878 = n8967 & ~n16049 ;
  assign n16879 = ( x0 & n8966 ) | ( x0 & n16047 ) | ( n8966 & n16047 ) ;
  assign n16880 = ( n8966 & n16878 ) | ( n8966 & ~n16879 ) | ( n16878 & ~n16879 ) ;
  assign n16881 = n35 & n16045 ;
  assign n16882 = ( n35 & n16880 ) | ( n35 & ~n16881 ) | ( n16880 & ~n16881 ) ;
  assign n16883 = ( ~x2 & n16877 ) | ( ~x2 & n16882 ) | ( n16877 & n16882 ) ;
  assign n16884 = ( n16877 & n16882 ) | ( n16877 & ~n16883 ) | ( n16882 & ~n16883 ) ;
  assign n16885 = ( x2 & n16883 ) | ( x2 & ~n16884 ) | ( n16883 & ~n16884 ) ;
  assign n16886 = ( n16811 & n16874 ) | ( n16811 & n16885 ) | ( n16874 & n16885 ) ;
  assign n16887 = n7296 & n16541 ;
  assign n16888 = n7879 & ~n16055 ;
  assign n16889 = n7300 & n16059 ;
  assign n16890 = n7299 & ~n16057 ;
  assign n16891 = n16889 | n16890 ;
  assign n16892 = ( ~n16887 & n16888 ) | ( ~n16887 & n16891 ) | ( n16888 & n16891 ) ;
  assign n16893 = ( ~x8 & n16887 ) | ( ~x8 & n16892 ) | ( n16887 & n16892 ) ;
  assign n16894 = ( n16887 & n16892 ) | ( n16887 & ~n16893 ) | ( n16892 & ~n16893 ) ;
  assign n16895 = ( x8 & n16893 ) | ( x8 & ~n16894 ) | ( n16893 & ~n16894 ) ;
  assign n16896 = n5966 & n16269 ;
  assign n16897 = n6464 & n16067 ;
  assign n16898 = n5970 & n16071 ;
  assign n16899 = n5969 & n16069 ;
  assign n16900 = n16898 | n16899 ;
  assign n16901 = ( ~n16896 & n16897 ) | ( ~n16896 & n16900 ) | ( n16897 & n16900 ) ;
  assign n16902 = ( ~x14 & n16896 ) | ( ~x14 & n16901 ) | ( n16896 & n16901 ) ;
  assign n16903 = ( n16896 & n16901 ) | ( n16896 & ~n16902 ) | ( n16901 & ~n16902 ) ;
  assign n16904 = ( x14 & n16902 ) | ( x14 & ~n16903 ) | ( n16902 & ~n16903 ) ;
  assign n16905 = n5508 & ~n16176 ;
  assign n16906 = n5507 & ~n16073 ;
  assign n16907 = n5504 & n16077 ;
  assign n16908 = n5666 & ~n16075 ;
  assign n16909 = n16907 | n16908 ;
  assign n16910 = ( ~n16905 & n16906 ) | ( ~n16905 & n16909 ) | ( n16906 & n16909 ) ;
  assign n16911 = ( ~x17 & n16905 ) | ( ~x17 & n16910 ) | ( n16905 & n16910 ) ;
  assign n16912 = ( n16905 & n16910 ) | ( n16905 & ~n16911 ) | ( n16910 & ~n16911 ) ;
  assign n16913 = ( x17 & n16911 ) | ( x17 & ~n16912 ) | ( n16911 & ~n16912 ) ;
  assign n16914 = x20 & n16832 ;
  assign n16915 = ( n4974 & n16155 ) | ( n4974 & n16187 ) | ( n16155 & n16187 ) ;
  assign n16916 = n4972 | n16081 ;
  assign n16917 = n5398 & ~n16079 ;
  assign n16918 = ( ~n16081 & n16916 ) | ( ~n16081 & n16917 ) | ( n16916 & n16917 ) ;
  assign n16919 = ( n16914 & n16915 ) | ( n16914 & n16918 ) | ( n16915 & n16918 ) ;
  assign n16920 = n16915 | n16918 ;
  assign n16921 = ~n16914 & n16920 ;
  assign n16922 = ( n16914 & ~n16919 ) | ( n16914 & n16921 ) | ( ~n16919 & n16921 ) ;
  assign n16923 = ( n16842 & n16913 ) | ( n16842 & n16922 ) | ( n16913 & n16922 ) ;
  assign n16924 = ( ~n16842 & n16913 ) | ( ~n16842 & n16922 ) | ( n16913 & n16922 ) ;
  assign n16925 = ( n16842 & ~n16923 ) | ( n16842 & n16924 ) | ( ~n16923 & n16924 ) ;
  assign n16926 = ( n16845 & n16904 ) | ( n16845 & n16925 ) | ( n16904 & n16925 ) ;
  assign n16927 = ( ~n16845 & n16904 ) | ( ~n16845 & n16925 ) | ( n16904 & n16925 ) ;
  assign n16928 = ( n16845 & ~n16926 ) | ( n16845 & n16927 ) | ( ~n16926 & n16927 ) ;
  assign n16929 = n6584 & ~n16354 ;
  assign n16930 = n7022 & ~n16061 ;
  assign n16931 = n6588 & n16065 ;
  assign n16932 = n6587 & n16063 ;
  assign n16933 = n16931 | n16932 ;
  assign n16934 = ( ~n16929 & n16930 ) | ( ~n16929 & n16933 ) | ( n16930 & n16933 ) ;
  assign n16935 = ( ~x11 & n16929 ) | ( ~x11 & n16934 ) | ( n16929 & n16934 ) ;
  assign n16936 = ( n16929 & n16934 ) | ( n16929 & ~n16935 ) | ( n16934 & ~n16935 ) ;
  assign n16937 = ( x11 & n16935 ) | ( x11 & ~n16936 ) | ( n16935 & ~n16936 ) ;
  assign n16938 = ( n16857 & n16928 ) | ( n16857 & n16937 ) | ( n16928 & n16937 ) ;
  assign n16939 = ( ~n16857 & n16928 ) | ( ~n16857 & n16937 ) | ( n16928 & n16937 ) ;
  assign n16940 = ( n16857 & ~n16938 ) | ( n16857 & n16939 ) | ( ~n16938 & n16939 ) ;
  assign n16941 = ( n16860 & n16895 ) | ( n16860 & n16940 ) | ( n16895 & n16940 ) ;
  assign n16942 = ( ~n16860 & n16895 ) | ( ~n16860 & n16940 ) | ( n16895 & n16940 ) ;
  assign n16943 = ( n16860 & ~n16941 ) | ( n16860 & n16942 ) | ( ~n16941 & n16942 ) ;
  assign n16944 = n8230 & ~n16674 ;
  assign n16945 = n8229 & ~n16049 ;
  assign n16946 = n8226 & n16053 ;
  assign n16947 = n8225 & ~n16051 ;
  assign n16948 = n16946 | n16947 ;
  assign n16949 = ( ~n16944 & n16945 ) | ( ~n16944 & n16948 ) | ( n16945 & n16948 ) ;
  assign n16950 = ( ~x5 & n16944 ) | ( ~x5 & n16949 ) | ( n16944 & n16949 ) ;
  assign n16951 = ( n16944 & n16949 ) | ( n16944 & ~n16950 ) | ( n16949 & ~n16950 ) ;
  assign n16952 = ( x5 & n16950 ) | ( x5 & ~n16951 ) | ( n16950 & ~n16951 ) ;
  assign n16953 = ( n16872 & n16943 ) | ( n16872 & n16952 ) | ( n16943 & n16952 ) ;
  assign n16954 = ( ~n16872 & n16943 ) | ( ~n16872 & n16952 ) | ( n16943 & n16952 ) ;
  assign n16955 = ( n16872 & ~n16953 ) | ( n16872 & n16954 ) | ( ~n16953 & n16954 ) ;
  assign n16956 = ( n16043 & ~n16045 ) | ( n16043 & n16100 ) | ( ~n16045 & n16100 ) ;
  assign n16957 = ( n16045 & ~n16101 ) | ( n16045 & n16956 ) | ( ~n16101 & n16956 ) ;
  assign n16958 = n36 & ~n16957 ;
  assign n16959 = n8967 & ~n16047 ;
  assign n16960 = ( x0 & n8966 ) | ( x0 & n16045 ) | ( n8966 & n16045 ) ;
  assign n16961 = ( n8966 & n16959 ) | ( n8966 & ~n16960 ) | ( n16959 & ~n16960 ) ;
  assign n16962 = n35 & n16043 ;
  assign n16963 = ( n35 & n16961 ) | ( n35 & ~n16962 ) | ( n16961 & ~n16962 ) ;
  assign n16964 = ( ~x2 & n16958 ) | ( ~x2 & n16963 ) | ( n16958 & n16963 ) ;
  assign n16965 = ( n16958 & n16963 ) | ( n16958 & ~n16964 ) | ( n16963 & ~n16964 ) ;
  assign n16966 = ( x2 & n16964 ) | ( x2 & ~n16965 ) | ( n16964 & ~n16965 ) ;
  assign n16967 = ( n16886 & n16955 ) | ( n16886 & n16966 ) | ( n16955 & n16966 ) ;
  assign n16968 = ( n16041 & ~n16043 ) | ( n16041 & n16101 ) | ( ~n16043 & n16101 ) ;
  assign n16969 = ( ~n16101 & n16102 ) | ( ~n16101 & n16968 ) | ( n16102 & n16968 ) ;
  assign n16970 = n36 & n16969 ;
  assign n16971 = n8967 & ~n16045 ;
  assign n16972 = ( x0 & n8966 ) | ( x0 & n16043 ) | ( n8966 & n16043 ) ;
  assign n16973 = ( n8966 & n16971 ) | ( n8966 & ~n16972 ) | ( n16971 & ~n16972 ) ;
  assign n16974 = n35 & ~n16041 ;
  assign n16975 = ( n35 & n16973 ) | ( n35 & ~n16974 ) | ( n16973 & ~n16974 ) ;
  assign n16976 = ( ~x2 & n16970 ) | ( ~x2 & n16975 ) | ( n16970 & n16975 ) ;
  assign n16977 = ( n16970 & n16975 ) | ( n16970 & ~n16976 ) | ( n16975 & ~n16976 ) ;
  assign n16978 = ( x2 & n16976 ) | ( x2 & ~n16977 ) | ( n16976 & ~n16977 ) ;
  assign n16979 = n8230 & ~n16801 ;
  assign n16980 = n8229 & ~n16047 ;
  assign n16981 = n8226 & ~n16051 ;
  assign n16982 = n8225 & ~n16049 ;
  assign n16983 = n16981 | n16982 ;
  assign n16984 = ( ~n16979 & n16980 ) | ( ~n16979 & n16983 ) | ( n16980 & n16983 ) ;
  assign n16985 = ( ~x5 & n16979 ) | ( ~x5 & n16984 ) | ( n16979 & n16984 ) ;
  assign n16986 = ( n16979 & n16984 ) | ( n16979 & ~n16985 ) | ( n16984 & ~n16985 ) ;
  assign n16987 = ( x5 & n16985 ) | ( x5 & ~n16986 ) | ( n16985 & ~n16986 ) ;
  assign n16988 = n6584 & ~n16433 ;
  assign n16989 = n7022 & n16059 ;
  assign n16990 = n6588 & n16063 ;
  assign n16991 = n6587 & ~n16061 ;
  assign n16992 = n16990 | n16991 ;
  assign n16993 = ( ~n16988 & n16989 ) | ( ~n16988 & n16992 ) | ( n16989 & n16992 ) ;
  assign n16994 = ( ~x11 & n16988 ) | ( ~x11 & n16993 ) | ( n16988 & n16993 ) ;
  assign n16995 = ( n16988 & n16993 ) | ( n16988 & ~n16994 ) | ( n16993 & ~n16994 ) ;
  assign n16996 = ( x11 & n16994 ) | ( x11 & ~n16995 ) | ( n16994 & ~n16995 ) ;
  assign n16997 = n5508 & n16209 ;
  assign n16998 = n5507 & n16071 ;
  assign n16999 = n5504 & ~n16075 ;
  assign n17000 = n5666 & ~n16073 ;
  assign n17001 = n16999 | n17000 ;
  assign n17002 = ( ~n16997 & n16998 ) | ( ~n16997 & n17001 ) | ( n16998 & n17001 ) ;
  assign n17003 = ( ~x17 & n16997 ) | ( ~x17 & n17002 ) | ( n16997 & n17002 ) ;
  assign n17004 = ( n16997 & n17002 ) | ( n16997 & ~n17003 ) | ( n17002 & ~n17003 ) ;
  assign n17005 = ( x17 & n17003 ) | ( x17 & ~n17004 ) | ( n17003 & ~n17004 ) ;
  assign n17006 = ( x20 & n16914 ) | ( x20 & n16920 ) | ( n16914 & n16920 ) ;
  assign n17007 = ( n4974 & n16083 ) | ( n4974 & n16198 ) | ( n16083 & n16198 ) ;
  assign n17008 = n4973 & ~n16081 ;
  assign n17009 = n4972 & ~n16079 ;
  assign n17010 = n17008 | n17009 ;
  assign n17011 = n5398 & ~n16077 ;
  assign n17012 = ( n5398 & n17010 ) | ( n5398 & ~n17011 ) | ( n17010 & ~n17011 ) ;
  assign n17013 = ( ~n17006 & n17007 ) | ( ~n17006 & n17012 ) | ( n17007 & n17012 ) ;
  assign n17014 = ( n17007 & n17012 ) | ( n17007 & ~n17013 ) | ( n17012 & ~n17013 ) ;
  assign n17015 = ( n17006 & n17013 ) | ( n17006 & ~n17014 ) | ( n17013 & ~n17014 ) ;
  assign n17016 = ( n16923 & n17005 ) | ( n16923 & n17015 ) | ( n17005 & n17015 ) ;
  assign n17017 = ( ~n16923 & n17005 ) | ( ~n16923 & n17015 ) | ( n17005 & n17015 ) ;
  assign n17018 = ( n16923 & ~n17016 ) | ( n16923 & n17017 ) | ( ~n17016 & n17017 ) ;
  assign n17019 = n5966 & n16281 ;
  assign n17020 = n6464 & n16065 ;
  assign n17021 = n5970 & n16069 ;
  assign n17022 = n5969 & n16067 ;
  assign n17023 = n17021 | n17022 ;
  assign n17024 = ( ~n17019 & n17020 ) | ( ~n17019 & n17023 ) | ( n17020 & n17023 ) ;
  assign n17025 = ( ~x14 & n17019 ) | ( ~x14 & n17024 ) | ( n17019 & n17024 ) ;
  assign n17026 = ( n17019 & n17024 ) | ( n17019 & ~n17025 ) | ( n17024 & ~n17025 ) ;
  assign n17027 = ( x14 & n17025 ) | ( x14 & ~n17026 ) | ( n17025 & ~n17026 ) ;
  assign n17028 = ( n16926 & n17018 ) | ( n16926 & n17027 ) | ( n17018 & n17027 ) ;
  assign n17029 = ( ~n16926 & n17018 ) | ( ~n16926 & n17027 ) | ( n17018 & n17027 ) ;
  assign n17030 = ( n16926 & ~n17028 ) | ( n16926 & n17029 ) | ( ~n17028 & n17029 ) ;
  assign n17031 = ( n16938 & n16996 ) | ( n16938 & n17030 ) | ( n16996 & n17030 ) ;
  assign n17032 = ( ~n16938 & n16996 ) | ( ~n16938 & n17030 ) | ( n16996 & n17030 ) ;
  assign n17033 = ( n16938 & ~n17031 ) | ( n16938 & n17032 ) | ( ~n17031 & n17032 ) ;
  assign n17034 = n7296 & n16553 ;
  assign n17035 = n7879 & n16053 ;
  assign n17036 = n7300 & ~n16057 ;
  assign n17037 = n7299 & ~n16055 ;
  assign n17038 = n17036 | n17037 ;
  assign n17039 = ( ~n17034 & n17035 ) | ( ~n17034 & n17038 ) | ( n17035 & n17038 ) ;
  assign n17040 = ( ~x8 & n17034 ) | ( ~x8 & n17039 ) | ( n17034 & n17039 ) ;
  assign n17041 = ( n17034 & n17039 ) | ( n17034 & ~n17040 ) | ( n17039 & ~n17040 ) ;
  assign n17042 = ( x8 & n17040 ) | ( x8 & ~n17041 ) | ( n17040 & ~n17041 ) ;
  assign n17043 = ( n16941 & n17033 ) | ( n16941 & n17042 ) | ( n17033 & n17042 ) ;
  assign n17044 = ( ~n16941 & n17033 ) | ( ~n16941 & n17042 ) | ( n17033 & n17042 ) ;
  assign n17045 = ( n16941 & ~n17043 ) | ( n16941 & n17044 ) | ( ~n17043 & n17044 ) ;
  assign n17046 = ( n16953 & n16987 ) | ( n16953 & n17045 ) | ( n16987 & n17045 ) ;
  assign n17047 = ( ~n16953 & n16987 ) | ( ~n16953 & n17045 ) | ( n16987 & n17045 ) ;
  assign n17048 = ( n16953 & ~n17046 ) | ( n16953 & n17047 ) | ( ~n17046 & n17047 ) ;
  assign n17049 = ( n16967 & n16978 ) | ( n16967 & n17048 ) | ( n16978 & n17048 ) ;
  assign n17050 = ( n16039 & n16041 ) | ( n16039 & ~n16103 ) | ( n16041 & ~n16103 ) ;
  assign n17051 = ( n16102 & n16103 ) | ( n16102 & ~n17050 ) | ( n16103 & ~n17050 ) ;
  assign n17052 = n36 & ~n17051 ;
  assign n17053 = n8967 & ~n16043 ;
  assign n17054 = ( x0 & n8966 ) | ( x0 & ~n16041 ) | ( n8966 & ~n16041 ) ;
  assign n17055 = ( n8966 & n17053 ) | ( n8966 & ~n17054 ) | ( n17053 & ~n17054 ) ;
  assign n17056 = n35 & ~n16039 ;
  assign n17057 = ( n35 & n17055 ) | ( n35 & ~n17056 ) | ( n17055 & ~n17056 ) ;
  assign n17058 = ( ~x2 & n17052 ) | ( ~x2 & n17057 ) | ( n17052 & n17057 ) ;
  assign n17059 = ( n17052 & n17057 ) | ( n17052 & ~n17058 ) | ( n17057 & ~n17058 ) ;
  assign n17060 = ( x2 & n17058 ) | ( x2 & ~n17059 ) | ( n17058 & ~n17059 ) ;
  assign n17061 = n8230 & ~n16876 ;
  assign n17062 = n8229 & ~n16045 ;
  assign n17063 = n8226 & ~n16049 ;
  assign n17064 = n8225 & ~n16047 ;
  assign n17065 = n17063 | n17064 ;
  assign n17066 = ( ~n17061 & n17062 ) | ( ~n17061 & n17065 ) | ( n17062 & n17065 ) ;
  assign n17067 = ( ~x5 & n17061 ) | ( ~x5 & n17066 ) | ( n17061 & n17066 ) ;
  assign n17068 = ( n17061 & n17066 ) | ( n17061 & ~n17067 ) | ( n17066 & ~n17067 ) ;
  assign n17069 = ( x5 & n17067 ) | ( x5 & ~n17068 ) | ( n17067 & ~n17068 ) ;
  assign n17070 = n6584 & ~n16484 ;
  assign n17071 = n7022 & ~n16057 ;
  assign n17072 = n6588 & ~n16061 ;
  assign n17073 = n6587 & n16059 ;
  assign n17074 = n17072 | n17073 ;
  assign n17075 = ( ~n17070 & n17071 ) | ( ~n17070 & n17074 ) | ( n17071 & n17074 ) ;
  assign n17076 = ( ~x11 & n17070 ) | ( ~x11 & n17075 ) | ( n17070 & n17075 ) ;
  assign n17077 = ( n17070 & n17075 ) | ( n17070 & ~n17076 ) | ( n17075 & ~n17076 ) ;
  assign n17078 = ( x11 & n17076 ) | ( x11 & ~n17077 ) | ( n17076 & ~n17077 ) ;
  assign n17079 = n5508 & ~n16221 ;
  assign n17080 = n5507 & n16069 ;
  assign n17081 = n5504 & ~n16073 ;
  assign n17082 = n5666 & n16071 ;
  assign n17083 = n17081 | n17082 ;
  assign n17084 = ( ~n17079 & n17080 ) | ( ~n17079 & n17083 ) | ( n17080 & n17083 ) ;
  assign n17085 = ( ~x17 & n17079 ) | ( ~x17 & n17084 ) | ( n17079 & n17084 ) ;
  assign n17086 = ( n17079 & n17084 ) | ( n17079 & ~n17085 ) | ( n17084 & ~n17085 ) ;
  assign n17087 = ( x17 & n17085 ) | ( x17 & ~n17086 ) | ( n17085 & ~n17086 ) ;
  assign n17088 = x20 & ~n17013 ;
  assign n17089 = ~n17006 & n17088 ;
  assign n17090 = n4711 & ~n16081 ;
  assign n17091 = n4974 & n16169 ;
  assign n17092 = n5398 & ~n16075 ;
  assign n17093 = n4973 & ~n16079 ;
  assign n17094 = n4972 & n16077 ;
  assign n17095 = n17093 | n17094 ;
  assign n17096 = ( ~n17091 & n17092 ) | ( ~n17091 & n17095 ) | ( n17092 & n17095 ) ;
  assign n17097 = ( ~x20 & n17091 ) | ( ~x20 & n17096 ) | ( n17091 & n17096 ) ;
  assign n17098 = ( n17091 & n17096 ) | ( n17091 & ~n17097 ) | ( n17096 & ~n17097 ) ;
  assign n17099 = ( x20 & n17097 ) | ( x20 & ~n17098 ) | ( n17097 & ~n17098 ) ;
  assign n17100 = ( n17089 & n17090 ) | ( n17089 & n17099 ) | ( n17090 & n17099 ) ;
  assign n17101 = ( ~n17089 & n17090 ) | ( ~n17089 & n17099 ) | ( n17090 & n17099 ) ;
  assign n17102 = ( n17089 & ~n17100 ) | ( n17089 & n17101 ) | ( ~n17100 & n17101 ) ;
  assign n17103 = ( n17016 & n17087 ) | ( n17016 & n17102 ) | ( n17087 & n17102 ) ;
  assign n17104 = ( ~n17016 & n17087 ) | ( ~n17016 & n17102 ) | ( n17087 & n17102 ) ;
  assign n17105 = ( n17016 & ~n17103 ) | ( n17016 & n17104 ) | ( ~n17103 & n17104 ) ;
  assign n17106 = n5966 & n16315 ;
  assign n17107 = n6464 & n16063 ;
  assign n17108 = n5970 & n16067 ;
  assign n17109 = n5969 & n16065 ;
  assign n17110 = n17108 | n17109 ;
  assign n17111 = ( ~n17106 & n17107 ) | ( ~n17106 & n17110 ) | ( n17107 & n17110 ) ;
  assign n17112 = ( ~x14 & n17106 ) | ( ~x14 & n17111 ) | ( n17106 & n17111 ) ;
  assign n17113 = ( n17106 & n17111 ) | ( n17106 & ~n17112 ) | ( n17111 & ~n17112 ) ;
  assign n17114 = ( x14 & n17112 ) | ( x14 & ~n17113 ) | ( n17112 & ~n17113 ) ;
  assign n17115 = ( n17028 & n17105 ) | ( n17028 & n17114 ) | ( n17105 & n17114 ) ;
  assign n17116 = ( ~n17028 & n17105 ) | ( ~n17028 & n17114 ) | ( n17105 & n17114 ) ;
  assign n17117 = ( n17028 & ~n17115 ) | ( n17028 & n17116 ) | ( ~n17115 & n17116 ) ;
  assign n17118 = ( n17031 & n17078 ) | ( n17031 & n17117 ) | ( n17078 & n17117 ) ;
  assign n17119 = ( ~n17031 & n17078 ) | ( ~n17031 & n17117 ) | ( n17078 & n17117 ) ;
  assign n17120 = ( n17031 & ~n17118 ) | ( n17031 & n17119 ) | ( ~n17118 & n17119 ) ;
  assign n17121 = n7296 & n16611 ;
  assign n17122 = n7879 & ~n16051 ;
  assign n17123 = n7300 & ~n16055 ;
  assign n17124 = n7299 & n16053 ;
  assign n17125 = n17123 | n17124 ;
  assign n17126 = ( ~n17121 & n17122 ) | ( ~n17121 & n17125 ) | ( n17122 & n17125 ) ;
  assign n17127 = ( ~x8 & n17121 ) | ( ~x8 & n17126 ) | ( n17121 & n17126 ) ;
  assign n17128 = ( n17121 & n17126 ) | ( n17121 & ~n17127 ) | ( n17126 & ~n17127 ) ;
  assign n17129 = ( x8 & n17127 ) | ( x8 & ~n17128 ) | ( n17127 & ~n17128 ) ;
  assign n17130 = ( n17043 & n17120 ) | ( n17043 & n17129 ) | ( n17120 & n17129 ) ;
  assign n17131 = ( ~n17043 & n17120 ) | ( ~n17043 & n17129 ) | ( n17120 & n17129 ) ;
  assign n17132 = ( n17043 & ~n17130 ) | ( n17043 & n17131 ) | ( ~n17130 & n17131 ) ;
  assign n17133 = ( n17046 & n17069 ) | ( n17046 & n17132 ) | ( n17069 & n17132 ) ;
  assign n17134 = ( ~n17046 & n17069 ) | ( ~n17046 & n17132 ) | ( n17069 & n17132 ) ;
  assign n17135 = ( n17046 & ~n17133 ) | ( n17046 & n17134 ) | ( ~n17133 & n17134 ) ;
  assign n17136 = ( n17049 & n17060 ) | ( n17049 & n17135 ) | ( n17060 & n17135 ) ;
  assign n17137 = ( n16037 & n16039 ) | ( n16037 & ~n16103 ) | ( n16039 & ~n16103 ) ;
  assign n17138 = ( ~n16039 & n16104 ) | ( ~n16039 & n17137 ) | ( n16104 & n17137 ) ;
  assign n17139 = n36 & ~n17138 ;
  assign n17140 = n8967 & n16041 ;
  assign n17141 = ( x0 & n8966 ) | ( x0 & ~n16039 ) | ( n8966 & ~n16039 ) ;
  assign n17142 = ( n8966 & n17140 ) | ( n8966 & ~n17141 ) | ( n17140 & ~n17141 ) ;
  assign n17143 = n35 & n16037 ;
  assign n17144 = ( n35 & n17142 ) | ( n35 & ~n17143 ) | ( n17142 & ~n17143 ) ;
  assign n17145 = ( ~x2 & n17139 ) | ( ~x2 & n17144 ) | ( n17139 & n17144 ) ;
  assign n17146 = ( n17139 & n17144 ) | ( n17139 & ~n17145 ) | ( n17144 & ~n17145 ) ;
  assign n17147 = ( x2 & n17145 ) | ( x2 & ~n17146 ) | ( n17145 & ~n17146 ) ;
  assign n17148 = n8230 & ~n16957 ;
  assign n17149 = n8229 & ~n16043 ;
  assign n17150 = n8226 & ~n16047 ;
  assign n17151 = n8225 & ~n16045 ;
  assign n17152 = n17150 | n17151 ;
  assign n17153 = ( ~n17148 & n17149 ) | ( ~n17148 & n17152 ) | ( n17149 & n17152 ) ;
  assign n17154 = ( ~x5 & n17148 ) | ( ~x5 & n17153 ) | ( n17148 & n17153 ) ;
  assign n17155 = ( n17148 & n17153 ) | ( n17148 & ~n17154 ) | ( n17153 & ~n17154 ) ;
  assign n17156 = ( x5 & n17154 ) | ( x5 & ~n17155 ) | ( n17154 & ~n17155 ) ;
  assign n17157 = n6584 & n16541 ;
  assign n17158 = n7022 & ~n16055 ;
  assign n17159 = n6588 & n16059 ;
  assign n17160 = n6587 & ~n16057 ;
  assign n17161 = n17159 | n17160 ;
  assign n17162 = ( ~n17157 & n17158 ) | ( ~n17157 & n17161 ) | ( n17158 & n17161 ) ;
  assign n17163 = ( ~x11 & n17157 ) | ( ~x11 & n17162 ) | ( n17157 & n17162 ) ;
  assign n17164 = ( n17157 & n17162 ) | ( n17157 & ~n17163 ) | ( n17162 & ~n17163 ) ;
  assign n17165 = ( x11 & n17163 ) | ( x11 & ~n17164 ) | ( n17163 & ~n17164 ) ;
  assign n17166 = n5508 & n16269 ;
  assign n17167 = n5507 & n16067 ;
  assign n17168 = n5504 & n16071 ;
  assign n17169 = n5666 & n16069 ;
  assign n17170 = n17168 | n17169 ;
  assign n17171 = ( ~n17166 & n17167 ) | ( ~n17166 & n17170 ) | ( n17167 & n17170 ) ;
  assign n17172 = ( ~x17 & n17166 ) | ( ~x17 & n17171 ) | ( n17166 & n17171 ) ;
  assign n17173 = ( n17166 & n17171 ) | ( n17166 & ~n17172 ) | ( n17171 & ~n17172 ) ;
  assign n17174 = ( x17 & n17172 ) | ( x17 & ~n17173 ) | ( n17172 & ~n17173 ) ;
  assign n17175 = n4974 & ~n16176 ;
  assign n17176 = n5398 & ~n16073 ;
  assign n17177 = n4973 & n16077 ;
  assign n17178 = n4972 & ~n16075 ;
  assign n17179 = n17177 | n17178 ;
  assign n17180 = ( ~n17175 & n17176 ) | ( ~n17175 & n17179 ) | ( n17176 & n17179 ) ;
  assign n17181 = ( ~x20 & n17175 ) | ( ~x20 & n17180 ) | ( n17175 & n17180 ) ;
  assign n17182 = ( n17175 & n17180 ) | ( n17175 & ~n17181 ) | ( n17180 & ~n17181 ) ;
  assign n17183 = ( x20 & n17181 ) | ( x20 & ~n17182 ) | ( n17181 & ~n17182 ) ;
  assign n17184 = x23 & n17090 ;
  assign n17185 = ( n4713 & n16155 ) | ( n4713 & n16187 ) | ( n16155 & n16187 ) ;
  assign n17186 = n4792 | n16081 ;
  assign n17187 = n4712 & ~n16079 ;
  assign n17188 = ( ~n16081 & n17186 ) | ( ~n16081 & n17187 ) | ( n17186 & n17187 ) ;
  assign n17189 = ( n17184 & n17185 ) | ( n17184 & n17188 ) | ( n17185 & n17188 ) ;
  assign n17190 = n17185 | n17188 ;
  assign n17191 = ~n17184 & n17190 ;
  assign n17192 = ( n17184 & ~n17189 ) | ( n17184 & n17191 ) | ( ~n17189 & n17191 ) ;
  assign n17193 = ( n17100 & n17183 ) | ( n17100 & n17192 ) | ( n17183 & n17192 ) ;
  assign n17194 = ( ~n17100 & n17183 ) | ( ~n17100 & n17192 ) | ( n17183 & n17192 ) ;
  assign n17195 = ( n17100 & ~n17193 ) | ( n17100 & n17194 ) | ( ~n17193 & n17194 ) ;
  assign n17196 = ( n17103 & n17174 ) | ( n17103 & n17195 ) | ( n17174 & n17195 ) ;
  assign n17197 = ( ~n17103 & n17174 ) | ( ~n17103 & n17195 ) | ( n17174 & n17195 ) ;
  assign n17198 = ( n17103 & ~n17196 ) | ( n17103 & n17197 ) | ( ~n17196 & n17197 ) ;
  assign n17199 = n5966 & ~n16354 ;
  assign n17200 = n6464 & ~n16061 ;
  assign n17201 = n5970 & n16065 ;
  assign n17202 = n5969 & n16063 ;
  assign n17203 = n17201 | n17202 ;
  assign n17204 = ( ~n17199 & n17200 ) | ( ~n17199 & n17203 ) | ( n17200 & n17203 ) ;
  assign n17205 = ( ~x14 & n17199 ) | ( ~x14 & n17204 ) | ( n17199 & n17204 ) ;
  assign n17206 = ( n17199 & n17204 ) | ( n17199 & ~n17205 ) | ( n17204 & ~n17205 ) ;
  assign n17207 = ( x14 & n17205 ) | ( x14 & ~n17206 ) | ( n17205 & ~n17206 ) ;
  assign n17208 = ( n17115 & n17198 ) | ( n17115 & n17207 ) | ( n17198 & n17207 ) ;
  assign n17209 = ( ~n17115 & n17198 ) | ( ~n17115 & n17207 ) | ( n17198 & n17207 ) ;
  assign n17210 = ( n17115 & ~n17208 ) | ( n17115 & n17209 ) | ( ~n17208 & n17209 ) ;
  assign n17211 = ( n17118 & n17165 ) | ( n17118 & n17210 ) | ( n17165 & n17210 ) ;
  assign n17212 = ( ~n17118 & n17165 ) | ( ~n17118 & n17210 ) | ( n17165 & n17210 ) ;
  assign n17213 = ( n17118 & ~n17211 ) | ( n17118 & n17212 ) | ( ~n17211 & n17212 ) ;
  assign n17214 = n7296 & ~n16674 ;
  assign n17215 = n7879 & ~n16049 ;
  assign n17216 = n7300 & n16053 ;
  assign n17217 = n7299 & ~n16051 ;
  assign n17218 = n17216 | n17217 ;
  assign n17219 = ( ~n17214 & n17215 ) | ( ~n17214 & n17218 ) | ( n17215 & n17218 ) ;
  assign n17220 = ( ~x8 & n17214 ) | ( ~x8 & n17219 ) | ( n17214 & n17219 ) ;
  assign n17221 = ( n17214 & n17219 ) | ( n17214 & ~n17220 ) | ( n17219 & ~n17220 ) ;
  assign n17222 = ( x8 & n17220 ) | ( x8 & ~n17221 ) | ( n17220 & ~n17221 ) ;
  assign n17223 = ( n17130 & n17213 ) | ( n17130 & n17222 ) | ( n17213 & n17222 ) ;
  assign n17224 = ( ~n17130 & n17213 ) | ( ~n17130 & n17222 ) | ( n17213 & n17222 ) ;
  assign n17225 = ( n17130 & ~n17223 ) | ( n17130 & n17224 ) | ( ~n17223 & n17224 ) ;
  assign n17226 = ( n17133 & n17156 ) | ( n17133 & n17225 ) | ( n17156 & n17225 ) ;
  assign n17227 = ( ~n17133 & n17156 ) | ( ~n17133 & n17225 ) | ( n17156 & n17225 ) ;
  assign n17228 = ( n17133 & ~n17226 ) | ( n17133 & n17227 ) | ( ~n17226 & n17227 ) ;
  assign n17229 = ( n17136 & n17147 ) | ( n17136 & n17228 ) | ( n17147 & n17228 ) ;
  assign n17230 = n7296 & ~n16801 ;
  assign n17231 = n7879 & ~n16047 ;
  assign n17232 = n7300 & ~n16051 ;
  assign n17233 = n7299 & ~n16049 ;
  assign n17234 = n17232 | n17233 ;
  assign n17235 = ( ~n17230 & n17231 ) | ( ~n17230 & n17234 ) | ( n17231 & n17234 ) ;
  assign n17236 = ( ~x8 & n17230 ) | ( ~x8 & n17235 ) | ( n17230 & n17235 ) ;
  assign n17237 = ( n17230 & n17235 ) | ( n17230 & ~n17236 ) | ( n17235 & ~n17236 ) ;
  assign n17238 = ( x8 & n17236 ) | ( x8 & ~n17237 ) | ( n17236 & ~n17237 ) ;
  assign n17239 = n5966 & ~n16433 ;
  assign n17240 = n6464 & n16059 ;
  assign n17241 = n5970 & n16063 ;
  assign n17242 = n5969 & ~n16061 ;
  assign n17243 = n17241 | n17242 ;
  assign n17244 = ( ~n17239 & n17240 ) | ( ~n17239 & n17243 ) | ( n17240 & n17243 ) ;
  assign n17245 = ( ~x14 & n17239 ) | ( ~x14 & n17244 ) | ( n17239 & n17244 ) ;
  assign n17246 = ( n17239 & n17244 ) | ( n17239 & ~n17245 ) | ( n17244 & ~n17245 ) ;
  assign n17247 = ( x14 & n17245 ) | ( x14 & ~n17246 ) | ( n17245 & ~n17246 ) ;
  assign n17248 = n4974 & n16209 ;
  assign n17249 = n5398 & n16071 ;
  assign n17250 = n4973 & ~n16075 ;
  assign n17251 = n4972 & ~n16073 ;
  assign n17252 = n17250 | n17251 ;
  assign n17253 = ( ~n17248 & n17249 ) | ( ~n17248 & n17252 ) | ( n17249 & n17252 ) ;
  assign n17254 = ( ~x20 & n17248 ) | ( ~x20 & n17253 ) | ( n17248 & n17253 ) ;
  assign n17255 = ( n17248 & n17253 ) | ( n17248 & ~n17254 ) | ( n17253 & ~n17254 ) ;
  assign n17256 = ( x20 & n17254 ) | ( x20 & ~n17255 ) | ( n17254 & ~n17255 ) ;
  assign n17257 = ( x23 & n17184 ) | ( x23 & n17190 ) | ( n17184 & n17190 ) ;
  assign n17258 = ( n4713 & n16083 ) | ( n4713 & n16198 ) | ( n16083 & n16198 ) ;
  assign n17259 = n4709 & ~n16081 ;
  assign n17260 = n4792 & ~n16079 ;
  assign n17261 = n17259 | n17260 ;
  assign n17262 = n4712 & ~n16077 ;
  assign n17263 = ( n4712 & n17261 ) | ( n4712 & ~n17262 ) | ( n17261 & ~n17262 ) ;
  assign n17264 = ( ~n17257 & n17258 ) | ( ~n17257 & n17263 ) | ( n17258 & n17263 ) ;
  assign n17265 = ( n17258 & n17263 ) | ( n17258 & ~n17264 ) | ( n17263 & ~n17264 ) ;
  assign n17266 = ( n17257 & n17264 ) | ( n17257 & ~n17265 ) | ( n17264 & ~n17265 ) ;
  assign n17267 = ( n17193 & n17256 ) | ( n17193 & n17266 ) | ( n17256 & n17266 ) ;
  assign n17268 = ( ~n17193 & n17256 ) | ( ~n17193 & n17266 ) | ( n17256 & n17266 ) ;
  assign n17269 = ( n17193 & ~n17267 ) | ( n17193 & n17268 ) | ( ~n17267 & n17268 ) ;
  assign n17270 = n5508 & n16281 ;
  assign n17271 = n5507 & n16065 ;
  assign n17272 = n5504 & n16069 ;
  assign n17273 = n5666 & n16067 ;
  assign n17274 = n17272 | n17273 ;
  assign n17275 = ( ~n17270 & n17271 ) | ( ~n17270 & n17274 ) | ( n17271 & n17274 ) ;
  assign n17276 = ( ~x17 & n17270 ) | ( ~x17 & n17275 ) | ( n17270 & n17275 ) ;
  assign n17277 = ( n17270 & n17275 ) | ( n17270 & ~n17276 ) | ( n17275 & ~n17276 ) ;
  assign n17278 = ( x17 & n17276 ) | ( x17 & ~n17277 ) | ( n17276 & ~n17277 ) ;
  assign n17279 = ( n17196 & n17269 ) | ( n17196 & n17278 ) | ( n17269 & n17278 ) ;
  assign n17280 = ( ~n17196 & n17269 ) | ( ~n17196 & n17278 ) | ( n17269 & n17278 ) ;
  assign n17281 = ( n17196 & ~n17279 ) | ( n17196 & n17280 ) | ( ~n17279 & n17280 ) ;
  assign n17282 = ( n17208 & n17247 ) | ( n17208 & n17281 ) | ( n17247 & n17281 ) ;
  assign n17283 = ( ~n17208 & n17247 ) | ( ~n17208 & n17281 ) | ( n17247 & n17281 ) ;
  assign n17284 = ( n17208 & ~n17282 ) | ( n17208 & n17283 ) | ( ~n17282 & n17283 ) ;
  assign n17285 = n6584 & n16553 ;
  assign n17286 = n7022 & n16053 ;
  assign n17287 = n6588 & ~n16057 ;
  assign n17288 = n6587 & ~n16055 ;
  assign n17289 = n17287 | n17288 ;
  assign n17290 = ( ~n17285 & n17286 ) | ( ~n17285 & n17289 ) | ( n17286 & n17289 ) ;
  assign n17291 = ( ~x11 & n17285 ) | ( ~x11 & n17290 ) | ( n17285 & n17290 ) ;
  assign n17292 = ( n17285 & n17290 ) | ( n17285 & ~n17291 ) | ( n17290 & ~n17291 ) ;
  assign n17293 = ( x11 & n17291 ) | ( x11 & ~n17292 ) | ( n17291 & ~n17292 ) ;
  assign n17294 = ( n17211 & n17284 ) | ( n17211 & n17293 ) | ( n17284 & n17293 ) ;
  assign n17295 = ( ~n17211 & n17284 ) | ( ~n17211 & n17293 ) | ( n17284 & n17293 ) ;
  assign n17296 = ( n17211 & ~n17294 ) | ( n17211 & n17295 ) | ( ~n17294 & n17295 ) ;
  assign n17297 = ( n17223 & n17238 ) | ( n17223 & n17296 ) | ( n17238 & n17296 ) ;
  assign n17298 = ( ~n17223 & n17238 ) | ( ~n17223 & n17296 ) | ( n17238 & n17296 ) ;
  assign n17299 = ( n17223 & ~n17297 ) | ( n17223 & n17298 ) | ( ~n17297 & n17298 ) ;
  assign n17300 = n8230 & n16969 ;
  assign n17301 = n8229 & n16041 ;
  assign n17302 = n8226 & ~n16045 ;
  assign n17303 = n8225 & ~n16043 ;
  assign n17304 = n17302 | n17303 ;
  assign n17305 = ( ~n17300 & n17301 ) | ( ~n17300 & n17304 ) | ( n17301 & n17304 ) ;
  assign n17306 = ( ~x5 & n17300 ) | ( ~x5 & n17305 ) | ( n17300 & n17305 ) ;
  assign n17307 = ( n17300 & n17305 ) | ( n17300 & ~n17306 ) | ( n17305 & ~n17306 ) ;
  assign n17308 = ( x5 & n17306 ) | ( x5 & ~n17307 ) | ( n17306 & ~n17307 ) ;
  assign n17309 = ( n17226 & n17299 ) | ( n17226 & n17308 ) | ( n17299 & n17308 ) ;
  assign n17310 = ( ~n17226 & n17299 ) | ( ~n17226 & n17308 ) | ( n17299 & n17308 ) ;
  assign n17311 = ( n17226 & ~n17309 ) | ( n17226 & n17310 ) | ( ~n17309 & n17310 ) ;
  assign n17312 = ( ~n16035 & n16037 ) | ( ~n16035 & n16104 ) | ( n16037 & n16104 ) ;
  assign n17313 = ( ~n16104 & n16105 ) | ( ~n16104 & n17312 ) | ( n16105 & n17312 ) ;
  assign n17314 = n36 & ~n17313 ;
  assign n17315 = n8967 & n16039 ;
  assign n17316 = ( x0 & n8966 ) | ( x0 & n16037 ) | ( n8966 & n16037 ) ;
  assign n17317 = ( n8966 & n17315 ) | ( n8966 & ~n17316 ) | ( n17315 & ~n17316 ) ;
  assign n17318 = n35 & ~n16035 ;
  assign n17319 = ( n35 & n17317 ) | ( n35 & ~n17318 ) | ( n17317 & ~n17318 ) ;
  assign n17320 = ( ~x2 & n17314 ) | ( ~x2 & n17319 ) | ( n17314 & n17319 ) ;
  assign n17321 = ( n17314 & n17319 ) | ( n17314 & ~n17320 ) | ( n17319 & ~n17320 ) ;
  assign n17322 = ( x2 & n17320 ) | ( x2 & ~n17321 ) | ( n17320 & ~n17321 ) ;
  assign n17323 = ( n17229 & n17311 ) | ( n17229 & n17322 ) | ( n17311 & n17322 ) ;
  assign n17324 = n7296 & ~n16876 ;
  assign n17325 = n7879 & ~n16045 ;
  assign n17326 = n7300 & ~n16049 ;
  assign n17327 = n7299 & ~n16047 ;
  assign n17328 = n17326 | n17327 ;
  assign n17329 = ( ~n17324 & n17325 ) | ( ~n17324 & n17328 ) | ( n17325 & n17328 ) ;
  assign n17330 = ( ~x8 & n17324 ) | ( ~x8 & n17329 ) | ( n17324 & n17329 ) ;
  assign n17331 = ( n17324 & n17329 ) | ( n17324 & ~n17330 ) | ( n17329 & ~n17330 ) ;
  assign n17332 = ( x8 & n17330 ) | ( x8 & ~n17331 ) | ( n17330 & ~n17331 ) ;
  assign n17333 = n5966 & ~n16484 ;
  assign n17334 = n6464 & ~n16057 ;
  assign n17335 = n5970 & ~n16061 ;
  assign n17336 = n5969 & n16059 ;
  assign n17337 = n17335 | n17336 ;
  assign n17338 = ( ~n17333 & n17334 ) | ( ~n17333 & n17337 ) | ( n17334 & n17337 ) ;
  assign n17339 = ( ~x14 & n17333 ) | ( ~x14 & n17338 ) | ( n17333 & n17338 ) ;
  assign n17340 = ( n17333 & n17338 ) | ( n17333 & ~n17339 ) | ( n17338 & ~n17339 ) ;
  assign n17341 = ( x14 & n17339 ) | ( x14 & ~n17340 ) | ( n17339 & ~n17340 ) ;
  assign n17342 = n4974 & ~n16221 ;
  assign n17343 = n5398 & n16069 ;
  assign n17344 = n4973 & ~n16073 ;
  assign n17345 = n4972 & n16071 ;
  assign n17346 = n17344 | n17345 ;
  assign n17347 = ( ~n17342 & n17343 ) | ( ~n17342 & n17346 ) | ( n17343 & n17346 ) ;
  assign n17348 = ( ~x20 & n17342 ) | ( ~x20 & n17347 ) | ( n17342 & n17347 ) ;
  assign n17349 = ( n17342 & n17347 ) | ( n17342 & ~n17348 ) | ( n17347 & ~n17348 ) ;
  assign n17350 = ( x20 & n17348 ) | ( x20 & ~n17349 ) | ( n17348 & ~n17349 ) ;
  assign n17351 = x23 & ~n17264 ;
  assign n17352 = ~n17257 & n17351 ;
  assign n17353 = n4195 & ~n16081 ;
  assign n17354 = n4713 & n16169 ;
  assign n17355 = n4712 & ~n16075 ;
  assign n17356 = n4709 & ~n16079 ;
  assign n17357 = n4792 & n16077 ;
  assign n17358 = n17356 | n17357 ;
  assign n17359 = ( ~n17354 & n17355 ) | ( ~n17354 & n17358 ) | ( n17355 & n17358 ) ;
  assign n17360 = ( ~x23 & n17354 ) | ( ~x23 & n17359 ) | ( n17354 & n17359 ) ;
  assign n17361 = ( n17354 & n17359 ) | ( n17354 & ~n17360 ) | ( n17359 & ~n17360 ) ;
  assign n17362 = ( x23 & n17360 ) | ( x23 & ~n17361 ) | ( n17360 & ~n17361 ) ;
  assign n17363 = ( n17352 & n17353 ) | ( n17352 & n17362 ) | ( n17353 & n17362 ) ;
  assign n17364 = ( ~n17352 & n17353 ) | ( ~n17352 & n17362 ) | ( n17353 & n17362 ) ;
  assign n17365 = ( n17352 & ~n17363 ) | ( n17352 & n17364 ) | ( ~n17363 & n17364 ) ;
  assign n17366 = ( n17267 & n17350 ) | ( n17267 & n17365 ) | ( n17350 & n17365 ) ;
  assign n17367 = ( ~n17267 & n17350 ) | ( ~n17267 & n17365 ) | ( n17350 & n17365 ) ;
  assign n17368 = ( n17267 & ~n17366 ) | ( n17267 & n17367 ) | ( ~n17366 & n17367 ) ;
  assign n17369 = n5508 & n16315 ;
  assign n17370 = n5507 & n16063 ;
  assign n17371 = n5504 & n16067 ;
  assign n17372 = n5666 & n16065 ;
  assign n17373 = n17371 | n17372 ;
  assign n17374 = ( ~n17369 & n17370 ) | ( ~n17369 & n17373 ) | ( n17370 & n17373 ) ;
  assign n17375 = ( ~x17 & n17369 ) | ( ~x17 & n17374 ) | ( n17369 & n17374 ) ;
  assign n17376 = ( n17369 & n17374 ) | ( n17369 & ~n17375 ) | ( n17374 & ~n17375 ) ;
  assign n17377 = ( x17 & n17375 ) | ( x17 & ~n17376 ) | ( n17375 & ~n17376 ) ;
  assign n17378 = ( n17279 & n17368 ) | ( n17279 & n17377 ) | ( n17368 & n17377 ) ;
  assign n17379 = ( ~n17279 & n17368 ) | ( ~n17279 & n17377 ) | ( n17368 & n17377 ) ;
  assign n17380 = ( n17279 & ~n17378 ) | ( n17279 & n17379 ) | ( ~n17378 & n17379 ) ;
  assign n17381 = ( n17282 & n17341 ) | ( n17282 & n17380 ) | ( n17341 & n17380 ) ;
  assign n17382 = ( ~n17282 & n17341 ) | ( ~n17282 & n17380 ) | ( n17341 & n17380 ) ;
  assign n17383 = ( n17282 & ~n17381 ) | ( n17282 & n17382 ) | ( ~n17381 & n17382 ) ;
  assign n17384 = n6584 & n16611 ;
  assign n17385 = n7022 & ~n16051 ;
  assign n17386 = n6588 & ~n16055 ;
  assign n17387 = n6587 & n16053 ;
  assign n17388 = n17386 | n17387 ;
  assign n17389 = ( ~n17384 & n17385 ) | ( ~n17384 & n17388 ) | ( n17385 & n17388 ) ;
  assign n17390 = ( ~x11 & n17384 ) | ( ~x11 & n17389 ) | ( n17384 & n17389 ) ;
  assign n17391 = ( n17384 & n17389 ) | ( n17384 & ~n17390 ) | ( n17389 & ~n17390 ) ;
  assign n17392 = ( x11 & n17390 ) | ( x11 & ~n17391 ) | ( n17390 & ~n17391 ) ;
  assign n17393 = ( n17294 & n17383 ) | ( n17294 & n17392 ) | ( n17383 & n17392 ) ;
  assign n17394 = ( ~n17294 & n17383 ) | ( ~n17294 & n17392 ) | ( n17383 & n17392 ) ;
  assign n17395 = ( n17294 & ~n17393 ) | ( n17294 & n17394 ) | ( ~n17393 & n17394 ) ;
  assign n17396 = ( n17297 & n17332 ) | ( n17297 & n17395 ) | ( n17332 & n17395 ) ;
  assign n17397 = ( ~n17297 & n17332 ) | ( ~n17297 & n17395 ) | ( n17332 & n17395 ) ;
  assign n17398 = ( n17297 & ~n17396 ) | ( n17297 & n17397 ) | ( ~n17396 & n17397 ) ;
  assign n17399 = n8230 & ~n17051 ;
  assign n17400 = n8229 & n16039 ;
  assign n17401 = n8226 & ~n16043 ;
  assign n17402 = n8225 & n16041 ;
  assign n17403 = n17401 | n17402 ;
  assign n17404 = ( ~n17399 & n17400 ) | ( ~n17399 & n17403 ) | ( n17400 & n17403 ) ;
  assign n17405 = ( ~x5 & n17399 ) | ( ~x5 & n17404 ) | ( n17399 & n17404 ) ;
  assign n17406 = ( n17399 & n17404 ) | ( n17399 & ~n17405 ) | ( n17404 & ~n17405 ) ;
  assign n17407 = ( x5 & n17405 ) | ( x5 & ~n17406 ) | ( n17405 & ~n17406 ) ;
  assign n17408 = ( n17309 & n17398 ) | ( n17309 & n17407 ) | ( n17398 & n17407 ) ;
  assign n17409 = ( ~n17309 & n17398 ) | ( ~n17309 & n17407 ) | ( n17398 & n17407 ) ;
  assign n17410 = ( n17309 & ~n17408 ) | ( n17309 & n17409 ) | ( ~n17408 & n17409 ) ;
  assign n17411 = ( n16033 & ~n16035 ) | ( n16033 & n16105 ) | ( ~n16035 & n16105 ) ;
  assign n17412 = ( ~n16105 & n16106 ) | ( ~n16105 & n17411 ) | ( n16106 & n17411 ) ;
  assign n17413 = n36 & ~n17412 ;
  assign n17414 = n8967 & ~n16037 ;
  assign n17415 = ( x0 & n8966 ) | ( x0 & ~n16035 ) | ( n8966 & ~n16035 ) ;
  assign n17416 = ( n8966 & n17414 ) | ( n8966 & ~n17415 ) | ( n17414 & ~n17415 ) ;
  assign n17417 = n35 & n16033 ;
  assign n17418 = ( n35 & n17416 ) | ( n35 & ~n17417 ) | ( n17416 & ~n17417 ) ;
  assign n17419 = ( ~x2 & n17413 ) | ( ~x2 & n17418 ) | ( n17413 & n17418 ) ;
  assign n17420 = ( n17413 & n17418 ) | ( n17413 & ~n17419 ) | ( n17418 & ~n17419 ) ;
  assign n17421 = ( x2 & n17419 ) | ( x2 & ~n17420 ) | ( n17419 & ~n17420 ) ;
  assign n17422 = ( n17323 & n17410 ) | ( n17323 & n17421 ) | ( n17410 & n17421 ) ;
  assign n17423 = n7296 & ~n16957 ;
  assign n17424 = n7879 & ~n16043 ;
  assign n17425 = n7300 & ~n16047 ;
  assign n17426 = n7299 & ~n16045 ;
  assign n17427 = n17425 | n17426 ;
  assign n17428 = ( ~n17423 & n17424 ) | ( ~n17423 & n17427 ) | ( n17424 & n17427 ) ;
  assign n17429 = ( ~x8 & n17423 ) | ( ~x8 & n17428 ) | ( n17423 & n17428 ) ;
  assign n17430 = ( n17423 & n17428 ) | ( n17423 & ~n17429 ) | ( n17428 & ~n17429 ) ;
  assign n17431 = ( x8 & n17429 ) | ( x8 & ~n17430 ) | ( n17429 & ~n17430 ) ;
  assign n17432 = n5966 & n16541 ;
  assign n17433 = n6464 & ~n16055 ;
  assign n17434 = n5970 & n16059 ;
  assign n17435 = n5969 & ~n16057 ;
  assign n17436 = n17434 | n17435 ;
  assign n17437 = ( ~n17432 & n17433 ) | ( ~n17432 & n17436 ) | ( n17433 & n17436 ) ;
  assign n17438 = ( ~x14 & n17432 ) | ( ~x14 & n17437 ) | ( n17432 & n17437 ) ;
  assign n17439 = ( n17432 & n17437 ) | ( n17432 & ~n17438 ) | ( n17437 & ~n17438 ) ;
  assign n17440 = ( x14 & n17438 ) | ( x14 & ~n17439 ) | ( n17438 & ~n17439 ) ;
  assign n17441 = n4974 & n16269 ;
  assign n17442 = n5398 & n16067 ;
  assign n17443 = n4973 & n16071 ;
  assign n17444 = n4972 & n16069 ;
  assign n17445 = n17443 | n17444 ;
  assign n17446 = ( ~n17441 & n17442 ) | ( ~n17441 & n17445 ) | ( n17442 & n17445 ) ;
  assign n17447 = ( ~x20 & n17441 ) | ( ~x20 & n17446 ) | ( n17441 & n17446 ) ;
  assign n17448 = ( n17441 & n17446 ) | ( n17441 & ~n17447 ) | ( n17446 & ~n17447 ) ;
  assign n17449 = ( x20 & n17447 ) | ( x20 & ~n17448 ) | ( n17447 & ~n17448 ) ;
  assign n17450 = n4713 & ~n16176 ;
  assign n17451 = n4712 & ~n16073 ;
  assign n17452 = n4709 & n16077 ;
  assign n17453 = n4792 & ~n16075 ;
  assign n17454 = n17452 | n17453 ;
  assign n17455 = ( ~n17450 & n17451 ) | ( ~n17450 & n17454 ) | ( n17451 & n17454 ) ;
  assign n17456 = ( ~x23 & n17450 ) | ( ~x23 & n17455 ) | ( n17450 & n17455 ) ;
  assign n17457 = ( n17450 & n17455 ) | ( n17450 & ~n17456 ) | ( n17455 & ~n17456 ) ;
  assign n17458 = ( x23 & n17456 ) | ( x23 & ~n17457 ) | ( n17456 & ~n17457 ) ;
  assign n17459 = x26 & n17353 ;
  assign n17460 = ( n4202 & n16155 ) | ( n4202 & n16187 ) | ( n16155 & n16187 ) ;
  assign n17461 = n4345 & ~n16081 ;
  assign n17462 = n4201 & ~n16079 ;
  assign n17463 = n17461 | n17462 ;
  assign n17464 = ( ~n17459 & n17460 ) | ( ~n17459 & n17463 ) | ( n17460 & n17463 ) ;
  assign n17465 = ( n17460 & n17463 ) | ( n17460 & ~n17464 ) | ( n17463 & ~n17464 ) ;
  assign n17466 = ( n17459 & n17464 ) | ( n17459 & ~n17465 ) | ( n17464 & ~n17465 ) ;
  assign n17467 = ( n17363 & n17458 ) | ( n17363 & n17466 ) | ( n17458 & n17466 ) ;
  assign n17468 = ( ~n17363 & n17458 ) | ( ~n17363 & n17466 ) | ( n17458 & n17466 ) ;
  assign n17469 = ( n17363 & ~n17467 ) | ( n17363 & n17468 ) | ( ~n17467 & n17468 ) ;
  assign n17470 = ( n17366 & n17449 ) | ( n17366 & n17469 ) | ( n17449 & n17469 ) ;
  assign n17471 = ( ~n17366 & n17449 ) | ( ~n17366 & n17469 ) | ( n17449 & n17469 ) ;
  assign n17472 = ( n17366 & ~n17470 ) | ( n17366 & n17471 ) | ( ~n17470 & n17471 ) ;
  assign n17473 = n5508 & ~n16354 ;
  assign n17474 = n5507 & ~n16061 ;
  assign n17475 = n5504 & n16065 ;
  assign n17476 = n5666 & n16063 ;
  assign n17477 = n17475 | n17476 ;
  assign n17478 = ( ~n17473 & n17474 ) | ( ~n17473 & n17477 ) | ( n17474 & n17477 ) ;
  assign n17479 = ( ~x17 & n17473 ) | ( ~x17 & n17478 ) | ( n17473 & n17478 ) ;
  assign n17480 = ( n17473 & n17478 ) | ( n17473 & ~n17479 ) | ( n17478 & ~n17479 ) ;
  assign n17481 = ( x17 & n17479 ) | ( x17 & ~n17480 ) | ( n17479 & ~n17480 ) ;
  assign n17482 = ( n17378 & n17472 ) | ( n17378 & n17481 ) | ( n17472 & n17481 ) ;
  assign n17483 = ( ~n17378 & n17472 ) | ( ~n17378 & n17481 ) | ( n17472 & n17481 ) ;
  assign n17484 = ( n17378 & ~n17482 ) | ( n17378 & n17483 ) | ( ~n17482 & n17483 ) ;
  assign n17485 = ( n17381 & n17440 ) | ( n17381 & n17484 ) | ( n17440 & n17484 ) ;
  assign n17486 = ( ~n17381 & n17440 ) | ( ~n17381 & n17484 ) | ( n17440 & n17484 ) ;
  assign n17487 = ( n17381 & ~n17485 ) | ( n17381 & n17486 ) | ( ~n17485 & n17486 ) ;
  assign n17488 = n6584 & ~n16674 ;
  assign n17489 = n7022 & ~n16049 ;
  assign n17490 = n6588 & n16053 ;
  assign n17491 = n6587 & ~n16051 ;
  assign n17492 = n17490 | n17491 ;
  assign n17493 = ( ~n17488 & n17489 ) | ( ~n17488 & n17492 ) | ( n17489 & n17492 ) ;
  assign n17494 = ( ~x11 & n17488 ) | ( ~x11 & n17493 ) | ( n17488 & n17493 ) ;
  assign n17495 = ( n17488 & n17493 ) | ( n17488 & ~n17494 ) | ( n17493 & ~n17494 ) ;
  assign n17496 = ( x11 & n17494 ) | ( x11 & ~n17495 ) | ( n17494 & ~n17495 ) ;
  assign n17497 = ( n17393 & n17487 ) | ( n17393 & n17496 ) | ( n17487 & n17496 ) ;
  assign n17498 = ( ~n17393 & n17487 ) | ( ~n17393 & n17496 ) | ( n17487 & n17496 ) ;
  assign n17499 = ( n17393 & ~n17497 ) | ( n17393 & n17498 ) | ( ~n17497 & n17498 ) ;
  assign n17500 = ( n17396 & n17431 ) | ( n17396 & n17499 ) | ( n17431 & n17499 ) ;
  assign n17501 = ( ~n17396 & n17431 ) | ( ~n17396 & n17499 ) | ( n17431 & n17499 ) ;
  assign n17502 = ( n17396 & ~n17500 ) | ( n17396 & n17501 ) | ( ~n17500 & n17501 ) ;
  assign n17503 = n8230 & ~n17138 ;
  assign n17504 = n8229 & ~n16037 ;
  assign n17505 = n8226 & n16041 ;
  assign n17506 = n8225 & n16039 ;
  assign n17507 = n17505 | n17506 ;
  assign n17508 = ( ~n17503 & n17504 ) | ( ~n17503 & n17507 ) | ( n17504 & n17507 ) ;
  assign n17509 = ( ~x5 & n17503 ) | ( ~x5 & n17508 ) | ( n17503 & n17508 ) ;
  assign n17510 = ( n17503 & n17508 ) | ( n17503 & ~n17509 ) | ( n17508 & ~n17509 ) ;
  assign n17511 = ( x5 & n17509 ) | ( x5 & ~n17510 ) | ( n17509 & ~n17510 ) ;
  assign n17512 = ( n17408 & n17502 ) | ( n17408 & n17511 ) | ( n17502 & n17511 ) ;
  assign n17513 = ( ~n17408 & n17502 ) | ( ~n17408 & n17511 ) | ( n17502 & n17511 ) ;
  assign n17514 = ( n17408 & ~n17512 ) | ( n17408 & n17513 ) | ( ~n17512 & n17513 ) ;
  assign n17515 = ( ~n16031 & n16033 ) | ( ~n16031 & n16106 ) | ( n16033 & n16106 ) ;
  assign n17516 = ( ~n16106 & n16107 ) | ( ~n16106 & n17515 ) | ( n16107 & n17515 ) ;
  assign n17517 = n36 & ~n17516 ;
  assign n17518 = n8967 & n16035 ;
  assign n17519 = ( x0 & n8966 ) | ( x0 & n16033 ) | ( n8966 & n16033 ) ;
  assign n17520 = ( n8966 & n17518 ) | ( n8966 & ~n17519 ) | ( n17518 & ~n17519 ) ;
  assign n17521 = n35 & ~n16031 ;
  assign n17522 = ( n35 & n17520 ) | ( n35 & ~n17521 ) | ( n17520 & ~n17521 ) ;
  assign n17523 = ( ~x2 & n17517 ) | ( ~x2 & n17522 ) | ( n17517 & n17522 ) ;
  assign n17524 = ( n17517 & n17522 ) | ( n17517 & ~n17523 ) | ( n17522 & ~n17523 ) ;
  assign n17525 = ( x2 & n17523 ) | ( x2 & ~n17524 ) | ( n17523 & ~n17524 ) ;
  assign n17526 = ( n17422 & n17514 ) | ( n17422 & n17525 ) | ( n17514 & n17525 ) ;
  assign n17527 = ( n16029 & ~n16031 ) | ( n16029 & n16107 ) | ( ~n16031 & n16107 ) ;
  assign n17528 = ( ~n16107 & n16108 ) | ( ~n16107 & n17527 ) | ( n16108 & n17527 ) ;
  assign n17529 = n36 & ~n17528 ;
  assign n17530 = n8967 & ~n16033 ;
  assign n17531 = ( x0 & n8966 ) | ( x0 & ~n16031 ) | ( n8966 & ~n16031 ) ;
  assign n17532 = ( n8966 & n17530 ) | ( n8966 & ~n17531 ) | ( n17530 & ~n17531 ) ;
  assign n17533 = n35 & n16029 ;
  assign n17534 = ( n35 & n17532 ) | ( n35 & ~n17533 ) | ( n17532 & ~n17533 ) ;
  assign n17535 = ( ~x2 & n17529 ) | ( ~x2 & n17534 ) | ( n17529 & n17534 ) ;
  assign n17536 = ( n17529 & n17534 ) | ( n17529 & ~n17535 ) | ( n17534 & ~n17535 ) ;
  assign n17537 = ( x2 & n17535 ) | ( x2 & ~n17536 ) | ( n17535 & ~n17536 ) ;
  assign n17538 = n8230 & ~n17313 ;
  assign n17539 = n8229 & n16035 ;
  assign n17540 = n8226 & n16039 ;
  assign n17541 = n8225 & ~n16037 ;
  assign n17542 = n17540 | n17541 ;
  assign n17543 = ( ~n17538 & n17539 ) | ( ~n17538 & n17542 ) | ( n17539 & n17542 ) ;
  assign n17544 = ( ~x5 & n17538 ) | ( ~x5 & n17543 ) | ( n17538 & n17543 ) ;
  assign n17545 = ( n17538 & n17543 ) | ( n17538 & ~n17544 ) | ( n17543 & ~n17544 ) ;
  assign n17546 = ( x5 & n17544 ) | ( x5 & ~n17545 ) | ( n17544 & ~n17545 ) ;
  assign n17547 = n6584 & ~n16801 ;
  assign n17548 = n7022 & ~n16047 ;
  assign n17549 = n6588 & ~n16051 ;
  assign n17550 = n6587 & ~n16049 ;
  assign n17551 = n17549 | n17550 ;
  assign n17552 = ( ~n17547 & n17548 ) | ( ~n17547 & n17551 ) | ( n17548 & n17551 ) ;
  assign n17553 = ( ~x11 & n17547 ) | ( ~x11 & n17552 ) | ( n17547 & n17552 ) ;
  assign n17554 = ( n17547 & n17552 ) | ( n17547 & ~n17553 ) | ( n17552 & ~n17553 ) ;
  assign n17555 = ( x11 & n17553 ) | ( x11 & ~n17554 ) | ( n17553 & ~n17554 ) ;
  assign n17556 = n5508 & ~n16433 ;
  assign n17557 = n5507 & n16059 ;
  assign n17558 = n5504 & n16063 ;
  assign n17559 = n5666 & ~n16061 ;
  assign n17560 = n17558 | n17559 ;
  assign n17561 = ( ~n17556 & n17557 ) | ( ~n17556 & n17560 ) | ( n17557 & n17560 ) ;
  assign n17562 = ( ~x17 & n17556 ) | ( ~x17 & n17561 ) | ( n17556 & n17561 ) ;
  assign n17563 = ( n17556 & n17561 ) | ( n17556 & ~n17562 ) | ( n17561 & ~n17562 ) ;
  assign n17564 = ( x17 & n17562 ) | ( x17 & ~n17563 ) | ( n17562 & ~n17563 ) ;
  assign n17565 = n4713 & n16209 ;
  assign n17566 = n4712 & n16071 ;
  assign n17567 = n4709 & ~n16075 ;
  assign n17568 = n4792 & ~n16073 ;
  assign n17569 = n17567 | n17568 ;
  assign n17570 = ( ~n17565 & n17566 ) | ( ~n17565 & n17569 ) | ( n17566 & n17569 ) ;
  assign n17571 = ( ~x23 & n17565 ) | ( ~x23 & n17570 ) | ( n17565 & n17570 ) ;
  assign n17572 = ( n17565 & n17570 ) | ( n17565 & ~n17571 ) | ( n17570 & ~n17571 ) ;
  assign n17573 = ( x23 & n17571 ) | ( x23 & ~n17572 ) | ( n17571 & ~n17572 ) ;
  assign n17574 = ( x26 & n17459 ) | ( x26 & n17464 ) | ( n17459 & n17464 ) ;
  assign n17575 = ( n4202 & n16083 ) | ( n4202 & n16198 ) | ( n16083 & n16198 ) ;
  assign n17576 = n4200 & ~n16081 ;
  assign n17577 = n4345 & ~n16079 ;
  assign n17578 = n17576 | n17577 ;
  assign n17579 = n4201 & ~n16077 ;
  assign n17580 = ( n4201 & n17578 ) | ( n4201 & ~n17579 ) | ( n17578 & ~n17579 ) ;
  assign n17581 = ( ~n17574 & n17575 ) | ( ~n17574 & n17580 ) | ( n17575 & n17580 ) ;
  assign n17582 = ( n17575 & n17580 ) | ( n17575 & ~n17581 ) | ( n17580 & ~n17581 ) ;
  assign n17583 = ( n17574 & n17581 ) | ( n17574 & ~n17582 ) | ( n17581 & ~n17582 ) ;
  assign n17584 = ( n17467 & n17573 ) | ( n17467 & n17583 ) | ( n17573 & n17583 ) ;
  assign n17585 = ( ~n17467 & n17573 ) | ( ~n17467 & n17583 ) | ( n17573 & n17583 ) ;
  assign n17586 = ( n17467 & ~n17584 ) | ( n17467 & n17585 ) | ( ~n17584 & n17585 ) ;
  assign n17587 = n4974 & n16281 ;
  assign n17588 = n5398 & n16065 ;
  assign n17589 = n4973 & n16069 ;
  assign n17590 = n4972 & n16067 ;
  assign n17591 = n17589 | n17590 ;
  assign n17592 = ( ~n17587 & n17588 ) | ( ~n17587 & n17591 ) | ( n17588 & n17591 ) ;
  assign n17593 = ( ~x20 & n17587 ) | ( ~x20 & n17592 ) | ( n17587 & n17592 ) ;
  assign n17594 = ( n17587 & n17592 ) | ( n17587 & ~n17593 ) | ( n17592 & ~n17593 ) ;
  assign n17595 = ( x20 & n17593 ) | ( x20 & ~n17594 ) | ( n17593 & ~n17594 ) ;
  assign n17596 = ( n17470 & n17586 ) | ( n17470 & n17595 ) | ( n17586 & n17595 ) ;
  assign n17597 = ( ~n17470 & n17586 ) | ( ~n17470 & n17595 ) | ( n17586 & n17595 ) ;
  assign n17598 = ( n17470 & ~n17596 ) | ( n17470 & n17597 ) | ( ~n17596 & n17597 ) ;
  assign n17599 = ( n17482 & n17564 ) | ( n17482 & n17598 ) | ( n17564 & n17598 ) ;
  assign n17600 = ( ~n17482 & n17564 ) | ( ~n17482 & n17598 ) | ( n17564 & n17598 ) ;
  assign n17601 = ( n17482 & ~n17599 ) | ( n17482 & n17600 ) | ( ~n17599 & n17600 ) ;
  assign n17602 = n5966 & n16553 ;
  assign n17603 = n6464 & n16053 ;
  assign n17604 = n5970 & ~n16057 ;
  assign n17605 = n5969 & ~n16055 ;
  assign n17606 = n17604 | n17605 ;
  assign n17607 = ( ~n17602 & n17603 ) | ( ~n17602 & n17606 ) | ( n17603 & n17606 ) ;
  assign n17608 = ( ~x14 & n17602 ) | ( ~x14 & n17607 ) | ( n17602 & n17607 ) ;
  assign n17609 = ( n17602 & n17607 ) | ( n17602 & ~n17608 ) | ( n17607 & ~n17608 ) ;
  assign n17610 = ( x14 & n17608 ) | ( x14 & ~n17609 ) | ( n17608 & ~n17609 ) ;
  assign n17611 = ( n17485 & n17601 ) | ( n17485 & n17610 ) | ( n17601 & n17610 ) ;
  assign n17612 = ( ~n17485 & n17601 ) | ( ~n17485 & n17610 ) | ( n17601 & n17610 ) ;
  assign n17613 = ( n17485 & ~n17611 ) | ( n17485 & n17612 ) | ( ~n17611 & n17612 ) ;
  assign n17614 = ( n17497 & n17555 ) | ( n17497 & n17613 ) | ( n17555 & n17613 ) ;
  assign n17615 = ( ~n17497 & n17555 ) | ( ~n17497 & n17613 ) | ( n17555 & n17613 ) ;
  assign n17616 = ( n17497 & ~n17614 ) | ( n17497 & n17615 ) | ( ~n17614 & n17615 ) ;
  assign n17617 = n7296 & n16969 ;
  assign n17618 = n7879 & n16041 ;
  assign n17619 = n7300 & ~n16045 ;
  assign n17620 = n7299 & ~n16043 ;
  assign n17621 = n17619 | n17620 ;
  assign n17622 = ( ~n17617 & n17618 ) | ( ~n17617 & n17621 ) | ( n17618 & n17621 ) ;
  assign n17623 = ( ~x8 & n17617 ) | ( ~x8 & n17622 ) | ( n17617 & n17622 ) ;
  assign n17624 = ( n17617 & n17622 ) | ( n17617 & ~n17623 ) | ( n17622 & ~n17623 ) ;
  assign n17625 = ( x8 & n17623 ) | ( x8 & ~n17624 ) | ( n17623 & ~n17624 ) ;
  assign n17626 = ( n17500 & n17616 ) | ( n17500 & n17625 ) | ( n17616 & n17625 ) ;
  assign n17627 = ( ~n17500 & n17616 ) | ( ~n17500 & n17625 ) | ( n17616 & n17625 ) ;
  assign n17628 = ( n17500 & ~n17626 ) | ( n17500 & n17627 ) | ( ~n17626 & n17627 ) ;
  assign n17629 = ( n17512 & n17546 ) | ( n17512 & n17628 ) | ( n17546 & n17628 ) ;
  assign n17630 = ( ~n17512 & n17546 ) | ( ~n17512 & n17628 ) | ( n17546 & n17628 ) ;
  assign n17631 = ( n17512 & ~n17629 ) | ( n17512 & n17630 ) | ( ~n17629 & n17630 ) ;
  assign n17632 = ( n17526 & n17537 ) | ( n17526 & n17631 ) | ( n17537 & n17631 ) ;
  assign n17633 = ( ~n16027 & n16031 ) | ( ~n16027 & n17527 ) | ( n16031 & n17527 ) ;
  assign n17634 = ( ~n16029 & n16109 ) | ( ~n16029 & n17633 ) | ( n16109 & n17633 ) ;
  assign n17635 = n36 & n17634 ;
  assign n17636 = n8967 & n16031 ;
  assign n17637 = ( x0 & n8966 ) | ( x0 & n16029 ) | ( n8966 & n16029 ) ;
  assign n17638 = ( n8966 & n17636 ) | ( n8966 & ~n17637 ) | ( n17636 & ~n17637 ) ;
  assign n17639 = n35 & n16027 ;
  assign n17640 = ( n35 & n17638 ) | ( n35 & ~n17639 ) | ( n17638 & ~n17639 ) ;
  assign n17641 = ( ~x2 & n17635 ) | ( ~x2 & n17640 ) | ( n17635 & n17640 ) ;
  assign n17642 = ( n17635 & n17640 ) | ( n17635 & ~n17641 ) | ( n17640 & ~n17641 ) ;
  assign n17643 = ( x2 & n17641 ) | ( x2 & ~n17642 ) | ( n17641 & ~n17642 ) ;
  assign n17644 = n8230 & ~n17412 ;
  assign n17645 = n8229 & ~n16033 ;
  assign n17646 = n8226 & ~n16037 ;
  assign n17647 = n8225 & n16035 ;
  assign n17648 = n17646 | n17647 ;
  assign n17649 = ( ~n17644 & n17645 ) | ( ~n17644 & n17648 ) | ( n17645 & n17648 ) ;
  assign n17650 = ( ~x5 & n17644 ) | ( ~x5 & n17649 ) | ( n17644 & n17649 ) ;
  assign n17651 = ( n17644 & n17649 ) | ( n17644 & ~n17650 ) | ( n17649 & ~n17650 ) ;
  assign n17652 = ( x5 & n17650 ) | ( x5 & ~n17651 ) | ( n17650 & ~n17651 ) ;
  assign n17653 = n6584 & ~n16876 ;
  assign n17654 = n7022 & ~n16045 ;
  assign n17655 = n6588 & ~n16049 ;
  assign n17656 = n6587 & ~n16047 ;
  assign n17657 = n17655 | n17656 ;
  assign n17658 = ( ~n17653 & n17654 ) | ( ~n17653 & n17657 ) | ( n17654 & n17657 ) ;
  assign n17659 = ( ~x11 & n17653 ) | ( ~x11 & n17658 ) | ( n17653 & n17658 ) ;
  assign n17660 = ( n17653 & n17658 ) | ( n17653 & ~n17659 ) | ( n17658 & ~n17659 ) ;
  assign n17661 = ( x11 & n17659 ) | ( x11 & ~n17660 ) | ( n17659 & ~n17660 ) ;
  assign n17662 = n5508 & ~n16484 ;
  assign n17663 = n5507 & ~n16057 ;
  assign n17664 = n5504 & ~n16061 ;
  assign n17665 = n5666 & n16059 ;
  assign n17666 = n17664 | n17665 ;
  assign n17667 = ( ~n17662 & n17663 ) | ( ~n17662 & n17666 ) | ( n17663 & n17666 ) ;
  assign n17668 = ( ~x17 & n17662 ) | ( ~x17 & n17667 ) | ( n17662 & n17667 ) ;
  assign n17669 = ( n17662 & n17667 ) | ( n17662 & ~n17668 ) | ( n17667 & ~n17668 ) ;
  assign n17670 = ( x17 & n17668 ) | ( x17 & ~n17669 ) | ( n17668 & ~n17669 ) ;
  assign n17671 = n4713 & ~n16221 ;
  assign n17672 = n4712 & n16069 ;
  assign n17673 = n4709 & ~n16073 ;
  assign n17674 = n4792 & n16071 ;
  assign n17675 = n17673 | n17674 ;
  assign n17676 = ( ~n17671 & n17672 ) | ( ~n17671 & n17675 ) | ( n17672 & n17675 ) ;
  assign n17677 = ( ~x23 & n17671 ) | ( ~x23 & n17676 ) | ( n17671 & n17676 ) ;
  assign n17678 = ( n17671 & n17676 ) | ( n17671 & ~n17677 ) | ( n17676 & ~n17677 ) ;
  assign n17679 = ( x23 & n17677 ) | ( x23 & ~n17678 ) | ( n17677 & ~n17678 ) ;
  assign n17680 = n3697 & ~n16081 ;
  assign n17681 = n4202 & n16169 ;
  assign n17682 = n4201 & ~n16075 ;
  assign n17683 = n4200 & ~n16079 ;
  assign n17684 = n4345 & n16077 ;
  assign n17685 = n17683 | n17684 ;
  assign n17686 = ( ~n17681 & n17682 ) | ( ~n17681 & n17685 ) | ( n17682 & n17685 ) ;
  assign n17687 = ( ~x26 & n17681 ) | ( ~x26 & n17686 ) | ( n17681 & n17686 ) ;
  assign n17688 = ( n17681 & n17686 ) | ( n17681 & ~n17687 ) | ( n17686 & ~n17687 ) ;
  assign n17689 = ( x26 & n17687 ) | ( x26 & ~n17688 ) | ( n17687 & ~n17688 ) ;
  assign n17690 = x26 & ~n17574 ;
  assign n17691 = ( ~n17575 & n17580 ) | ( ~n17575 & n17690 ) | ( n17580 & n17690 ) ;
  assign n17692 = ~n17580 & n17691 ;
  assign n17693 = ( n17680 & n17689 ) | ( n17680 & n17692 ) | ( n17689 & n17692 ) ;
  assign n17694 = ( ~n17680 & n17689 ) | ( ~n17680 & n17692 ) | ( n17689 & n17692 ) ;
  assign n17695 = ( n17680 & ~n17693 ) | ( n17680 & n17694 ) | ( ~n17693 & n17694 ) ;
  assign n17696 = ( n17584 & n17679 ) | ( n17584 & n17695 ) | ( n17679 & n17695 ) ;
  assign n17697 = ( ~n17584 & n17679 ) | ( ~n17584 & n17695 ) | ( n17679 & n17695 ) ;
  assign n17698 = ( n17584 & ~n17696 ) | ( n17584 & n17697 ) | ( ~n17696 & n17697 ) ;
  assign n17699 = n4974 & n16315 ;
  assign n17700 = n5398 & n16063 ;
  assign n17701 = n4973 & n16067 ;
  assign n17702 = n4972 & n16065 ;
  assign n17703 = n17701 | n17702 ;
  assign n17704 = ( ~n17699 & n17700 ) | ( ~n17699 & n17703 ) | ( n17700 & n17703 ) ;
  assign n17705 = ( ~x20 & n17699 ) | ( ~x20 & n17704 ) | ( n17699 & n17704 ) ;
  assign n17706 = ( n17699 & n17704 ) | ( n17699 & ~n17705 ) | ( n17704 & ~n17705 ) ;
  assign n17707 = ( x20 & n17705 ) | ( x20 & ~n17706 ) | ( n17705 & ~n17706 ) ;
  assign n17708 = ( n17596 & n17698 ) | ( n17596 & n17707 ) | ( n17698 & n17707 ) ;
  assign n17709 = ( ~n17596 & n17698 ) | ( ~n17596 & n17707 ) | ( n17698 & n17707 ) ;
  assign n17710 = ( n17596 & ~n17708 ) | ( n17596 & n17709 ) | ( ~n17708 & n17709 ) ;
  assign n17711 = ( n17599 & n17670 ) | ( n17599 & n17710 ) | ( n17670 & n17710 ) ;
  assign n17712 = ( ~n17599 & n17670 ) | ( ~n17599 & n17710 ) | ( n17670 & n17710 ) ;
  assign n17713 = ( n17599 & ~n17711 ) | ( n17599 & n17712 ) | ( ~n17711 & n17712 ) ;
  assign n17714 = n5966 & n16611 ;
  assign n17715 = n6464 & ~n16051 ;
  assign n17716 = n5970 & ~n16055 ;
  assign n17717 = n5969 & n16053 ;
  assign n17718 = n17716 | n17717 ;
  assign n17719 = ( ~n17714 & n17715 ) | ( ~n17714 & n17718 ) | ( n17715 & n17718 ) ;
  assign n17720 = ( ~x14 & n17714 ) | ( ~x14 & n17719 ) | ( n17714 & n17719 ) ;
  assign n17721 = ( n17714 & n17719 ) | ( n17714 & ~n17720 ) | ( n17719 & ~n17720 ) ;
  assign n17722 = ( x14 & n17720 ) | ( x14 & ~n17721 ) | ( n17720 & ~n17721 ) ;
  assign n17723 = ( n17611 & n17713 ) | ( n17611 & n17722 ) | ( n17713 & n17722 ) ;
  assign n17724 = ( ~n17611 & n17713 ) | ( ~n17611 & n17722 ) | ( n17713 & n17722 ) ;
  assign n17725 = ( n17611 & ~n17723 ) | ( n17611 & n17724 ) | ( ~n17723 & n17724 ) ;
  assign n17726 = ( n17614 & n17661 ) | ( n17614 & n17725 ) | ( n17661 & n17725 ) ;
  assign n17727 = ( ~n17614 & n17661 ) | ( ~n17614 & n17725 ) | ( n17661 & n17725 ) ;
  assign n17728 = ( n17614 & ~n17726 ) | ( n17614 & n17727 ) | ( ~n17726 & n17727 ) ;
  assign n17729 = n7296 & ~n17051 ;
  assign n17730 = n7879 & n16039 ;
  assign n17731 = n7300 & ~n16043 ;
  assign n17732 = n7299 & n16041 ;
  assign n17733 = n17731 | n17732 ;
  assign n17734 = ( ~n17729 & n17730 ) | ( ~n17729 & n17733 ) | ( n17730 & n17733 ) ;
  assign n17735 = ( ~x8 & n17729 ) | ( ~x8 & n17734 ) | ( n17729 & n17734 ) ;
  assign n17736 = ( n17729 & n17734 ) | ( n17729 & ~n17735 ) | ( n17734 & ~n17735 ) ;
  assign n17737 = ( x8 & n17735 ) | ( x8 & ~n17736 ) | ( n17735 & ~n17736 ) ;
  assign n17738 = ( n17626 & n17728 ) | ( n17626 & n17737 ) | ( n17728 & n17737 ) ;
  assign n17739 = ( ~n17626 & n17728 ) | ( ~n17626 & n17737 ) | ( n17728 & n17737 ) ;
  assign n17740 = ( n17626 & ~n17738 ) | ( n17626 & n17739 ) | ( ~n17738 & n17739 ) ;
  assign n17741 = ( n17629 & n17652 ) | ( n17629 & n17740 ) | ( n17652 & n17740 ) ;
  assign n17742 = ( ~n17629 & n17652 ) | ( ~n17629 & n17740 ) | ( n17652 & n17740 ) ;
  assign n17743 = ( n17629 & ~n17741 ) | ( n17629 & n17742 ) | ( ~n17741 & n17742 ) ;
  assign n17744 = ( n17632 & n17643 ) | ( n17632 & n17743 ) | ( n17643 & n17743 ) ;
  assign n17745 = ( n16025 & n16108 ) | ( n16025 & ~n17633 ) | ( n16108 & ~n17633 ) ;
  assign n17746 = ( n16109 & ~n16110 ) | ( n16109 & n17745 ) | ( ~n16110 & n17745 ) ;
  assign n17747 = n36 & ~n17746 ;
  assign n17748 = n8967 & ~n16029 ;
  assign n17749 = ( x0 & n8966 ) | ( x0 & n16027 ) | ( n8966 & n16027 ) ;
  assign n17750 = ( n8966 & n17748 ) | ( n8966 & ~n17749 ) | ( n17748 & ~n17749 ) ;
  assign n17751 = n35 & n16025 ;
  assign n17752 = ( n35 & n17750 ) | ( n35 & ~n17751 ) | ( n17750 & ~n17751 ) ;
  assign n17753 = ( ~x2 & n17747 ) | ( ~x2 & n17752 ) | ( n17747 & n17752 ) ;
  assign n17754 = ( n17747 & n17752 ) | ( n17747 & ~n17753 ) | ( n17752 & ~n17753 ) ;
  assign n17755 = ( x2 & n17753 ) | ( x2 & ~n17754 ) | ( n17753 & ~n17754 ) ;
  assign n17756 = n8230 & ~n17516 ;
  assign n17757 = n8229 & n16031 ;
  assign n17758 = n8226 & n16035 ;
  assign n17759 = n8225 & ~n16033 ;
  assign n17760 = n17758 | n17759 ;
  assign n17761 = ( ~n17756 & n17757 ) | ( ~n17756 & n17760 ) | ( n17757 & n17760 ) ;
  assign n17762 = ( ~x5 & n17756 ) | ( ~x5 & n17761 ) | ( n17756 & n17761 ) ;
  assign n17763 = ( n17756 & n17761 ) | ( n17756 & ~n17762 ) | ( n17761 & ~n17762 ) ;
  assign n17764 = ( x5 & n17762 ) | ( x5 & ~n17763 ) | ( n17762 & ~n17763 ) ;
  assign n17765 = n6584 & ~n16957 ;
  assign n17766 = n7022 & ~n16043 ;
  assign n17767 = n6588 & ~n16047 ;
  assign n17768 = n6587 & ~n16045 ;
  assign n17769 = n17767 | n17768 ;
  assign n17770 = ( ~n17765 & n17766 ) | ( ~n17765 & n17769 ) | ( n17766 & n17769 ) ;
  assign n17771 = ( ~x11 & n17765 ) | ( ~x11 & n17770 ) | ( n17765 & n17770 ) ;
  assign n17772 = ( n17765 & n17770 ) | ( n17765 & ~n17771 ) | ( n17770 & ~n17771 ) ;
  assign n17773 = ( x11 & n17771 ) | ( x11 & ~n17772 ) | ( n17771 & ~n17772 ) ;
  assign n17774 = n5508 & n16541 ;
  assign n17775 = n5507 & ~n16055 ;
  assign n17776 = n5504 & n16059 ;
  assign n17777 = n5666 & ~n16057 ;
  assign n17778 = n17776 | n17777 ;
  assign n17779 = ( ~n17774 & n17775 ) | ( ~n17774 & n17778 ) | ( n17775 & n17778 ) ;
  assign n17780 = ( ~x17 & n17774 ) | ( ~x17 & n17779 ) | ( n17774 & n17779 ) ;
  assign n17781 = ( n17774 & n17779 ) | ( n17774 & ~n17780 ) | ( n17779 & ~n17780 ) ;
  assign n17782 = ( x17 & n17780 ) | ( x17 & ~n17781 ) | ( n17780 & ~n17781 ) ;
  assign n17783 = n4713 & n16269 ;
  assign n17784 = n4712 & n16067 ;
  assign n17785 = n4709 & n16071 ;
  assign n17786 = n4792 & n16069 ;
  assign n17787 = n17785 | n17786 ;
  assign n17788 = ( ~n17783 & n17784 ) | ( ~n17783 & n17787 ) | ( n17784 & n17787 ) ;
  assign n17789 = ( ~x23 & n17783 ) | ( ~x23 & n17788 ) | ( n17783 & n17788 ) ;
  assign n17790 = ( n17783 & n17788 ) | ( n17783 & ~n17789 ) | ( n17788 & ~n17789 ) ;
  assign n17791 = ( x23 & n17789 ) | ( x23 & ~n17790 ) | ( n17789 & ~n17790 ) ;
  assign n17792 = x29 & n17680 ;
  assign n17793 = ( n3800 & n16155 ) | ( n3800 & n16187 ) | ( n16155 & n16187 ) ;
  assign n17794 = n3802 | n16081 ;
  assign n17795 = n3799 & ~n16079 ;
  assign n17796 = ( ~n16081 & n17794 ) | ( ~n16081 & n17795 ) | ( n17794 & n17795 ) ;
  assign n17797 = ( ~n17792 & n17793 ) | ( ~n17792 & n17796 ) | ( n17793 & n17796 ) ;
  assign n17798 = ( n17793 & n17796 ) | ( n17793 & ~n17797 ) | ( n17796 & ~n17797 ) ;
  assign n17799 = ( n17792 & n17797 ) | ( n17792 & ~n17798 ) | ( n17797 & ~n17798 ) ;
  assign n17800 = n4202 & ~n16176 ;
  assign n17801 = n4201 & ~n16073 ;
  assign n17802 = n4200 & n16077 ;
  assign n17803 = n4345 & ~n16075 ;
  assign n17804 = n17802 | n17803 ;
  assign n17805 = ( ~n17800 & n17801 ) | ( ~n17800 & n17804 ) | ( n17801 & n17804 ) ;
  assign n17806 = ( ~x26 & n17800 ) | ( ~x26 & n17805 ) | ( n17800 & n17805 ) ;
  assign n17807 = ( n17800 & n17805 ) | ( n17800 & ~n17806 ) | ( n17805 & ~n17806 ) ;
  assign n17808 = ( x26 & n17806 ) | ( x26 & ~n17807 ) | ( n17806 & ~n17807 ) ;
  assign n17809 = ( n17693 & n17799 ) | ( n17693 & n17808 ) | ( n17799 & n17808 ) ;
  assign n17810 = ( n17693 & ~n17799 ) | ( n17693 & n17808 ) | ( ~n17799 & n17808 ) ;
  assign n17811 = ( n17799 & ~n17809 ) | ( n17799 & n17810 ) | ( ~n17809 & n17810 ) ;
  assign n17812 = ( n17696 & n17791 ) | ( n17696 & n17811 ) | ( n17791 & n17811 ) ;
  assign n17813 = ( n17696 & ~n17791 ) | ( n17696 & n17811 ) | ( ~n17791 & n17811 ) ;
  assign n17814 = ( n17791 & ~n17812 ) | ( n17791 & n17813 ) | ( ~n17812 & n17813 ) ;
  assign n17815 = n4974 & ~n16354 ;
  assign n17816 = n5398 & ~n16061 ;
  assign n17817 = n4973 & n16065 ;
  assign n17818 = n4972 & n16063 ;
  assign n17819 = n17817 | n17818 ;
  assign n17820 = ( ~n17815 & n17816 ) | ( ~n17815 & n17819 ) | ( n17816 & n17819 ) ;
  assign n17821 = ( ~x20 & n17815 ) | ( ~x20 & n17820 ) | ( n17815 & n17820 ) ;
  assign n17822 = ( n17815 & n17820 ) | ( n17815 & ~n17821 ) | ( n17820 & ~n17821 ) ;
  assign n17823 = ( x20 & n17821 ) | ( x20 & ~n17822 ) | ( n17821 & ~n17822 ) ;
  assign n17824 = ( n17708 & n17814 ) | ( n17708 & n17823 ) | ( n17814 & n17823 ) ;
  assign n17825 = ( ~n17708 & n17814 ) | ( ~n17708 & n17823 ) | ( n17814 & n17823 ) ;
  assign n17826 = ( n17708 & ~n17824 ) | ( n17708 & n17825 ) | ( ~n17824 & n17825 ) ;
  assign n17827 = ( n17711 & n17782 ) | ( n17711 & n17826 ) | ( n17782 & n17826 ) ;
  assign n17828 = ( ~n17711 & n17782 ) | ( ~n17711 & n17826 ) | ( n17782 & n17826 ) ;
  assign n17829 = ( n17711 & ~n17827 ) | ( n17711 & n17828 ) | ( ~n17827 & n17828 ) ;
  assign n17830 = n5966 & ~n16674 ;
  assign n17831 = n6464 & ~n16049 ;
  assign n17832 = n5970 & n16053 ;
  assign n17833 = n5969 & ~n16051 ;
  assign n17834 = n17832 | n17833 ;
  assign n17835 = ( ~n17830 & n17831 ) | ( ~n17830 & n17834 ) | ( n17831 & n17834 ) ;
  assign n17836 = ( ~x14 & n17830 ) | ( ~x14 & n17835 ) | ( n17830 & n17835 ) ;
  assign n17837 = ( n17830 & n17835 ) | ( n17830 & ~n17836 ) | ( n17835 & ~n17836 ) ;
  assign n17838 = ( x14 & n17836 ) | ( x14 & ~n17837 ) | ( n17836 & ~n17837 ) ;
  assign n17839 = ( n17723 & n17829 ) | ( n17723 & n17838 ) | ( n17829 & n17838 ) ;
  assign n17840 = ( ~n17723 & n17829 ) | ( ~n17723 & n17838 ) | ( n17829 & n17838 ) ;
  assign n17841 = ( n17723 & ~n17839 ) | ( n17723 & n17840 ) | ( ~n17839 & n17840 ) ;
  assign n17842 = ( n17726 & n17773 ) | ( n17726 & n17841 ) | ( n17773 & n17841 ) ;
  assign n17843 = ( ~n17726 & n17773 ) | ( ~n17726 & n17841 ) | ( n17773 & n17841 ) ;
  assign n17844 = ( n17726 & ~n17842 ) | ( n17726 & n17843 ) | ( ~n17842 & n17843 ) ;
  assign n17845 = n7296 & ~n17138 ;
  assign n17846 = n7879 & ~n16037 ;
  assign n17847 = n7300 & n16041 ;
  assign n17848 = n7299 & n16039 ;
  assign n17849 = n17847 | n17848 ;
  assign n17850 = ( ~n17845 & n17846 ) | ( ~n17845 & n17849 ) | ( n17846 & n17849 ) ;
  assign n17851 = ( ~x8 & n17845 ) | ( ~x8 & n17850 ) | ( n17845 & n17850 ) ;
  assign n17852 = ( n17845 & n17850 ) | ( n17845 & ~n17851 ) | ( n17850 & ~n17851 ) ;
  assign n17853 = ( x8 & n17851 ) | ( x8 & ~n17852 ) | ( n17851 & ~n17852 ) ;
  assign n17854 = ( n17738 & n17844 ) | ( n17738 & n17853 ) | ( n17844 & n17853 ) ;
  assign n17855 = ( ~n17738 & n17844 ) | ( ~n17738 & n17853 ) | ( n17844 & n17853 ) ;
  assign n17856 = ( n17738 & ~n17854 ) | ( n17738 & n17855 ) | ( ~n17854 & n17855 ) ;
  assign n17857 = ( n17741 & n17764 ) | ( n17741 & n17856 ) | ( n17764 & n17856 ) ;
  assign n17858 = ( ~n17741 & n17764 ) | ( ~n17741 & n17856 ) | ( n17764 & n17856 ) ;
  assign n17859 = ( n17741 & ~n17857 ) | ( n17741 & n17858 ) | ( ~n17857 & n17858 ) ;
  assign n17860 = ( n17744 & n17755 ) | ( n17744 & n17859 ) | ( n17755 & n17859 ) ;
  assign n17861 = n7296 & ~n17313 ;
  assign n17862 = n7879 & n16035 ;
  assign n17863 = n7300 & n16039 ;
  assign n17864 = n7299 & ~n16037 ;
  assign n17865 = n17863 | n17864 ;
  assign n17866 = ( ~n17861 & n17862 ) | ( ~n17861 & n17865 ) | ( n17862 & n17865 ) ;
  assign n17867 = ( ~x8 & n17861 ) | ( ~x8 & n17866 ) | ( n17861 & n17866 ) ;
  assign n17868 = ( n17861 & n17866 ) | ( n17861 & ~n17867 ) | ( n17866 & ~n17867 ) ;
  assign n17869 = ( x8 & n17867 ) | ( x8 & ~n17868 ) | ( n17867 & ~n17868 ) ;
  assign n17870 = n5966 & ~n16801 ;
  assign n17871 = n6464 & ~n16047 ;
  assign n17872 = n5970 & ~n16051 ;
  assign n17873 = n5969 & ~n16049 ;
  assign n17874 = n17872 | n17873 ;
  assign n17875 = ( ~n17870 & n17871 ) | ( ~n17870 & n17874 ) | ( n17871 & n17874 ) ;
  assign n17876 = ( ~x14 & n17870 ) | ( ~x14 & n17875 ) | ( n17870 & n17875 ) ;
  assign n17877 = ( n17870 & n17875 ) | ( n17870 & ~n17876 ) | ( n17875 & ~n17876 ) ;
  assign n17878 = ( x14 & n17876 ) | ( x14 & ~n17877 ) | ( n17876 & ~n17877 ) ;
  assign n17879 = n4974 & ~n16433 ;
  assign n17880 = n5398 & n16059 ;
  assign n17881 = n4973 & n16063 ;
  assign n17882 = n4972 & ~n16061 ;
  assign n17883 = n17881 | n17882 ;
  assign n17884 = ( ~n17879 & n17880 ) | ( ~n17879 & n17883 ) | ( n17880 & n17883 ) ;
  assign n17885 = ( ~x20 & n17879 ) | ( ~x20 & n17884 ) | ( n17879 & n17884 ) ;
  assign n17886 = ( n17879 & n17884 ) | ( n17879 & ~n17885 ) | ( n17884 & ~n17885 ) ;
  assign n17887 = ( x20 & n17885 ) | ( x20 & ~n17886 ) | ( n17885 & ~n17886 ) ;
  assign n17888 = n4202 & n16209 ;
  assign n17889 = n4201 & n16071 ;
  assign n17890 = n4200 & ~n16075 ;
  assign n17891 = n4345 & ~n16073 ;
  assign n17892 = n17890 | n17891 ;
  assign n17893 = ( ~n17888 & n17889 ) | ( ~n17888 & n17892 ) | ( n17889 & n17892 ) ;
  assign n17894 = ( ~x26 & n17888 ) | ( ~x26 & n17893 ) | ( n17888 & n17893 ) ;
  assign n17895 = ( n17888 & n17893 ) | ( n17888 & ~n17894 ) | ( n17893 & ~n17894 ) ;
  assign n17896 = ( x26 & n17894 ) | ( x26 & ~n17895 ) | ( n17894 & ~n17895 ) ;
  assign n17897 = ( x29 & n17792 ) | ( x29 & n17797 ) | ( n17792 & n17797 ) ;
  assign n17898 = ( n3800 & n16083 ) | ( n3800 & n16198 ) | ( n16083 & n16198 ) ;
  assign n17899 = n3700 & ~n16081 ;
  assign n17900 = n3802 & ~n16079 ;
  assign n17901 = n17899 | n17900 ;
  assign n17902 = n3799 & ~n16077 ;
  assign n17903 = ( n3799 & n17901 ) | ( n3799 & ~n17902 ) | ( n17901 & ~n17902 ) ;
  assign n17904 = ( ~n17897 & n17898 ) | ( ~n17897 & n17903 ) | ( n17898 & n17903 ) ;
  assign n17905 = ( n17898 & n17903 ) | ( n17898 & ~n17904 ) | ( n17903 & ~n17904 ) ;
  assign n17906 = ( n17897 & n17904 ) | ( n17897 & ~n17905 ) | ( n17904 & ~n17905 ) ;
  assign n17907 = ( n17809 & n17896 ) | ( n17809 & n17906 ) | ( n17896 & n17906 ) ;
  assign n17908 = ( n17809 & ~n17896 ) | ( n17809 & n17906 ) | ( ~n17896 & n17906 ) ;
  assign n17909 = ( n17896 & ~n17907 ) | ( n17896 & n17908 ) | ( ~n17907 & n17908 ) ;
  assign n17910 = n4713 & n16281 ;
  assign n17911 = n4712 & n16065 ;
  assign n17912 = n4709 & n16069 ;
  assign n17913 = n4792 & n16067 ;
  assign n17914 = n17912 | n17913 ;
  assign n17915 = ( ~n17910 & n17911 ) | ( ~n17910 & n17914 ) | ( n17911 & n17914 ) ;
  assign n17916 = ( ~x23 & n17910 ) | ( ~x23 & n17915 ) | ( n17910 & n17915 ) ;
  assign n17917 = ( n17910 & n17915 ) | ( n17910 & ~n17916 ) | ( n17915 & ~n17916 ) ;
  assign n17918 = ( x23 & n17916 ) | ( x23 & ~n17917 ) | ( n17916 & ~n17917 ) ;
  assign n17919 = ( n17812 & n17909 ) | ( n17812 & n17918 ) | ( n17909 & n17918 ) ;
  assign n17920 = ( n17812 & ~n17909 ) | ( n17812 & n17918 ) | ( ~n17909 & n17918 ) ;
  assign n17921 = ( n17909 & ~n17919 ) | ( n17909 & n17920 ) | ( ~n17919 & n17920 ) ;
  assign n17922 = ( n17824 & n17887 ) | ( n17824 & n17921 ) | ( n17887 & n17921 ) ;
  assign n17923 = ( n17824 & ~n17887 ) | ( n17824 & n17921 ) | ( ~n17887 & n17921 ) ;
  assign n17924 = ( n17887 & ~n17922 ) | ( n17887 & n17923 ) | ( ~n17922 & n17923 ) ;
  assign n17925 = n5508 & n16553 ;
  assign n17926 = n5507 & n16053 ;
  assign n17927 = n5504 & ~n16057 ;
  assign n17928 = n5666 & ~n16055 ;
  assign n17929 = n17927 | n17928 ;
  assign n17930 = ( ~n17925 & n17926 ) | ( ~n17925 & n17929 ) | ( n17926 & n17929 ) ;
  assign n17931 = ( ~x17 & n17925 ) | ( ~x17 & n17930 ) | ( n17925 & n17930 ) ;
  assign n17932 = ( n17925 & n17930 ) | ( n17925 & ~n17931 ) | ( n17930 & ~n17931 ) ;
  assign n17933 = ( x17 & n17931 ) | ( x17 & ~n17932 ) | ( n17931 & ~n17932 ) ;
  assign n17934 = ( n17827 & n17924 ) | ( n17827 & n17933 ) | ( n17924 & n17933 ) ;
  assign n17935 = ( ~n17827 & n17924 ) | ( ~n17827 & n17933 ) | ( n17924 & n17933 ) ;
  assign n17936 = ( n17827 & ~n17934 ) | ( n17827 & n17935 ) | ( ~n17934 & n17935 ) ;
  assign n17937 = ( n17839 & n17878 ) | ( n17839 & n17936 ) | ( n17878 & n17936 ) ;
  assign n17938 = ( ~n17839 & n17878 ) | ( ~n17839 & n17936 ) | ( n17878 & n17936 ) ;
  assign n17939 = ( n17839 & ~n17937 ) | ( n17839 & n17938 ) | ( ~n17937 & n17938 ) ;
  assign n17940 = n6584 & n16969 ;
  assign n17941 = n7022 & n16041 ;
  assign n17942 = n6588 & ~n16045 ;
  assign n17943 = n6587 & ~n16043 ;
  assign n17944 = n17942 | n17943 ;
  assign n17945 = ( ~n17940 & n17941 ) | ( ~n17940 & n17944 ) | ( n17941 & n17944 ) ;
  assign n17946 = ( ~x11 & n17940 ) | ( ~x11 & n17945 ) | ( n17940 & n17945 ) ;
  assign n17947 = ( n17940 & n17945 ) | ( n17940 & ~n17946 ) | ( n17945 & ~n17946 ) ;
  assign n17948 = ( x11 & n17946 ) | ( x11 & ~n17947 ) | ( n17946 & ~n17947 ) ;
  assign n17949 = ( n17842 & n17939 ) | ( n17842 & n17948 ) | ( n17939 & n17948 ) ;
  assign n17950 = ( ~n17842 & n17939 ) | ( ~n17842 & n17948 ) | ( n17939 & n17948 ) ;
  assign n17951 = ( n17842 & ~n17949 ) | ( n17842 & n17950 ) | ( ~n17949 & n17950 ) ;
  assign n17952 = ( n17854 & n17869 ) | ( n17854 & n17951 ) | ( n17869 & n17951 ) ;
  assign n17953 = ( ~n17854 & n17869 ) | ( ~n17854 & n17951 ) | ( n17869 & n17951 ) ;
  assign n17954 = ( n17854 & ~n17952 ) | ( n17854 & n17953 ) | ( ~n17952 & n17953 ) ;
  assign n17955 = n8230 & ~n17528 ;
  assign n17956 = n8229 & ~n16029 ;
  assign n17957 = n8226 & ~n16033 ;
  assign n17958 = n8225 & n16031 ;
  assign n17959 = n17957 | n17958 ;
  assign n17960 = ( ~n17955 & n17956 ) | ( ~n17955 & n17959 ) | ( n17956 & n17959 ) ;
  assign n17961 = ( ~x5 & n17955 ) | ( ~x5 & n17960 ) | ( n17955 & n17960 ) ;
  assign n17962 = ( n17955 & n17960 ) | ( n17955 & ~n17961 ) | ( n17960 & ~n17961 ) ;
  assign n17963 = ( x5 & n17961 ) | ( x5 & ~n17962 ) | ( n17961 & ~n17962 ) ;
  assign n17964 = ( n17857 & n17954 ) | ( n17857 & n17963 ) | ( n17954 & n17963 ) ;
  assign n17965 = ( ~n17857 & n17954 ) | ( ~n17857 & n17963 ) | ( n17954 & n17963 ) ;
  assign n17966 = ( n17857 & ~n17964 ) | ( n17857 & n17965 ) | ( ~n17964 & n17965 ) ;
  assign n17967 = ( n16023 & n16025 ) | ( n16023 & ~n16110 ) | ( n16025 & ~n16110 ) ;
  assign n17968 = ( ~n16025 & n16111 ) | ( ~n16025 & n17967 ) | ( n16111 & n17967 ) ;
  assign n17969 = n36 & n17968 ;
  assign n17970 = n8967 & ~n16027 ;
  assign n17971 = ( x0 & n8966 ) | ( x0 & n16025 ) | ( n8966 & n16025 ) ;
  assign n17972 = ( n8966 & n17970 ) | ( n8966 & ~n17971 ) | ( n17970 & ~n17971 ) ;
  assign n17973 = n35 & ~n16023 ;
  assign n17974 = ( n35 & n17972 ) | ( n35 & ~n17973 ) | ( n17972 & ~n17973 ) ;
  assign n17975 = ( ~x2 & n17969 ) | ( ~x2 & n17974 ) | ( n17969 & n17974 ) ;
  assign n17976 = ( n17969 & n17974 ) | ( n17969 & ~n17975 ) | ( n17974 & ~n17975 ) ;
  assign n17977 = ( x2 & n17975 ) | ( x2 & ~n17976 ) | ( n17975 & ~n17976 ) ;
  assign n17978 = ( n17860 & n17966 ) | ( n17860 & n17977 ) | ( n17966 & n17977 ) ;
  assign n17979 = n7296 & ~n17412 ;
  assign n17980 = n7879 & ~n16033 ;
  assign n17981 = n7300 & ~n16037 ;
  assign n17982 = n7299 & n16035 ;
  assign n17983 = n17981 | n17982 ;
  assign n17984 = ( ~n17979 & n17980 ) | ( ~n17979 & n17983 ) | ( n17980 & n17983 ) ;
  assign n17985 = ( ~x8 & n17979 ) | ( ~x8 & n17984 ) | ( n17979 & n17984 ) ;
  assign n17986 = ( n17979 & n17984 ) | ( n17979 & ~n17985 ) | ( n17984 & ~n17985 ) ;
  assign n17987 = ( x8 & n17985 ) | ( x8 & ~n17986 ) | ( n17985 & ~n17986 ) ;
  assign n17988 = n5966 & ~n16876 ;
  assign n17989 = n6464 & ~n16045 ;
  assign n17990 = n5970 & ~n16049 ;
  assign n17991 = n5969 & ~n16047 ;
  assign n17992 = n17990 | n17991 ;
  assign n17993 = ( ~n17988 & n17989 ) | ( ~n17988 & n17992 ) | ( n17989 & n17992 ) ;
  assign n17994 = ( ~x14 & n17988 ) | ( ~x14 & n17993 ) | ( n17988 & n17993 ) ;
  assign n17995 = ( n17988 & n17993 ) | ( n17988 & ~n17994 ) | ( n17993 & ~n17994 ) ;
  assign n17996 = ( x14 & n17994 ) | ( x14 & ~n17995 ) | ( n17994 & ~n17995 ) ;
  assign n17997 = n4974 & ~n16484 ;
  assign n17998 = n5398 & ~n16057 ;
  assign n17999 = n4973 & ~n16061 ;
  assign n18000 = n4972 & n16059 ;
  assign n18001 = n17999 | n18000 ;
  assign n18002 = ( ~n17997 & n17998 ) | ( ~n17997 & n18001 ) | ( n17998 & n18001 ) ;
  assign n18003 = ( ~x20 & n17997 ) | ( ~x20 & n18002 ) | ( n17997 & n18002 ) ;
  assign n18004 = ( n17997 & n18002 ) | ( n17997 & ~n18003 ) | ( n18002 & ~n18003 ) ;
  assign n18005 = ( x20 & n18003 ) | ( x20 & ~n18004 ) | ( n18003 & ~n18004 ) ;
  assign n18006 = n4202 & ~n16221 ;
  assign n18007 = n4201 & n16069 ;
  assign n18008 = n4200 & ~n16073 ;
  assign n18009 = n4345 & n16071 ;
  assign n18010 = n18008 | n18009 ;
  assign n18011 = ( ~n18006 & n18007 ) | ( ~n18006 & n18010 ) | ( n18007 & n18010 ) ;
  assign n18012 = ( ~x26 & n18006 ) | ( ~x26 & n18011 ) | ( n18006 & n18011 ) ;
  assign n18013 = ( n18006 & n18011 ) | ( n18006 & ~n18012 ) | ( n18011 & ~n18012 ) ;
  assign n18014 = ( x26 & n18012 ) | ( x26 & ~n18013 ) | ( n18012 & ~n18013 ) ;
  assign n18015 = ( n58 & n96 ) | ( n58 & ~n16081 ) | ( n96 & ~n16081 ) ;
  assign n18016 = n3800 & n16169 ;
  assign n18017 = n3799 & ~n16075 ;
  assign n18018 = n3700 & ~n16079 ;
  assign n18019 = n3802 & n16077 ;
  assign n18020 = n18018 | n18019 ;
  assign n18021 = ( ~n18016 & n18017 ) | ( ~n18016 & n18020 ) | ( n18017 & n18020 ) ;
  assign n18022 = ( ~x29 & n18016 ) | ( ~x29 & n18021 ) | ( n18016 & n18021 ) ;
  assign n18023 = ( n18016 & n18021 ) | ( n18016 & ~n18022 ) | ( n18021 & ~n18022 ) ;
  assign n18024 = ( x29 & n18022 ) | ( x29 & ~n18023 ) | ( n18022 & ~n18023 ) ;
  assign n18025 = x29 & ~n17897 ;
  assign n18026 = ~n17904 & n18025 ;
  assign n18027 = ( n18015 & n18024 ) | ( n18015 & n18026 ) | ( n18024 & n18026 ) ;
  assign n18028 = ( ~n18015 & n18024 ) | ( ~n18015 & n18026 ) | ( n18024 & n18026 ) ;
  assign n18029 = ( n18015 & ~n18027 ) | ( n18015 & n18028 ) | ( ~n18027 & n18028 ) ;
  assign n18030 = ( n17907 & n18014 ) | ( n17907 & n18029 ) | ( n18014 & n18029 ) ;
  assign n18031 = ( n17907 & ~n18014 ) | ( n17907 & n18029 ) | ( ~n18014 & n18029 ) ;
  assign n18032 = ( n18014 & ~n18030 ) | ( n18014 & n18031 ) | ( ~n18030 & n18031 ) ;
  assign n18033 = n4713 & n16315 ;
  assign n18034 = n4712 & n16063 ;
  assign n18035 = n4709 & n16067 ;
  assign n18036 = n4792 & n16065 ;
  assign n18037 = n18035 | n18036 ;
  assign n18038 = ( ~n18033 & n18034 ) | ( ~n18033 & n18037 ) | ( n18034 & n18037 ) ;
  assign n18039 = ( ~x23 & n18033 ) | ( ~x23 & n18038 ) | ( n18033 & n18038 ) ;
  assign n18040 = ( n18033 & n18038 ) | ( n18033 & ~n18039 ) | ( n18038 & ~n18039 ) ;
  assign n18041 = ( x23 & n18039 ) | ( x23 & ~n18040 ) | ( n18039 & ~n18040 ) ;
  assign n18042 = ( n17919 & n18032 ) | ( n17919 & n18041 ) | ( n18032 & n18041 ) ;
  assign n18043 = ( n17919 & ~n18032 ) | ( n17919 & n18041 ) | ( ~n18032 & n18041 ) ;
  assign n18044 = ( n18032 & ~n18042 ) | ( n18032 & n18043 ) | ( ~n18042 & n18043 ) ;
  assign n18045 = ( n17922 & n18005 ) | ( n17922 & n18044 ) | ( n18005 & n18044 ) ;
  assign n18046 = ( n17922 & ~n18005 ) | ( n17922 & n18044 ) | ( ~n18005 & n18044 ) ;
  assign n18047 = ( n18005 & ~n18045 ) | ( n18005 & n18046 ) | ( ~n18045 & n18046 ) ;
  assign n18048 = n5508 & n16611 ;
  assign n18049 = n5507 & ~n16051 ;
  assign n18050 = n5504 & ~n16055 ;
  assign n18051 = n5666 & n16053 ;
  assign n18052 = n18050 | n18051 ;
  assign n18053 = ( ~n18048 & n18049 ) | ( ~n18048 & n18052 ) | ( n18049 & n18052 ) ;
  assign n18054 = ( ~x17 & n18048 ) | ( ~x17 & n18053 ) | ( n18048 & n18053 ) ;
  assign n18055 = ( n18048 & n18053 ) | ( n18048 & ~n18054 ) | ( n18053 & ~n18054 ) ;
  assign n18056 = ( x17 & n18054 ) | ( x17 & ~n18055 ) | ( n18054 & ~n18055 ) ;
  assign n18057 = ( n17934 & n18047 ) | ( n17934 & n18056 ) | ( n18047 & n18056 ) ;
  assign n18058 = ( n17934 & ~n18047 ) | ( n17934 & n18056 ) | ( ~n18047 & n18056 ) ;
  assign n18059 = ( n18047 & ~n18057 ) | ( n18047 & n18058 ) | ( ~n18057 & n18058 ) ;
  assign n18060 = ( n17937 & n17996 ) | ( n17937 & n18059 ) | ( n17996 & n18059 ) ;
  assign n18061 = ( ~n17937 & n17996 ) | ( ~n17937 & n18059 ) | ( n17996 & n18059 ) ;
  assign n18062 = ( n17937 & ~n18060 ) | ( n17937 & n18061 ) | ( ~n18060 & n18061 ) ;
  assign n18063 = n6584 & ~n17051 ;
  assign n18064 = n7022 & n16039 ;
  assign n18065 = n6588 & ~n16043 ;
  assign n18066 = n6587 & n16041 ;
  assign n18067 = n18065 | n18066 ;
  assign n18068 = ( ~n18063 & n18064 ) | ( ~n18063 & n18067 ) | ( n18064 & n18067 ) ;
  assign n18069 = ( ~x11 & n18063 ) | ( ~x11 & n18068 ) | ( n18063 & n18068 ) ;
  assign n18070 = ( n18063 & n18068 ) | ( n18063 & ~n18069 ) | ( n18068 & ~n18069 ) ;
  assign n18071 = ( x11 & n18069 ) | ( x11 & ~n18070 ) | ( n18069 & ~n18070 ) ;
  assign n18072 = ( n17949 & n18062 ) | ( n17949 & n18071 ) | ( n18062 & n18071 ) ;
  assign n18073 = ( ~n17949 & n18062 ) | ( ~n17949 & n18071 ) | ( n18062 & n18071 ) ;
  assign n18074 = ( n17949 & ~n18072 ) | ( n17949 & n18073 ) | ( ~n18072 & n18073 ) ;
  assign n18075 = ( n17952 & n17987 ) | ( n17952 & n18074 ) | ( n17987 & n18074 ) ;
  assign n18076 = ( ~n17952 & n17987 ) | ( ~n17952 & n18074 ) | ( n17987 & n18074 ) ;
  assign n18077 = ( n17952 & ~n18075 ) | ( n17952 & n18076 ) | ( ~n18075 & n18076 ) ;
  assign n18078 = n8230 & n17634 ;
  assign n18079 = n8229 & ~n16027 ;
  assign n18080 = n8226 & n16031 ;
  assign n18081 = n8225 & ~n16029 ;
  assign n18082 = n18080 | n18081 ;
  assign n18083 = ( ~n18078 & n18079 ) | ( ~n18078 & n18082 ) | ( n18079 & n18082 ) ;
  assign n18084 = ( ~x5 & n18078 ) | ( ~x5 & n18083 ) | ( n18078 & n18083 ) ;
  assign n18085 = ( n18078 & n18083 ) | ( n18078 & ~n18084 ) | ( n18083 & ~n18084 ) ;
  assign n18086 = ( x5 & n18084 ) | ( x5 & ~n18085 ) | ( n18084 & ~n18085 ) ;
  assign n18087 = ( n17964 & n18077 ) | ( n17964 & n18086 ) | ( n18077 & n18086 ) ;
  assign n18088 = ( ~n17964 & n18077 ) | ( ~n17964 & n18086 ) | ( n18077 & n18086 ) ;
  assign n18089 = ( n17964 & ~n18087 ) | ( n17964 & n18088 ) | ( ~n18087 & n18088 ) ;
  assign n18090 = ( n16021 & n16023 ) | ( n16021 & ~n16112 ) | ( n16023 & ~n16112 ) ;
  assign n18091 = ( n16111 & n16112 ) | ( n16111 & ~n18090 ) | ( n16112 & ~n18090 ) ;
  assign n18092 = n36 & ~n18091 ;
  assign n18093 = n8967 & ~n16025 ;
  assign n18094 = ( x0 & n8966 ) | ( x0 & ~n16023 ) | ( n8966 & ~n16023 ) ;
  assign n18095 = ( n8966 & n18093 ) | ( n8966 & ~n18094 ) | ( n18093 & ~n18094 ) ;
  assign n18096 = n35 & ~n16021 ;
  assign n18097 = ( n35 & n18095 ) | ( n35 & ~n18096 ) | ( n18095 & ~n18096 ) ;
  assign n18098 = ( ~x2 & n18092 ) | ( ~x2 & n18097 ) | ( n18092 & n18097 ) ;
  assign n18099 = ( n18092 & n18097 ) | ( n18092 & ~n18098 ) | ( n18097 & ~n18098 ) ;
  assign n18100 = ( x2 & n18098 ) | ( x2 & ~n18099 ) | ( n18098 & ~n18099 ) ;
  assign n18101 = ( n17978 & n18089 ) | ( n17978 & n18100 ) | ( n18089 & n18100 ) ;
  assign n18102 = ( n16019 & n16021 ) | ( n16019 & ~n16112 ) | ( n16021 & ~n16112 ) ;
  assign n18103 = ( n16112 & ~n16113 ) | ( n16112 & n18102 ) | ( ~n16113 & n18102 ) ;
  assign n18104 = n36 & n18103 ;
  assign n18105 = n8967 & n16023 ;
  assign n18106 = ( x0 & n8966 ) | ( x0 & ~n16021 ) | ( n8966 & ~n16021 ) ;
  assign n18107 = ( n8966 & n18105 ) | ( n8966 & ~n18106 ) | ( n18105 & ~n18106 ) ;
  assign n18108 = n35 & ~n16019 ;
  assign n18109 = ( n35 & n18107 ) | ( n35 & ~n18108 ) | ( n18107 & ~n18108 ) ;
  assign n18110 = ( ~x2 & n18104 ) | ( ~x2 & n18109 ) | ( n18104 & n18109 ) ;
  assign n18111 = ( n18104 & n18109 ) | ( n18104 & ~n18110 ) | ( n18109 & ~n18110 ) ;
  assign n18112 = ( x2 & n18110 ) | ( x2 & ~n18111 ) | ( n18110 & ~n18111 ) ;
  assign n18113 = n8230 & ~n17746 ;
  assign n18114 = n8229 & ~n16025 ;
  assign n18115 = n8226 & ~n16029 ;
  assign n18116 = n8225 & ~n16027 ;
  assign n18117 = n18115 | n18116 ;
  assign n18118 = ( ~n18113 & n18114 ) | ( ~n18113 & n18117 ) | ( n18114 & n18117 ) ;
  assign n18119 = ( ~x5 & n18113 ) | ( ~x5 & n18118 ) | ( n18113 & n18118 ) ;
  assign n18120 = ( n18113 & n18118 ) | ( n18113 & ~n18119 ) | ( n18118 & ~n18119 ) ;
  assign n18121 = ( x5 & n18119 ) | ( x5 & ~n18120 ) | ( n18119 & ~n18120 ) ;
  assign n18122 = n7296 & ~n17516 ;
  assign n18123 = n7879 & n16031 ;
  assign n18124 = n7300 & n16035 ;
  assign n18125 = n7299 & ~n16033 ;
  assign n18126 = n18124 | n18125 ;
  assign n18127 = ( ~n18122 & n18123 ) | ( ~n18122 & n18126 ) | ( n18123 & n18126 ) ;
  assign n18128 = ( ~x8 & n18122 ) | ( ~x8 & n18127 ) | ( n18122 & n18127 ) ;
  assign n18129 = ( n18122 & n18127 ) | ( n18122 & ~n18128 ) | ( n18127 & ~n18128 ) ;
  assign n18130 = ( x8 & n18128 ) | ( x8 & ~n18129 ) | ( n18128 & ~n18129 ) ;
  assign n18131 = n6584 & ~n17138 ;
  assign n18132 = n7022 & ~n16037 ;
  assign n18133 = n6588 & n16041 ;
  assign n18134 = n6587 & n16039 ;
  assign n18135 = n18133 | n18134 ;
  assign n18136 = ( ~n18131 & n18132 ) | ( ~n18131 & n18135 ) | ( n18132 & n18135 ) ;
  assign n18137 = ( ~x11 & n18131 ) | ( ~x11 & n18136 ) | ( n18131 & n18136 ) ;
  assign n18138 = ( n18131 & n18136 ) | ( n18131 & ~n18137 ) | ( n18136 & ~n18137 ) ;
  assign n18139 = ( x11 & n18137 ) | ( x11 & ~n18138 ) | ( n18137 & ~n18138 ) ;
  assign n18140 = n146 | n2434 ;
  assign n18141 = ( n72 & n109 ) | ( n72 & n116 ) | ( n109 & n116 ) ;
  assign n18142 = ( n3042 & ~n18140 ) | ( n3042 & n18141 ) | ( ~n18140 & n18141 ) ;
  assign n18143 = n18140 | n18142 ;
  assign n18144 = n5996 | n11901 ;
  assign n18145 = ( n838 & ~n947 ) | ( n838 & n1494 ) | ( ~n947 & n1494 ) ;
  assign n18146 = n947 | n18145 ;
  assign n18147 = n712 | n1720 ;
  assign n18148 = ( n2161 & ~n18146 ) | ( n2161 & n18147 ) | ( ~n18146 & n18147 ) ;
  assign n18149 = n18146 | n18148 ;
  assign n18150 = ( ~n18143 & n18144 ) | ( ~n18143 & n18149 ) | ( n18144 & n18149 ) ;
  assign n18151 = n18143 | n18150 ;
  assign n18152 = n340 | n386 ;
  assign n18153 = n1024 | n1589 ;
  assign n18154 = n256 | n978 ;
  assign n18155 = ( n3568 & ~n3879 ) | ( n3568 & n18154 ) | ( ~n3879 & n18154 ) ;
  assign n18156 = ~n18154 & n18155 ;
  assign n18157 = ( n18152 & ~n18153 ) | ( n18152 & n18156 ) | ( ~n18153 & n18156 ) ;
  assign n18158 = ~n18152 & n18157 ;
  assign n18159 = ( n41 & n44 ) | ( n41 & n80 ) | ( n44 & n80 ) ;
  assign n18160 = ( n211 & n544 ) | ( n211 & ~n18159 ) | ( n544 & ~n18159 ) ;
  assign n18161 = n18159 | n18160 ;
  assign n18162 = n404 | n4391 ;
  assign n18163 = n18161 | n18162 ;
  assign n18164 = ( n10816 & n18158 ) | ( n10816 & n18163 ) | ( n18158 & n18163 ) ;
  assign n18165 = n18158 & ~n18164 ;
  assign n18166 = ~n11990 & n18165 ;
  assign n18167 = n1145 | n1737 ;
  assign n18168 = n76 | n123 ;
  assign n18169 = n253 | n1533 ;
  assign n18170 = ( n1523 & n1653 ) | ( n1523 & ~n18169 ) | ( n1653 & ~n18169 ) ;
  assign n18171 = n18169 | n18170 ;
  assign n18172 = ( n545 & ~n18168 ) | ( n545 & n18171 ) | ( ~n18168 & n18171 ) ;
  assign n18173 = n18168 | n18172 ;
  assign n18174 = ( n4849 & ~n18167 ) | ( n4849 & n18173 ) | ( ~n18167 & n18173 ) ;
  assign n18175 = n18167 | n18174 ;
  assign n18176 = ( n18151 & n18166 ) | ( n18151 & ~n18175 ) | ( n18166 & ~n18175 ) ;
  assign n18177 = ~n18151 & n18176 ;
  assign n18178 = ( n1248 & n16155 ) | ( n1248 & n16187 ) | ( n16155 & n16187 ) ;
  assign n18179 = ( n606 & ~n16079 ) | ( n606 & n18178 ) | ( ~n16079 & n18178 ) ;
  assign n18180 = ( n1250 & ~n16081 ) | ( n1250 & n18178 ) | ( ~n16081 & n18178 ) ;
  assign n18181 = n18179 | n18180 ;
  assign n18182 = ~n18177 & n18181 ;
  assign n18183 = n18177 & n18181 ;
  assign n18184 = ( n18177 & n18182 ) | ( n18177 & ~n18183 ) | ( n18182 & ~n18183 ) ;
  assign n18185 = n3800 & ~n16176 ;
  assign n18186 = n3799 & ~n16073 ;
  assign n18187 = n3700 & n16077 ;
  assign n18188 = n3802 & ~n16075 ;
  assign n18189 = n18187 | n18188 ;
  assign n18190 = ( ~n18185 & n18186 ) | ( ~n18185 & n18189 ) | ( n18186 & n18189 ) ;
  assign n18191 = ( ~x29 & n18185 ) | ( ~x29 & n18190 ) | ( n18185 & n18190 ) ;
  assign n18192 = ( n18185 & n18190 ) | ( n18185 & ~n18191 ) | ( n18190 & ~n18191 ) ;
  assign n18193 = ( x29 & n18191 ) | ( x29 & ~n18192 ) | ( n18191 & ~n18192 ) ;
  assign n18194 = ( n18027 & ~n18184 ) | ( n18027 & n18193 ) | ( ~n18184 & n18193 ) ;
  assign n18195 = ( n18027 & n18184 ) | ( n18027 & n18193 ) | ( n18184 & n18193 ) ;
  assign n18196 = ( n18184 & n18194 ) | ( n18184 & ~n18195 ) | ( n18194 & ~n18195 ) ;
  assign n18197 = n4202 & n16269 ;
  assign n18198 = n4201 & n16067 ;
  assign n18199 = n4200 & n16071 ;
  assign n18200 = n4345 & n16069 ;
  assign n18201 = n18199 | n18200 ;
  assign n18202 = ( ~n18197 & n18198 ) | ( ~n18197 & n18201 ) | ( n18198 & n18201 ) ;
  assign n18203 = ( ~x26 & n18197 ) | ( ~x26 & n18202 ) | ( n18197 & n18202 ) ;
  assign n18204 = ( n18197 & n18202 ) | ( n18197 & ~n18203 ) | ( n18202 & ~n18203 ) ;
  assign n18205 = ( x26 & n18203 ) | ( x26 & ~n18204 ) | ( n18203 & ~n18204 ) ;
  assign n18206 = ( n18030 & ~n18196 ) | ( n18030 & n18205 ) | ( ~n18196 & n18205 ) ;
  assign n18207 = ( n18030 & n18196 ) | ( n18030 & n18205 ) | ( n18196 & n18205 ) ;
  assign n18208 = ( n18196 & n18206 ) | ( n18196 & ~n18207 ) | ( n18206 & ~n18207 ) ;
  assign n18209 = n4713 & ~n16354 ;
  assign n18210 = n4712 & ~n16061 ;
  assign n18211 = n4709 & n16065 ;
  assign n18212 = n4792 & n16063 ;
  assign n18213 = n18211 | n18212 ;
  assign n18214 = ( ~n18209 & n18210 ) | ( ~n18209 & n18213 ) | ( n18210 & n18213 ) ;
  assign n18215 = ( ~x23 & n18209 ) | ( ~x23 & n18214 ) | ( n18209 & n18214 ) ;
  assign n18216 = ( n18209 & n18214 ) | ( n18209 & ~n18215 ) | ( n18214 & ~n18215 ) ;
  assign n18217 = ( x23 & n18215 ) | ( x23 & ~n18216 ) | ( n18215 & ~n18216 ) ;
  assign n18218 = ( n18042 & ~n18208 ) | ( n18042 & n18217 ) | ( ~n18208 & n18217 ) ;
  assign n18219 = ( n18042 & n18208 ) | ( n18042 & n18217 ) | ( n18208 & n18217 ) ;
  assign n18220 = ( n18208 & n18218 ) | ( n18208 & ~n18219 ) | ( n18218 & ~n18219 ) ;
  assign n18221 = n4974 & n16541 ;
  assign n18222 = n5398 & ~n16055 ;
  assign n18223 = n4973 & n16059 ;
  assign n18224 = n4972 & ~n16057 ;
  assign n18225 = n18223 | n18224 ;
  assign n18226 = ( ~n18221 & n18222 ) | ( ~n18221 & n18225 ) | ( n18222 & n18225 ) ;
  assign n18227 = ( ~x20 & n18221 ) | ( ~x20 & n18226 ) | ( n18221 & n18226 ) ;
  assign n18228 = ( n18221 & n18226 ) | ( n18221 & ~n18227 ) | ( n18226 & ~n18227 ) ;
  assign n18229 = ( x20 & n18227 ) | ( x20 & ~n18228 ) | ( n18227 & ~n18228 ) ;
  assign n18230 = ( n18045 & ~n18220 ) | ( n18045 & n18229 ) | ( ~n18220 & n18229 ) ;
  assign n18231 = ( n18045 & n18220 ) | ( n18045 & n18229 ) | ( n18220 & n18229 ) ;
  assign n18232 = ( n18220 & n18230 ) | ( n18220 & ~n18231 ) | ( n18230 & ~n18231 ) ;
  assign n18233 = n5508 & ~n16674 ;
  assign n18234 = n5507 & ~n16049 ;
  assign n18235 = n5504 & n16053 ;
  assign n18236 = n5666 & ~n16051 ;
  assign n18237 = n18235 | n18236 ;
  assign n18238 = ( ~n18233 & n18234 ) | ( ~n18233 & n18237 ) | ( n18234 & n18237 ) ;
  assign n18239 = ( ~x17 & n18233 ) | ( ~x17 & n18238 ) | ( n18233 & n18238 ) ;
  assign n18240 = ( n18233 & n18238 ) | ( n18233 & ~n18239 ) | ( n18238 & ~n18239 ) ;
  assign n18241 = ( x17 & n18239 ) | ( x17 & ~n18240 ) | ( n18239 & ~n18240 ) ;
  assign n18242 = ( n18057 & ~n18232 ) | ( n18057 & n18241 ) | ( ~n18232 & n18241 ) ;
  assign n18243 = ( n18057 & n18232 ) | ( n18057 & n18241 ) | ( n18232 & n18241 ) ;
  assign n18244 = ( n18232 & n18242 ) | ( n18232 & ~n18243 ) | ( n18242 & ~n18243 ) ;
  assign n18245 = n5966 & ~n16957 ;
  assign n18246 = n6464 & ~n16043 ;
  assign n18247 = n5970 & ~n16047 ;
  assign n18248 = n5969 & ~n16045 ;
  assign n18249 = n18247 | n18248 ;
  assign n18250 = ( ~n18245 & n18246 ) | ( ~n18245 & n18249 ) | ( n18246 & n18249 ) ;
  assign n18251 = ( ~x14 & n18245 ) | ( ~x14 & n18250 ) | ( n18245 & n18250 ) ;
  assign n18252 = ( n18245 & n18250 ) | ( n18245 & ~n18251 ) | ( n18250 & ~n18251 ) ;
  assign n18253 = ( x14 & n18251 ) | ( x14 & ~n18252 ) | ( n18251 & ~n18252 ) ;
  assign n18254 = ( n18060 & ~n18244 ) | ( n18060 & n18253 ) | ( ~n18244 & n18253 ) ;
  assign n18255 = ( n18060 & n18244 ) | ( n18060 & n18253 ) | ( n18244 & n18253 ) ;
  assign n18256 = ( n18244 & n18254 ) | ( n18244 & ~n18255 ) | ( n18254 & ~n18255 ) ;
  assign n18257 = ( n18072 & n18139 ) | ( n18072 & ~n18256 ) | ( n18139 & ~n18256 ) ;
  assign n18258 = ( ~n18072 & n18139 ) | ( ~n18072 & n18256 ) | ( n18139 & n18256 ) ;
  assign n18259 = ( ~n18139 & n18257 ) | ( ~n18139 & n18258 ) | ( n18257 & n18258 ) ;
  assign n18260 = ( n18075 & n18130 ) | ( n18075 & ~n18259 ) | ( n18130 & ~n18259 ) ;
  assign n18261 = ( ~n18075 & n18130 ) | ( ~n18075 & n18259 ) | ( n18130 & n18259 ) ;
  assign n18262 = ( ~n18130 & n18260 ) | ( ~n18130 & n18261 ) | ( n18260 & n18261 ) ;
  assign n18263 = ( n18087 & n18121 ) | ( n18087 & ~n18262 ) | ( n18121 & ~n18262 ) ;
  assign n18264 = ( n18087 & ~n18121 ) | ( n18087 & n18262 ) | ( ~n18121 & n18262 ) ;
  assign n18265 = ( ~n18087 & n18263 ) | ( ~n18087 & n18264 ) | ( n18263 & n18264 ) ;
  assign n18266 = ( n18101 & n18112 ) | ( n18101 & ~n18265 ) | ( n18112 & ~n18265 ) ;
  assign n18267 = ( ~n16019 & n16114 ) | ( ~n16019 & n16140 ) | ( n16114 & n16140 ) ;
  assign n18268 = n36 & ~n18267 ;
  assign n18269 = n8967 & n16021 ;
  assign n18270 = ( x0 & n8966 ) | ( x0 & ~n16019 ) | ( n8966 & ~n16019 ) ;
  assign n18271 = ( n8966 & n18269 ) | ( n8966 & ~n18270 ) | ( n18269 & ~n18270 ) ;
  assign n18272 = n35 & n16017 ;
  assign n18273 = ( n35 & n18271 ) | ( n35 & ~n18272 ) | ( n18271 & ~n18272 ) ;
  assign n18274 = ( ~x2 & n18268 ) | ( ~x2 & n18273 ) | ( n18268 & n18273 ) ;
  assign n18275 = ( n18268 & n18273 ) | ( n18268 & ~n18274 ) | ( n18273 & ~n18274 ) ;
  assign n18276 = ( x2 & n18274 ) | ( x2 & ~n18275 ) | ( n18274 & ~n18275 ) ;
  assign n18277 = n8230 & n17968 ;
  assign n18278 = n8229 & n16023 ;
  assign n18279 = n8226 & ~n16027 ;
  assign n18280 = n8225 & ~n16025 ;
  assign n18281 = n18279 | n18280 ;
  assign n18282 = ( ~n18277 & n18278 ) | ( ~n18277 & n18281 ) | ( n18278 & n18281 ) ;
  assign n18283 = ( ~x5 & n18277 ) | ( ~x5 & n18282 ) | ( n18277 & n18282 ) ;
  assign n18284 = ( n18277 & n18282 ) | ( n18277 & ~n18283 ) | ( n18282 & ~n18283 ) ;
  assign n18285 = ( x5 & n18283 ) | ( x5 & ~n18284 ) | ( n18283 & ~n18284 ) ;
  assign n18286 = n7296 & ~n17528 ;
  assign n18287 = n7879 & ~n16029 ;
  assign n18288 = n7300 & ~n16033 ;
  assign n18289 = n7299 & n16031 ;
  assign n18290 = n18288 | n18289 ;
  assign n18291 = ( ~n18286 & n18287 ) | ( ~n18286 & n18290 ) | ( n18287 & n18290 ) ;
  assign n18292 = ( ~x8 & n18286 ) | ( ~x8 & n18291 ) | ( n18286 & n18291 ) ;
  assign n18293 = ( n18286 & n18291 ) | ( n18286 & ~n18292 ) | ( n18291 & ~n18292 ) ;
  assign n18294 = ( x8 & n18292 ) | ( x8 & ~n18293 ) | ( n18292 & ~n18293 ) ;
  assign n18295 = n1680 | n2011 ;
  assign n18296 = n1185 | n1205 ;
  assign n18297 = n76 | n148 ;
  assign n18298 = ( n217 & ~n356 ) | ( n217 & n435 ) | ( ~n356 & n435 ) ;
  assign n18299 = n356 | n18298 ;
  assign n18300 = ( ~n54 & n129 ) | ( ~n54 & n1031 ) | ( n129 & n1031 ) ;
  assign n18301 = ( ~n18297 & n18299 ) | ( ~n18297 & n18300 ) | ( n18299 & n18300 ) ;
  assign n18302 = n18297 | n18301 ;
  assign n18303 = ( ~n18295 & n18296 ) | ( ~n18295 & n18302 ) | ( n18296 & n18302 ) ;
  assign n18304 = n18295 | n18303 ;
  assign n18305 = n781 | n4569 ;
  assign n18306 = ( n2169 & n10120 ) | ( n2169 & ~n18305 ) | ( n10120 & ~n18305 ) ;
  assign n18307 = n18305 | n18306 ;
  assign n18308 = ( n3904 & n4267 ) | ( n3904 & ~n18307 ) | ( n4267 & ~n18307 ) ;
  assign n18309 = n18307 | n18308 ;
  assign n18310 = ( ~n6124 & n18304 ) | ( ~n6124 & n18309 ) | ( n18304 & n18309 ) ;
  assign n18311 = n5129 & ~n18310 ;
  assign n18312 = ( n6124 & n11990 ) | ( n6124 & n18311 ) | ( n11990 & n18311 ) ;
  assign n18313 = n18311 & ~n18312 ;
  assign n18314 = ( n1248 & n16077 ) | ( n1248 & ~n16082 ) | ( n16077 & ~n16082 ) ;
  assign n18315 = ~n16198 & n18314 ;
  assign n18316 = n607 & ~n16081 ;
  assign n18317 = n1250 & ~n16079 ;
  assign n18318 = n18316 | n18317 ;
  assign n18319 = n606 & ~n16077 ;
  assign n18320 = ( n606 & n18318 ) | ( n606 & ~n18319 ) | ( n18318 & ~n18319 ) ;
  assign n18321 = ( n1248 & ~n18315 ) | ( n1248 & n18320 ) | ( ~n18315 & n18320 ) ;
  assign n18322 = ( n18182 & ~n18313 ) | ( n18182 & n18321 ) | ( ~n18313 & n18321 ) ;
  assign n18323 = ( n18182 & n18313 ) | ( n18182 & n18321 ) | ( n18313 & n18321 ) ;
  assign n18324 = ( n18313 & n18322 ) | ( n18313 & ~n18323 ) | ( n18322 & ~n18323 ) ;
  assign n18325 = n3800 & n16209 ;
  assign n18326 = n3799 & n16071 ;
  assign n18327 = n3700 & ~n16075 ;
  assign n18328 = n3802 & ~n16073 ;
  assign n18329 = n18327 | n18328 ;
  assign n18330 = ( ~n18325 & n18326 ) | ( ~n18325 & n18329 ) | ( n18326 & n18329 ) ;
  assign n18331 = ( ~x29 & n18325 ) | ( ~x29 & n18330 ) | ( n18325 & n18330 ) ;
  assign n18332 = ( n18325 & n18330 ) | ( n18325 & ~n18331 ) | ( n18330 & ~n18331 ) ;
  assign n18333 = ( x29 & n18331 ) | ( x29 & ~n18332 ) | ( n18331 & ~n18332 ) ;
  assign n18334 = ( n18194 & ~n18324 ) | ( n18194 & n18333 ) | ( ~n18324 & n18333 ) ;
  assign n18335 = ( n18194 & n18324 ) | ( n18194 & n18333 ) | ( n18324 & n18333 ) ;
  assign n18336 = ( n18324 & n18334 ) | ( n18324 & ~n18335 ) | ( n18334 & ~n18335 ) ;
  assign n18337 = n4202 & n16281 ;
  assign n18338 = n4201 & n16065 ;
  assign n18339 = n4200 & n16069 ;
  assign n18340 = n4345 & n16067 ;
  assign n18341 = n18339 | n18340 ;
  assign n18342 = ( ~n18337 & n18338 ) | ( ~n18337 & n18341 ) | ( n18338 & n18341 ) ;
  assign n18343 = ( ~x26 & n18337 ) | ( ~x26 & n18342 ) | ( n18337 & n18342 ) ;
  assign n18344 = ( n18337 & n18342 ) | ( n18337 & ~n18343 ) | ( n18342 & ~n18343 ) ;
  assign n18345 = ( x26 & n18343 ) | ( x26 & ~n18344 ) | ( n18343 & ~n18344 ) ;
  assign n18346 = ( n18206 & ~n18336 ) | ( n18206 & n18345 ) | ( ~n18336 & n18345 ) ;
  assign n18347 = ( n18206 & n18336 ) | ( n18206 & n18345 ) | ( n18336 & n18345 ) ;
  assign n18348 = ( n18336 & n18346 ) | ( n18336 & ~n18347 ) | ( n18346 & ~n18347 ) ;
  assign n18349 = n4713 & ~n16433 ;
  assign n18350 = n4712 & n16059 ;
  assign n18351 = n4709 & n16063 ;
  assign n18352 = n4792 & ~n16061 ;
  assign n18353 = n18351 | n18352 ;
  assign n18354 = ( ~n18349 & n18350 ) | ( ~n18349 & n18353 ) | ( n18350 & n18353 ) ;
  assign n18355 = ( ~x23 & n18349 ) | ( ~x23 & n18354 ) | ( n18349 & n18354 ) ;
  assign n18356 = ( n18349 & n18354 ) | ( n18349 & ~n18355 ) | ( n18354 & ~n18355 ) ;
  assign n18357 = ( x23 & n18355 ) | ( x23 & ~n18356 ) | ( n18355 & ~n18356 ) ;
  assign n18358 = ( n18218 & ~n18348 ) | ( n18218 & n18357 ) | ( ~n18348 & n18357 ) ;
  assign n18359 = ( n18218 & n18348 ) | ( n18218 & n18357 ) | ( n18348 & n18357 ) ;
  assign n18360 = ( n18348 & n18358 ) | ( n18348 & ~n18359 ) | ( n18358 & ~n18359 ) ;
  assign n18361 = n4974 & n16553 ;
  assign n18362 = n5398 & n16053 ;
  assign n18363 = n4973 & ~n16057 ;
  assign n18364 = n4972 & ~n16055 ;
  assign n18365 = n18363 | n18364 ;
  assign n18366 = ( ~n18361 & n18362 ) | ( ~n18361 & n18365 ) | ( n18362 & n18365 ) ;
  assign n18367 = ( ~x20 & n18361 ) | ( ~x20 & n18366 ) | ( n18361 & n18366 ) ;
  assign n18368 = ( n18361 & n18366 ) | ( n18361 & ~n18367 ) | ( n18366 & ~n18367 ) ;
  assign n18369 = ( x20 & n18367 ) | ( x20 & ~n18368 ) | ( n18367 & ~n18368 ) ;
  assign n18370 = ( n18230 & ~n18360 ) | ( n18230 & n18369 ) | ( ~n18360 & n18369 ) ;
  assign n18371 = ( n18230 & n18360 ) | ( n18230 & n18369 ) | ( n18360 & n18369 ) ;
  assign n18372 = ( n18360 & n18370 ) | ( n18360 & ~n18371 ) | ( n18370 & ~n18371 ) ;
  assign n18373 = n5508 & ~n16801 ;
  assign n18374 = n5507 & ~n16047 ;
  assign n18375 = n5504 & ~n16051 ;
  assign n18376 = n5666 & ~n16049 ;
  assign n18377 = n18375 | n18376 ;
  assign n18378 = ( ~n18373 & n18374 ) | ( ~n18373 & n18377 ) | ( n18374 & n18377 ) ;
  assign n18379 = ( ~x17 & n18373 ) | ( ~x17 & n18378 ) | ( n18373 & n18378 ) ;
  assign n18380 = ( n18373 & n18378 ) | ( n18373 & ~n18379 ) | ( n18378 & ~n18379 ) ;
  assign n18381 = ( x17 & n18379 ) | ( x17 & ~n18380 ) | ( n18379 & ~n18380 ) ;
  assign n18382 = ( n18242 & ~n18372 ) | ( n18242 & n18381 ) | ( ~n18372 & n18381 ) ;
  assign n18383 = ( n18242 & n18372 ) | ( n18242 & n18381 ) | ( n18372 & n18381 ) ;
  assign n18384 = ( n18372 & n18382 ) | ( n18372 & ~n18383 ) | ( n18382 & ~n18383 ) ;
  assign n18385 = n5966 & n16969 ;
  assign n18386 = n6464 & n16041 ;
  assign n18387 = n5970 & ~n16045 ;
  assign n18388 = n5969 & ~n16043 ;
  assign n18389 = n18387 | n18388 ;
  assign n18390 = ( ~n18385 & n18386 ) | ( ~n18385 & n18389 ) | ( n18386 & n18389 ) ;
  assign n18391 = ( ~x14 & n18385 ) | ( ~x14 & n18390 ) | ( n18385 & n18390 ) ;
  assign n18392 = ( n18385 & n18390 ) | ( n18385 & ~n18391 ) | ( n18390 & ~n18391 ) ;
  assign n18393 = ( x14 & n18391 ) | ( x14 & ~n18392 ) | ( n18391 & ~n18392 ) ;
  assign n18394 = ( n18254 & ~n18384 ) | ( n18254 & n18393 ) | ( ~n18384 & n18393 ) ;
  assign n18395 = ( n18254 & n18384 ) | ( n18254 & n18393 ) | ( n18384 & n18393 ) ;
  assign n18396 = ( n18384 & n18394 ) | ( n18384 & ~n18395 ) | ( n18394 & ~n18395 ) ;
  assign n18397 = n6584 & ~n17313 ;
  assign n18398 = n7022 & n16035 ;
  assign n18399 = n6588 & n16039 ;
  assign n18400 = n6587 & ~n16037 ;
  assign n18401 = n18399 | n18400 ;
  assign n18402 = ( ~n18397 & n18398 ) | ( ~n18397 & n18401 ) | ( n18398 & n18401 ) ;
  assign n18403 = ( ~x11 & n18397 ) | ( ~x11 & n18402 ) | ( n18397 & n18402 ) ;
  assign n18404 = ( n18397 & n18402 ) | ( n18397 & ~n18403 ) | ( n18402 & ~n18403 ) ;
  assign n18405 = ( x11 & n18403 ) | ( x11 & ~n18404 ) | ( n18403 & ~n18404 ) ;
  assign n18406 = ( n18257 & ~n18396 ) | ( n18257 & n18405 ) | ( ~n18396 & n18405 ) ;
  assign n18407 = ( n18257 & n18396 ) | ( n18257 & n18405 ) | ( n18396 & n18405 ) ;
  assign n18408 = ( n18396 & n18406 ) | ( n18396 & ~n18407 ) | ( n18406 & ~n18407 ) ;
  assign n18409 = ( n18260 & n18294 ) | ( n18260 & ~n18408 ) | ( n18294 & ~n18408 ) ;
  assign n18410 = ( ~n18260 & n18294 ) | ( ~n18260 & n18408 ) | ( n18294 & n18408 ) ;
  assign n18411 = ( ~n18294 & n18409 ) | ( ~n18294 & n18410 ) | ( n18409 & n18410 ) ;
  assign n18412 = ( n18263 & n18285 ) | ( n18263 & ~n18411 ) | ( n18285 & ~n18411 ) ;
  assign n18413 = ( n18263 & ~n18285 ) | ( n18263 & n18411 ) | ( ~n18285 & n18411 ) ;
  assign n18414 = ( ~n18263 & n18412 ) | ( ~n18263 & n18413 ) | ( n18412 & n18413 ) ;
  assign n18415 = ( n18266 & n18276 ) | ( n18266 & ~n18414 ) | ( n18276 & ~n18414 ) ;
  assign n18416 = ( ~n16114 & n16115 ) | ( ~n16114 & n16141 ) | ( n16115 & n16141 ) ;
  assign n18417 = n36 & ~n18416 ;
  assign n18418 = n8967 & n16019 ;
  assign n18419 = ( x0 & n8966 ) | ( x0 & n16017 ) | ( n8966 & n16017 ) ;
  assign n18420 = ( n8966 & n18418 ) | ( n8966 & ~n18419 ) | ( n18418 & ~n18419 ) ;
  assign n18421 = n35 & ~n16015 ;
  assign n18422 = ( n35 & n18420 ) | ( n35 & ~n18421 ) | ( n18420 & ~n18421 ) ;
  assign n18423 = ( ~x2 & n18417 ) | ( ~x2 & n18422 ) | ( n18417 & n18422 ) ;
  assign n18424 = ( n18417 & n18422 ) | ( n18417 & ~n18423 ) | ( n18422 & ~n18423 ) ;
  assign n18425 = ( x2 & n18423 ) | ( x2 & ~n18424 ) | ( n18423 & ~n18424 ) ;
  assign n18426 = n8230 & ~n18091 ;
  assign n18427 = n8229 & n16021 ;
  assign n18428 = n8226 & ~n16025 ;
  assign n18429 = n8225 & n16023 ;
  assign n18430 = n18428 | n18429 ;
  assign n18431 = ( ~n18426 & n18427 ) | ( ~n18426 & n18430 ) | ( n18427 & n18430 ) ;
  assign n18432 = ( ~x5 & n18426 ) | ( ~x5 & n18431 ) | ( n18426 & n18431 ) ;
  assign n18433 = ( n18426 & n18431 ) | ( n18426 & ~n18432 ) | ( n18431 & ~n18432 ) ;
  assign n18434 = ( x5 & n18432 ) | ( x5 & ~n18433 ) | ( n18432 & ~n18433 ) ;
  assign n18435 = n6584 & ~n17412 ;
  assign n18436 = n7022 & ~n16033 ;
  assign n18437 = n6588 & ~n16037 ;
  assign n18438 = n6587 & n16035 ;
  assign n18439 = n18437 | n18438 ;
  assign n18440 = ( ~n18435 & n18436 ) | ( ~n18435 & n18439 ) | ( n18436 & n18439 ) ;
  assign n18441 = ( ~x11 & n18435 ) | ( ~x11 & n18440 ) | ( n18435 & n18440 ) ;
  assign n18442 = ( n18435 & n18440 ) | ( n18435 & ~n18441 ) | ( n18440 & ~n18441 ) ;
  assign n18443 = ( x11 & n18441 ) | ( x11 & ~n18442 ) | ( n18441 & ~n18442 ) ;
  assign n18444 = n5508 & ~n16876 ;
  assign n18445 = n5507 & ~n16045 ;
  assign n18446 = n5504 & ~n16049 ;
  assign n18447 = n5666 & ~n16047 ;
  assign n18448 = n18446 | n18447 ;
  assign n18449 = ( ~n18444 & n18445 ) | ( ~n18444 & n18448 ) | ( n18445 & n18448 ) ;
  assign n18450 = ( ~x17 & n18444 ) | ( ~x17 & n18449 ) | ( n18444 & n18449 ) ;
  assign n18451 = ( n18444 & n18449 ) | ( n18444 & ~n18450 ) | ( n18449 & ~n18450 ) ;
  assign n18452 = ( x17 & n18450 ) | ( x17 & ~n18451 ) | ( n18450 & ~n18451 ) ;
  assign n18453 = n4713 & ~n16484 ;
  assign n18454 = n4712 & ~n16057 ;
  assign n18455 = n4709 & ~n16061 ;
  assign n18456 = n4792 & n16059 ;
  assign n18457 = n18455 | n18456 ;
  assign n18458 = ( ~n18453 & n18454 ) | ( ~n18453 & n18457 ) | ( n18454 & n18457 ) ;
  assign n18459 = ( ~x23 & n18453 ) | ( ~x23 & n18458 ) | ( n18453 & n18458 ) ;
  assign n18460 = ( n18453 & n18458 ) | ( n18453 & ~n18459 ) | ( n18458 & ~n18459 ) ;
  assign n18461 = ( x23 & n18459 ) | ( x23 & ~n18460 ) | ( n18459 & ~n18460 ) ;
  assign n18462 = n3800 & ~n16221 ;
  assign n18463 = n3799 & n16069 ;
  assign n18464 = n3700 & ~n16073 ;
  assign n18465 = n3802 & n16071 ;
  assign n18466 = n18464 | n18465 ;
  assign n18467 = ( ~n18462 & n18463 ) | ( ~n18462 & n18466 ) | ( n18463 & n18466 ) ;
  assign n18468 = ( ~x29 & n18462 ) | ( ~x29 & n18467 ) | ( n18462 & n18467 ) ;
  assign n18469 = ( n18462 & n18467 ) | ( n18462 & ~n18468 ) | ( n18467 & ~n18468 ) ;
  assign n18470 = ( x29 & n18468 ) | ( x29 & ~n18469 ) | ( n18468 & ~n18469 ) ;
  assign n18471 = n2569 | n5002 ;
  assign n18472 = n226 | n1002 ;
  assign n18473 = n782 | n1032 ;
  assign n18474 = n138 | n689 ;
  assign n18475 = ( n73 & n109 ) | ( n73 & n129 ) | ( n109 & n129 ) ;
  assign n18476 = n133 | n18475 ;
  assign n18477 = ( n865 & ~n18474 ) | ( n865 & n18476 ) | ( ~n18474 & n18476 ) ;
  assign n18478 = n18474 | n18477 ;
  assign n18479 = ( ~n18472 & n18473 ) | ( ~n18472 & n18478 ) | ( n18473 & n18478 ) ;
  assign n18480 = n18472 | n18479 ;
  assign n18481 = n702 | n2898 ;
  assign n18482 = ( ~n18471 & n18480 ) | ( ~n18471 & n18481 ) | ( n18480 & n18481 ) ;
  assign n18483 = n18471 | n18482 ;
  assign n18484 = ( ~n4226 & n5177 ) | ( ~n4226 & n18483 ) | ( n5177 & n18483 ) ;
  assign n18485 = ( n2042 & ~n2880 ) | ( n2042 & n4226 ) | ( ~n2880 & n4226 ) ;
  assign n18486 = ( n2880 & ~n18484 ) | ( n2880 & n18485 ) | ( ~n18484 & n18485 ) ;
  assign n18487 = n18484 | n18486 ;
  assign n18488 = n607 & ~n16079 ;
  assign n18489 = n1250 & n16077 ;
  assign n18490 = n18488 | n18489 ;
  assign n18491 = n606 & n16075 ;
  assign n18492 = ( n606 & n18490 ) | ( n606 & ~n18491 ) | ( n18490 & ~n18491 ) ;
  assign n18493 = n1248 & n16169 ;
  assign n18494 = n18492 | n18493 ;
  assign n18495 = ( n18322 & n18487 ) | ( n18322 & n18494 ) | ( n18487 & n18494 ) ;
  assign n18496 = ( n18322 & ~n18487 ) | ( n18322 & n18494 ) | ( ~n18487 & n18494 ) ;
  assign n18497 = ( n18487 & ~n18495 ) | ( n18487 & n18496 ) | ( ~n18495 & n18496 ) ;
  assign n18498 = ( n18334 & n18470 ) | ( n18334 & n18497 ) | ( n18470 & n18497 ) ;
  assign n18499 = ( n18334 & ~n18470 ) | ( n18334 & n18497 ) | ( ~n18470 & n18497 ) ;
  assign n18500 = ( n18470 & ~n18498 ) | ( n18470 & n18499 ) | ( ~n18498 & n18499 ) ;
  assign n18501 = n4202 & n16315 ;
  assign n18502 = n4201 & n16063 ;
  assign n18503 = n4200 & n16067 ;
  assign n18504 = n4345 & n16065 ;
  assign n18505 = n18503 | n18504 ;
  assign n18506 = ( ~n18501 & n18502 ) | ( ~n18501 & n18505 ) | ( n18502 & n18505 ) ;
  assign n18507 = ( ~x26 & n18501 ) | ( ~x26 & n18506 ) | ( n18501 & n18506 ) ;
  assign n18508 = ( n18501 & n18506 ) | ( n18501 & ~n18507 ) | ( n18506 & ~n18507 ) ;
  assign n18509 = ( x26 & n18507 ) | ( x26 & ~n18508 ) | ( n18507 & ~n18508 ) ;
  assign n18510 = ( n18346 & n18500 ) | ( n18346 & n18509 ) | ( n18500 & n18509 ) ;
  assign n18511 = ( n18346 & ~n18500 ) | ( n18346 & n18509 ) | ( ~n18500 & n18509 ) ;
  assign n18512 = ( n18500 & ~n18510 ) | ( n18500 & n18511 ) | ( ~n18510 & n18511 ) ;
  assign n18513 = ( n18358 & n18461 ) | ( n18358 & n18512 ) | ( n18461 & n18512 ) ;
  assign n18514 = ( n18358 & ~n18461 ) | ( n18358 & n18512 ) | ( ~n18461 & n18512 ) ;
  assign n18515 = ( n18461 & ~n18513 ) | ( n18461 & n18514 ) | ( ~n18513 & n18514 ) ;
  assign n18516 = n4974 & n16611 ;
  assign n18517 = n5398 & ~n16051 ;
  assign n18518 = n4973 & ~n16055 ;
  assign n18519 = n4972 & n16053 ;
  assign n18520 = n18518 | n18519 ;
  assign n18521 = ( ~n18516 & n18517 ) | ( ~n18516 & n18520 ) | ( n18517 & n18520 ) ;
  assign n18522 = ( ~x20 & n18516 ) | ( ~x20 & n18521 ) | ( n18516 & n18521 ) ;
  assign n18523 = ( n18516 & n18521 ) | ( n18516 & ~n18522 ) | ( n18521 & ~n18522 ) ;
  assign n18524 = ( x20 & n18522 ) | ( x20 & ~n18523 ) | ( n18522 & ~n18523 ) ;
  assign n18525 = ( n18370 & n18515 ) | ( n18370 & n18524 ) | ( n18515 & n18524 ) ;
  assign n18526 = ( n18370 & ~n18515 ) | ( n18370 & n18524 ) | ( ~n18515 & n18524 ) ;
  assign n18527 = ( n18515 & ~n18525 ) | ( n18515 & n18526 ) | ( ~n18525 & n18526 ) ;
  assign n18528 = ( n18382 & n18452 ) | ( n18382 & n18527 ) | ( n18452 & n18527 ) ;
  assign n18529 = ( n18382 & ~n18452 ) | ( n18382 & n18527 ) | ( ~n18452 & n18527 ) ;
  assign n18530 = ( n18452 & ~n18528 ) | ( n18452 & n18529 ) | ( ~n18528 & n18529 ) ;
  assign n18531 = n5966 & ~n17051 ;
  assign n18532 = n6464 & n16039 ;
  assign n18533 = n5970 & ~n16043 ;
  assign n18534 = n5969 & n16041 ;
  assign n18535 = n18533 | n18534 ;
  assign n18536 = ( ~n18531 & n18532 ) | ( ~n18531 & n18535 ) | ( n18532 & n18535 ) ;
  assign n18537 = ( ~x14 & n18531 ) | ( ~x14 & n18536 ) | ( n18531 & n18536 ) ;
  assign n18538 = ( n18531 & n18536 ) | ( n18531 & ~n18537 ) | ( n18536 & ~n18537 ) ;
  assign n18539 = ( x14 & n18537 ) | ( x14 & ~n18538 ) | ( n18537 & ~n18538 ) ;
  assign n18540 = ( n18394 & n18530 ) | ( n18394 & n18539 ) | ( n18530 & n18539 ) ;
  assign n18541 = ( n18394 & ~n18530 ) | ( n18394 & n18539 ) | ( ~n18530 & n18539 ) ;
  assign n18542 = ( n18530 & ~n18540 ) | ( n18530 & n18541 ) | ( ~n18540 & n18541 ) ;
  assign n18543 = ( n18406 & n18443 ) | ( n18406 & n18542 ) | ( n18443 & n18542 ) ;
  assign n18544 = ( n18406 & ~n18443 ) | ( n18406 & n18542 ) | ( ~n18443 & n18542 ) ;
  assign n18545 = ( n18443 & ~n18543 ) | ( n18443 & n18544 ) | ( ~n18543 & n18544 ) ;
  assign n18546 = n7296 & n17634 ;
  assign n18547 = n7879 & ~n16027 ;
  assign n18548 = n7300 & n16031 ;
  assign n18549 = n7299 & ~n16029 ;
  assign n18550 = n18548 | n18549 ;
  assign n18551 = ( ~n18546 & n18547 ) | ( ~n18546 & n18550 ) | ( n18547 & n18550 ) ;
  assign n18552 = ( ~x8 & n18546 ) | ( ~x8 & n18551 ) | ( n18546 & n18551 ) ;
  assign n18553 = ( n18546 & n18551 ) | ( n18546 & ~n18552 ) | ( n18551 & ~n18552 ) ;
  assign n18554 = ( x8 & n18552 ) | ( x8 & ~n18553 ) | ( n18552 & ~n18553 ) ;
  assign n18555 = ( n18409 & n18545 ) | ( n18409 & n18554 ) | ( n18545 & n18554 ) ;
  assign n18556 = ( n18409 & ~n18545 ) | ( n18409 & n18554 ) | ( ~n18545 & n18554 ) ;
  assign n18557 = ( n18545 & ~n18555 ) | ( n18545 & n18556 ) | ( ~n18555 & n18556 ) ;
  assign n18558 = ( n18412 & n18434 ) | ( n18412 & n18557 ) | ( n18434 & n18557 ) ;
  assign n18559 = ( ~n18412 & n18434 ) | ( ~n18412 & n18557 ) | ( n18434 & n18557 ) ;
  assign n18560 = ( n18412 & ~n18558 ) | ( n18412 & n18559 ) | ( ~n18558 & n18559 ) ;
  assign n18561 = ( n18415 & n18425 ) | ( n18415 & n18560 ) | ( n18425 & n18560 ) ;
  assign n18562 = n1380 | n5554 ;
  assign n18563 = ( n66 & n80 ) | ( n66 & n149 ) | ( n80 & n149 ) ;
  assign n18564 = n995 | n18563 ;
  assign n18565 = ( ~n130 & n689 ) | ( ~n130 & n18564 ) | ( n689 & n18564 ) ;
  assign n18566 = ( n130 & n146 ) | ( n130 & ~n18565 ) | ( n146 & ~n18565 ) ;
  assign n18567 = n18565 | n18566 ;
  assign n18568 = n847 | n1893 ;
  assign n18569 = ( n4463 & n10207 ) | ( n4463 & ~n18568 ) | ( n10207 & ~n18568 ) ;
  assign n18570 = n18568 | n18569 ;
  assign n18571 = ( n10092 & ~n18567 ) | ( n10092 & n18570 ) | ( ~n18567 & n18570 ) ;
  assign n18572 = ( ~n18562 & n18567 ) | ( ~n18562 & n18571 ) | ( n18567 & n18571 ) ;
  assign n18573 = n10078 | n18562 ;
  assign n18574 = ( n11962 & n18572 ) | ( n11962 & ~n18573 ) | ( n18572 & ~n18573 ) ;
  assign n18575 = ~n18572 & n18574 ;
  assign n18576 = n607 & n16077 ;
  assign n18577 = n1250 & ~n16075 ;
  assign n18578 = n18576 | n18577 ;
  assign n18579 = n606 & n16073 ;
  assign n18580 = ( n606 & n18578 ) | ( n606 & ~n18579 ) | ( n18578 & ~n18579 ) ;
  assign n18581 = n1248 & ~n16176 ;
  assign n18582 = n18580 | n18581 ;
  assign n18583 = ( n18495 & ~n18575 ) | ( n18495 & n18582 ) | ( ~n18575 & n18582 ) ;
  assign n18584 = ( n18495 & n18575 ) | ( n18495 & n18582 ) | ( n18575 & n18582 ) ;
  assign n18585 = ( n18575 & n18583 ) | ( n18575 & ~n18584 ) | ( n18583 & ~n18584 ) ;
  assign n18586 = n3800 & n16269 ;
  assign n18587 = n3799 & n16067 ;
  assign n18588 = n3700 & n16071 ;
  assign n18589 = n3802 & n16069 ;
  assign n18590 = n18588 | n18589 ;
  assign n18591 = ( ~n18586 & n18587 ) | ( ~n18586 & n18590 ) | ( n18587 & n18590 ) ;
  assign n18592 = ( ~x29 & n18586 ) | ( ~x29 & n18591 ) | ( n18586 & n18591 ) ;
  assign n18593 = ( n18586 & n18591 ) | ( n18586 & ~n18592 ) | ( n18591 & ~n18592 ) ;
  assign n18594 = ( x29 & n18592 ) | ( x29 & ~n18593 ) | ( n18592 & ~n18593 ) ;
  assign n18595 = ( n18498 & ~n18585 ) | ( n18498 & n18594 ) | ( ~n18585 & n18594 ) ;
  assign n18596 = ( n18498 & n18585 ) | ( n18498 & n18594 ) | ( n18585 & n18594 ) ;
  assign n18597 = ( n18585 & n18595 ) | ( n18585 & ~n18596 ) | ( n18595 & ~n18596 ) ;
  assign n18598 = n4202 & ~n16354 ;
  assign n18599 = n4201 & ~n16061 ;
  assign n18600 = n4200 & n16065 ;
  assign n18601 = n4345 & n16063 ;
  assign n18602 = n18600 | n18601 ;
  assign n18603 = ( ~n18598 & n18599 ) | ( ~n18598 & n18602 ) | ( n18599 & n18602 ) ;
  assign n18604 = ( ~x26 & n18598 ) | ( ~x26 & n18603 ) | ( n18598 & n18603 ) ;
  assign n18605 = ( n18598 & n18603 ) | ( n18598 & ~n18604 ) | ( n18603 & ~n18604 ) ;
  assign n18606 = ( x26 & n18604 ) | ( x26 & ~n18605 ) | ( n18604 & ~n18605 ) ;
  assign n18607 = ( n18510 & ~n18597 ) | ( n18510 & n18606 ) | ( ~n18597 & n18606 ) ;
  assign n18608 = ( n18510 & n18597 ) | ( n18510 & n18606 ) | ( n18597 & n18606 ) ;
  assign n18609 = ( n18597 & n18607 ) | ( n18597 & ~n18608 ) | ( n18607 & ~n18608 ) ;
  assign n18610 = n4713 & n16541 ;
  assign n18611 = n4712 & ~n16055 ;
  assign n18612 = n4709 & n16059 ;
  assign n18613 = n4792 & ~n16057 ;
  assign n18614 = n18612 | n18613 ;
  assign n18615 = ( ~n18610 & n18611 ) | ( ~n18610 & n18614 ) | ( n18611 & n18614 ) ;
  assign n18616 = ( ~x23 & n18610 ) | ( ~x23 & n18615 ) | ( n18610 & n18615 ) ;
  assign n18617 = ( n18610 & n18615 ) | ( n18610 & ~n18616 ) | ( n18615 & ~n18616 ) ;
  assign n18618 = ( x23 & n18616 ) | ( x23 & ~n18617 ) | ( n18616 & ~n18617 ) ;
  assign n18619 = ( n18513 & ~n18609 ) | ( n18513 & n18618 ) | ( ~n18609 & n18618 ) ;
  assign n18620 = ( n18513 & n18609 ) | ( n18513 & n18618 ) | ( n18609 & n18618 ) ;
  assign n18621 = ( n18609 & n18619 ) | ( n18609 & ~n18620 ) | ( n18619 & ~n18620 ) ;
  assign n18622 = n4974 & ~n16674 ;
  assign n18623 = n5398 & ~n16049 ;
  assign n18624 = n4973 & n16053 ;
  assign n18625 = n4972 & ~n16051 ;
  assign n18626 = n18624 | n18625 ;
  assign n18627 = ( ~n18622 & n18623 ) | ( ~n18622 & n18626 ) | ( n18623 & n18626 ) ;
  assign n18628 = ( ~x20 & n18622 ) | ( ~x20 & n18627 ) | ( n18622 & n18627 ) ;
  assign n18629 = ( n18622 & n18627 ) | ( n18622 & ~n18628 ) | ( n18627 & ~n18628 ) ;
  assign n18630 = ( x20 & n18628 ) | ( x20 & ~n18629 ) | ( n18628 & ~n18629 ) ;
  assign n18631 = ( n18525 & ~n18621 ) | ( n18525 & n18630 ) | ( ~n18621 & n18630 ) ;
  assign n18632 = ( n18525 & n18621 ) | ( n18525 & n18630 ) | ( n18621 & n18630 ) ;
  assign n18633 = ( n18621 & n18631 ) | ( n18621 & ~n18632 ) | ( n18631 & ~n18632 ) ;
  assign n18634 = n5508 & ~n16957 ;
  assign n18635 = n5507 & ~n16043 ;
  assign n18636 = n5504 & ~n16047 ;
  assign n18637 = n5666 & ~n16045 ;
  assign n18638 = n18636 | n18637 ;
  assign n18639 = ( ~n18634 & n18635 ) | ( ~n18634 & n18638 ) | ( n18635 & n18638 ) ;
  assign n18640 = ( ~x17 & n18634 ) | ( ~x17 & n18639 ) | ( n18634 & n18639 ) ;
  assign n18641 = ( n18634 & n18639 ) | ( n18634 & ~n18640 ) | ( n18639 & ~n18640 ) ;
  assign n18642 = ( x17 & n18640 ) | ( x17 & ~n18641 ) | ( n18640 & ~n18641 ) ;
  assign n18643 = ( n18528 & ~n18633 ) | ( n18528 & n18642 ) | ( ~n18633 & n18642 ) ;
  assign n18644 = ( n18528 & n18633 ) | ( n18528 & n18642 ) | ( n18633 & n18642 ) ;
  assign n18645 = ( n18633 & n18643 ) | ( n18633 & ~n18644 ) | ( n18643 & ~n18644 ) ;
  assign n18646 = n5966 & ~n17138 ;
  assign n18647 = n6464 & ~n16037 ;
  assign n18648 = n5970 & n16041 ;
  assign n18649 = n5969 & n16039 ;
  assign n18650 = n18648 | n18649 ;
  assign n18651 = ( ~n18646 & n18647 ) | ( ~n18646 & n18650 ) | ( n18647 & n18650 ) ;
  assign n18652 = ( ~x14 & n18646 ) | ( ~x14 & n18651 ) | ( n18646 & n18651 ) ;
  assign n18653 = ( n18646 & n18651 ) | ( n18646 & ~n18652 ) | ( n18651 & ~n18652 ) ;
  assign n18654 = ( x14 & n18652 ) | ( x14 & ~n18653 ) | ( n18652 & ~n18653 ) ;
  assign n18655 = ( n18540 & ~n18645 ) | ( n18540 & n18654 ) | ( ~n18645 & n18654 ) ;
  assign n18656 = ( n18540 & n18645 ) | ( n18540 & n18654 ) | ( n18645 & n18654 ) ;
  assign n18657 = ( n18645 & n18655 ) | ( n18645 & ~n18656 ) | ( n18655 & ~n18656 ) ;
  assign n18658 = n6584 & ~n17516 ;
  assign n18659 = n7022 & n16031 ;
  assign n18660 = n6588 & n16035 ;
  assign n18661 = n6587 & ~n16033 ;
  assign n18662 = n18660 | n18661 ;
  assign n18663 = ( ~n18658 & n18659 ) | ( ~n18658 & n18662 ) | ( n18659 & n18662 ) ;
  assign n18664 = ( ~x11 & n18658 ) | ( ~x11 & n18663 ) | ( n18658 & n18663 ) ;
  assign n18665 = ( n18658 & n18663 ) | ( n18658 & ~n18664 ) | ( n18663 & ~n18664 ) ;
  assign n18666 = ( x11 & n18664 ) | ( x11 & ~n18665 ) | ( n18664 & ~n18665 ) ;
  assign n18667 = ( n18543 & ~n18657 ) | ( n18543 & n18666 ) | ( ~n18657 & n18666 ) ;
  assign n18668 = ( n18543 & n18657 ) | ( n18543 & n18666 ) | ( n18657 & n18666 ) ;
  assign n18669 = ( n18657 & n18667 ) | ( n18657 & ~n18668 ) | ( n18667 & ~n18668 ) ;
  assign n18670 = n7296 & ~n17746 ;
  assign n18671 = n7879 & ~n16025 ;
  assign n18672 = n7300 & ~n16029 ;
  assign n18673 = n7299 & ~n16027 ;
  assign n18674 = n18672 | n18673 ;
  assign n18675 = ( ~n18670 & n18671 ) | ( ~n18670 & n18674 ) | ( n18671 & n18674 ) ;
  assign n18676 = ( ~x8 & n18670 ) | ( ~x8 & n18675 ) | ( n18670 & n18675 ) ;
  assign n18677 = ( n18670 & n18675 ) | ( n18670 & ~n18676 ) | ( n18675 & ~n18676 ) ;
  assign n18678 = ( x8 & n18676 ) | ( x8 & ~n18677 ) | ( n18676 & ~n18677 ) ;
  assign n18679 = ( n18555 & ~n18669 ) | ( n18555 & n18678 ) | ( ~n18669 & n18678 ) ;
  assign n18680 = ( n18555 & n18669 ) | ( n18555 & n18678 ) | ( n18669 & n18678 ) ;
  assign n18681 = ( n18669 & n18679 ) | ( n18669 & ~n18680 ) | ( n18679 & ~n18680 ) ;
  assign n18682 = n8230 & n18103 ;
  assign n18683 = n8229 & n16019 ;
  assign n18684 = n8226 & n16023 ;
  assign n18685 = n8225 & n16021 ;
  assign n18686 = n18684 | n18685 ;
  assign n18687 = ( ~n18682 & n18683 ) | ( ~n18682 & n18686 ) | ( n18683 & n18686 ) ;
  assign n18688 = ( ~x5 & n18682 ) | ( ~x5 & n18687 ) | ( n18682 & n18687 ) ;
  assign n18689 = ( n18682 & n18687 ) | ( n18682 & ~n18688 ) | ( n18687 & ~n18688 ) ;
  assign n18690 = ( x5 & n18688 ) | ( x5 & ~n18689 ) | ( n18688 & ~n18689 ) ;
  assign n18691 = ( n18558 & ~n18681 ) | ( n18558 & n18690 ) | ( ~n18681 & n18690 ) ;
  assign n18692 = ( n18558 & n18681 ) | ( n18558 & n18690 ) | ( n18681 & n18690 ) ;
  assign n18693 = ( n18681 & n18691 ) | ( n18681 & ~n18692 ) | ( n18691 & ~n18692 ) ;
  assign n18694 = ( ~n16115 & n16116 ) | ( ~n16115 & n16142 ) | ( n16116 & n16142 ) ;
  assign n18695 = n36 & ~n18694 ;
  assign n18696 = n8967 & ~n16017 ;
  assign n18697 = ( x0 & n8966 ) | ( x0 & ~n16015 ) | ( n8966 & ~n16015 ) ;
  assign n18698 = ( n8966 & n18696 ) | ( n8966 & ~n18697 ) | ( n18696 & ~n18697 ) ;
  assign n18699 = n35 & n16013 ;
  assign n18700 = ( n35 & n18698 ) | ( n35 & ~n18699 ) | ( n18698 & ~n18699 ) ;
  assign n18701 = ( ~x2 & n18695 ) | ( ~x2 & n18700 ) | ( n18695 & n18700 ) ;
  assign n18702 = ( n18695 & n18700 ) | ( n18695 & ~n18701 ) | ( n18700 & ~n18701 ) ;
  assign n18703 = ( x2 & n18701 ) | ( x2 & ~n18702 ) | ( n18701 & ~n18702 ) ;
  assign n18704 = ( n18561 & ~n18693 ) | ( n18561 & n18703 ) | ( ~n18693 & n18703 ) ;
  assign n18705 = ~n4525 & n10516 ;
  assign n18706 = n1600 | n2067 ;
  assign n18707 = n133 | n1435 ;
  assign n18708 = ( n2833 & n18706 ) | ( n2833 & ~n18707 ) | ( n18706 & ~n18707 ) ;
  assign n18709 = ( n4121 & n18707 ) | ( n4121 & ~n18708 ) | ( n18707 & ~n18708 ) ;
  assign n18710 = n18708 | n18709 ;
  assign n18711 = n703 | n10202 ;
  assign n18712 = n807 | n2647 ;
  assign n18713 = ( n4837 & ~n18711 ) | ( n4837 & n18712 ) | ( ~n18711 & n18712 ) ;
  assign n18714 = n18711 | n18713 ;
  assign n18715 = ( n10516 & n18710 ) | ( n10516 & n18714 ) | ( n18710 & n18714 ) ;
  assign n18716 = ( n10571 & n18705 ) | ( n10571 & ~n18715 ) | ( n18705 & ~n18715 ) ;
  assign n18717 = ~n10571 & n18716 ;
  assign n18718 = n607 & ~n16075 ;
  assign n18719 = n1250 & ~n16073 ;
  assign n18720 = n18718 | n18719 ;
  assign n18721 = n606 & ~n16071 ;
  assign n18722 = ( n606 & n18720 ) | ( n606 & ~n18721 ) | ( n18720 & ~n18721 ) ;
  assign n18723 = n1248 & n16209 ;
  assign n18724 = n18722 | n18723 ;
  assign n18725 = ( n18583 & ~n18717 ) | ( n18583 & n18724 ) | ( ~n18717 & n18724 ) ;
  assign n18726 = ( n18583 & n18717 ) | ( n18583 & n18724 ) | ( n18717 & n18724 ) ;
  assign n18727 = ( n18717 & n18725 ) | ( n18717 & ~n18726 ) | ( n18725 & ~n18726 ) ;
  assign n18728 = n3800 & n16281 ;
  assign n18729 = n3799 & n16065 ;
  assign n18730 = n3700 & n16069 ;
  assign n18731 = n3802 & n16067 ;
  assign n18732 = n18730 | n18731 ;
  assign n18733 = ( ~n18728 & n18729 ) | ( ~n18728 & n18732 ) | ( n18729 & n18732 ) ;
  assign n18734 = ( ~x29 & n18728 ) | ( ~x29 & n18733 ) | ( n18728 & n18733 ) ;
  assign n18735 = ( n18728 & n18733 ) | ( n18728 & ~n18734 ) | ( n18733 & ~n18734 ) ;
  assign n18736 = ( x29 & n18734 ) | ( x29 & ~n18735 ) | ( n18734 & ~n18735 ) ;
  assign n18737 = ( n18595 & ~n18727 ) | ( n18595 & n18736 ) | ( ~n18727 & n18736 ) ;
  assign n18738 = ( n18595 & n18727 ) | ( n18595 & n18736 ) | ( n18727 & n18736 ) ;
  assign n18739 = ( n18727 & n18737 ) | ( n18727 & ~n18738 ) | ( n18737 & ~n18738 ) ;
  assign n18740 = n4202 & ~n16433 ;
  assign n18741 = n4201 & n16059 ;
  assign n18742 = n4200 & n16063 ;
  assign n18743 = n4345 & ~n16061 ;
  assign n18744 = n18742 | n18743 ;
  assign n18745 = ( ~n18740 & n18741 ) | ( ~n18740 & n18744 ) | ( n18741 & n18744 ) ;
  assign n18746 = ( ~x26 & n18740 ) | ( ~x26 & n18745 ) | ( n18740 & n18745 ) ;
  assign n18747 = ( n18740 & n18745 ) | ( n18740 & ~n18746 ) | ( n18745 & ~n18746 ) ;
  assign n18748 = ( x26 & n18746 ) | ( x26 & ~n18747 ) | ( n18746 & ~n18747 ) ;
  assign n18749 = ( n18607 & ~n18739 ) | ( n18607 & n18748 ) | ( ~n18739 & n18748 ) ;
  assign n18750 = ( n18607 & n18739 ) | ( n18607 & n18748 ) | ( n18739 & n18748 ) ;
  assign n18751 = ( n18739 & n18749 ) | ( n18739 & ~n18750 ) | ( n18749 & ~n18750 ) ;
  assign n18752 = n4713 & n16553 ;
  assign n18753 = n4712 & n16053 ;
  assign n18754 = n4709 & ~n16057 ;
  assign n18755 = n4792 & ~n16055 ;
  assign n18756 = n18754 | n18755 ;
  assign n18757 = ( ~n18752 & n18753 ) | ( ~n18752 & n18756 ) | ( n18753 & n18756 ) ;
  assign n18758 = ( ~x23 & n18752 ) | ( ~x23 & n18757 ) | ( n18752 & n18757 ) ;
  assign n18759 = ( n18752 & n18757 ) | ( n18752 & ~n18758 ) | ( n18757 & ~n18758 ) ;
  assign n18760 = ( x23 & n18758 ) | ( x23 & ~n18759 ) | ( n18758 & ~n18759 ) ;
  assign n18761 = ( n18619 & ~n18751 ) | ( n18619 & n18760 ) | ( ~n18751 & n18760 ) ;
  assign n18762 = ( n18619 & n18751 ) | ( n18619 & n18760 ) | ( n18751 & n18760 ) ;
  assign n18763 = ( n18751 & n18761 ) | ( n18751 & ~n18762 ) | ( n18761 & ~n18762 ) ;
  assign n18764 = n4974 & ~n16801 ;
  assign n18765 = n5398 & ~n16047 ;
  assign n18766 = n4973 & ~n16051 ;
  assign n18767 = n4972 & ~n16049 ;
  assign n18768 = n18766 | n18767 ;
  assign n18769 = ( ~n18764 & n18765 ) | ( ~n18764 & n18768 ) | ( n18765 & n18768 ) ;
  assign n18770 = ( ~x20 & n18764 ) | ( ~x20 & n18769 ) | ( n18764 & n18769 ) ;
  assign n18771 = ( n18764 & n18769 ) | ( n18764 & ~n18770 ) | ( n18769 & ~n18770 ) ;
  assign n18772 = ( x20 & n18770 ) | ( x20 & ~n18771 ) | ( n18770 & ~n18771 ) ;
  assign n18773 = ( n18631 & ~n18763 ) | ( n18631 & n18772 ) | ( ~n18763 & n18772 ) ;
  assign n18774 = ( n18631 & n18763 ) | ( n18631 & n18772 ) | ( n18763 & n18772 ) ;
  assign n18775 = ( n18763 & n18773 ) | ( n18763 & ~n18774 ) | ( n18773 & ~n18774 ) ;
  assign n18776 = n5508 & n16969 ;
  assign n18777 = n5507 & n16041 ;
  assign n18778 = n5504 & ~n16045 ;
  assign n18779 = n5666 & ~n16043 ;
  assign n18780 = n18778 | n18779 ;
  assign n18781 = ( ~n18776 & n18777 ) | ( ~n18776 & n18780 ) | ( n18777 & n18780 ) ;
  assign n18782 = ( ~x17 & n18776 ) | ( ~x17 & n18781 ) | ( n18776 & n18781 ) ;
  assign n18783 = ( n18776 & n18781 ) | ( n18776 & ~n18782 ) | ( n18781 & ~n18782 ) ;
  assign n18784 = ( x17 & n18782 ) | ( x17 & ~n18783 ) | ( n18782 & ~n18783 ) ;
  assign n18785 = ( n18643 & ~n18775 ) | ( n18643 & n18784 ) | ( ~n18775 & n18784 ) ;
  assign n18786 = ( n18643 & n18775 ) | ( n18643 & n18784 ) | ( n18775 & n18784 ) ;
  assign n18787 = ( n18775 & n18785 ) | ( n18775 & ~n18786 ) | ( n18785 & ~n18786 ) ;
  assign n18788 = n5966 & ~n17313 ;
  assign n18789 = n6464 & n16035 ;
  assign n18790 = n5970 & n16039 ;
  assign n18791 = n5969 & ~n16037 ;
  assign n18792 = n18790 | n18791 ;
  assign n18793 = ( ~n18788 & n18789 ) | ( ~n18788 & n18792 ) | ( n18789 & n18792 ) ;
  assign n18794 = ( ~x14 & n18788 ) | ( ~x14 & n18793 ) | ( n18788 & n18793 ) ;
  assign n18795 = ( n18788 & n18793 ) | ( n18788 & ~n18794 ) | ( n18793 & ~n18794 ) ;
  assign n18796 = ( x14 & n18794 ) | ( x14 & ~n18795 ) | ( n18794 & ~n18795 ) ;
  assign n18797 = ( n18655 & ~n18787 ) | ( n18655 & n18796 ) | ( ~n18787 & n18796 ) ;
  assign n18798 = ( n18655 & n18787 ) | ( n18655 & n18796 ) | ( n18787 & n18796 ) ;
  assign n18799 = ( n18787 & n18797 ) | ( n18787 & ~n18798 ) | ( n18797 & ~n18798 ) ;
  assign n18800 = n6584 & ~n17528 ;
  assign n18801 = n7022 & ~n16029 ;
  assign n18802 = n6588 & ~n16033 ;
  assign n18803 = n6587 & n16031 ;
  assign n18804 = n18802 | n18803 ;
  assign n18805 = ( ~n18800 & n18801 ) | ( ~n18800 & n18804 ) | ( n18801 & n18804 ) ;
  assign n18806 = ( ~x11 & n18800 ) | ( ~x11 & n18805 ) | ( n18800 & n18805 ) ;
  assign n18807 = ( n18800 & n18805 ) | ( n18800 & ~n18806 ) | ( n18805 & ~n18806 ) ;
  assign n18808 = ( x11 & n18806 ) | ( x11 & ~n18807 ) | ( n18806 & ~n18807 ) ;
  assign n18809 = ( n18667 & ~n18799 ) | ( n18667 & n18808 ) | ( ~n18799 & n18808 ) ;
  assign n18810 = ( n18667 & n18799 ) | ( n18667 & n18808 ) | ( n18799 & n18808 ) ;
  assign n18811 = ( n18799 & n18809 ) | ( n18799 & ~n18810 ) | ( n18809 & ~n18810 ) ;
  assign n18812 = n7296 & n17968 ;
  assign n18813 = n7879 & n16023 ;
  assign n18814 = n7300 & ~n16027 ;
  assign n18815 = n7299 & ~n16025 ;
  assign n18816 = n18814 | n18815 ;
  assign n18817 = ( ~n18812 & n18813 ) | ( ~n18812 & n18816 ) | ( n18813 & n18816 ) ;
  assign n18818 = ( ~x8 & n18812 ) | ( ~x8 & n18817 ) | ( n18812 & n18817 ) ;
  assign n18819 = ( n18812 & n18817 ) | ( n18812 & ~n18818 ) | ( n18817 & ~n18818 ) ;
  assign n18820 = ( x8 & n18818 ) | ( x8 & ~n18819 ) | ( n18818 & ~n18819 ) ;
  assign n18821 = ( n18679 & ~n18811 ) | ( n18679 & n18820 ) | ( ~n18811 & n18820 ) ;
  assign n18822 = ( n18679 & n18811 ) | ( n18679 & n18820 ) | ( n18811 & n18820 ) ;
  assign n18823 = ( n18811 & n18821 ) | ( n18811 & ~n18822 ) | ( n18821 & ~n18822 ) ;
  assign n18824 = n8230 & ~n18267 ;
  assign n18825 = n8229 & ~n16017 ;
  assign n18826 = n8226 & n16021 ;
  assign n18827 = n8225 & n16019 ;
  assign n18828 = n18826 | n18827 ;
  assign n18829 = ( ~n18824 & n18825 ) | ( ~n18824 & n18828 ) | ( n18825 & n18828 ) ;
  assign n18830 = ( ~x5 & n18824 ) | ( ~x5 & n18829 ) | ( n18824 & n18829 ) ;
  assign n18831 = ( n18824 & n18829 ) | ( n18824 & ~n18830 ) | ( n18829 & ~n18830 ) ;
  assign n18832 = ( x5 & n18830 ) | ( x5 & ~n18831 ) | ( n18830 & ~n18831 ) ;
  assign n18833 = ( n18691 & ~n18823 ) | ( n18691 & n18832 ) | ( ~n18823 & n18832 ) ;
  assign n18834 = ( n18691 & n18823 ) | ( n18691 & n18832 ) | ( n18823 & n18832 ) ;
  assign n18835 = ( n18823 & n18833 ) | ( n18823 & ~n18834 ) | ( n18833 & ~n18834 ) ;
  assign n18836 = ( n16153 & n18704 ) | ( n16153 & ~n18835 ) | ( n18704 & ~n18835 ) ;
  assign n18837 = ( n16153 & ~n18704 ) | ( n16153 & n18835 ) | ( ~n18704 & n18835 ) ;
  assign n18838 = ( ~n16153 & n18836 ) | ( ~n16153 & n18837 ) | ( n18836 & n18837 ) ;
  assign n18839 = ( ~n18561 & n18693 ) | ( ~n18561 & n18703 ) | ( n18693 & n18703 ) ;
  assign n18840 = ( ~n18703 & n18704 ) | ( ~n18703 & n18839 ) | ( n18704 & n18839 ) ;
  assign n18841 = n18838 | n18840 ;
  assign n18842 = ( n18838 & n18840 ) | ( n18838 & ~n18841 ) | ( n18840 & ~n18841 ) ;
  assign n18843 = n18841 & ~n18842 ;
  assign n18844 = ( ~n1667 & n3255 ) | ( ~n1667 & n11030 ) | ( n3255 & n11030 ) ;
  assign n18845 = n1235 | n1459 ;
  assign n18846 = n267 | n613 ;
  assign n18847 = ( n2926 & n18845 ) | ( n2926 & ~n18846 ) | ( n18845 & ~n18846 ) ;
  assign n18848 = ( n5985 & n18846 ) | ( n5985 & ~n18847 ) | ( n18846 & ~n18847 ) ;
  assign n18849 = n18847 | n18848 ;
  assign n18850 = ( n148 & n2628 ) | ( n148 & ~n11978 ) | ( n2628 & ~n11978 ) ;
  assign n18851 = n11978 | n18850 ;
  assign n18852 = n916 | n2363 ;
  assign n18853 = ( ~n807 & n2439 ) | ( ~n807 & n18852 ) | ( n2439 & n18852 ) ;
  assign n18854 = ~n18852 & n18853 ;
  assign n18855 = ( ~n6132 & n18851 ) | ( ~n6132 & n18854 ) | ( n18851 & n18854 ) ;
  assign n18856 = ~n18851 & n18855 ;
  assign n18857 = ( n11030 & ~n18849 ) | ( n11030 & n18856 ) | ( ~n18849 & n18856 ) ;
  assign n18858 = ( n1667 & ~n18844 ) | ( n1667 & n18857 ) | ( ~n18844 & n18857 ) ;
  assign n18859 = ~n1667 & n18858 ;
  assign n18860 = n607 & ~n16073 ;
  assign n18861 = n1250 & n16071 ;
  assign n18862 = n18860 | n18861 ;
  assign n18863 = n606 & ~n16069 ;
  assign n18864 = ( n606 & n18862 ) | ( n606 & ~n18863 ) | ( n18862 & ~n18863 ) ;
  assign n18865 = n1248 & ~n16221 ;
  assign n18866 = n18864 | n18865 ;
  assign n18867 = ( n18725 & ~n18859 ) | ( n18725 & n18866 ) | ( ~n18859 & n18866 ) ;
  assign n18868 = ( n18725 & n18859 ) | ( n18725 & n18866 ) | ( n18859 & n18866 ) ;
  assign n18869 = ( n18859 & n18867 ) | ( n18859 & ~n18868 ) | ( n18867 & ~n18868 ) ;
  assign n18870 = n3800 & n16315 ;
  assign n18871 = n3799 & n16063 ;
  assign n18872 = n3700 & n16067 ;
  assign n18873 = n3802 & n16065 ;
  assign n18874 = n18872 | n18873 ;
  assign n18875 = ( ~n18870 & n18871 ) | ( ~n18870 & n18874 ) | ( n18871 & n18874 ) ;
  assign n18876 = ( ~x29 & n18870 ) | ( ~x29 & n18875 ) | ( n18870 & n18875 ) ;
  assign n18877 = ( n18870 & n18875 ) | ( n18870 & ~n18876 ) | ( n18875 & ~n18876 ) ;
  assign n18878 = ( x29 & n18876 ) | ( x29 & ~n18877 ) | ( n18876 & ~n18877 ) ;
  assign n18879 = ( n18737 & ~n18869 ) | ( n18737 & n18878 ) | ( ~n18869 & n18878 ) ;
  assign n18880 = ( n18737 & n18869 ) | ( n18737 & n18878 ) | ( n18869 & n18878 ) ;
  assign n18881 = ( n18869 & n18879 ) | ( n18869 & ~n18880 ) | ( n18879 & ~n18880 ) ;
  assign n18882 = n4202 & ~n16484 ;
  assign n18883 = n4201 & ~n16057 ;
  assign n18884 = n4200 & ~n16061 ;
  assign n18885 = n4345 & n16059 ;
  assign n18886 = n18884 | n18885 ;
  assign n18887 = ( ~n18882 & n18883 ) | ( ~n18882 & n18886 ) | ( n18883 & n18886 ) ;
  assign n18888 = ( ~x26 & n18882 ) | ( ~x26 & n18887 ) | ( n18882 & n18887 ) ;
  assign n18889 = ( n18882 & n18887 ) | ( n18882 & ~n18888 ) | ( n18887 & ~n18888 ) ;
  assign n18890 = ( x26 & n18888 ) | ( x26 & ~n18889 ) | ( n18888 & ~n18889 ) ;
  assign n18891 = ( n18749 & ~n18881 ) | ( n18749 & n18890 ) | ( ~n18881 & n18890 ) ;
  assign n18892 = ( n18749 & n18881 ) | ( n18749 & n18890 ) | ( n18881 & n18890 ) ;
  assign n18893 = ( n18881 & n18891 ) | ( n18881 & ~n18892 ) | ( n18891 & ~n18892 ) ;
  assign n18894 = n4713 & n16611 ;
  assign n18895 = n4712 & ~n16051 ;
  assign n18896 = n4709 & ~n16055 ;
  assign n18897 = n4792 & n16053 ;
  assign n18898 = n18896 | n18897 ;
  assign n18899 = ( ~n18894 & n18895 ) | ( ~n18894 & n18898 ) | ( n18895 & n18898 ) ;
  assign n18900 = ( ~x23 & n18894 ) | ( ~x23 & n18899 ) | ( n18894 & n18899 ) ;
  assign n18901 = ( n18894 & n18899 ) | ( n18894 & ~n18900 ) | ( n18899 & ~n18900 ) ;
  assign n18902 = ( x23 & n18900 ) | ( x23 & ~n18901 ) | ( n18900 & ~n18901 ) ;
  assign n18903 = ( n18761 & ~n18893 ) | ( n18761 & n18902 ) | ( ~n18893 & n18902 ) ;
  assign n18904 = ( n18761 & n18893 ) | ( n18761 & n18902 ) | ( n18893 & n18902 ) ;
  assign n18905 = ( n18893 & n18903 ) | ( n18893 & ~n18904 ) | ( n18903 & ~n18904 ) ;
  assign n18906 = n4974 & ~n16876 ;
  assign n18907 = n5398 & ~n16045 ;
  assign n18908 = n4973 & ~n16049 ;
  assign n18909 = n4972 & ~n16047 ;
  assign n18910 = n18908 | n18909 ;
  assign n18911 = ( ~n18906 & n18907 ) | ( ~n18906 & n18910 ) | ( n18907 & n18910 ) ;
  assign n18912 = ( ~x20 & n18906 ) | ( ~x20 & n18911 ) | ( n18906 & n18911 ) ;
  assign n18913 = ( n18906 & n18911 ) | ( n18906 & ~n18912 ) | ( n18911 & ~n18912 ) ;
  assign n18914 = ( x20 & n18912 ) | ( x20 & ~n18913 ) | ( n18912 & ~n18913 ) ;
  assign n18915 = ( n18773 & ~n18905 ) | ( n18773 & n18914 ) | ( ~n18905 & n18914 ) ;
  assign n18916 = ( n18773 & n18905 ) | ( n18773 & n18914 ) | ( n18905 & n18914 ) ;
  assign n18917 = ( n18905 & n18915 ) | ( n18905 & ~n18916 ) | ( n18915 & ~n18916 ) ;
  assign n18918 = n5508 & ~n17051 ;
  assign n18919 = n5507 & n16039 ;
  assign n18920 = n5504 & ~n16043 ;
  assign n18921 = n5666 & n16041 ;
  assign n18922 = n18920 | n18921 ;
  assign n18923 = ( ~n18918 & n18919 ) | ( ~n18918 & n18922 ) | ( n18919 & n18922 ) ;
  assign n18924 = ( ~x17 & n18918 ) | ( ~x17 & n18923 ) | ( n18918 & n18923 ) ;
  assign n18925 = ( n18918 & n18923 ) | ( n18918 & ~n18924 ) | ( n18923 & ~n18924 ) ;
  assign n18926 = ( x17 & n18924 ) | ( x17 & ~n18925 ) | ( n18924 & ~n18925 ) ;
  assign n18927 = ( n18785 & ~n18917 ) | ( n18785 & n18926 ) | ( ~n18917 & n18926 ) ;
  assign n18928 = ( n18785 & n18917 ) | ( n18785 & n18926 ) | ( n18917 & n18926 ) ;
  assign n18929 = ( n18917 & n18927 ) | ( n18917 & ~n18928 ) | ( n18927 & ~n18928 ) ;
  assign n18930 = n5966 & ~n17412 ;
  assign n18931 = n6464 & ~n16033 ;
  assign n18932 = n5970 & ~n16037 ;
  assign n18933 = n5969 & n16035 ;
  assign n18934 = n18932 | n18933 ;
  assign n18935 = ( ~n18930 & n18931 ) | ( ~n18930 & n18934 ) | ( n18931 & n18934 ) ;
  assign n18936 = ( ~x14 & n18930 ) | ( ~x14 & n18935 ) | ( n18930 & n18935 ) ;
  assign n18937 = ( n18930 & n18935 ) | ( n18930 & ~n18936 ) | ( n18935 & ~n18936 ) ;
  assign n18938 = ( x14 & n18936 ) | ( x14 & ~n18937 ) | ( n18936 & ~n18937 ) ;
  assign n18939 = ( n18797 & ~n18929 ) | ( n18797 & n18938 ) | ( ~n18929 & n18938 ) ;
  assign n18940 = ( n18797 & n18929 ) | ( n18797 & n18938 ) | ( n18929 & n18938 ) ;
  assign n18941 = ( n18929 & n18939 ) | ( n18929 & ~n18940 ) | ( n18939 & ~n18940 ) ;
  assign n18942 = n6584 & n17634 ;
  assign n18943 = n7022 & ~n16027 ;
  assign n18944 = n6588 & n16031 ;
  assign n18945 = n6587 & ~n16029 ;
  assign n18946 = n18944 | n18945 ;
  assign n18947 = ( ~n18942 & n18943 ) | ( ~n18942 & n18946 ) | ( n18943 & n18946 ) ;
  assign n18948 = ( ~x11 & n18942 ) | ( ~x11 & n18947 ) | ( n18942 & n18947 ) ;
  assign n18949 = ( n18942 & n18947 ) | ( n18942 & ~n18948 ) | ( n18947 & ~n18948 ) ;
  assign n18950 = ( x11 & n18948 ) | ( x11 & ~n18949 ) | ( n18948 & ~n18949 ) ;
  assign n18951 = ( n18809 & ~n18941 ) | ( n18809 & n18950 ) | ( ~n18941 & n18950 ) ;
  assign n18952 = ( n18809 & n18941 ) | ( n18809 & n18950 ) | ( n18941 & n18950 ) ;
  assign n18953 = ( n18941 & n18951 ) | ( n18941 & ~n18952 ) | ( n18951 & ~n18952 ) ;
  assign n18954 = n7296 & ~n18091 ;
  assign n18955 = n7879 & n16021 ;
  assign n18956 = n7300 & ~n16025 ;
  assign n18957 = n7299 & n16023 ;
  assign n18958 = n18956 | n18957 ;
  assign n18959 = ( ~n18954 & n18955 ) | ( ~n18954 & n18958 ) | ( n18955 & n18958 ) ;
  assign n18960 = ( ~x8 & n18954 ) | ( ~x8 & n18959 ) | ( n18954 & n18959 ) ;
  assign n18961 = ( n18954 & n18959 ) | ( n18954 & ~n18960 ) | ( n18959 & ~n18960 ) ;
  assign n18962 = ( x8 & n18960 ) | ( x8 & ~n18961 ) | ( n18960 & ~n18961 ) ;
  assign n18963 = ( n18821 & ~n18953 ) | ( n18821 & n18962 ) | ( ~n18953 & n18962 ) ;
  assign n18964 = ( n18821 & n18953 ) | ( n18821 & n18962 ) | ( n18953 & n18962 ) ;
  assign n18965 = ( n18953 & n18963 ) | ( n18953 & ~n18964 ) | ( n18963 & ~n18964 ) ;
  assign n18966 = n8230 & ~n18416 ;
  assign n18967 = n8229 & n16015 ;
  assign n18968 = n8226 & n16019 ;
  assign n18969 = n8225 & ~n16017 ;
  assign n18970 = n18968 | n18969 ;
  assign n18971 = ( ~n18966 & n18967 ) | ( ~n18966 & n18970 ) | ( n18967 & n18970 ) ;
  assign n18972 = ( ~x5 & n18966 ) | ( ~x5 & n18971 ) | ( n18966 & n18971 ) ;
  assign n18973 = ( n18966 & n18971 ) | ( n18966 & ~n18972 ) | ( n18971 & ~n18972 ) ;
  assign n18974 = ( x5 & n18972 ) | ( x5 & ~n18973 ) | ( n18972 & ~n18973 ) ;
  assign n18975 = ( n18833 & ~n18965 ) | ( n18833 & n18974 ) | ( ~n18965 & n18974 ) ;
  assign n18976 = ( n18833 & n18965 ) | ( n18833 & n18974 ) | ( n18965 & n18974 ) ;
  assign n18977 = ( n18965 & n18975 ) | ( n18965 & ~n18976 ) | ( n18975 & ~n18976 ) ;
  assign n18978 = n3655 | n3689 ;
  assign n18979 = ( n460 & ~n16127 ) | ( n460 & n18978 ) | ( ~n16127 & n18978 ) ;
  assign n18980 = ( ~n460 & n16127 ) | ( ~n460 & n18978 ) | ( n16127 & n18978 ) ;
  assign n18981 = ( ~n18978 & n18979 ) | ( ~n18978 & n18980 ) | ( n18979 & n18980 ) ;
  assign n18982 = n1248 & ~n10362 ;
  assign n18983 = n1250 & ~n10302 ;
  assign n18984 = n606 | n607 ;
  assign n18985 = ( n606 & ~n10056 ) | ( n606 & n18984 ) | ( ~n10056 & n18984 ) ;
  assign n18986 = n18983 | n18985 ;
  assign n18987 = ( n1248 & ~n18982 ) | ( n1248 & n18986 ) | ( ~n18982 & n18986 ) ;
  assign n18988 = ( n16132 & n18981 ) | ( n16132 & n18987 ) | ( n18981 & n18987 ) ;
  assign n18989 = ( ~n16132 & n18981 ) | ( ~n16132 & n18987 ) | ( n18981 & n18987 ) ;
  assign n18990 = ( n16132 & ~n18988 ) | ( n16132 & n18989 ) | ( ~n18988 & n18989 ) ;
  assign n18991 = ( n16133 & n16136 ) | ( n16133 & n18990 ) | ( n16136 & n18990 ) ;
  assign n18992 = ( ~n16133 & n16136 ) | ( ~n16133 & n18990 ) | ( n16136 & n18990 ) ;
  assign n18993 = ( n16133 & ~n18991 ) | ( n16133 & n18992 ) | ( ~n18991 & n18992 ) ;
  assign n18994 = ( n16138 & n16139 ) | ( n16138 & n18993 ) | ( n16139 & n18993 ) ;
  assign n18995 = ( n16138 & ~n16139 ) | ( n16138 & n18993 ) | ( ~n16139 & n18993 ) ;
  assign n18996 = ( n16139 & ~n18994 ) | ( n16139 & n18995 ) | ( ~n18994 & n18995 ) ;
  assign n18997 = n36 & n18996 ;
  assign n18998 = n8967 & ~n16013 ;
  assign n18999 = ( x0 & n8966 ) | ( x0 & ~n16138 ) | ( n8966 & ~n16138 ) ;
  assign n19000 = ( n8966 & n18998 ) | ( n8966 & ~n18999 ) | ( n18998 & ~n18999 ) ;
  assign n19001 = n35 & ~n18993 ;
  assign n19002 = ( n35 & n19000 ) | ( n35 & ~n19001 ) | ( n19000 & ~n19001 ) ;
  assign n19003 = ( ~x2 & n18997 ) | ( ~x2 & n19002 ) | ( n18997 & n19002 ) ;
  assign n19004 = ( n18997 & n19002 ) | ( n18997 & ~n19003 ) | ( n19002 & ~n19003 ) ;
  assign n19005 = ( x2 & n19003 ) | ( x2 & ~n19004 ) | ( n19003 & ~n19004 ) ;
  assign n19006 = ( n18836 & ~n18977 ) | ( n18836 & n19005 ) | ( ~n18977 & n19005 ) ;
  assign n19007 = ( n18836 & n18977 ) | ( n18836 & n19005 ) | ( n18977 & n19005 ) ;
  assign n19008 = ( n18977 & n19006 ) | ( n18977 & ~n19007 ) | ( n19006 & ~n19007 ) ;
  assign n19009 = n18841 | n19008 ;
  assign n19010 = ( n18841 & n19008 ) | ( n18841 & ~n19009 ) | ( n19008 & ~n19009 ) ;
  assign n19011 = n19009 & ~n19010 ;
  assign n19012 = n8230 & ~n18694 ;
  assign n19013 = n8229 & ~n16013 ;
  assign n19014 = n8226 & ~n16017 ;
  assign n19015 = n8225 & n16015 ;
  assign n19016 = n19014 | n19015 ;
  assign n19017 = ( ~n19012 & n19013 ) | ( ~n19012 & n19016 ) | ( n19013 & n19016 ) ;
  assign n19018 = ( ~x5 & n19012 ) | ( ~x5 & n19017 ) | ( n19012 & n19017 ) ;
  assign n19019 = ( n19012 & n19017 ) | ( n19012 & ~n19018 ) | ( n19017 & ~n19018 ) ;
  assign n19020 = ( x5 & n19018 ) | ( x5 & ~n19019 ) | ( n19018 & ~n19019 ) ;
  assign n19021 = n6584 & ~n17746 ;
  assign n19022 = n7022 & ~n16025 ;
  assign n19023 = n6588 & ~n16029 ;
  assign n19024 = n6587 & ~n16027 ;
  assign n19025 = n19023 | n19024 ;
  assign n19026 = ( ~n19021 & n19022 ) | ( ~n19021 & n19025 ) | ( n19022 & n19025 ) ;
  assign n19027 = ( ~x11 & n19021 ) | ( ~x11 & n19026 ) | ( n19021 & n19026 ) ;
  assign n19028 = ( n19021 & n19026 ) | ( n19021 & ~n19027 ) | ( n19026 & ~n19027 ) ;
  assign n19029 = ( x11 & n19027 ) | ( x11 & ~n19028 ) | ( n19027 & ~n19028 ) ;
  assign n19030 = n5508 & ~n17138 ;
  assign n19031 = n5507 & ~n16037 ;
  assign n19032 = n5504 & n16041 ;
  assign n19033 = n5666 & n16039 ;
  assign n19034 = n19032 | n19033 ;
  assign n19035 = ( ~n19030 & n19031 ) | ( ~n19030 & n19034 ) | ( n19031 & n19034 ) ;
  assign n19036 = ( ~x17 & n19030 ) | ( ~x17 & n19035 ) | ( n19030 & n19035 ) ;
  assign n19037 = ( n19030 & n19035 ) | ( n19030 & ~n19036 ) | ( n19035 & ~n19036 ) ;
  assign n19038 = ( x17 & n19036 ) | ( x17 & ~n19037 ) | ( n19036 & ~n19037 ) ;
  assign n19039 = n4713 & ~n16674 ;
  assign n19040 = n4712 & ~n16049 ;
  assign n19041 = n4709 & n16053 ;
  assign n19042 = n4792 & ~n16051 ;
  assign n19043 = n19041 | n19042 ;
  assign n19044 = ( ~n19039 & n19040 ) | ( ~n19039 & n19043 ) | ( n19040 & n19043 ) ;
  assign n19045 = ( ~x23 & n19039 ) | ( ~x23 & n19044 ) | ( n19039 & n19044 ) ;
  assign n19046 = ( n19039 & n19044 ) | ( n19039 & ~n19045 ) | ( n19044 & ~n19045 ) ;
  assign n19047 = ( x23 & n19045 ) | ( x23 & ~n19046 ) | ( n19045 & ~n19046 ) ;
  assign n19048 = n3800 & ~n16354 ;
  assign n19049 = n3799 & ~n16061 ;
  assign n19050 = n3700 & n16065 ;
  assign n19051 = n3802 & n16063 ;
  assign n19052 = n19050 | n19051 ;
  assign n19053 = ( ~n19048 & n19049 ) | ( ~n19048 & n19052 ) | ( n19049 & n19052 ) ;
  assign n19054 = ( ~x29 & n19048 ) | ( ~x29 & n19053 ) | ( n19048 & n19053 ) ;
  assign n19055 = ( n19048 & n19053 ) | ( n19048 & ~n19054 ) | ( n19053 & ~n19054 ) ;
  assign n19056 = ( x29 & n19054 ) | ( x29 & ~n19055 ) | ( n19054 & ~n19055 ) ;
  assign n19057 = n2749 | n6041 ;
  assign n19058 = n2605 | n19057 ;
  assign n19059 = n1879 | n10626 ;
  assign n19060 = ( n4099 & n11053 ) | ( n4099 & ~n19059 ) | ( n11053 & ~n19059 ) ;
  assign n19061 = n19059 | n19060 ;
  assign n19062 = n1481 | n3273 ;
  assign n19063 = n130 | n1494 ;
  assign n19064 = n544 | n719 ;
  assign n19065 = n1116 | n19064 ;
  assign n19066 = ( n77 & n1173 ) | ( n77 & ~n19065 ) | ( n1173 & ~n19065 ) ;
  assign n19067 = n19065 | n19066 ;
  assign n19068 = ( ~n19062 & n19063 ) | ( ~n19062 & n19067 ) | ( n19063 & n19067 ) ;
  assign n19069 = n19062 | n19068 ;
  assign n19070 = ( ~n19057 & n19061 ) | ( ~n19057 & n19069 ) | ( n19061 & n19069 ) ;
  assign n19071 = ( ~n4080 & n19058 ) | ( ~n4080 & n19070 ) | ( n19058 & n19070 ) ;
  assign n19072 = n4080 | n19071 ;
  assign n19073 = n607 & n16071 ;
  assign n19074 = n1250 & n16069 ;
  assign n19075 = n19073 | n19074 ;
  assign n19076 = n606 & ~n16067 ;
  assign n19077 = ( n606 & n19075 ) | ( n606 & ~n19076 ) | ( n19075 & ~n19076 ) ;
  assign n19078 = n1248 & n16269 ;
  assign n19079 = n19077 | n19078 ;
  assign n19080 = ( n18867 & n19072 ) | ( n18867 & n19079 ) | ( n19072 & n19079 ) ;
  assign n19081 = ( n18867 & ~n19072 ) | ( n18867 & n19079 ) | ( ~n19072 & n19079 ) ;
  assign n19082 = ( n19072 & ~n19080 ) | ( n19072 & n19081 ) | ( ~n19080 & n19081 ) ;
  assign n19083 = ( n18879 & n19056 ) | ( n18879 & n19082 ) | ( n19056 & n19082 ) ;
  assign n19084 = ( n18879 & ~n19056 ) | ( n18879 & n19082 ) | ( ~n19056 & n19082 ) ;
  assign n19085 = ( n19056 & ~n19083 ) | ( n19056 & n19084 ) | ( ~n19083 & n19084 ) ;
  assign n19086 = n4202 & n16541 ;
  assign n19087 = n4201 & ~n16055 ;
  assign n19088 = n4200 & n16059 ;
  assign n19089 = n4345 & ~n16057 ;
  assign n19090 = n19088 | n19089 ;
  assign n19091 = ( ~n19086 & n19087 ) | ( ~n19086 & n19090 ) | ( n19087 & n19090 ) ;
  assign n19092 = ( ~x26 & n19086 ) | ( ~x26 & n19091 ) | ( n19086 & n19091 ) ;
  assign n19093 = ( n19086 & n19091 ) | ( n19086 & ~n19092 ) | ( n19091 & ~n19092 ) ;
  assign n19094 = ( x26 & n19092 ) | ( x26 & ~n19093 ) | ( n19092 & ~n19093 ) ;
  assign n19095 = ( n18891 & n19085 ) | ( n18891 & n19094 ) | ( n19085 & n19094 ) ;
  assign n19096 = ( n18891 & ~n19085 ) | ( n18891 & n19094 ) | ( ~n19085 & n19094 ) ;
  assign n19097 = ( n19085 & ~n19095 ) | ( n19085 & n19096 ) | ( ~n19095 & n19096 ) ;
  assign n19098 = ( n18903 & n19047 ) | ( n18903 & n19097 ) | ( n19047 & n19097 ) ;
  assign n19099 = ( n18903 & ~n19047 ) | ( n18903 & n19097 ) | ( ~n19047 & n19097 ) ;
  assign n19100 = ( n19047 & ~n19098 ) | ( n19047 & n19099 ) | ( ~n19098 & n19099 ) ;
  assign n19101 = n4974 & ~n16957 ;
  assign n19102 = n5398 & ~n16043 ;
  assign n19103 = n4973 & ~n16047 ;
  assign n19104 = n4972 & ~n16045 ;
  assign n19105 = n19103 | n19104 ;
  assign n19106 = ( ~n19101 & n19102 ) | ( ~n19101 & n19105 ) | ( n19102 & n19105 ) ;
  assign n19107 = ( ~x20 & n19101 ) | ( ~x20 & n19106 ) | ( n19101 & n19106 ) ;
  assign n19108 = ( n19101 & n19106 ) | ( n19101 & ~n19107 ) | ( n19106 & ~n19107 ) ;
  assign n19109 = ( x20 & n19107 ) | ( x20 & ~n19108 ) | ( n19107 & ~n19108 ) ;
  assign n19110 = ( n18915 & n19100 ) | ( n18915 & n19109 ) | ( n19100 & n19109 ) ;
  assign n19111 = ( n18915 & ~n19100 ) | ( n18915 & n19109 ) | ( ~n19100 & n19109 ) ;
  assign n19112 = ( n19100 & ~n19110 ) | ( n19100 & n19111 ) | ( ~n19110 & n19111 ) ;
  assign n19113 = ( n18927 & n19038 ) | ( n18927 & n19112 ) | ( n19038 & n19112 ) ;
  assign n19114 = ( n18927 & ~n19038 ) | ( n18927 & n19112 ) | ( ~n19038 & n19112 ) ;
  assign n19115 = ( n19038 & ~n19113 ) | ( n19038 & n19114 ) | ( ~n19113 & n19114 ) ;
  assign n19116 = n5966 & ~n17516 ;
  assign n19117 = n6464 & n16031 ;
  assign n19118 = n5970 & n16035 ;
  assign n19119 = n5969 & ~n16033 ;
  assign n19120 = n19118 | n19119 ;
  assign n19121 = ( ~n19116 & n19117 ) | ( ~n19116 & n19120 ) | ( n19117 & n19120 ) ;
  assign n19122 = ( ~x14 & n19116 ) | ( ~x14 & n19121 ) | ( n19116 & n19121 ) ;
  assign n19123 = ( n19116 & n19121 ) | ( n19116 & ~n19122 ) | ( n19121 & ~n19122 ) ;
  assign n19124 = ( x14 & n19122 ) | ( x14 & ~n19123 ) | ( n19122 & ~n19123 ) ;
  assign n19125 = ( n18939 & n19115 ) | ( n18939 & n19124 ) | ( n19115 & n19124 ) ;
  assign n19126 = ( n18939 & ~n19115 ) | ( n18939 & n19124 ) | ( ~n19115 & n19124 ) ;
  assign n19127 = ( n19115 & ~n19125 ) | ( n19115 & n19126 ) | ( ~n19125 & n19126 ) ;
  assign n19128 = ( n18951 & n19029 ) | ( n18951 & n19127 ) | ( n19029 & n19127 ) ;
  assign n19129 = ( n18951 & ~n19029 ) | ( n18951 & n19127 ) | ( ~n19029 & n19127 ) ;
  assign n19130 = ( n19029 & ~n19128 ) | ( n19029 & n19129 ) | ( ~n19128 & n19129 ) ;
  assign n19131 = n7296 & n18103 ;
  assign n19132 = n7879 & n16019 ;
  assign n19133 = n7300 & n16023 ;
  assign n19134 = n7299 & n16021 ;
  assign n19135 = n19133 | n19134 ;
  assign n19136 = ( ~n19131 & n19132 ) | ( ~n19131 & n19135 ) | ( n19132 & n19135 ) ;
  assign n19137 = ( ~x8 & n19131 ) | ( ~x8 & n19136 ) | ( n19131 & n19136 ) ;
  assign n19138 = ( n19131 & n19136 ) | ( n19131 & ~n19137 ) | ( n19136 & ~n19137 ) ;
  assign n19139 = ( x8 & n19137 ) | ( x8 & ~n19138 ) | ( n19137 & ~n19138 ) ;
  assign n19140 = ( n18963 & n19130 ) | ( n18963 & n19139 ) | ( n19130 & n19139 ) ;
  assign n19141 = ( n18963 & ~n19130 ) | ( n18963 & n19139 ) | ( ~n19130 & n19139 ) ;
  assign n19142 = ( n19130 & ~n19140 ) | ( n19130 & n19141 ) | ( ~n19140 & n19141 ) ;
  assign n19143 = ( n18975 & n19020 ) | ( n18975 & n19142 ) | ( n19020 & n19142 ) ;
  assign n19144 = ( n18975 & ~n19020 ) | ( n18975 & n19142 ) | ( ~n19020 & n19142 ) ;
  assign n19145 = ( n19020 & ~n19143 ) | ( n19020 & n19144 ) | ( ~n19143 & n19144 ) ;
  assign n19146 = ( ~n1248 & n10346 ) | ( ~n1248 & n10347 ) | ( n10346 & n10347 ) ;
  assign n19147 = n1250 | n18984 ;
  assign n19148 = ( n10346 & ~n19146 ) | ( n10346 & n19147 ) | ( ~n19146 & n19147 ) ;
  assign n19149 = ( n10343 & ~n16132 ) | ( n10343 & n18978 ) | ( ~n16132 & n18978 ) ;
  assign n19150 = ( n10343 & n16132 ) | ( n10343 & n18978 ) | ( n16132 & n18978 ) ;
  assign n19151 = ( n16132 & n19149 ) | ( n16132 & ~n19150 ) | ( n19149 & ~n19150 ) ;
  assign n19152 = ( n18979 & ~n19148 ) | ( n18979 & n19151 ) | ( ~n19148 & n19151 ) ;
  assign n19153 = ( n18979 & n19151 ) | ( n18979 & ~n19152 ) | ( n19151 & ~n19152 ) ;
  assign n19154 = ( n19148 & n19152 ) | ( n19148 & ~n19153 ) | ( n19152 & ~n19153 ) ;
  assign n19155 = ( n18988 & n18991 ) | ( n18988 & n19154 ) | ( n18991 & n19154 ) ;
  assign n19156 = ( ~n18988 & n18991 ) | ( ~n18988 & n19154 ) | ( n18991 & n19154 ) ;
  assign n19157 = ( n18988 & ~n19155 ) | ( n18988 & n19156 ) | ( ~n19155 & n19156 ) ;
  assign n19158 = ( n18993 & n18994 ) | ( n18993 & n19157 ) | ( n18994 & n19157 ) ;
  assign n19159 = ( ~n18993 & n18994 ) | ( ~n18993 & n19157 ) | ( n18994 & n19157 ) ;
  assign n19160 = ( n18993 & ~n19158 ) | ( n18993 & n19159 ) | ( ~n19158 & n19159 ) ;
  assign n19161 = n36 & n19160 ;
  assign n19162 = n8967 & n16138 ;
  assign n19163 = ( x0 & n8966 ) | ( x0 & ~n18993 ) | ( n8966 & ~n18993 ) ;
  assign n19164 = ( n8966 & n19162 ) | ( n8966 & ~n19163 ) | ( n19162 & ~n19163 ) ;
  assign n19165 = n35 & ~n19157 ;
  assign n19166 = ( n35 & n19164 ) | ( n35 & ~n19165 ) | ( n19164 & ~n19165 ) ;
  assign n19167 = ( ~x2 & n19161 ) | ( ~x2 & n19166 ) | ( n19161 & n19166 ) ;
  assign n19168 = ( n19161 & n19166 ) | ( n19161 & ~n19167 ) | ( n19166 & ~n19167 ) ;
  assign n19169 = ( x2 & n19167 ) | ( x2 & ~n19168 ) | ( n19167 & ~n19168 ) ;
  assign n19170 = ( n19006 & n19145 ) | ( n19006 & n19169 ) | ( n19145 & n19169 ) ;
  assign n19171 = ( ~n19006 & n19145 ) | ( ~n19006 & n19169 ) | ( n19145 & n19169 ) ;
  assign n19172 = ( n19006 & ~n19170 ) | ( n19006 & n19171 ) | ( ~n19170 & n19171 ) ;
  assign n19173 = ~n19009 & n19172 ;
  assign n19174 = n19009 & n19172 ;
  assign n19175 = ( n19009 & n19173 ) | ( n19009 & ~n19174 ) | ( n19173 & ~n19174 ) ;
  assign n19176 = n1023 | n1838 ;
  assign n19177 = ( n369 & ~n684 ) | ( n369 & n959 ) | ( ~n684 & n959 ) ;
  assign n19178 = n684 | n19177 ;
  assign n19179 = ( n3273 & ~n19176 ) | ( n3273 & n19178 ) | ( ~n19176 & n19178 ) ;
  assign n19180 = n19176 | n19179 ;
  assign n19181 = ( n2688 & n4829 ) | ( n2688 & ~n12119 ) | ( n4829 & ~n12119 ) ;
  assign n19182 = n12119 | n19181 ;
  assign n19183 = n124 | n159 ;
  assign n19184 = ( n1477 & n2721 ) | ( n1477 & ~n19183 ) | ( n2721 & ~n19183 ) ;
  assign n19185 = n19183 | n19184 ;
  assign n19186 = ( ~n19180 & n19182 ) | ( ~n19180 & n19185 ) | ( n19182 & n19185 ) ;
  assign n19187 = n19180 | n19186 ;
  assign n19188 = n3096 | n3943 ;
  assign n19189 = ( n6052 & n19187 ) | ( n6052 & ~n19188 ) | ( n19187 & ~n19188 ) ;
  assign n19190 = ~n19187 & n19189 ;
  assign n19191 = n607 & n16069 ;
  assign n19192 = n1250 & n16067 ;
  assign n19193 = n19191 | n19192 ;
  assign n19194 = n606 & ~n16065 ;
  assign n19195 = ( n606 & n19193 ) | ( n606 & ~n19194 ) | ( n19193 & ~n19194 ) ;
  assign n19196 = n1248 & n16281 ;
  assign n19197 = n19195 | n19196 ;
  assign n19198 = ( n19080 & ~n19190 ) | ( n19080 & n19197 ) | ( ~n19190 & n19197 ) ;
  assign n19199 = ( n19080 & n19190 ) | ( n19080 & n19197 ) | ( n19190 & n19197 ) ;
  assign n19200 = ( n19190 & n19198 ) | ( n19190 & ~n19199 ) | ( n19198 & ~n19199 ) ;
  assign n19201 = n3800 & ~n16433 ;
  assign n19202 = n3799 & n16059 ;
  assign n19203 = n3700 & n16063 ;
  assign n19204 = n3802 & ~n16061 ;
  assign n19205 = n19203 | n19204 ;
  assign n19206 = ( ~n19201 & n19202 ) | ( ~n19201 & n19205 ) | ( n19202 & n19205 ) ;
  assign n19207 = ( ~x29 & n19201 ) | ( ~x29 & n19206 ) | ( n19201 & n19206 ) ;
  assign n19208 = ( n19201 & n19206 ) | ( n19201 & ~n19207 ) | ( n19206 & ~n19207 ) ;
  assign n19209 = ( x29 & n19207 ) | ( x29 & ~n19208 ) | ( n19207 & ~n19208 ) ;
  assign n19210 = ( n19083 & ~n19200 ) | ( n19083 & n19209 ) | ( ~n19200 & n19209 ) ;
  assign n19211 = ( n19083 & n19200 ) | ( n19083 & n19209 ) | ( n19200 & n19209 ) ;
  assign n19212 = ( n19200 & n19210 ) | ( n19200 & ~n19211 ) | ( n19210 & ~n19211 ) ;
  assign n19213 = n4202 & n16553 ;
  assign n19214 = n4201 & n16053 ;
  assign n19215 = n4200 & ~n16057 ;
  assign n19216 = n4345 & ~n16055 ;
  assign n19217 = n19215 | n19216 ;
  assign n19218 = ( ~n19213 & n19214 ) | ( ~n19213 & n19217 ) | ( n19214 & n19217 ) ;
  assign n19219 = ( ~x26 & n19213 ) | ( ~x26 & n19218 ) | ( n19213 & n19218 ) ;
  assign n19220 = ( n19213 & n19218 ) | ( n19213 & ~n19219 ) | ( n19218 & ~n19219 ) ;
  assign n19221 = ( x26 & n19219 ) | ( x26 & ~n19220 ) | ( n19219 & ~n19220 ) ;
  assign n19222 = ( n19095 & ~n19212 ) | ( n19095 & n19221 ) | ( ~n19212 & n19221 ) ;
  assign n19223 = ( n19095 & n19212 ) | ( n19095 & n19221 ) | ( n19212 & n19221 ) ;
  assign n19224 = ( n19212 & n19222 ) | ( n19212 & ~n19223 ) | ( n19222 & ~n19223 ) ;
  assign n19225 = n4713 & ~n16801 ;
  assign n19226 = n4712 & ~n16047 ;
  assign n19227 = n4709 & ~n16051 ;
  assign n19228 = n4792 & ~n16049 ;
  assign n19229 = n19227 | n19228 ;
  assign n19230 = ( ~n19225 & n19226 ) | ( ~n19225 & n19229 ) | ( n19226 & n19229 ) ;
  assign n19231 = ( ~x23 & n19225 ) | ( ~x23 & n19230 ) | ( n19225 & n19230 ) ;
  assign n19232 = ( n19225 & n19230 ) | ( n19225 & ~n19231 ) | ( n19230 & ~n19231 ) ;
  assign n19233 = ( x23 & n19231 ) | ( x23 & ~n19232 ) | ( n19231 & ~n19232 ) ;
  assign n19234 = ( n19098 & ~n19224 ) | ( n19098 & n19233 ) | ( ~n19224 & n19233 ) ;
  assign n19235 = ( n19098 & n19224 ) | ( n19098 & n19233 ) | ( n19224 & n19233 ) ;
  assign n19236 = ( n19224 & n19234 ) | ( n19224 & ~n19235 ) | ( n19234 & ~n19235 ) ;
  assign n19237 = n4974 & n16969 ;
  assign n19238 = n5398 & n16041 ;
  assign n19239 = n4973 & ~n16045 ;
  assign n19240 = n4972 & ~n16043 ;
  assign n19241 = n19239 | n19240 ;
  assign n19242 = ( ~n19237 & n19238 ) | ( ~n19237 & n19241 ) | ( n19238 & n19241 ) ;
  assign n19243 = ( ~x20 & n19237 ) | ( ~x20 & n19242 ) | ( n19237 & n19242 ) ;
  assign n19244 = ( n19237 & n19242 ) | ( n19237 & ~n19243 ) | ( n19242 & ~n19243 ) ;
  assign n19245 = ( x20 & n19243 ) | ( x20 & ~n19244 ) | ( n19243 & ~n19244 ) ;
  assign n19246 = ( n19110 & ~n19236 ) | ( n19110 & n19245 ) | ( ~n19236 & n19245 ) ;
  assign n19247 = ( n19110 & n19236 ) | ( n19110 & n19245 ) | ( n19236 & n19245 ) ;
  assign n19248 = ( n19236 & n19246 ) | ( n19236 & ~n19247 ) | ( n19246 & ~n19247 ) ;
  assign n19249 = n5508 & ~n17313 ;
  assign n19250 = n5507 & n16035 ;
  assign n19251 = n5504 & n16039 ;
  assign n19252 = n5666 & ~n16037 ;
  assign n19253 = n19251 | n19252 ;
  assign n19254 = ( ~n19249 & n19250 ) | ( ~n19249 & n19253 ) | ( n19250 & n19253 ) ;
  assign n19255 = ( ~x17 & n19249 ) | ( ~x17 & n19254 ) | ( n19249 & n19254 ) ;
  assign n19256 = ( n19249 & n19254 ) | ( n19249 & ~n19255 ) | ( n19254 & ~n19255 ) ;
  assign n19257 = ( x17 & n19255 ) | ( x17 & ~n19256 ) | ( n19255 & ~n19256 ) ;
  assign n19258 = ( n19113 & ~n19248 ) | ( n19113 & n19257 ) | ( ~n19248 & n19257 ) ;
  assign n19259 = ( n19113 & n19248 ) | ( n19113 & n19257 ) | ( n19248 & n19257 ) ;
  assign n19260 = ( n19248 & n19258 ) | ( n19248 & ~n19259 ) | ( n19258 & ~n19259 ) ;
  assign n19261 = n5966 & ~n17528 ;
  assign n19262 = n6464 & ~n16029 ;
  assign n19263 = n5970 & ~n16033 ;
  assign n19264 = n5969 & n16031 ;
  assign n19265 = n19263 | n19264 ;
  assign n19266 = ( ~n19261 & n19262 ) | ( ~n19261 & n19265 ) | ( n19262 & n19265 ) ;
  assign n19267 = ( ~x14 & n19261 ) | ( ~x14 & n19266 ) | ( n19261 & n19266 ) ;
  assign n19268 = ( n19261 & n19266 ) | ( n19261 & ~n19267 ) | ( n19266 & ~n19267 ) ;
  assign n19269 = ( x14 & n19267 ) | ( x14 & ~n19268 ) | ( n19267 & ~n19268 ) ;
  assign n19270 = ( n19125 & ~n19260 ) | ( n19125 & n19269 ) | ( ~n19260 & n19269 ) ;
  assign n19271 = ( n19125 & n19260 ) | ( n19125 & n19269 ) | ( n19260 & n19269 ) ;
  assign n19272 = ( n19260 & n19270 ) | ( n19260 & ~n19271 ) | ( n19270 & ~n19271 ) ;
  assign n19273 = n6584 & n17968 ;
  assign n19274 = n7022 & n16023 ;
  assign n19275 = n6588 & ~n16027 ;
  assign n19276 = n6587 & ~n16025 ;
  assign n19277 = n19275 | n19276 ;
  assign n19278 = ( ~n19273 & n19274 ) | ( ~n19273 & n19277 ) | ( n19274 & n19277 ) ;
  assign n19279 = ( ~x11 & n19273 ) | ( ~x11 & n19278 ) | ( n19273 & n19278 ) ;
  assign n19280 = ( n19273 & n19278 ) | ( n19273 & ~n19279 ) | ( n19278 & ~n19279 ) ;
  assign n19281 = ( x11 & n19279 ) | ( x11 & ~n19280 ) | ( n19279 & ~n19280 ) ;
  assign n19282 = ( n19128 & ~n19272 ) | ( n19128 & n19281 ) | ( ~n19272 & n19281 ) ;
  assign n19283 = ( n19128 & n19272 ) | ( n19128 & n19281 ) | ( n19272 & n19281 ) ;
  assign n19284 = ( n19272 & n19282 ) | ( n19272 & ~n19283 ) | ( n19282 & ~n19283 ) ;
  assign n19285 = n7296 & ~n18267 ;
  assign n19286 = n7879 & ~n16017 ;
  assign n19287 = n7300 & n16021 ;
  assign n19288 = n7299 & n16019 ;
  assign n19289 = n19287 | n19288 ;
  assign n19290 = ( ~n19285 & n19286 ) | ( ~n19285 & n19289 ) | ( n19286 & n19289 ) ;
  assign n19291 = ( ~x8 & n19285 ) | ( ~x8 & n19290 ) | ( n19285 & n19290 ) ;
  assign n19292 = ( n19285 & n19290 ) | ( n19285 & ~n19291 ) | ( n19290 & ~n19291 ) ;
  assign n19293 = ( x8 & n19291 ) | ( x8 & ~n19292 ) | ( n19291 & ~n19292 ) ;
  assign n19294 = ( n19140 & ~n19284 ) | ( n19140 & n19293 ) | ( ~n19284 & n19293 ) ;
  assign n19295 = ( n19140 & n19284 ) | ( n19140 & n19293 ) | ( n19284 & n19293 ) ;
  assign n19296 = ( n19284 & n19294 ) | ( n19284 & ~n19295 ) | ( n19294 & ~n19295 ) ;
  assign n19297 = n8230 & ~n16144 ;
  assign n19298 = n8229 & n16138 ;
  assign n19299 = n8226 & n16015 ;
  assign n19300 = n8225 & ~n16013 ;
  assign n19301 = n19299 | n19300 ;
  assign n19302 = ( ~n19297 & n19298 ) | ( ~n19297 & n19301 ) | ( n19298 & n19301 ) ;
  assign n19303 = ( ~x5 & n19297 ) | ( ~x5 & n19302 ) | ( n19297 & n19302 ) ;
  assign n19304 = ( n19297 & n19302 ) | ( n19297 & ~n19303 ) | ( n19302 & ~n19303 ) ;
  assign n19305 = ( x5 & n19303 ) | ( x5 & ~n19304 ) | ( n19303 & ~n19304 ) ;
  assign n19306 = ( n19143 & ~n19296 ) | ( n19143 & n19305 ) | ( ~n19296 & n19305 ) ;
  assign n19307 = ( n19143 & n19296 ) | ( n19143 & n19305 ) | ( n19296 & n19305 ) ;
  assign n19308 = ( n19296 & n19306 ) | ( n19296 & ~n19307 ) | ( n19306 & ~n19307 ) ;
  assign n19309 = n19148 | n19157 ;
  assign n19310 = ( n19157 & n19158 ) | ( n19157 & ~n19309 ) | ( n19158 & ~n19309 ) ;
  assign n19311 = ( ~n19157 & n19158 ) | ( ~n19157 & n19309 ) | ( n19158 & n19309 ) ;
  assign n19312 = ( ~n19158 & n19310 ) | ( ~n19158 & n19311 ) | ( n19310 & n19311 ) ;
  assign n19313 = n36 & ~n19312 ;
  assign n19314 = n8967 & n18993 ;
  assign n19315 = ( x0 & n8966 ) | ( x0 & ~n19157 ) | ( n8966 & ~n19157 ) ;
  assign n19316 = ( n8966 & n19314 ) | ( n8966 & ~n19315 ) | ( n19314 & ~n19315 ) ;
  assign n19317 = n35 & n19309 ;
  assign n19318 = ( n35 & n19316 ) | ( n35 & ~n19317 ) | ( n19316 & ~n19317 ) ;
  assign n19319 = ( ~x2 & n19313 ) | ( ~x2 & n19318 ) | ( n19313 & n19318 ) ;
  assign n19320 = ( n19313 & n19318 ) | ( n19313 & ~n19319 ) | ( n19318 & ~n19319 ) ;
  assign n19321 = ( x2 & n19319 ) | ( x2 & ~n19320 ) | ( n19319 & ~n19320 ) ;
  assign n19322 = ( n19170 & ~n19308 ) | ( n19170 & n19321 ) | ( ~n19308 & n19321 ) ;
  assign n19323 = ( n19170 & n19308 ) | ( n19170 & n19321 ) | ( n19308 & n19321 ) ;
  assign n19324 = ( n19308 & n19322 ) | ( n19308 & ~n19323 ) | ( n19322 & ~n19323 ) ;
  assign n19325 = n19173 & ~n19324 ;
  assign n19326 = ~n19173 & n19324 ;
  assign n19327 = n19325 | n19326 ;
  assign n19328 = n2952 & ~n4042 ;
  assign n19329 = n2182 | n2390 ;
  assign n19330 = n5725 | n10965 ;
  assign n19331 = n2628 | n2966 ;
  assign n19332 = n132 | n544 ;
  assign n19333 = ( n142 & n890 ) | ( n142 & ~n19332 ) | ( n890 & ~n19332 ) ;
  assign n19334 = n19332 | n19333 ;
  assign n19335 = ( n916 & n1646 ) | ( n916 & ~n19334 ) | ( n1646 & ~n19334 ) ;
  assign n19336 = n19334 | n19335 ;
  assign n19337 = ( ~n19330 & n19331 ) | ( ~n19330 & n19336 ) | ( n19331 & n19336 ) ;
  assign n19338 = n19330 | n19337 ;
  assign n19339 = n233 | n1225 ;
  assign n19340 = ( n1116 & n1442 ) | ( n1116 & ~n19339 ) | ( n1442 & ~n19339 ) ;
  assign n19341 = n19339 | n19340 ;
  assign n19342 = ( ~n19329 & n19338 ) | ( ~n19329 & n19341 ) | ( n19338 & n19341 ) ;
  assign n19343 = n19329 | n19342 ;
  assign n19344 = n2975 | n5156 ;
  assign n19345 = n866 | n2636 ;
  assign n19346 = n679 | n1423 ;
  assign n19347 = ( n1253 & n1510 ) | ( n1253 & ~n19346 ) | ( n1510 & ~n19346 ) ;
  assign n19348 = n19346 | n19347 ;
  assign n19349 = ( ~n19344 & n19345 ) | ( ~n19344 & n19348 ) | ( n19345 & n19348 ) ;
  assign n19350 = n19344 | n19349 ;
  assign n19351 = ( ~n4042 & n19343 ) | ( ~n4042 & n19350 ) | ( n19343 & n19350 ) ;
  assign n19352 = ( n4581 & n19328 ) | ( n4581 & ~n19351 ) | ( n19328 & ~n19351 ) ;
  assign n19353 = ~n4581 & n19352 ;
  assign n19354 = n607 & n16067 ;
  assign n19355 = n1250 & n16065 ;
  assign n19356 = n19354 | n19355 ;
  assign n19357 = n606 & ~n16063 ;
  assign n19358 = ( n606 & n19356 ) | ( n606 & ~n19357 ) | ( n19356 & ~n19357 ) ;
  assign n19359 = n1248 & n16315 ;
  assign n19360 = n19358 | n19359 ;
  assign n19361 = ( n19198 & ~n19353 ) | ( n19198 & n19360 ) | ( ~n19353 & n19360 ) ;
  assign n19362 = ( n19198 & n19353 ) | ( n19198 & n19360 ) | ( n19353 & n19360 ) ;
  assign n19363 = ( n19353 & n19361 ) | ( n19353 & ~n19362 ) | ( n19361 & ~n19362 ) ;
  assign n19364 = n3800 & ~n16484 ;
  assign n19365 = n3799 & ~n16057 ;
  assign n19366 = n3700 & ~n16061 ;
  assign n19367 = n3802 & n16059 ;
  assign n19368 = n19366 | n19367 ;
  assign n19369 = ( ~n19364 & n19365 ) | ( ~n19364 & n19368 ) | ( n19365 & n19368 ) ;
  assign n19370 = ( ~x29 & n19364 ) | ( ~x29 & n19369 ) | ( n19364 & n19369 ) ;
  assign n19371 = ( n19364 & n19369 ) | ( n19364 & ~n19370 ) | ( n19369 & ~n19370 ) ;
  assign n19372 = ( x29 & n19370 ) | ( x29 & ~n19371 ) | ( n19370 & ~n19371 ) ;
  assign n19373 = ( n19210 & ~n19363 ) | ( n19210 & n19372 ) | ( ~n19363 & n19372 ) ;
  assign n19374 = ( n19210 & n19363 ) | ( n19210 & n19372 ) | ( n19363 & n19372 ) ;
  assign n19375 = ( n19363 & n19373 ) | ( n19363 & ~n19374 ) | ( n19373 & ~n19374 ) ;
  assign n19376 = n4202 & n16611 ;
  assign n19377 = n4201 & ~n16051 ;
  assign n19378 = n4200 & ~n16055 ;
  assign n19379 = n4345 & n16053 ;
  assign n19380 = n19378 | n19379 ;
  assign n19381 = ( ~n19376 & n19377 ) | ( ~n19376 & n19380 ) | ( n19377 & n19380 ) ;
  assign n19382 = ( ~x26 & n19376 ) | ( ~x26 & n19381 ) | ( n19376 & n19381 ) ;
  assign n19383 = ( n19376 & n19381 ) | ( n19376 & ~n19382 ) | ( n19381 & ~n19382 ) ;
  assign n19384 = ( x26 & n19382 ) | ( x26 & ~n19383 ) | ( n19382 & ~n19383 ) ;
  assign n19385 = ( n19222 & ~n19375 ) | ( n19222 & n19384 ) | ( ~n19375 & n19384 ) ;
  assign n19386 = ( n19222 & n19375 ) | ( n19222 & n19384 ) | ( n19375 & n19384 ) ;
  assign n19387 = ( n19375 & n19385 ) | ( n19375 & ~n19386 ) | ( n19385 & ~n19386 ) ;
  assign n19388 = n4713 & ~n16876 ;
  assign n19389 = n4712 & ~n16045 ;
  assign n19390 = n4709 & ~n16049 ;
  assign n19391 = n4792 & ~n16047 ;
  assign n19392 = n19390 | n19391 ;
  assign n19393 = ( ~n19388 & n19389 ) | ( ~n19388 & n19392 ) | ( n19389 & n19392 ) ;
  assign n19394 = ( ~x23 & n19388 ) | ( ~x23 & n19393 ) | ( n19388 & n19393 ) ;
  assign n19395 = ( n19388 & n19393 ) | ( n19388 & ~n19394 ) | ( n19393 & ~n19394 ) ;
  assign n19396 = ( x23 & n19394 ) | ( x23 & ~n19395 ) | ( n19394 & ~n19395 ) ;
  assign n19397 = ( n19234 & ~n19387 ) | ( n19234 & n19396 ) | ( ~n19387 & n19396 ) ;
  assign n19398 = ( n19234 & n19387 ) | ( n19234 & n19396 ) | ( n19387 & n19396 ) ;
  assign n19399 = ( n19387 & n19397 ) | ( n19387 & ~n19398 ) | ( n19397 & ~n19398 ) ;
  assign n19400 = n4974 & ~n17051 ;
  assign n19401 = n5398 & n16039 ;
  assign n19402 = n4973 & ~n16043 ;
  assign n19403 = n4972 & n16041 ;
  assign n19404 = n19402 | n19403 ;
  assign n19405 = ( ~n19400 & n19401 ) | ( ~n19400 & n19404 ) | ( n19401 & n19404 ) ;
  assign n19406 = ( ~x20 & n19400 ) | ( ~x20 & n19405 ) | ( n19400 & n19405 ) ;
  assign n19407 = ( n19400 & n19405 ) | ( n19400 & ~n19406 ) | ( n19405 & ~n19406 ) ;
  assign n19408 = ( x20 & n19406 ) | ( x20 & ~n19407 ) | ( n19406 & ~n19407 ) ;
  assign n19409 = ( n19246 & ~n19399 ) | ( n19246 & n19408 ) | ( ~n19399 & n19408 ) ;
  assign n19410 = ( n19246 & n19399 ) | ( n19246 & n19408 ) | ( n19399 & n19408 ) ;
  assign n19411 = ( n19399 & n19409 ) | ( n19399 & ~n19410 ) | ( n19409 & ~n19410 ) ;
  assign n19412 = n5508 & ~n17412 ;
  assign n19413 = n5507 & ~n16033 ;
  assign n19414 = n5504 & ~n16037 ;
  assign n19415 = n5666 & n16035 ;
  assign n19416 = n19414 | n19415 ;
  assign n19417 = ( ~n19412 & n19413 ) | ( ~n19412 & n19416 ) | ( n19413 & n19416 ) ;
  assign n19418 = ( ~x17 & n19412 ) | ( ~x17 & n19417 ) | ( n19412 & n19417 ) ;
  assign n19419 = ( n19412 & n19417 ) | ( n19412 & ~n19418 ) | ( n19417 & ~n19418 ) ;
  assign n19420 = ( x17 & n19418 ) | ( x17 & ~n19419 ) | ( n19418 & ~n19419 ) ;
  assign n19421 = ( n19258 & ~n19411 ) | ( n19258 & n19420 ) | ( ~n19411 & n19420 ) ;
  assign n19422 = ( n19258 & n19411 ) | ( n19258 & n19420 ) | ( n19411 & n19420 ) ;
  assign n19423 = ( n19411 & n19421 ) | ( n19411 & ~n19422 ) | ( n19421 & ~n19422 ) ;
  assign n19424 = n5966 & n17634 ;
  assign n19425 = n6464 & ~n16027 ;
  assign n19426 = n5970 & n16031 ;
  assign n19427 = n5969 & ~n16029 ;
  assign n19428 = n19426 | n19427 ;
  assign n19429 = ( ~n19424 & n19425 ) | ( ~n19424 & n19428 ) | ( n19425 & n19428 ) ;
  assign n19430 = ( ~x14 & n19424 ) | ( ~x14 & n19429 ) | ( n19424 & n19429 ) ;
  assign n19431 = ( n19424 & n19429 ) | ( n19424 & ~n19430 ) | ( n19429 & ~n19430 ) ;
  assign n19432 = ( x14 & n19430 ) | ( x14 & ~n19431 ) | ( n19430 & ~n19431 ) ;
  assign n19433 = ( n19270 & ~n19423 ) | ( n19270 & n19432 ) | ( ~n19423 & n19432 ) ;
  assign n19434 = ( n19270 & n19423 ) | ( n19270 & n19432 ) | ( n19423 & n19432 ) ;
  assign n19435 = ( n19423 & n19433 ) | ( n19423 & ~n19434 ) | ( n19433 & ~n19434 ) ;
  assign n19436 = n6584 & ~n18091 ;
  assign n19437 = n7022 & n16021 ;
  assign n19438 = n6588 & ~n16025 ;
  assign n19439 = n6587 & n16023 ;
  assign n19440 = n19438 | n19439 ;
  assign n19441 = ( ~n19436 & n19437 ) | ( ~n19436 & n19440 ) | ( n19437 & n19440 ) ;
  assign n19442 = ( ~x11 & n19436 ) | ( ~x11 & n19441 ) | ( n19436 & n19441 ) ;
  assign n19443 = ( n19436 & n19441 ) | ( n19436 & ~n19442 ) | ( n19441 & ~n19442 ) ;
  assign n19444 = ( x11 & n19442 ) | ( x11 & ~n19443 ) | ( n19442 & ~n19443 ) ;
  assign n19445 = ( n19282 & ~n19435 ) | ( n19282 & n19444 ) | ( ~n19435 & n19444 ) ;
  assign n19446 = ( n19282 & n19435 ) | ( n19282 & n19444 ) | ( n19435 & n19444 ) ;
  assign n19447 = ( n19435 & n19445 ) | ( n19435 & ~n19446 ) | ( n19445 & ~n19446 ) ;
  assign n19448 = n7296 & ~n18416 ;
  assign n19449 = n7879 & n16015 ;
  assign n19450 = n7300 & n16019 ;
  assign n19451 = n7299 & ~n16017 ;
  assign n19452 = n19450 | n19451 ;
  assign n19453 = ( ~n19448 & n19449 ) | ( ~n19448 & n19452 ) | ( n19449 & n19452 ) ;
  assign n19454 = ( ~x8 & n19448 ) | ( ~x8 & n19453 ) | ( n19448 & n19453 ) ;
  assign n19455 = ( n19448 & n19453 ) | ( n19448 & ~n19454 ) | ( n19453 & ~n19454 ) ;
  assign n19456 = ( x8 & n19454 ) | ( x8 & ~n19455 ) | ( n19454 & ~n19455 ) ;
  assign n19457 = ( n19294 & ~n19447 ) | ( n19294 & n19456 ) | ( ~n19447 & n19456 ) ;
  assign n19458 = ( n19294 & n19447 ) | ( n19294 & n19456 ) | ( n19447 & n19456 ) ;
  assign n19459 = ( n19447 & n19457 ) | ( n19447 & ~n19458 ) | ( n19457 & ~n19458 ) ;
  assign n19460 = n8230 & n18996 ;
  assign n19461 = n8229 & n18993 ;
  assign n19462 = n8226 & ~n16013 ;
  assign n19463 = n8225 & n16138 ;
  assign n19464 = n19462 | n19463 ;
  assign n19465 = ( ~n19460 & n19461 ) | ( ~n19460 & n19464 ) | ( n19461 & n19464 ) ;
  assign n19466 = ( ~x5 & n19460 ) | ( ~x5 & n19465 ) | ( n19460 & n19465 ) ;
  assign n19467 = ( n19460 & n19465 ) | ( n19460 & ~n19466 ) | ( n19465 & ~n19466 ) ;
  assign n19468 = ( x5 & n19466 ) | ( x5 & ~n19467 ) | ( n19466 & ~n19467 ) ;
  assign n19469 = ( n19306 & ~n19459 ) | ( n19306 & n19468 ) | ( ~n19459 & n19468 ) ;
  assign n19470 = ( n19306 & n19459 ) | ( n19306 & n19468 ) | ( n19459 & n19468 ) ;
  assign n19471 = ( n19459 & n19469 ) | ( n19459 & ~n19470 ) | ( n19469 & ~n19470 ) ;
  assign n19472 = n19309 & ~n19310 ;
  assign n19473 = n36 & ~n19472 ;
  assign n19474 = n8967 & n19157 ;
  assign n19475 = ( x0 & n8966 ) | ( x0 & n19309 ) | ( n8966 & n19309 ) ;
  assign n19476 = ( n8966 & n19474 ) | ( n8966 & ~n19475 ) | ( n19474 & ~n19475 ) ;
  assign n19477 = ( ~x2 & n19473 ) | ( ~x2 & n19476 ) | ( n19473 & n19476 ) ;
  assign n19478 = ( n19473 & n19476 ) | ( n19473 & ~n19477 ) | ( n19476 & ~n19477 ) ;
  assign n19479 = ( x2 & n19477 ) | ( x2 & ~n19478 ) | ( n19477 & ~n19478 ) ;
  assign n19480 = ( n19322 & ~n19471 ) | ( n19322 & n19479 ) | ( ~n19471 & n19479 ) ;
  assign n19481 = ( n19322 & n19471 ) | ( n19322 & n19479 ) | ( n19471 & n19479 ) ;
  assign n19482 = ( n19471 & n19480 ) | ( n19471 & ~n19481 ) | ( n19480 & ~n19481 ) ;
  assign n19483 = n19325 & ~n19482 ;
  assign n19484 = n19325 & n19482 ;
  assign n19485 = ( n19482 & n19483 ) | ( n19482 & ~n19484 ) | ( n19483 & ~n19484 ) ;
  assign n19486 = n1891 | n5061 ;
  assign n19487 = n132 | n254 ;
  assign n19488 = ( n1407 & ~n19486 ) | ( n1407 & n19487 ) | ( ~n19486 & n19487 ) ;
  assign n19489 = n19486 | n19488 ;
  assign n19490 = n3840 | n3918 ;
  assign n19491 = n586 | n1048 ;
  assign n19492 = ( n50 & n97 ) | ( n50 & n810 ) | ( n97 & n810 ) ;
  assign n19493 = ( n171 & n873 ) | ( n171 & ~n19492 ) | ( n873 & ~n19492 ) ;
  assign n19494 = n19492 | n19493 ;
  assign n19495 = ( n450 & n1377 ) | ( n450 & ~n19494 ) | ( n1377 & ~n19494 ) ;
  assign n19496 = n19494 | n19495 ;
  assign n19497 = ( n1556 & ~n19491 ) | ( n1556 & n19496 ) | ( ~n19491 & n19496 ) ;
  assign n19498 = n19491 | n19497 ;
  assign n19499 = ( ~n19489 & n19490 ) | ( ~n19489 & n19498 ) | ( n19490 & n19498 ) ;
  assign n19500 = n19489 | n19499 ;
  assign n19501 = ~n5220 & n11913 ;
  assign n19502 = ~n19500 & n19501 ;
  assign n19503 = n607 & n16065 ;
  assign n19504 = n1250 & n16063 ;
  assign n19505 = n19503 | n19504 ;
  assign n19506 = n606 & ~n16061 ;
  assign n19507 = n19505 | n19506 ;
  assign n19508 = n1248 & ~n16354 ;
  assign n19509 = n19507 | n19508 ;
  assign n19510 = ( n19361 & ~n19502 ) | ( n19361 & n19509 ) | ( ~n19502 & n19509 ) ;
  assign n19511 = ( n19361 & n19502 ) | ( n19361 & n19509 ) | ( n19502 & n19509 ) ;
  assign n19512 = ( n19502 & n19510 ) | ( n19502 & ~n19511 ) | ( n19510 & ~n19511 ) ;
  assign n19513 = n3800 & n16541 ;
  assign n19514 = n3799 & ~n16055 ;
  assign n19515 = n3700 & n16059 ;
  assign n19516 = n3802 & ~n16057 ;
  assign n19517 = n19515 | n19516 ;
  assign n19518 = ( ~n19513 & n19514 ) | ( ~n19513 & n19517 ) | ( n19514 & n19517 ) ;
  assign n19519 = ( ~x29 & n19513 ) | ( ~x29 & n19518 ) | ( n19513 & n19518 ) ;
  assign n19520 = ( n19513 & n19518 ) | ( n19513 & ~n19519 ) | ( n19518 & ~n19519 ) ;
  assign n19521 = ( x29 & n19519 ) | ( x29 & ~n19520 ) | ( n19519 & ~n19520 ) ;
  assign n19522 = ( n19373 & ~n19512 ) | ( n19373 & n19521 ) | ( ~n19512 & n19521 ) ;
  assign n19523 = ( n19373 & n19512 ) | ( n19373 & n19521 ) | ( n19512 & n19521 ) ;
  assign n19524 = ( n19512 & n19522 ) | ( n19512 & ~n19523 ) | ( n19522 & ~n19523 ) ;
  assign n19525 = n4202 & ~n16674 ;
  assign n19526 = n4201 & ~n16049 ;
  assign n19527 = n4200 & n16053 ;
  assign n19528 = n4345 & ~n16051 ;
  assign n19529 = n19527 | n19528 ;
  assign n19530 = ( ~n19525 & n19526 ) | ( ~n19525 & n19529 ) | ( n19526 & n19529 ) ;
  assign n19531 = ( ~x26 & n19525 ) | ( ~x26 & n19530 ) | ( n19525 & n19530 ) ;
  assign n19532 = ( n19525 & n19530 ) | ( n19525 & ~n19531 ) | ( n19530 & ~n19531 ) ;
  assign n19533 = ( x26 & n19531 ) | ( x26 & ~n19532 ) | ( n19531 & ~n19532 ) ;
  assign n19534 = ( n19385 & ~n19524 ) | ( n19385 & n19533 ) | ( ~n19524 & n19533 ) ;
  assign n19535 = ( n19385 & n19524 ) | ( n19385 & n19533 ) | ( n19524 & n19533 ) ;
  assign n19536 = ( n19524 & n19534 ) | ( n19524 & ~n19535 ) | ( n19534 & ~n19535 ) ;
  assign n19537 = n4713 & ~n16957 ;
  assign n19538 = n4712 & ~n16043 ;
  assign n19539 = n4709 & ~n16047 ;
  assign n19540 = n4792 & ~n16045 ;
  assign n19541 = n19539 | n19540 ;
  assign n19542 = ( ~n19537 & n19538 ) | ( ~n19537 & n19541 ) | ( n19538 & n19541 ) ;
  assign n19543 = ( ~x23 & n19537 ) | ( ~x23 & n19542 ) | ( n19537 & n19542 ) ;
  assign n19544 = ( n19537 & n19542 ) | ( n19537 & ~n19543 ) | ( n19542 & ~n19543 ) ;
  assign n19545 = ( x23 & n19543 ) | ( x23 & ~n19544 ) | ( n19543 & ~n19544 ) ;
  assign n19546 = ( n19397 & ~n19536 ) | ( n19397 & n19545 ) | ( ~n19536 & n19545 ) ;
  assign n19547 = ( n19397 & n19536 ) | ( n19397 & n19545 ) | ( n19536 & n19545 ) ;
  assign n19548 = ( n19536 & n19546 ) | ( n19536 & ~n19547 ) | ( n19546 & ~n19547 ) ;
  assign n19549 = n4974 & ~n17138 ;
  assign n19550 = n5398 & ~n16037 ;
  assign n19551 = n4973 & n16041 ;
  assign n19552 = n4972 & n16039 ;
  assign n19553 = n19551 | n19552 ;
  assign n19554 = ( ~n19549 & n19550 ) | ( ~n19549 & n19553 ) | ( n19550 & n19553 ) ;
  assign n19555 = ( ~x20 & n19549 ) | ( ~x20 & n19554 ) | ( n19549 & n19554 ) ;
  assign n19556 = ( n19549 & n19554 ) | ( n19549 & ~n19555 ) | ( n19554 & ~n19555 ) ;
  assign n19557 = ( x20 & n19555 ) | ( x20 & ~n19556 ) | ( n19555 & ~n19556 ) ;
  assign n19558 = ( n19409 & ~n19548 ) | ( n19409 & n19557 ) | ( ~n19548 & n19557 ) ;
  assign n19559 = ( n19409 & n19548 ) | ( n19409 & n19557 ) | ( n19548 & n19557 ) ;
  assign n19560 = ( n19548 & n19558 ) | ( n19548 & ~n19559 ) | ( n19558 & ~n19559 ) ;
  assign n19561 = n5508 & ~n17516 ;
  assign n19562 = n5507 & n16031 ;
  assign n19563 = n5504 & n16035 ;
  assign n19564 = n5666 & ~n16033 ;
  assign n19565 = n19563 | n19564 ;
  assign n19566 = ( ~n19561 & n19562 ) | ( ~n19561 & n19565 ) | ( n19562 & n19565 ) ;
  assign n19567 = ( ~x17 & n19561 ) | ( ~x17 & n19566 ) | ( n19561 & n19566 ) ;
  assign n19568 = ( n19561 & n19566 ) | ( n19561 & ~n19567 ) | ( n19566 & ~n19567 ) ;
  assign n19569 = ( x17 & n19567 ) | ( x17 & ~n19568 ) | ( n19567 & ~n19568 ) ;
  assign n19570 = ( n19421 & ~n19560 ) | ( n19421 & n19569 ) | ( ~n19560 & n19569 ) ;
  assign n19571 = ( n19421 & n19560 ) | ( n19421 & n19569 ) | ( n19560 & n19569 ) ;
  assign n19572 = ( n19560 & n19570 ) | ( n19560 & ~n19571 ) | ( n19570 & ~n19571 ) ;
  assign n19573 = n5966 & ~n17746 ;
  assign n19574 = n6464 & ~n16025 ;
  assign n19575 = n5970 & ~n16029 ;
  assign n19576 = n5969 & ~n16027 ;
  assign n19577 = n19575 | n19576 ;
  assign n19578 = ( ~n19573 & n19574 ) | ( ~n19573 & n19577 ) | ( n19574 & n19577 ) ;
  assign n19579 = ( ~x14 & n19573 ) | ( ~x14 & n19578 ) | ( n19573 & n19578 ) ;
  assign n19580 = ( n19573 & n19578 ) | ( n19573 & ~n19579 ) | ( n19578 & ~n19579 ) ;
  assign n19581 = ( x14 & n19579 ) | ( x14 & ~n19580 ) | ( n19579 & ~n19580 ) ;
  assign n19582 = ( n19433 & ~n19572 ) | ( n19433 & n19581 ) | ( ~n19572 & n19581 ) ;
  assign n19583 = ( n19433 & n19572 ) | ( n19433 & n19581 ) | ( n19572 & n19581 ) ;
  assign n19584 = ( n19572 & n19582 ) | ( n19572 & ~n19583 ) | ( n19582 & ~n19583 ) ;
  assign n19585 = n6584 & n18103 ;
  assign n19586 = n7022 & n16019 ;
  assign n19587 = n6588 & n16023 ;
  assign n19588 = n6587 & n16021 ;
  assign n19589 = n19587 | n19588 ;
  assign n19590 = ( ~n19585 & n19586 ) | ( ~n19585 & n19589 ) | ( n19586 & n19589 ) ;
  assign n19591 = ( ~x11 & n19585 ) | ( ~x11 & n19590 ) | ( n19585 & n19590 ) ;
  assign n19592 = ( n19585 & n19590 ) | ( n19585 & ~n19591 ) | ( n19590 & ~n19591 ) ;
  assign n19593 = ( x11 & n19591 ) | ( x11 & ~n19592 ) | ( n19591 & ~n19592 ) ;
  assign n19594 = ( n19445 & ~n19584 ) | ( n19445 & n19593 ) | ( ~n19584 & n19593 ) ;
  assign n19595 = ( n19445 & n19584 ) | ( n19445 & n19593 ) | ( n19584 & n19593 ) ;
  assign n19596 = ( n19584 & n19594 ) | ( n19584 & ~n19595 ) | ( n19594 & ~n19595 ) ;
  assign n19597 = n7296 & ~n18694 ;
  assign n19598 = n7879 & ~n16013 ;
  assign n19599 = n7300 & ~n16017 ;
  assign n19600 = n7299 & n16015 ;
  assign n19601 = n19599 | n19600 ;
  assign n19602 = ( ~n19597 & n19598 ) | ( ~n19597 & n19601 ) | ( n19598 & n19601 ) ;
  assign n19603 = ( ~x8 & n19597 ) | ( ~x8 & n19602 ) | ( n19597 & n19602 ) ;
  assign n19604 = ( n19597 & n19602 ) | ( n19597 & ~n19603 ) | ( n19602 & ~n19603 ) ;
  assign n19605 = ( x8 & n19603 ) | ( x8 & ~n19604 ) | ( n19603 & ~n19604 ) ;
  assign n19606 = ( n19457 & ~n19596 ) | ( n19457 & n19605 ) | ( ~n19596 & n19605 ) ;
  assign n19607 = ( n19457 & n19596 ) | ( n19457 & n19605 ) | ( n19596 & n19605 ) ;
  assign n19608 = ( n19596 & n19606 ) | ( n19596 & ~n19607 ) | ( n19606 & ~n19607 ) ;
  assign n19609 = n8230 & n19160 ;
  assign n19610 = n8229 & n19157 ;
  assign n19611 = n8226 & n16138 ;
  assign n19612 = n8225 & n18993 ;
  assign n19613 = n19611 | n19612 ;
  assign n19614 = ( ~n19609 & n19610 ) | ( ~n19609 & n19613 ) | ( n19610 & n19613 ) ;
  assign n19615 = ( ~x5 & n19609 ) | ( ~x5 & n19614 ) | ( n19609 & n19614 ) ;
  assign n19616 = ( n19609 & n19614 ) | ( n19609 & ~n19615 ) | ( n19614 & ~n19615 ) ;
  assign n19617 = ( x5 & n19615 ) | ( x5 & ~n19616 ) | ( n19615 & ~n19616 ) ;
  assign n19618 = ( n19469 & ~n19608 ) | ( n19469 & n19617 ) | ( ~n19608 & n19617 ) ;
  assign n19619 = ( n19469 & n19608 ) | ( n19469 & n19617 ) | ( n19608 & n19617 ) ;
  assign n19620 = ( n19608 & n19618 ) | ( n19608 & ~n19619 ) | ( n19618 & ~n19619 ) ;
  assign n19621 = n8967 & ~n19309 ;
  assign n19622 = x2 & ~n19621 ;
  assign n19623 = ( n19480 & ~n19620 ) | ( n19480 & n19622 ) | ( ~n19620 & n19622 ) ;
  assign n19624 = ( n19480 & n19620 ) | ( n19480 & n19622 ) | ( n19620 & n19622 ) ;
  assign n19625 = ( n19620 & n19623 ) | ( n19620 & ~n19624 ) | ( n19623 & ~n19624 ) ;
  assign n19626 = n19483 & ~n19625 ;
  assign n19627 = ~n19483 & n19625 ;
  assign n19628 = n19626 | n19627 ;
  assign n19629 = n3255 | n5012 ;
  assign n19630 = n837 | n1009 ;
  assign n19631 = ( n2325 & n19178 ) | ( n2325 & ~n19630 ) | ( n19178 & ~n19630 ) ;
  assign n19632 = n19630 | n19631 ;
  assign n19633 = n1132 | n2661 ;
  assign n19634 = n541 | n3445 ;
  assign n19635 = ( n4993 & ~n19633 ) | ( n4993 & n19634 ) | ( ~n19633 & n19634 ) ;
  assign n19636 = n19633 | n19635 ;
  assign n19637 = n11055 | n19636 ;
  assign n19638 = n1523 | n1679 ;
  assign n19639 = n133 | n1253 ;
  assign n19640 = n218 & ~n679 ;
  assign n19641 = ( n66 & n84 ) | ( n66 & n136 ) | ( n84 & n136 ) ;
  assign n19642 = ( n123 & n697 ) | ( n123 & ~n19641 ) | ( n697 & ~n19641 ) ;
  assign n19643 = n19641 | n19642 ;
  assign n19644 = ( n753 & n19640 ) | ( n753 & n19643 ) | ( n19640 & n19643 ) ;
  assign n19645 = n19640 & ~n19644 ;
  assign n19646 = ( n19638 & ~n19639 ) | ( n19638 & n19645 ) | ( ~n19639 & n19645 ) ;
  assign n19647 = ~n19638 & n19646 ;
  assign n19648 = ( n19632 & ~n19637 ) | ( n19632 & n19647 ) | ( ~n19637 & n19647 ) ;
  assign n19649 = ~n19632 & n19648 ;
  assign n19650 = ( ~n11370 & n19629 ) | ( ~n11370 & n19649 ) | ( n19629 & n19649 ) ;
  assign n19651 = ~n19629 & n19650 ;
  assign n19652 = n607 & n16063 ;
  assign n19653 = n1250 & ~n16061 ;
  assign n19654 = n19652 | n19653 ;
  assign n19655 = n606 & ~n16059 ;
  assign n19656 = ( n606 & n19654 ) | ( n606 & ~n19655 ) | ( n19654 & ~n19655 ) ;
  assign n19657 = n1248 & n16433 ;
  assign n19658 = ( n1248 & n19656 ) | ( n1248 & ~n19657 ) | ( n19656 & ~n19657 ) ;
  assign n19659 = ( n19510 & ~n19651 ) | ( n19510 & n19658 ) | ( ~n19651 & n19658 ) ;
  assign n19660 = ( n19510 & n19651 ) | ( n19510 & n19658 ) | ( n19651 & n19658 ) ;
  assign n19661 = ( n19651 & n19659 ) | ( n19651 & ~n19660 ) | ( n19659 & ~n19660 ) ;
  assign n19662 = n3800 & n16553 ;
  assign n19663 = n3799 & n16053 ;
  assign n19664 = n3700 & ~n16057 ;
  assign n19665 = n3802 & ~n16055 ;
  assign n19666 = n19664 | n19665 ;
  assign n19667 = ( ~n19662 & n19663 ) | ( ~n19662 & n19666 ) | ( n19663 & n19666 ) ;
  assign n19668 = ( ~x29 & n19662 ) | ( ~x29 & n19667 ) | ( n19662 & n19667 ) ;
  assign n19669 = ( n19662 & n19667 ) | ( n19662 & ~n19668 ) | ( n19667 & ~n19668 ) ;
  assign n19670 = ( x29 & n19668 ) | ( x29 & ~n19669 ) | ( n19668 & ~n19669 ) ;
  assign n19671 = ( n19522 & ~n19661 ) | ( n19522 & n19670 ) | ( ~n19661 & n19670 ) ;
  assign n19672 = ( n19522 & n19661 ) | ( n19522 & n19670 ) | ( n19661 & n19670 ) ;
  assign n19673 = ( n19661 & n19671 ) | ( n19661 & ~n19672 ) | ( n19671 & ~n19672 ) ;
  assign n19674 = n4202 & ~n16801 ;
  assign n19675 = n4201 & ~n16047 ;
  assign n19676 = n4200 & ~n16051 ;
  assign n19677 = n4345 & ~n16049 ;
  assign n19678 = n19676 | n19677 ;
  assign n19679 = ( ~n19674 & n19675 ) | ( ~n19674 & n19678 ) | ( n19675 & n19678 ) ;
  assign n19680 = ( ~x26 & n19674 ) | ( ~x26 & n19679 ) | ( n19674 & n19679 ) ;
  assign n19681 = ( n19674 & n19679 ) | ( n19674 & ~n19680 ) | ( n19679 & ~n19680 ) ;
  assign n19682 = ( x26 & n19680 ) | ( x26 & ~n19681 ) | ( n19680 & ~n19681 ) ;
  assign n19683 = ( n19534 & ~n19673 ) | ( n19534 & n19682 ) | ( ~n19673 & n19682 ) ;
  assign n19684 = ( n19534 & n19673 ) | ( n19534 & n19682 ) | ( n19673 & n19682 ) ;
  assign n19685 = ( n19673 & n19683 ) | ( n19673 & ~n19684 ) | ( n19683 & ~n19684 ) ;
  assign n19686 = n4713 & n16969 ;
  assign n19687 = n4712 & n16041 ;
  assign n19688 = n4709 & ~n16045 ;
  assign n19689 = n4792 & ~n16043 ;
  assign n19690 = n19688 | n19689 ;
  assign n19691 = ( ~n19686 & n19687 ) | ( ~n19686 & n19690 ) | ( n19687 & n19690 ) ;
  assign n19692 = ( ~x23 & n19686 ) | ( ~x23 & n19691 ) | ( n19686 & n19691 ) ;
  assign n19693 = ( n19686 & n19691 ) | ( n19686 & ~n19692 ) | ( n19691 & ~n19692 ) ;
  assign n19694 = ( x23 & n19692 ) | ( x23 & ~n19693 ) | ( n19692 & ~n19693 ) ;
  assign n19695 = ( n19546 & ~n19685 ) | ( n19546 & n19694 ) | ( ~n19685 & n19694 ) ;
  assign n19696 = ( n19546 & n19685 ) | ( n19546 & n19694 ) | ( n19685 & n19694 ) ;
  assign n19697 = ( n19685 & n19695 ) | ( n19685 & ~n19696 ) | ( n19695 & ~n19696 ) ;
  assign n19698 = n4974 & ~n17313 ;
  assign n19699 = n5398 & n16035 ;
  assign n19700 = n4973 & n16039 ;
  assign n19701 = n4972 & ~n16037 ;
  assign n19702 = n19700 | n19701 ;
  assign n19703 = ( ~n19698 & n19699 ) | ( ~n19698 & n19702 ) | ( n19699 & n19702 ) ;
  assign n19704 = ( ~x20 & n19698 ) | ( ~x20 & n19703 ) | ( n19698 & n19703 ) ;
  assign n19705 = ( n19698 & n19703 ) | ( n19698 & ~n19704 ) | ( n19703 & ~n19704 ) ;
  assign n19706 = ( x20 & n19704 ) | ( x20 & ~n19705 ) | ( n19704 & ~n19705 ) ;
  assign n19707 = ( n19558 & ~n19697 ) | ( n19558 & n19706 ) | ( ~n19697 & n19706 ) ;
  assign n19708 = ( n19558 & n19697 ) | ( n19558 & n19706 ) | ( n19697 & n19706 ) ;
  assign n19709 = ( n19697 & n19707 ) | ( n19697 & ~n19708 ) | ( n19707 & ~n19708 ) ;
  assign n19710 = n5508 & ~n17528 ;
  assign n19711 = n5507 & ~n16029 ;
  assign n19712 = n5504 & ~n16033 ;
  assign n19713 = n5666 & n16031 ;
  assign n19714 = n19712 | n19713 ;
  assign n19715 = ( ~n19710 & n19711 ) | ( ~n19710 & n19714 ) | ( n19711 & n19714 ) ;
  assign n19716 = ( ~x17 & n19710 ) | ( ~x17 & n19715 ) | ( n19710 & n19715 ) ;
  assign n19717 = ( n19710 & n19715 ) | ( n19710 & ~n19716 ) | ( n19715 & ~n19716 ) ;
  assign n19718 = ( x17 & n19716 ) | ( x17 & ~n19717 ) | ( n19716 & ~n19717 ) ;
  assign n19719 = ( n19570 & ~n19709 ) | ( n19570 & n19718 ) | ( ~n19709 & n19718 ) ;
  assign n19720 = ( n19570 & n19709 ) | ( n19570 & n19718 ) | ( n19709 & n19718 ) ;
  assign n19721 = ( n19709 & n19719 ) | ( n19709 & ~n19720 ) | ( n19719 & ~n19720 ) ;
  assign n19722 = n5966 & n17968 ;
  assign n19723 = n6464 & n16023 ;
  assign n19724 = n5970 & ~n16027 ;
  assign n19725 = n5969 & ~n16025 ;
  assign n19726 = n19724 | n19725 ;
  assign n19727 = ( ~n19722 & n19723 ) | ( ~n19722 & n19726 ) | ( n19723 & n19726 ) ;
  assign n19728 = ( ~x14 & n19722 ) | ( ~x14 & n19727 ) | ( n19722 & n19727 ) ;
  assign n19729 = ( n19722 & n19727 ) | ( n19722 & ~n19728 ) | ( n19727 & ~n19728 ) ;
  assign n19730 = ( x14 & n19728 ) | ( x14 & ~n19729 ) | ( n19728 & ~n19729 ) ;
  assign n19731 = ( n19582 & ~n19721 ) | ( n19582 & n19730 ) | ( ~n19721 & n19730 ) ;
  assign n19732 = ( n19582 & n19721 ) | ( n19582 & n19730 ) | ( n19721 & n19730 ) ;
  assign n19733 = ( n19721 & n19731 ) | ( n19721 & ~n19732 ) | ( n19731 & ~n19732 ) ;
  assign n19734 = n6584 & ~n18267 ;
  assign n19735 = n7022 & ~n16017 ;
  assign n19736 = n6588 & n16021 ;
  assign n19737 = n6587 & n16019 ;
  assign n19738 = n19736 | n19737 ;
  assign n19739 = ( ~n19734 & n19735 ) | ( ~n19734 & n19738 ) | ( n19735 & n19738 ) ;
  assign n19740 = ( ~x11 & n19734 ) | ( ~x11 & n19739 ) | ( n19734 & n19739 ) ;
  assign n19741 = ( n19734 & n19739 ) | ( n19734 & ~n19740 ) | ( n19739 & ~n19740 ) ;
  assign n19742 = ( x11 & n19740 ) | ( x11 & ~n19741 ) | ( n19740 & ~n19741 ) ;
  assign n19743 = ( n19594 & ~n19733 ) | ( n19594 & n19742 ) | ( ~n19733 & n19742 ) ;
  assign n19744 = ( n19594 & n19733 ) | ( n19594 & n19742 ) | ( n19733 & n19742 ) ;
  assign n19745 = ( n19733 & n19743 ) | ( n19733 & ~n19744 ) | ( n19743 & ~n19744 ) ;
  assign n19746 = n7296 & ~n16144 ;
  assign n19747 = n7879 & n16138 ;
  assign n19748 = n7300 & n16015 ;
  assign n19749 = n7299 & ~n16013 ;
  assign n19750 = n19748 | n19749 ;
  assign n19751 = ( ~n19746 & n19747 ) | ( ~n19746 & n19750 ) | ( n19747 & n19750 ) ;
  assign n19752 = ( ~x8 & n19746 ) | ( ~x8 & n19751 ) | ( n19746 & n19751 ) ;
  assign n19753 = ( n19746 & n19751 ) | ( n19746 & ~n19752 ) | ( n19751 & ~n19752 ) ;
  assign n19754 = ( x8 & n19752 ) | ( x8 & ~n19753 ) | ( n19752 & ~n19753 ) ;
  assign n19755 = ( n19606 & ~n19745 ) | ( n19606 & n19754 ) | ( ~n19745 & n19754 ) ;
  assign n19756 = ( n19606 & n19745 ) | ( n19606 & n19754 ) | ( n19745 & n19754 ) ;
  assign n19757 = ( n19745 & n19755 ) | ( n19745 & ~n19756 ) | ( n19755 & ~n19756 ) ;
  assign n19758 = n8230 & ~n19312 ;
  assign n19759 = n8229 & ~n19309 ;
  assign n19760 = n8226 & n18993 ;
  assign n19761 = n8225 & n19157 ;
  assign n19762 = n19760 | n19761 ;
  assign n19763 = ( ~n19758 & n19759 ) | ( ~n19758 & n19762 ) | ( n19759 & n19762 ) ;
  assign n19764 = ( ~x5 & n19758 ) | ( ~x5 & n19763 ) | ( n19758 & n19763 ) ;
  assign n19765 = ( n19758 & n19763 ) | ( n19758 & ~n19764 ) | ( n19763 & ~n19764 ) ;
  assign n19766 = ( x5 & n19764 ) | ( x5 & ~n19765 ) | ( n19764 & ~n19765 ) ;
  assign n19767 = ( x2 & ~n19757 ) | ( x2 & n19766 ) | ( ~n19757 & n19766 ) ;
  assign n19768 = ( x2 & n19766 ) | ( x2 & ~n19767 ) | ( n19766 & ~n19767 ) ;
  assign n19769 = ( n19757 & n19767 ) | ( n19757 & ~n19768 ) | ( n19767 & ~n19768 ) ;
  assign n19770 = ( n19618 & n19623 ) | ( n19618 & ~n19769 ) | ( n19623 & ~n19769 ) ;
  assign n19771 = ( n19618 & ~n19623 ) | ( n19618 & n19769 ) | ( ~n19623 & n19769 ) ;
  assign n19772 = ( ~n19618 & n19770 ) | ( ~n19618 & n19771 ) | ( n19770 & n19771 ) ;
  assign n19773 = n19626 & ~n19772 ;
  assign n19774 = n19626 & n19772 ;
  assign n19775 = ( n19772 & n19773 ) | ( n19772 & ~n19774 ) | ( n19773 & ~n19774 ) ;
  assign n19776 = n4713 & ~n17051 ;
  assign n19777 = n4712 & n16039 ;
  assign n19778 = n4709 & ~n16043 ;
  assign n19779 = n4792 & n16041 ;
  assign n19780 = n19778 | n19779 ;
  assign n19781 = ( ~n19776 & n19777 ) | ( ~n19776 & n19780 ) | ( n19777 & n19780 ) ;
  assign n19782 = ( ~x23 & n19776 ) | ( ~x23 & n19781 ) | ( n19776 & n19781 ) ;
  assign n19783 = ( n19776 & n19781 ) | ( n19776 & ~n19782 ) | ( n19781 & ~n19782 ) ;
  assign n19784 = ( x23 & n19782 ) | ( x23 & ~n19783 ) | ( n19782 & ~n19783 ) ;
  assign n19785 = n254 | n992 ;
  assign n19786 = ( n732 & n1346 ) | ( n732 & ~n19785 ) | ( n1346 & ~n19785 ) ;
  assign n19787 = n19785 | n19786 ;
  assign n19788 = ( n10534 & ~n10941 ) | ( n10534 & n19787 ) | ( ~n10941 & n19787 ) ;
  assign n19789 = ( ~n3011 & n10941 ) | ( ~n3011 & n19788 ) | ( n10941 & n19788 ) ;
  assign n19790 = n3284 | n6026 ;
  assign n19791 = n434 | n1356 ;
  assign n19792 = ( n10973 & ~n19790 ) | ( n10973 & n19791 ) | ( ~n19790 & n19791 ) ;
  assign n19793 = n19790 | n19792 ;
  assign n19794 = ( n3011 & ~n19789 ) | ( n3011 & n19793 ) | ( ~n19789 & n19793 ) ;
  assign n19795 = n19789 | n19794 ;
  assign n19796 = n90 | n2815 ;
  assign n19797 = ( n10191 & n19795 ) | ( n10191 & ~n19796 ) | ( n19795 & ~n19796 ) ;
  assign n19798 = ~n19795 & n19797 ;
  assign n19799 = ( n573 & n3353 ) | ( n573 & n19798 ) | ( n3353 & n19798 ) ;
  assign n19800 = n19798 & ~n19799 ;
  assign n19801 = n607 & ~n16061 ;
  assign n19802 = n1250 & n16059 ;
  assign n19803 = n19801 | n19802 ;
  assign n19804 = n606 & n16057 ;
  assign n19805 = ( n606 & n19803 ) | ( n606 & ~n19804 ) | ( n19803 & ~n19804 ) ;
  assign n19806 = n1248 & n16484 ;
  assign n19807 = ( n1248 & n19805 ) | ( n1248 & ~n19806 ) | ( n19805 & ~n19806 ) ;
  assign n19808 = ( x2 & ~n19800 ) | ( x2 & n19807 ) | ( ~n19800 & n19807 ) ;
  assign n19809 = ( x2 & n19807 ) | ( x2 & ~n19808 ) | ( n19807 & ~n19808 ) ;
  assign n19810 = ( n19800 & n19808 ) | ( n19800 & ~n19809 ) | ( n19808 & ~n19809 ) ;
  assign n19811 = n3800 & n16611 ;
  assign n19812 = n3799 & ~n16051 ;
  assign n19813 = n3700 & ~n16055 ;
  assign n19814 = n3802 & n16053 ;
  assign n19815 = n19813 | n19814 ;
  assign n19816 = ( ~n19811 & n19812 ) | ( ~n19811 & n19815 ) | ( n19812 & n19815 ) ;
  assign n19817 = ( ~x29 & n19811 ) | ( ~x29 & n19816 ) | ( n19811 & n19816 ) ;
  assign n19818 = ( n19811 & n19816 ) | ( n19811 & ~n19817 ) | ( n19816 & ~n19817 ) ;
  assign n19819 = ( x29 & n19817 ) | ( x29 & ~n19818 ) | ( n19817 & ~n19818 ) ;
  assign n19820 = ( n19659 & ~n19810 ) | ( n19659 & n19819 ) | ( ~n19810 & n19819 ) ;
  assign n19821 = ( n19659 & n19810 ) | ( n19659 & n19819 ) | ( n19810 & n19819 ) ;
  assign n19822 = ( n19810 & n19820 ) | ( n19810 & ~n19821 ) | ( n19820 & ~n19821 ) ;
  assign n19823 = n4202 & ~n16876 ;
  assign n19824 = n4201 & ~n16045 ;
  assign n19825 = n4200 & ~n16049 ;
  assign n19826 = n4345 & ~n16047 ;
  assign n19827 = n19825 | n19826 ;
  assign n19828 = ( ~n19823 & n19824 ) | ( ~n19823 & n19827 ) | ( n19824 & n19827 ) ;
  assign n19829 = ( ~x26 & n19823 ) | ( ~x26 & n19828 ) | ( n19823 & n19828 ) ;
  assign n19830 = ( n19823 & n19828 ) | ( n19823 & ~n19829 ) | ( n19828 & ~n19829 ) ;
  assign n19831 = ( x26 & n19829 ) | ( x26 & ~n19830 ) | ( n19829 & ~n19830 ) ;
  assign n19832 = ( n19671 & ~n19822 ) | ( n19671 & n19831 ) | ( ~n19822 & n19831 ) ;
  assign n19833 = ( n19671 & n19822 ) | ( n19671 & n19831 ) | ( n19822 & n19831 ) ;
  assign n19834 = ( n19822 & n19832 ) | ( n19822 & ~n19833 ) | ( n19832 & ~n19833 ) ;
  assign n19835 = ( n19683 & n19784 ) | ( n19683 & ~n19834 ) | ( n19784 & ~n19834 ) ;
  assign n19836 = ( ~n19683 & n19784 ) | ( ~n19683 & n19834 ) | ( n19784 & n19834 ) ;
  assign n19837 = ( ~n19784 & n19835 ) | ( ~n19784 & n19836 ) | ( n19835 & n19836 ) ;
  assign n19838 = n4974 & ~n17412 ;
  assign n19839 = n5398 & ~n16033 ;
  assign n19840 = n4973 & ~n16037 ;
  assign n19841 = n4972 & n16035 ;
  assign n19842 = n19840 | n19841 ;
  assign n19843 = ( ~n19838 & n19839 ) | ( ~n19838 & n19842 ) | ( n19839 & n19842 ) ;
  assign n19844 = ( ~x20 & n19838 ) | ( ~x20 & n19843 ) | ( n19838 & n19843 ) ;
  assign n19845 = ( n19838 & n19843 ) | ( n19838 & ~n19844 ) | ( n19843 & ~n19844 ) ;
  assign n19846 = ( x20 & n19844 ) | ( x20 & ~n19845 ) | ( n19844 & ~n19845 ) ;
  assign n19847 = ( n19695 & ~n19837 ) | ( n19695 & n19846 ) | ( ~n19837 & n19846 ) ;
  assign n19848 = ( n19695 & n19837 ) | ( n19695 & n19846 ) | ( n19837 & n19846 ) ;
  assign n19849 = ( n19837 & n19847 ) | ( n19837 & ~n19848 ) | ( n19847 & ~n19848 ) ;
  assign n19850 = n5508 & n17634 ;
  assign n19851 = n5507 & ~n16027 ;
  assign n19852 = n5504 & n16031 ;
  assign n19853 = n5666 & ~n16029 ;
  assign n19854 = n19852 | n19853 ;
  assign n19855 = ( ~n19850 & n19851 ) | ( ~n19850 & n19854 ) | ( n19851 & n19854 ) ;
  assign n19856 = ( ~x17 & n19850 ) | ( ~x17 & n19855 ) | ( n19850 & n19855 ) ;
  assign n19857 = ( n19850 & n19855 ) | ( n19850 & ~n19856 ) | ( n19855 & ~n19856 ) ;
  assign n19858 = ( x17 & n19856 ) | ( x17 & ~n19857 ) | ( n19856 & ~n19857 ) ;
  assign n19859 = ( n19707 & ~n19849 ) | ( n19707 & n19858 ) | ( ~n19849 & n19858 ) ;
  assign n19860 = ( n19707 & n19849 ) | ( n19707 & n19858 ) | ( n19849 & n19858 ) ;
  assign n19861 = ( n19849 & n19859 ) | ( n19849 & ~n19860 ) | ( n19859 & ~n19860 ) ;
  assign n19862 = n5966 & ~n18091 ;
  assign n19863 = n6464 & n16021 ;
  assign n19864 = n5970 & ~n16025 ;
  assign n19865 = n5969 & n16023 ;
  assign n19866 = n19864 | n19865 ;
  assign n19867 = ( ~n19862 & n19863 ) | ( ~n19862 & n19866 ) | ( n19863 & n19866 ) ;
  assign n19868 = ( ~x14 & n19862 ) | ( ~x14 & n19867 ) | ( n19862 & n19867 ) ;
  assign n19869 = ( n19862 & n19867 ) | ( n19862 & ~n19868 ) | ( n19867 & ~n19868 ) ;
  assign n19870 = ( x14 & n19868 ) | ( x14 & ~n19869 ) | ( n19868 & ~n19869 ) ;
  assign n19871 = ( n19719 & ~n19861 ) | ( n19719 & n19870 ) | ( ~n19861 & n19870 ) ;
  assign n19872 = ( n19719 & n19861 ) | ( n19719 & n19870 ) | ( n19861 & n19870 ) ;
  assign n19873 = ( n19861 & n19871 ) | ( n19861 & ~n19872 ) | ( n19871 & ~n19872 ) ;
  assign n19874 = n6584 & ~n18416 ;
  assign n19875 = n7022 & n16015 ;
  assign n19876 = n6588 & n16019 ;
  assign n19877 = n6587 & ~n16017 ;
  assign n19878 = n19876 | n19877 ;
  assign n19879 = ( ~n19874 & n19875 ) | ( ~n19874 & n19878 ) | ( n19875 & n19878 ) ;
  assign n19880 = ( ~x11 & n19874 ) | ( ~x11 & n19879 ) | ( n19874 & n19879 ) ;
  assign n19881 = ( n19874 & n19879 ) | ( n19874 & ~n19880 ) | ( n19879 & ~n19880 ) ;
  assign n19882 = ( x11 & n19880 ) | ( x11 & ~n19881 ) | ( n19880 & ~n19881 ) ;
  assign n19883 = ( n19731 & ~n19873 ) | ( n19731 & n19882 ) | ( ~n19873 & n19882 ) ;
  assign n19884 = ( n19731 & n19873 ) | ( n19731 & n19882 ) | ( n19873 & n19882 ) ;
  assign n19885 = ( n19873 & n19883 ) | ( n19873 & ~n19884 ) | ( n19883 & ~n19884 ) ;
  assign n19886 = n7296 & n18996 ;
  assign n19887 = n7879 & n18993 ;
  assign n19888 = n7300 & ~n16013 ;
  assign n19889 = n7299 & n16138 ;
  assign n19890 = n19888 | n19889 ;
  assign n19891 = ( ~n19886 & n19887 ) | ( ~n19886 & n19890 ) | ( n19887 & n19890 ) ;
  assign n19892 = ( ~x8 & n19886 ) | ( ~x8 & n19891 ) | ( n19886 & n19891 ) ;
  assign n19893 = ( n19886 & n19891 ) | ( n19886 & ~n19892 ) | ( n19891 & ~n19892 ) ;
  assign n19894 = ( x8 & n19892 ) | ( x8 & ~n19893 ) | ( n19892 & ~n19893 ) ;
  assign n19895 = ( n19743 & ~n19885 ) | ( n19743 & n19894 ) | ( ~n19885 & n19894 ) ;
  assign n19896 = ( n19743 & n19885 ) | ( n19743 & n19894 ) | ( n19885 & n19894 ) ;
  assign n19897 = ( n19885 & n19895 ) | ( n19885 & ~n19896 ) | ( n19895 & ~n19896 ) ;
  assign n19898 = n8230 & ~n19472 ;
  assign n19899 = n8226 & n19157 ;
  assign n19900 = n8225 & ~n19309 ;
  assign n19901 = n19899 | n19900 ;
  assign n19902 = ~n19898 & n19901 ;
  assign n19903 = ( ~x5 & n19898 ) | ( ~x5 & n19902 ) | ( n19898 & n19902 ) ;
  assign n19904 = ( n19898 & n19902 ) | ( n19898 & ~n19903 ) | ( n19902 & ~n19903 ) ;
  assign n19905 = ( x5 & n19903 ) | ( x5 & ~n19904 ) | ( n19903 & ~n19904 ) ;
  assign n19906 = ( n19755 & ~n19897 ) | ( n19755 & n19905 ) | ( ~n19897 & n19905 ) ;
  assign n19907 = ( n19755 & n19897 ) | ( n19755 & n19905 ) | ( n19897 & n19905 ) ;
  assign n19908 = ( n19897 & n19906 ) | ( n19897 & ~n19907 ) | ( n19906 & ~n19907 ) ;
  assign n19909 = ( n19767 & n19770 ) | ( n19767 & ~n19908 ) | ( n19770 & ~n19908 ) ;
  assign n19910 = ( n19767 & ~n19770 ) | ( n19767 & n19908 ) | ( ~n19770 & n19908 ) ;
  assign n19911 = ( ~n19767 & n19909 ) | ( ~n19767 & n19910 ) | ( n19909 & n19910 ) ;
  assign n19912 = n19773 & ~n19911 ;
  assign n19913 = ~n19773 & n19911 ;
  assign n19914 = n19912 | n19913 ;
  assign n19915 = n2305 | n11830 ;
  assign n19916 = n172 | n185 ;
  assign n19917 = n519 | n1313 ;
  assign n19918 = ( n10141 & ~n19916 ) | ( n10141 & n19917 ) | ( ~n19916 & n19917 ) ;
  assign n19919 = n19916 | n19918 ;
  assign n19920 = n1144 | n2078 ;
  assign n19921 = n383 | n963 ;
  assign n19922 = n2414 | n2791 ;
  assign n19923 = ( n3273 & n3879 ) | ( n3273 & ~n19922 ) | ( n3879 & ~n19922 ) ;
  assign n19924 = n19922 | n19923 ;
  assign n19925 = ( n19920 & ~n19921 ) | ( n19920 & n19924 ) | ( ~n19921 & n19924 ) ;
  assign n19926 = n135 | n168 ;
  assign n19927 = ( n912 & n933 ) | ( n912 & ~n19926 ) | ( n933 & ~n19926 ) ;
  assign n19928 = n19926 | n19927 ;
  assign n19929 = n327 | n1235 ;
  assign n19930 = ( n18299 & ~n19928 ) | ( n18299 & n19929 ) | ( ~n19928 & n19929 ) ;
  assign n19931 = n19928 | n19930 ;
  assign n19932 = ( n19921 & ~n19925 ) | ( n19921 & n19931 ) | ( ~n19925 & n19931 ) ;
  assign n19933 = n19925 | n19932 ;
  assign n19934 = ( ~n19915 & n19919 ) | ( ~n19915 & n19933 ) | ( n19919 & n19933 ) ;
  assign n19935 = ( ~n3044 & n19915 ) | ( ~n3044 & n19934 ) | ( n19915 & n19934 ) ;
  assign n19936 = n3044 | n19935 ;
  assign n19937 = ( x2 & n19808 ) | ( x2 & n19936 ) | ( n19808 & n19936 ) ;
  assign n19938 = ( x2 & ~n19808 ) | ( x2 & n19936 ) | ( ~n19808 & n19936 ) ;
  assign n19939 = ( n19808 & ~n19937 ) | ( n19808 & n19938 ) | ( ~n19937 & n19938 ) ;
  assign n19940 = n607 & n16059 ;
  assign n19941 = n1250 & ~n16057 ;
  assign n19942 = n19940 | n19941 ;
  assign n19943 = n606 & n16055 ;
  assign n19944 = ( n606 & n19942 ) | ( n606 & ~n19943 ) | ( n19942 & ~n19943 ) ;
  assign n19945 = n1248 & n16541 ;
  assign n19946 = n19944 | n19945 ;
  assign n19947 = ( n19820 & n19939 ) | ( n19820 & n19946 ) | ( n19939 & n19946 ) ;
  assign n19948 = ( n19820 & ~n19939 ) | ( n19820 & n19946 ) | ( ~n19939 & n19946 ) ;
  assign n19949 = ( n19939 & ~n19947 ) | ( n19939 & n19948 ) | ( ~n19947 & n19948 ) ;
  assign n19950 = n4202 & ~n16957 ;
  assign n19951 = n4201 & ~n16043 ;
  assign n19952 = n4200 & ~n16047 ;
  assign n19953 = n4345 & ~n16045 ;
  assign n19954 = n19952 | n19953 ;
  assign n19955 = ( ~n19950 & n19951 ) | ( ~n19950 & n19954 ) | ( n19951 & n19954 ) ;
  assign n19956 = ( ~x26 & n19950 ) | ( ~x26 & n19955 ) | ( n19950 & n19955 ) ;
  assign n19957 = ( n19950 & n19955 ) | ( n19950 & ~n19956 ) | ( n19955 & ~n19956 ) ;
  assign n19958 = ( x26 & n19956 ) | ( x26 & ~n19957 ) | ( n19956 & ~n19957 ) ;
  assign n19959 = n3800 & ~n16674 ;
  assign n19960 = n3799 & ~n16049 ;
  assign n19961 = n3700 & n16053 ;
  assign n19962 = n3802 & ~n16051 ;
  assign n19963 = n19961 | n19962 ;
  assign n19964 = ( ~n19959 & n19960 ) | ( ~n19959 & n19963 ) | ( n19960 & n19963 ) ;
  assign n19965 = ( ~x29 & n19959 ) | ( ~x29 & n19964 ) | ( n19959 & n19964 ) ;
  assign n19966 = ( n19959 & n19964 ) | ( n19959 & ~n19965 ) | ( n19964 & ~n19965 ) ;
  assign n19967 = ( x29 & n19965 ) | ( x29 & ~n19966 ) | ( n19965 & ~n19966 ) ;
  assign n19968 = ( n19949 & n19958 ) | ( n19949 & n19967 ) | ( n19958 & n19967 ) ;
  assign n19969 = ( ~n19949 & n19958 ) | ( ~n19949 & n19967 ) | ( n19958 & n19967 ) ;
  assign n19970 = ( n19949 & ~n19968 ) | ( n19949 & n19969 ) | ( ~n19968 & n19969 ) ;
  assign n19971 = n4713 & ~n17138 ;
  assign n19972 = n4712 & ~n16037 ;
  assign n19973 = n4709 & n16041 ;
  assign n19974 = n4792 & n16039 ;
  assign n19975 = n19973 | n19974 ;
  assign n19976 = ( ~n19971 & n19972 ) | ( ~n19971 & n19975 ) | ( n19972 & n19975 ) ;
  assign n19977 = ( ~x23 & n19971 ) | ( ~x23 & n19976 ) | ( n19971 & n19976 ) ;
  assign n19978 = ( n19971 & n19976 ) | ( n19971 & ~n19977 ) | ( n19976 & ~n19977 ) ;
  assign n19979 = ( x23 & n19977 ) | ( x23 & ~n19978 ) | ( n19977 & ~n19978 ) ;
  assign n19980 = ( n19832 & n19970 ) | ( n19832 & n19979 ) | ( n19970 & n19979 ) ;
  assign n19981 = ( ~n19832 & n19970 ) | ( ~n19832 & n19979 ) | ( n19970 & n19979 ) ;
  assign n19982 = ( n19832 & ~n19980 ) | ( n19832 & n19981 ) | ( ~n19980 & n19981 ) ;
  assign n19983 = n4974 & ~n17516 ;
  assign n19984 = n5398 & n16031 ;
  assign n19985 = n4973 & n16035 ;
  assign n19986 = n4972 & ~n16033 ;
  assign n19987 = n19985 | n19986 ;
  assign n19988 = ( ~n19983 & n19984 ) | ( ~n19983 & n19987 ) | ( n19984 & n19987 ) ;
  assign n19989 = ( ~x20 & n19983 ) | ( ~x20 & n19988 ) | ( n19983 & n19988 ) ;
  assign n19990 = ( n19983 & n19988 ) | ( n19983 & ~n19989 ) | ( n19988 & ~n19989 ) ;
  assign n19991 = ( x20 & n19989 ) | ( x20 & ~n19990 ) | ( n19989 & ~n19990 ) ;
  assign n19992 = ( n19835 & n19982 ) | ( n19835 & n19991 ) | ( n19982 & n19991 ) ;
  assign n19993 = ( n19835 & ~n19982 ) | ( n19835 & n19991 ) | ( ~n19982 & n19991 ) ;
  assign n19994 = ( n19982 & ~n19992 ) | ( n19982 & n19993 ) | ( ~n19992 & n19993 ) ;
  assign n19995 = n5508 & ~n17746 ;
  assign n19996 = n5507 & ~n16025 ;
  assign n19997 = n5504 & ~n16029 ;
  assign n19998 = n5666 & ~n16027 ;
  assign n19999 = n19997 | n19998 ;
  assign n20000 = ( ~n19995 & n19996 ) | ( ~n19995 & n19999 ) | ( n19996 & n19999 ) ;
  assign n20001 = ( ~x17 & n19995 ) | ( ~x17 & n20000 ) | ( n19995 & n20000 ) ;
  assign n20002 = ( n19995 & n20000 ) | ( n19995 & ~n20001 ) | ( n20000 & ~n20001 ) ;
  assign n20003 = ( x17 & n20001 ) | ( x17 & ~n20002 ) | ( n20001 & ~n20002 ) ;
  assign n20004 = ( n19847 & n19994 ) | ( n19847 & n20003 ) | ( n19994 & n20003 ) ;
  assign n20005 = ( n19847 & ~n19994 ) | ( n19847 & n20003 ) | ( ~n19994 & n20003 ) ;
  assign n20006 = ( n19994 & ~n20004 ) | ( n19994 & n20005 ) | ( ~n20004 & n20005 ) ;
  assign n20007 = n5966 & n18103 ;
  assign n20008 = n6464 & n16019 ;
  assign n20009 = n5970 & n16023 ;
  assign n20010 = n5969 & n16021 ;
  assign n20011 = n20009 | n20010 ;
  assign n20012 = ( ~n20007 & n20008 ) | ( ~n20007 & n20011 ) | ( n20008 & n20011 ) ;
  assign n20013 = ( ~x14 & n20007 ) | ( ~x14 & n20012 ) | ( n20007 & n20012 ) ;
  assign n20014 = ( n20007 & n20012 ) | ( n20007 & ~n20013 ) | ( n20012 & ~n20013 ) ;
  assign n20015 = ( x14 & n20013 ) | ( x14 & ~n20014 ) | ( n20013 & ~n20014 ) ;
  assign n20016 = ( n19859 & n20006 ) | ( n19859 & n20015 ) | ( n20006 & n20015 ) ;
  assign n20017 = ( n19859 & ~n20006 ) | ( n19859 & n20015 ) | ( ~n20006 & n20015 ) ;
  assign n20018 = ( n20006 & ~n20016 ) | ( n20006 & n20017 ) | ( ~n20016 & n20017 ) ;
  assign n20019 = n6584 & ~n18694 ;
  assign n20020 = n7022 & ~n16013 ;
  assign n20021 = n6588 & ~n16017 ;
  assign n20022 = n6587 & n16015 ;
  assign n20023 = n20021 | n20022 ;
  assign n20024 = ( ~n20019 & n20020 ) | ( ~n20019 & n20023 ) | ( n20020 & n20023 ) ;
  assign n20025 = ( ~x11 & n20019 ) | ( ~x11 & n20024 ) | ( n20019 & n20024 ) ;
  assign n20026 = ( n20019 & n20024 ) | ( n20019 & ~n20025 ) | ( n20024 & ~n20025 ) ;
  assign n20027 = ( x11 & n20025 ) | ( x11 & ~n20026 ) | ( n20025 & ~n20026 ) ;
  assign n20028 = ( n19871 & n20018 ) | ( n19871 & n20027 ) | ( n20018 & n20027 ) ;
  assign n20029 = ( n19871 & ~n20018 ) | ( n19871 & n20027 ) | ( ~n20018 & n20027 ) ;
  assign n20030 = ( n20018 & ~n20028 ) | ( n20018 & n20029 ) | ( ~n20028 & n20029 ) ;
  assign n20031 = n7296 & n19160 ;
  assign n20032 = n7879 & n19157 ;
  assign n20033 = n7300 & n16138 ;
  assign n20034 = n7299 & n18993 ;
  assign n20035 = n20033 | n20034 ;
  assign n20036 = ( ~n20031 & n20032 ) | ( ~n20031 & n20035 ) | ( n20032 & n20035 ) ;
  assign n20037 = ( ~x8 & n20031 ) | ( ~x8 & n20036 ) | ( n20031 & n20036 ) ;
  assign n20038 = ( n20031 & n20036 ) | ( n20031 & ~n20037 ) | ( n20036 & ~n20037 ) ;
  assign n20039 = ( x8 & n20037 ) | ( x8 & ~n20038 ) | ( n20037 & ~n20038 ) ;
  assign n20040 = ( n19883 & n20030 ) | ( n19883 & n20039 ) | ( n20030 & n20039 ) ;
  assign n20041 = ( n19883 & ~n20030 ) | ( n19883 & n20039 ) | ( ~n20030 & n20039 ) ;
  assign n20042 = ( n20030 & ~n20040 ) | ( n20030 & n20041 ) | ( ~n20040 & n20041 ) ;
  assign n20043 = n8226 & ~n19309 ;
  assign n20044 = ~x5 & n20043 ;
  assign n20045 = n20043 & ~n20044 ;
  assign n20046 = ( x5 & n20044 ) | ( x5 & ~n20045 ) | ( n20044 & ~n20045 ) ;
  assign n20047 = ( n19895 & n20042 ) | ( n19895 & n20046 ) | ( n20042 & n20046 ) ;
  assign n20048 = ( n19895 & ~n20042 ) | ( n19895 & n20046 ) | ( ~n20042 & n20046 ) ;
  assign n20049 = ( n20042 & ~n20047 ) | ( n20042 & n20048 ) | ( ~n20047 & n20048 ) ;
  assign n20050 = ( n19906 & n19909 ) | ( n19906 & n20049 ) | ( n19909 & n20049 ) ;
  assign n20051 = ( n19906 & ~n19909 ) | ( n19906 & n20049 ) | ( ~n19909 & n20049 ) ;
  assign n20052 = ( n19909 & ~n20050 ) | ( n19909 & n20051 ) | ( ~n20050 & n20051 ) ;
  assign n20053 = n19912 & n20052 ;
  assign n20054 = n19912 & ~n20052 ;
  assign n20055 = ( n20052 & ~n20053 ) | ( n20052 & n20054 ) | ( ~n20053 & n20054 ) ;
  assign n20056 = n3285 | n3830 ;
  assign n20057 = n2232 | n3522 ;
  assign n20058 = n4848 | n20057 ;
  assign n20059 = ( ~n11579 & n20056 ) | ( ~n11579 & n20058 ) | ( n20056 & n20058 ) ;
  assign n20060 = n394 | n1237 ;
  assign n20061 = n514 | n20060 ;
  assign n20062 = n159 | n208 ;
  assign n20063 = ( n969 & ~n20061 ) | ( n969 & n20062 ) | ( ~n20061 & n20062 ) ;
  assign n20064 = n20061 | n20063 ;
  assign n20065 = n11579 | n20064 ;
  assign n20066 = ( n1769 & n5107 ) | ( n1769 & ~n20064 ) | ( n5107 & ~n20064 ) ;
  assign n20067 = ( ~n20059 & n20065 ) | ( ~n20059 & n20066 ) | ( n20065 & n20066 ) ;
  assign n20068 = n20059 | n20067 ;
  assign n20069 = ( n2021 & n3057 ) | ( n2021 & ~n20068 ) | ( n3057 & ~n20068 ) ;
  assign n20070 = n20068 | n20069 ;
  assign n20071 = ( x2 & n19937 ) | ( x2 & n20070 ) | ( n19937 & n20070 ) ;
  assign n20072 = ( ~x2 & n19937 ) | ( ~x2 & n20070 ) | ( n19937 & n20070 ) ;
  assign n20073 = ( x2 & ~n20071 ) | ( x2 & n20072 ) | ( ~n20071 & n20072 ) ;
  assign n20074 = n607 & ~n16057 ;
  assign n20075 = n1250 & ~n16055 ;
  assign n20076 = n20074 | n20075 ;
  assign n20077 = n606 & ~n16053 ;
  assign n20078 = ( n606 & n20076 ) | ( n606 & ~n20077 ) | ( n20076 & ~n20077 ) ;
  assign n20079 = n1248 & ~n16553 ;
  assign n20080 = ( n1248 & n20078 ) | ( n1248 & ~n20079 ) | ( n20078 & ~n20079 ) ;
  assign n20081 = ( n19947 & n20073 ) | ( n19947 & n20080 ) | ( n20073 & n20080 ) ;
  assign n20082 = ( n19947 & ~n20073 ) | ( n19947 & n20080 ) | ( ~n20073 & n20080 ) ;
  assign n20083 = ( n20073 & ~n20081 ) | ( n20073 & n20082 ) | ( ~n20081 & n20082 ) ;
  assign n20084 = n4202 & n16969 ;
  assign n20085 = n4201 & n16041 ;
  assign n20086 = n4200 & ~n16045 ;
  assign n20087 = n4345 & ~n16043 ;
  assign n20088 = n20086 | n20087 ;
  assign n20089 = ( ~n20084 & n20085 ) | ( ~n20084 & n20088 ) | ( n20085 & n20088 ) ;
  assign n20090 = ( ~x26 & n20084 ) | ( ~x26 & n20089 ) | ( n20084 & n20089 ) ;
  assign n20091 = ( n20084 & n20089 ) | ( n20084 & ~n20090 ) | ( n20089 & ~n20090 ) ;
  assign n20092 = ( x26 & n20090 ) | ( x26 & ~n20091 ) | ( n20090 & ~n20091 ) ;
  assign n20093 = n3800 & ~n16801 ;
  assign n20094 = n3799 & ~n16047 ;
  assign n20095 = n3700 & ~n16051 ;
  assign n20096 = n3802 & ~n16049 ;
  assign n20097 = n20095 | n20096 ;
  assign n20098 = ( ~n20093 & n20094 ) | ( ~n20093 & n20097 ) | ( n20094 & n20097 ) ;
  assign n20099 = ( ~x29 & n20093 ) | ( ~x29 & n20098 ) | ( n20093 & n20098 ) ;
  assign n20100 = ( n20093 & n20098 ) | ( n20093 & ~n20099 ) | ( n20098 & ~n20099 ) ;
  assign n20101 = ( x29 & n20099 ) | ( x29 & ~n20100 ) | ( n20099 & ~n20100 ) ;
  assign n20102 = ( n20083 & n20092 ) | ( n20083 & n20101 ) | ( n20092 & n20101 ) ;
  assign n20103 = ( ~n20083 & n20092 ) | ( ~n20083 & n20101 ) | ( n20092 & n20101 ) ;
  assign n20104 = ( n20083 & ~n20102 ) | ( n20083 & n20103 ) | ( ~n20102 & n20103 ) ;
  assign n20105 = n4713 & ~n17313 ;
  assign n20106 = n4712 & n16035 ;
  assign n20107 = n4709 & n16039 ;
  assign n20108 = n4792 & ~n16037 ;
  assign n20109 = n20107 | n20108 ;
  assign n20110 = ( ~n20105 & n20106 ) | ( ~n20105 & n20109 ) | ( n20106 & n20109 ) ;
  assign n20111 = ( ~x23 & n20105 ) | ( ~x23 & n20110 ) | ( n20105 & n20110 ) ;
  assign n20112 = ( n20105 & n20110 ) | ( n20105 & ~n20111 ) | ( n20110 & ~n20111 ) ;
  assign n20113 = ( x23 & n20111 ) | ( x23 & ~n20112 ) | ( n20111 & ~n20112 ) ;
  assign n20114 = ( n19968 & n20104 ) | ( n19968 & n20113 ) | ( n20104 & n20113 ) ;
  assign n20115 = ( n19968 & ~n20104 ) | ( n19968 & n20113 ) | ( ~n20104 & n20113 ) ;
  assign n20116 = ( n20104 & ~n20114 ) | ( n20104 & n20115 ) | ( ~n20114 & n20115 ) ;
  assign n20117 = n4974 & ~n17528 ;
  assign n20118 = n5398 & ~n16029 ;
  assign n20119 = n4973 & ~n16033 ;
  assign n20120 = n4972 & n16031 ;
  assign n20121 = n20119 | n20120 ;
  assign n20122 = ( ~n20117 & n20118 ) | ( ~n20117 & n20121 ) | ( n20118 & n20121 ) ;
  assign n20123 = ( ~x20 & n20117 ) | ( ~x20 & n20122 ) | ( n20117 & n20122 ) ;
  assign n20124 = ( n20117 & n20122 ) | ( n20117 & ~n20123 ) | ( n20122 & ~n20123 ) ;
  assign n20125 = ( x20 & n20123 ) | ( x20 & ~n20124 ) | ( n20123 & ~n20124 ) ;
  assign n20126 = ( n19980 & n20116 ) | ( n19980 & n20125 ) | ( n20116 & n20125 ) ;
  assign n20127 = ( n19980 & ~n20116 ) | ( n19980 & n20125 ) | ( ~n20116 & n20125 ) ;
  assign n20128 = ( n20116 & ~n20126 ) | ( n20116 & n20127 ) | ( ~n20126 & n20127 ) ;
  assign n20129 = n5508 & n17968 ;
  assign n20130 = n5507 & n16023 ;
  assign n20131 = n5504 & ~n16027 ;
  assign n20132 = n5666 & ~n16025 ;
  assign n20133 = n20131 | n20132 ;
  assign n20134 = ( ~n20129 & n20130 ) | ( ~n20129 & n20133 ) | ( n20130 & n20133 ) ;
  assign n20135 = ( ~x17 & n20129 ) | ( ~x17 & n20134 ) | ( n20129 & n20134 ) ;
  assign n20136 = ( n20129 & n20134 ) | ( n20129 & ~n20135 ) | ( n20134 & ~n20135 ) ;
  assign n20137 = ( x17 & n20135 ) | ( x17 & ~n20136 ) | ( n20135 & ~n20136 ) ;
  assign n20138 = ( n19992 & n20128 ) | ( n19992 & n20137 ) | ( n20128 & n20137 ) ;
  assign n20139 = ( n19992 & ~n20128 ) | ( n19992 & n20137 ) | ( ~n20128 & n20137 ) ;
  assign n20140 = ( n20128 & ~n20138 ) | ( n20128 & n20139 ) | ( ~n20138 & n20139 ) ;
  assign n20141 = n5966 & ~n18267 ;
  assign n20142 = n6464 & ~n16017 ;
  assign n20143 = n5970 & n16021 ;
  assign n20144 = n5969 & n16019 ;
  assign n20145 = n20143 | n20144 ;
  assign n20146 = ( ~n20141 & n20142 ) | ( ~n20141 & n20145 ) | ( n20142 & n20145 ) ;
  assign n20147 = ( ~x14 & n20141 ) | ( ~x14 & n20146 ) | ( n20141 & n20146 ) ;
  assign n20148 = ( n20141 & n20146 ) | ( n20141 & ~n20147 ) | ( n20146 & ~n20147 ) ;
  assign n20149 = ( x14 & n20147 ) | ( x14 & ~n20148 ) | ( n20147 & ~n20148 ) ;
  assign n20150 = ( n20004 & n20140 ) | ( n20004 & n20149 ) | ( n20140 & n20149 ) ;
  assign n20151 = ( n20004 & ~n20140 ) | ( n20004 & n20149 ) | ( ~n20140 & n20149 ) ;
  assign n20152 = ( n20140 & ~n20150 ) | ( n20140 & n20151 ) | ( ~n20150 & n20151 ) ;
  assign n20153 = n6584 & ~n16144 ;
  assign n20154 = n7022 & n16138 ;
  assign n20155 = n6588 & n16015 ;
  assign n20156 = n6587 & ~n16013 ;
  assign n20157 = n20155 | n20156 ;
  assign n20158 = ( ~n20153 & n20154 ) | ( ~n20153 & n20157 ) | ( n20154 & n20157 ) ;
  assign n20159 = ( ~x11 & n20153 ) | ( ~x11 & n20158 ) | ( n20153 & n20158 ) ;
  assign n20160 = ( n20153 & n20158 ) | ( n20153 & ~n20159 ) | ( n20158 & ~n20159 ) ;
  assign n20161 = ( x11 & n20159 ) | ( x11 & ~n20160 ) | ( n20159 & ~n20160 ) ;
  assign n20162 = ( n20016 & n20152 ) | ( n20016 & n20161 ) | ( n20152 & n20161 ) ;
  assign n20163 = ( n20016 & ~n20152 ) | ( n20016 & n20161 ) | ( ~n20152 & n20161 ) ;
  assign n20164 = ( n20152 & ~n20162 ) | ( n20152 & n20163 ) | ( ~n20162 & n20163 ) ;
  assign n20165 = n7296 & ~n19312 ;
  assign n20166 = n7879 & ~n19309 ;
  assign n20167 = n7300 & n18993 ;
  assign n20168 = n7299 & n19157 ;
  assign n20169 = n20167 | n20168 ;
  assign n20170 = ( ~n20165 & n20166 ) | ( ~n20165 & n20169 ) | ( n20166 & n20169 ) ;
  assign n20171 = ( ~x8 & n20165 ) | ( ~x8 & n20170 ) | ( n20165 & n20170 ) ;
  assign n20172 = ( n20165 & n20170 ) | ( n20165 & ~n20171 ) | ( n20170 & ~n20171 ) ;
  assign n20173 = ( x8 & n20171 ) | ( x8 & ~n20172 ) | ( n20171 & ~n20172 ) ;
  assign n20174 = ( n20028 & n20164 ) | ( n20028 & n20173 ) | ( n20164 & n20173 ) ;
  assign n20175 = ( n20028 & ~n20164 ) | ( n20028 & n20173 ) | ( ~n20164 & n20173 ) ;
  assign n20176 = ( n20164 & ~n20174 ) | ( n20164 & n20175 ) | ( ~n20174 & n20175 ) ;
  assign n20177 = ( x5 & n20040 ) | ( x5 & n20176 ) | ( n20040 & n20176 ) ;
  assign n20178 = ( ~x5 & n20040 ) | ( ~x5 & n20176 ) | ( n20040 & n20176 ) ;
  assign n20179 = ( x5 & ~n20177 ) | ( x5 & n20178 ) | ( ~n20177 & n20178 ) ;
  assign n20180 = ( n20047 & n20050 ) | ( n20047 & n20179 ) | ( n20050 & n20179 ) ;
  assign n20181 = ( n20047 & ~n20050 ) | ( n20047 & n20179 ) | ( ~n20050 & n20179 ) ;
  assign n20182 = ( n20050 & ~n20180 ) | ( n20050 & n20181 ) | ( ~n20180 & n20181 ) ;
  assign n20183 = n20053 & n20182 ;
  assign n20184 = n20053 | n20182 ;
  assign n20185 = ~n20183 & n20184 ;
  assign n20186 = n4202 & ~n17051 ;
  assign n20187 = n4201 & n16039 ;
  assign n20188 = n4200 & ~n16043 ;
  assign n20189 = n4345 & n16041 ;
  assign n20190 = n20188 | n20189 ;
  assign n20191 = ( ~n20186 & n20187 ) | ( ~n20186 & n20190 ) | ( n20187 & n20190 ) ;
  assign n20192 = ( ~x26 & n20186 ) | ( ~x26 & n20191 ) | ( n20186 & n20191 ) ;
  assign n20193 = ( n20186 & n20191 ) | ( n20186 & ~n20192 ) | ( n20191 & ~n20192 ) ;
  assign n20194 = ( x26 & n20192 ) | ( x26 & ~n20193 ) | ( n20192 & ~n20193 ) ;
  assign n20195 = ( n72 & n129 ) | ( n72 & n136 ) | ( n129 & n136 ) ;
  assign n20196 = ( n83 & n109 ) | ( n83 & n116 ) | ( n109 & n116 ) ;
  assign n20197 = n20195 | n20196 ;
  assign n20198 = n1254 | n1423 ;
  assign n20199 = ( n5008 & ~n20197 ) | ( n5008 & n20198 ) | ( ~n20197 & n20198 ) ;
  assign n20200 = n20197 | n20199 ;
  assign n20201 = n2167 | n2205 ;
  assign n20202 = ( n3339 & n4495 ) | ( n3339 & ~n20201 ) | ( n4495 & ~n20201 ) ;
  assign n20203 = n20201 | n20202 ;
  assign n20204 = ( n10622 & ~n20200 ) | ( n10622 & n20203 ) | ( ~n20200 & n20203 ) ;
  assign n20205 = n20200 | n20204 ;
  assign n20206 = ( ~n2757 & n4001 ) | ( ~n2757 & n18175 ) | ( n4001 & n18175 ) ;
  assign n20207 = ( n2757 & ~n20205 ) | ( n2757 & n20206 ) | ( ~n20205 & n20206 ) ;
  assign n20208 = n20205 | n20207 ;
  assign n20209 = ( x2 & x5 ) | ( x2 & ~n20208 ) | ( x5 & ~n20208 ) ;
  assign n20210 = ( x2 & x5 ) | ( x2 & n20208 ) | ( x5 & n20208 ) ;
  assign n20211 = ( n20208 & n20209 ) | ( n20208 & ~n20210 ) | ( n20209 & ~n20210 ) ;
  assign n20212 = n607 & ~n16055 ;
  assign n20213 = n1250 & n16053 ;
  assign n20214 = n20212 | n20213 ;
  assign n20215 = n606 & n16051 ;
  assign n20216 = ( n606 & n20214 ) | ( n606 & ~n20215 ) | ( n20214 & ~n20215 ) ;
  assign n20217 = n1248 & ~n16611 ;
  assign n20218 = ( n1248 & n20216 ) | ( n1248 & ~n20217 ) | ( n20216 & ~n20217 ) ;
  assign n20219 = ( n20071 & n20211 ) | ( n20071 & n20218 ) | ( n20211 & n20218 ) ;
  assign n20220 = ( n20071 & ~n20211 ) | ( n20071 & n20218 ) | ( ~n20211 & n20218 ) ;
  assign n20221 = ( n20211 & ~n20219 ) | ( n20211 & n20220 ) | ( ~n20219 & n20220 ) ;
  assign n20222 = n3800 & ~n16876 ;
  assign n20223 = n3799 & ~n16045 ;
  assign n20224 = n3700 & ~n16049 ;
  assign n20225 = n3802 & ~n16047 ;
  assign n20226 = n20224 | n20225 ;
  assign n20227 = ( ~n20222 & n20223 ) | ( ~n20222 & n20226 ) | ( n20223 & n20226 ) ;
  assign n20228 = ( ~x29 & n20222 ) | ( ~x29 & n20227 ) | ( n20222 & n20227 ) ;
  assign n20229 = ( n20222 & n20227 ) | ( n20222 & ~n20228 ) | ( n20227 & ~n20228 ) ;
  assign n20230 = ( x29 & n20228 ) | ( x29 & ~n20229 ) | ( n20228 & ~n20229 ) ;
  assign n20231 = ( n20081 & n20221 ) | ( n20081 & n20230 ) | ( n20221 & n20230 ) ;
  assign n20232 = ( n20081 & ~n20221 ) | ( n20081 & n20230 ) | ( ~n20221 & n20230 ) ;
  assign n20233 = ( n20221 & ~n20231 ) | ( n20221 & n20232 ) | ( ~n20231 & n20232 ) ;
  assign n20234 = ( n20102 & n20194 ) | ( n20102 & n20233 ) | ( n20194 & n20233 ) ;
  assign n20235 = ( n20102 & ~n20194 ) | ( n20102 & n20233 ) | ( ~n20194 & n20233 ) ;
  assign n20236 = ( n20194 & ~n20234 ) | ( n20194 & n20235 ) | ( ~n20234 & n20235 ) ;
  assign n20237 = n4713 & ~n17412 ;
  assign n20238 = n4712 & ~n16033 ;
  assign n20239 = n4709 & ~n16037 ;
  assign n20240 = n4792 & n16035 ;
  assign n20241 = n20239 | n20240 ;
  assign n20242 = ( ~n20237 & n20238 ) | ( ~n20237 & n20241 ) | ( n20238 & n20241 ) ;
  assign n20243 = ( ~x23 & n20237 ) | ( ~x23 & n20242 ) | ( n20237 & n20242 ) ;
  assign n20244 = ( n20237 & n20242 ) | ( n20237 & ~n20243 ) | ( n20242 & ~n20243 ) ;
  assign n20245 = ( x23 & n20243 ) | ( x23 & ~n20244 ) | ( n20243 & ~n20244 ) ;
  assign n20246 = ( n20114 & n20236 ) | ( n20114 & n20245 ) | ( n20236 & n20245 ) ;
  assign n20247 = ( n20114 & ~n20236 ) | ( n20114 & n20245 ) | ( ~n20236 & n20245 ) ;
  assign n20248 = ( n20236 & ~n20246 ) | ( n20236 & n20247 ) | ( ~n20246 & n20247 ) ;
  assign n20249 = n4974 & n17634 ;
  assign n20250 = n5398 & ~n16027 ;
  assign n20251 = n4973 & n16031 ;
  assign n20252 = n4972 & ~n16029 ;
  assign n20253 = n20251 | n20252 ;
  assign n20254 = ( ~n20249 & n20250 ) | ( ~n20249 & n20253 ) | ( n20250 & n20253 ) ;
  assign n20255 = ( ~x20 & n20249 ) | ( ~x20 & n20254 ) | ( n20249 & n20254 ) ;
  assign n20256 = ( n20249 & n20254 ) | ( n20249 & ~n20255 ) | ( n20254 & ~n20255 ) ;
  assign n20257 = ( x20 & n20255 ) | ( x20 & ~n20256 ) | ( n20255 & ~n20256 ) ;
  assign n20258 = ( n20126 & n20248 ) | ( n20126 & n20257 ) | ( n20248 & n20257 ) ;
  assign n20259 = ( n20126 & ~n20248 ) | ( n20126 & n20257 ) | ( ~n20248 & n20257 ) ;
  assign n20260 = ( n20248 & ~n20258 ) | ( n20248 & n20259 ) | ( ~n20258 & n20259 ) ;
  assign n20261 = n5508 & ~n18091 ;
  assign n20262 = n5507 & n16021 ;
  assign n20263 = n5504 & ~n16025 ;
  assign n20264 = n5666 & n16023 ;
  assign n20265 = n20263 | n20264 ;
  assign n20266 = ( ~n20261 & n20262 ) | ( ~n20261 & n20265 ) | ( n20262 & n20265 ) ;
  assign n20267 = ( ~x17 & n20261 ) | ( ~x17 & n20266 ) | ( n20261 & n20266 ) ;
  assign n20268 = ( n20261 & n20266 ) | ( n20261 & ~n20267 ) | ( n20266 & ~n20267 ) ;
  assign n20269 = ( x17 & n20267 ) | ( x17 & ~n20268 ) | ( n20267 & ~n20268 ) ;
  assign n20270 = ( n20138 & n20260 ) | ( n20138 & n20269 ) | ( n20260 & n20269 ) ;
  assign n20271 = ( n20138 & ~n20260 ) | ( n20138 & n20269 ) | ( ~n20260 & n20269 ) ;
  assign n20272 = ( n20260 & ~n20270 ) | ( n20260 & n20271 ) | ( ~n20270 & n20271 ) ;
  assign n20273 = n5966 & ~n18416 ;
  assign n20274 = n6464 & n16015 ;
  assign n20275 = n5970 & n16019 ;
  assign n20276 = n5969 & ~n16017 ;
  assign n20277 = n20275 | n20276 ;
  assign n20278 = ( ~n20273 & n20274 ) | ( ~n20273 & n20277 ) | ( n20274 & n20277 ) ;
  assign n20279 = ( ~x14 & n20273 ) | ( ~x14 & n20278 ) | ( n20273 & n20278 ) ;
  assign n20280 = ( n20273 & n20278 ) | ( n20273 & ~n20279 ) | ( n20278 & ~n20279 ) ;
  assign n20281 = ( x14 & n20279 ) | ( x14 & ~n20280 ) | ( n20279 & ~n20280 ) ;
  assign n20282 = ( n20150 & n20272 ) | ( n20150 & n20281 ) | ( n20272 & n20281 ) ;
  assign n20283 = ( ~n20150 & n20272 ) | ( ~n20150 & n20281 ) | ( n20272 & n20281 ) ;
  assign n20284 = ( n20150 & ~n20282 ) | ( n20150 & n20283 ) | ( ~n20282 & n20283 ) ;
  assign n20285 = n6584 & n18996 ;
  assign n20286 = n7022 & n18993 ;
  assign n20287 = n6588 & ~n16013 ;
  assign n20288 = n6587 & n16138 ;
  assign n20289 = n20287 | n20288 ;
  assign n20290 = ( ~n20285 & n20286 ) | ( ~n20285 & n20289 ) | ( n20286 & n20289 ) ;
  assign n20291 = ( ~x11 & n20285 ) | ( ~x11 & n20290 ) | ( n20285 & n20290 ) ;
  assign n20292 = ( n20285 & n20290 ) | ( n20285 & ~n20291 ) | ( n20290 & ~n20291 ) ;
  assign n20293 = ( x11 & n20291 ) | ( x11 & ~n20292 ) | ( n20291 & ~n20292 ) ;
  assign n20294 = ( n20162 & n20284 ) | ( n20162 & n20293 ) | ( n20284 & n20293 ) ;
  assign n20295 = ( n20162 & ~n20284 ) | ( n20162 & n20293 ) | ( ~n20284 & n20293 ) ;
  assign n20296 = ( n20284 & ~n20294 ) | ( n20284 & n20295 ) | ( ~n20294 & n20295 ) ;
  assign n20297 = n7296 & ~n19472 ;
  assign n20298 = n7300 & n19157 ;
  assign n20299 = n7299 & ~n19309 ;
  assign n20300 = n20298 | n20299 ;
  assign n20301 = ~n20297 & n20300 ;
  assign n20302 = ( ~x8 & n20297 ) | ( ~x8 & n20301 ) | ( n20297 & n20301 ) ;
  assign n20303 = ( n20297 & n20301 ) | ( n20297 & ~n20302 ) | ( n20301 & ~n20302 ) ;
  assign n20304 = ( x8 & n20302 ) | ( x8 & ~n20303 ) | ( n20302 & ~n20303 ) ;
  assign n20305 = ( n20174 & n20296 ) | ( n20174 & n20304 ) | ( n20296 & n20304 ) ;
  assign n20306 = ( ~n20174 & n20296 ) | ( ~n20174 & n20304 ) | ( n20296 & n20304 ) ;
  assign n20307 = ( n20174 & ~n20305 ) | ( n20174 & n20306 ) | ( ~n20305 & n20306 ) ;
  assign n20308 = ( n20177 & n20180 ) | ( n20177 & n20307 ) | ( n20180 & n20307 ) ;
  assign n20309 = ( ~n20177 & n20180 ) | ( ~n20177 & n20307 ) | ( n20180 & n20307 ) ;
  assign n20310 = ( n20177 & ~n20308 ) | ( n20177 & n20309 ) | ( ~n20308 & n20309 ) ;
  assign n20311 = n20183 & n20310 ;
  assign n20312 = n20183 & ~n20310 ;
  assign n20313 = ( n20310 & ~n20311 ) | ( n20310 & n20312 ) | ( ~n20311 & n20312 ) ;
  assign n20314 = ( n810 & n1237 ) | ( n810 & ~n1588 ) | ( n1237 & ~n1588 ) ;
  assign n20315 = n1588 | n20314 ;
  assign n20316 = n931 | n1652 ;
  assign n20317 = n92 | n890 ;
  assign n20318 = ( n888 & n3514 ) | ( n888 & ~n20317 ) | ( n3514 & ~n20317 ) ;
  assign n20319 = n20317 | n20318 ;
  assign n20320 = ( ~n20315 & n20316 ) | ( ~n20315 & n20319 ) | ( n20316 & n20319 ) ;
  assign n20321 = n20315 | n20320 ;
  assign n20322 = ( ~n1822 & n2488 ) | ( ~n1822 & n20321 ) | ( n2488 & n20321 ) ;
  assign n20323 = n5723 | n6023 ;
  assign n20324 = n2324 | n2380 ;
  assign n20325 = n11079 | n20324 ;
  assign n20326 = n169 | n551 ;
  assign n20327 = n1711 | n2078 ;
  assign n20328 = ( n2274 & ~n20326 ) | ( n2274 & n20327 ) | ( ~n20326 & n20327 ) ;
  assign n20329 = ( ~n1538 & n20326 ) | ( ~n1538 & n20328 ) | ( n20326 & n20328 ) ;
  assign n20330 = n1538 | n20329 ;
  assign n20331 = ( ~n20323 & n20325 ) | ( ~n20323 & n20330 ) | ( n20325 & n20330 ) ;
  assign n20332 = n20323 | n20331 ;
  assign n20333 = n676 | n792 ;
  assign n20334 = ( n3983 & n4069 ) | ( n3983 & ~n5991 ) | ( n4069 & ~n5991 ) ;
  assign n20335 = n5991 | n20334 ;
  assign n20336 = ( n1889 & ~n20333 ) | ( n1889 & n20335 ) | ( ~n20333 & n20335 ) ;
  assign n20337 = n20333 | n20336 ;
  assign n20338 = ( ~n20321 & n20332 ) | ( ~n20321 & n20337 ) | ( n20332 & n20337 ) ;
  assign n20339 = ( ~n1822 & n20322 ) | ( ~n1822 & n20338 ) | ( n20322 & n20338 ) ;
  assign n20340 = n1822 | n20339 ;
  assign n20341 = n607 & n16053 ;
  assign n20342 = n1250 & ~n16051 ;
  assign n20343 = n20341 | n20342 ;
  assign n20344 = n606 & n16049 ;
  assign n20345 = ( n606 & n20343 ) | ( n606 & ~n20344 ) | ( n20343 & ~n20344 ) ;
  assign n20346 = n1248 & n16674 ;
  assign n20347 = ( n1248 & n20345 ) | ( n1248 & ~n20346 ) | ( n20345 & ~n20346 ) ;
  assign n20348 = ( n20209 & n20340 ) | ( n20209 & ~n20347 ) | ( n20340 & ~n20347 ) ;
  assign n20349 = ( ~n20209 & n20340 ) | ( ~n20209 & n20347 ) | ( n20340 & n20347 ) ;
  assign n20350 = ( ~n20340 & n20348 ) | ( ~n20340 & n20349 ) | ( n20348 & n20349 ) ;
  assign n20351 = n3800 & ~n16957 ;
  assign n20352 = n3799 & ~n16043 ;
  assign n20353 = n3700 & ~n16047 ;
  assign n20354 = n3802 & ~n16045 ;
  assign n20355 = n20353 | n20354 ;
  assign n20356 = ( ~n20351 & n20352 ) | ( ~n20351 & n20355 ) | ( n20352 & n20355 ) ;
  assign n20357 = ( ~x29 & n20351 ) | ( ~x29 & n20356 ) | ( n20351 & n20356 ) ;
  assign n20358 = ( n20351 & n20356 ) | ( n20351 & ~n20357 ) | ( n20356 & ~n20357 ) ;
  assign n20359 = ( x29 & n20357 ) | ( x29 & ~n20358 ) | ( n20357 & ~n20358 ) ;
  assign n20360 = ( n20219 & n20350 ) | ( n20219 & n20359 ) | ( n20350 & n20359 ) ;
  assign n20361 = ( n20219 & ~n20350 ) | ( n20219 & n20359 ) | ( ~n20350 & n20359 ) ;
  assign n20362 = ( n20350 & ~n20360 ) | ( n20350 & n20361 ) | ( ~n20360 & n20361 ) ;
  assign n20363 = n4202 & ~n17138 ;
  assign n20364 = n4201 & ~n16037 ;
  assign n20365 = n4200 & n16041 ;
  assign n20366 = n4345 & n16039 ;
  assign n20367 = n20365 | n20366 ;
  assign n20368 = ( ~n20363 & n20364 ) | ( ~n20363 & n20367 ) | ( n20364 & n20367 ) ;
  assign n20369 = ( ~x26 & n20363 ) | ( ~x26 & n20368 ) | ( n20363 & n20368 ) ;
  assign n20370 = ( n20363 & n20368 ) | ( n20363 & ~n20369 ) | ( n20368 & ~n20369 ) ;
  assign n20371 = ( x26 & n20369 ) | ( x26 & ~n20370 ) | ( n20369 & ~n20370 ) ;
  assign n20372 = ( n20231 & n20362 ) | ( n20231 & n20371 ) | ( n20362 & n20371 ) ;
  assign n20373 = ( n20231 & ~n20362 ) | ( n20231 & n20371 ) | ( ~n20362 & n20371 ) ;
  assign n20374 = ( n20362 & ~n20372 ) | ( n20362 & n20373 ) | ( ~n20372 & n20373 ) ;
  assign n20375 = n4713 & ~n17516 ;
  assign n20376 = n4712 & n16031 ;
  assign n20377 = n4709 & n16035 ;
  assign n20378 = n4792 & ~n16033 ;
  assign n20379 = n20377 | n20378 ;
  assign n20380 = ( ~n20375 & n20376 ) | ( ~n20375 & n20379 ) | ( n20376 & n20379 ) ;
  assign n20381 = ( ~x23 & n20375 ) | ( ~x23 & n20380 ) | ( n20375 & n20380 ) ;
  assign n20382 = ( n20375 & n20380 ) | ( n20375 & ~n20381 ) | ( n20380 & ~n20381 ) ;
  assign n20383 = ( x23 & n20381 ) | ( x23 & ~n20382 ) | ( n20381 & ~n20382 ) ;
  assign n20384 = ( n20234 & n20374 ) | ( n20234 & n20383 ) | ( n20374 & n20383 ) ;
  assign n20385 = ( n20234 & ~n20374 ) | ( n20234 & n20383 ) | ( ~n20374 & n20383 ) ;
  assign n20386 = ( n20374 & ~n20384 ) | ( n20374 & n20385 ) | ( ~n20384 & n20385 ) ;
  assign n20387 = n4974 & ~n17746 ;
  assign n20388 = n5398 & ~n16025 ;
  assign n20389 = n4973 & ~n16029 ;
  assign n20390 = n4972 & ~n16027 ;
  assign n20391 = n20389 | n20390 ;
  assign n20392 = ( ~n20387 & n20388 ) | ( ~n20387 & n20391 ) | ( n20388 & n20391 ) ;
  assign n20393 = ( ~x20 & n20387 ) | ( ~x20 & n20392 ) | ( n20387 & n20392 ) ;
  assign n20394 = ( n20387 & n20392 ) | ( n20387 & ~n20393 ) | ( n20392 & ~n20393 ) ;
  assign n20395 = ( x20 & n20393 ) | ( x20 & ~n20394 ) | ( n20393 & ~n20394 ) ;
  assign n20396 = ( n20246 & n20386 ) | ( n20246 & n20395 ) | ( n20386 & n20395 ) ;
  assign n20397 = ( n20246 & ~n20386 ) | ( n20246 & n20395 ) | ( ~n20386 & n20395 ) ;
  assign n20398 = ( n20386 & ~n20396 ) | ( n20386 & n20397 ) | ( ~n20396 & n20397 ) ;
  assign n20399 = n5508 & n18103 ;
  assign n20400 = n5507 & n16019 ;
  assign n20401 = n5504 & n16023 ;
  assign n20402 = n5666 & n16021 ;
  assign n20403 = n20401 | n20402 ;
  assign n20404 = ( ~n20399 & n20400 ) | ( ~n20399 & n20403 ) | ( n20400 & n20403 ) ;
  assign n20405 = ( ~x17 & n20399 ) | ( ~x17 & n20404 ) | ( n20399 & n20404 ) ;
  assign n20406 = ( n20399 & n20404 ) | ( n20399 & ~n20405 ) | ( n20404 & ~n20405 ) ;
  assign n20407 = ( x17 & n20405 ) | ( x17 & ~n20406 ) | ( n20405 & ~n20406 ) ;
  assign n20408 = ( n20258 & n20398 ) | ( n20258 & n20407 ) | ( n20398 & n20407 ) ;
  assign n20409 = ( n20258 & ~n20398 ) | ( n20258 & n20407 ) | ( ~n20398 & n20407 ) ;
  assign n20410 = ( n20398 & ~n20408 ) | ( n20398 & n20409 ) | ( ~n20408 & n20409 ) ;
  assign n20411 = n5966 & ~n18694 ;
  assign n20412 = n6464 & ~n16013 ;
  assign n20413 = n5970 & ~n16017 ;
  assign n20414 = n5969 & n16015 ;
  assign n20415 = n20413 | n20414 ;
  assign n20416 = ( ~n20411 & n20412 ) | ( ~n20411 & n20415 ) | ( n20412 & n20415 ) ;
  assign n20417 = ( ~x14 & n20411 ) | ( ~x14 & n20416 ) | ( n20411 & n20416 ) ;
  assign n20418 = ( n20411 & n20416 ) | ( n20411 & ~n20417 ) | ( n20416 & ~n20417 ) ;
  assign n20419 = ( x14 & n20417 ) | ( x14 & ~n20418 ) | ( n20417 & ~n20418 ) ;
  assign n20420 = ( n20270 & n20410 ) | ( n20270 & n20419 ) | ( n20410 & n20419 ) ;
  assign n20421 = ( n20270 & ~n20410 ) | ( n20270 & n20419 ) | ( ~n20410 & n20419 ) ;
  assign n20422 = ( n20410 & ~n20420 ) | ( n20410 & n20421 ) | ( ~n20420 & n20421 ) ;
  assign n20423 = n6584 & n19160 ;
  assign n20424 = n7022 & n19157 ;
  assign n20425 = n6588 & n16138 ;
  assign n20426 = n6587 & n18993 ;
  assign n20427 = n20425 | n20426 ;
  assign n20428 = ( ~n20423 & n20424 ) | ( ~n20423 & n20427 ) | ( n20424 & n20427 ) ;
  assign n20429 = ( ~x11 & n20423 ) | ( ~x11 & n20428 ) | ( n20423 & n20428 ) ;
  assign n20430 = ( n20423 & n20428 ) | ( n20423 & ~n20429 ) | ( n20428 & ~n20429 ) ;
  assign n20431 = ( x11 & n20429 ) | ( x11 & ~n20430 ) | ( n20429 & ~n20430 ) ;
  assign n20432 = ( n20282 & n20422 ) | ( n20282 & n20431 ) | ( n20422 & n20431 ) ;
  assign n20433 = ( n20282 & ~n20422 ) | ( n20282 & n20431 ) | ( ~n20422 & n20431 ) ;
  assign n20434 = ( n20422 & ~n20432 ) | ( n20422 & n20433 ) | ( ~n20432 & n20433 ) ;
  assign n20435 = n7300 & ~n19309 ;
  assign n20436 = ~x8 & n20435 ;
  assign n20437 = n20435 & ~n20436 ;
  assign n20438 = ( x8 & n20436 ) | ( x8 & ~n20437 ) | ( n20436 & ~n20437 ) ;
  assign n20439 = ( n20294 & n20434 ) | ( n20294 & n20438 ) | ( n20434 & n20438 ) ;
  assign n20440 = ( n20294 & ~n20434 ) | ( n20294 & n20438 ) | ( ~n20434 & n20438 ) ;
  assign n20441 = ( n20434 & ~n20439 ) | ( n20434 & n20440 ) | ( ~n20439 & n20440 ) ;
  assign n20442 = ( n20305 & n20308 ) | ( n20305 & n20441 ) | ( n20308 & n20441 ) ;
  assign n20443 = ( ~n20305 & n20308 ) | ( ~n20305 & n20441 ) | ( n20308 & n20441 ) ;
  assign n20444 = ( n20305 & ~n20442 ) | ( n20305 & n20443 ) | ( ~n20442 & n20443 ) ;
  assign n20445 = n20311 & n20444 ;
  assign n20446 = n20311 | n20444 ;
  assign n20447 = ~n20445 & n20446 ;
  assign n20448 = n170 | n328 ;
  assign n20449 = n124 | n20448 ;
  assign n20450 = ( n450 & n1145 ) | ( n450 & ~n20449 ) | ( n1145 & ~n20449 ) ;
  assign n20451 = n20449 | n20450 ;
  assign n20452 = ( n863 & n4510 ) | ( n863 & ~n20451 ) | ( n4510 & ~n20451 ) ;
  assign n20453 = n20451 | n20452 ;
  assign n20454 = n968 | n2638 ;
  assign n20455 = ( n943 & n2082 ) | ( n943 & ~n20454 ) | ( n2082 & ~n20454 ) ;
  assign n20456 = n20454 | n20455 ;
  assign n20457 = ( n3277 & n20453 ) | ( n3277 & ~n20456 ) | ( n20453 & ~n20456 ) ;
  assign n20458 = ~n20453 & n20457 ;
  assign n20459 = n890 | n5140 ;
  assign n20460 = ( n59 & n119 ) | ( n59 & n129 ) | ( n119 & n129 ) ;
  assign n20461 = ( n74 & n641 ) | ( n74 & ~n1170 ) | ( n641 & ~n1170 ) ;
  assign n20462 = n1170 | n20461 ;
  assign n20463 = ( ~n20459 & n20460 ) | ( ~n20459 & n20462 ) | ( n20460 & n20462 ) ;
  assign n20464 = n20459 | n20463 ;
  assign n20465 = n217 | n493 ;
  assign n20466 = ( n483 & n1346 ) | ( n483 & ~n20465 ) | ( n1346 & ~n20465 ) ;
  assign n20467 = n20465 | n20466 ;
  assign n20468 = ( n3053 & n3677 ) | ( n3053 & ~n10182 ) | ( n3677 & ~n10182 ) ;
  assign n20469 = n10182 | n20468 ;
  assign n20470 = ( n6179 & ~n20467 ) | ( n6179 & n20469 ) | ( ~n20467 & n20469 ) ;
  assign n20471 = n20467 | n20470 ;
  assign n20472 = ( ~n3906 & n3977 ) | ( ~n3906 & n20471 ) | ( n3977 & n20471 ) ;
  assign n20473 = ( n3906 & ~n20464 ) | ( n3906 & n20472 ) | ( ~n20464 & n20472 ) ;
  assign n20474 = n20464 | n20473 ;
  assign n20475 = ( n10597 & n20458 ) | ( n10597 & n20474 ) | ( n20458 & n20474 ) ;
  assign n20476 = n20458 & ~n20475 ;
  assign n20477 = ( n20340 & n20348 ) | ( n20340 & n20476 ) | ( n20348 & n20476 ) ;
  assign n20478 = ( ~n20340 & n20348 ) | ( ~n20340 & n20476 ) | ( n20348 & n20476 ) ;
  assign n20479 = ( n20340 & ~n20477 ) | ( n20340 & n20478 ) | ( ~n20477 & n20478 ) ;
  assign n20480 = n607 & ~n16051 ;
  assign n20481 = n1250 & ~n16049 ;
  assign n20482 = n20480 | n20481 ;
  assign n20483 = n606 & n16047 ;
  assign n20484 = ( n606 & n20482 ) | ( n606 & ~n20483 ) | ( n20482 & ~n20483 ) ;
  assign n20485 = n1248 & n16801 ;
  assign n20486 = ( n1248 & n20484 ) | ( n1248 & ~n20485 ) | ( n20484 & ~n20485 ) ;
  assign n20487 = ( n20360 & ~n20479 ) | ( n20360 & n20486 ) | ( ~n20479 & n20486 ) ;
  assign n20488 = ( n20360 & n20479 ) | ( n20360 & n20486 ) | ( n20479 & n20486 ) ;
  assign n20489 = ( n20479 & n20487 ) | ( n20479 & ~n20488 ) | ( n20487 & ~n20488 ) ;
  assign n20490 = n4202 & ~n17313 ;
  assign n20491 = n4201 & n16035 ;
  assign n20492 = n4200 & n16039 ;
  assign n20493 = n4345 & ~n16037 ;
  assign n20494 = n20492 | n20493 ;
  assign n20495 = ( ~n20490 & n20491 ) | ( ~n20490 & n20494 ) | ( n20491 & n20494 ) ;
  assign n20496 = ( ~x26 & n20490 ) | ( ~x26 & n20495 ) | ( n20490 & n20495 ) ;
  assign n20497 = ( n20490 & n20495 ) | ( n20490 & ~n20496 ) | ( n20495 & ~n20496 ) ;
  assign n20498 = ( x26 & n20496 ) | ( x26 & ~n20497 ) | ( n20496 & ~n20497 ) ;
  assign n20499 = n3800 & n16969 ;
  assign n20500 = n3799 & n16041 ;
  assign n20501 = n3700 & ~n16045 ;
  assign n20502 = n3802 & ~n16043 ;
  assign n20503 = n20501 | n20502 ;
  assign n20504 = ( ~n20499 & n20500 ) | ( ~n20499 & n20503 ) | ( n20500 & n20503 ) ;
  assign n20505 = ( ~x29 & n20499 ) | ( ~x29 & n20504 ) | ( n20499 & n20504 ) ;
  assign n20506 = ( n20499 & n20504 ) | ( n20499 & ~n20505 ) | ( n20504 & ~n20505 ) ;
  assign n20507 = ( x29 & n20505 ) | ( x29 & ~n20506 ) | ( n20505 & ~n20506 ) ;
  assign n20508 = ( ~n20489 & n20498 ) | ( ~n20489 & n20507 ) | ( n20498 & n20507 ) ;
  assign n20509 = ( n20498 & n20507 ) | ( n20498 & ~n20508 ) | ( n20507 & ~n20508 ) ;
  assign n20510 = ( n20489 & n20508 ) | ( n20489 & ~n20509 ) | ( n20508 & ~n20509 ) ;
  assign n20511 = n4713 & ~n17528 ;
  assign n20512 = n4712 & ~n16029 ;
  assign n20513 = n4709 & ~n16033 ;
  assign n20514 = n4792 & n16031 ;
  assign n20515 = n20513 | n20514 ;
  assign n20516 = ( ~n20511 & n20512 ) | ( ~n20511 & n20515 ) | ( n20512 & n20515 ) ;
  assign n20517 = ( ~x23 & n20511 ) | ( ~x23 & n20516 ) | ( n20511 & n20516 ) ;
  assign n20518 = ( n20511 & n20516 ) | ( n20511 & ~n20517 ) | ( n20516 & ~n20517 ) ;
  assign n20519 = ( x23 & n20517 ) | ( x23 & ~n20518 ) | ( n20517 & ~n20518 ) ;
  assign n20520 = ( n20372 & ~n20510 ) | ( n20372 & n20519 ) | ( ~n20510 & n20519 ) ;
  assign n20521 = ( n20372 & n20510 ) | ( n20372 & n20519 ) | ( n20510 & n20519 ) ;
  assign n20522 = ( n20510 & n20520 ) | ( n20510 & ~n20521 ) | ( n20520 & ~n20521 ) ;
  assign n20523 = n4974 & n17968 ;
  assign n20524 = n5398 & n16023 ;
  assign n20525 = n4973 & ~n16027 ;
  assign n20526 = n4972 & ~n16025 ;
  assign n20527 = n20525 | n20526 ;
  assign n20528 = ( ~n20523 & n20524 ) | ( ~n20523 & n20527 ) | ( n20524 & n20527 ) ;
  assign n20529 = ( ~x20 & n20523 ) | ( ~x20 & n20528 ) | ( n20523 & n20528 ) ;
  assign n20530 = ( n20523 & n20528 ) | ( n20523 & ~n20529 ) | ( n20528 & ~n20529 ) ;
  assign n20531 = ( x20 & n20529 ) | ( x20 & ~n20530 ) | ( n20529 & ~n20530 ) ;
  assign n20532 = ( n20384 & ~n20522 ) | ( n20384 & n20531 ) | ( ~n20522 & n20531 ) ;
  assign n20533 = ( n20384 & n20522 ) | ( n20384 & n20531 ) | ( n20522 & n20531 ) ;
  assign n20534 = ( n20522 & n20532 ) | ( n20522 & ~n20533 ) | ( n20532 & ~n20533 ) ;
  assign n20535 = n5508 & ~n18267 ;
  assign n20536 = n5507 & ~n16017 ;
  assign n20537 = n5504 & n16021 ;
  assign n20538 = n5666 & n16019 ;
  assign n20539 = n20537 | n20538 ;
  assign n20540 = ( ~n20535 & n20536 ) | ( ~n20535 & n20539 ) | ( n20536 & n20539 ) ;
  assign n20541 = ( ~x17 & n20535 ) | ( ~x17 & n20540 ) | ( n20535 & n20540 ) ;
  assign n20542 = ( n20535 & n20540 ) | ( n20535 & ~n20541 ) | ( n20540 & ~n20541 ) ;
  assign n20543 = ( x17 & n20541 ) | ( x17 & ~n20542 ) | ( n20541 & ~n20542 ) ;
  assign n20544 = ( n20396 & ~n20534 ) | ( n20396 & n20543 ) | ( ~n20534 & n20543 ) ;
  assign n20545 = ( n20396 & n20534 ) | ( n20396 & n20543 ) | ( n20534 & n20543 ) ;
  assign n20546 = ( n20534 & n20544 ) | ( n20534 & ~n20545 ) | ( n20544 & ~n20545 ) ;
  assign n20547 = n5966 & ~n16144 ;
  assign n20548 = n6464 & n16138 ;
  assign n20549 = n5970 & n16015 ;
  assign n20550 = n5969 & ~n16013 ;
  assign n20551 = n20549 | n20550 ;
  assign n20552 = ( ~n20547 & n20548 ) | ( ~n20547 & n20551 ) | ( n20548 & n20551 ) ;
  assign n20553 = ( ~x14 & n20547 ) | ( ~x14 & n20552 ) | ( n20547 & n20552 ) ;
  assign n20554 = ( n20547 & n20552 ) | ( n20547 & ~n20553 ) | ( n20552 & ~n20553 ) ;
  assign n20555 = ( x14 & n20553 ) | ( x14 & ~n20554 ) | ( n20553 & ~n20554 ) ;
  assign n20556 = ( n20408 & ~n20546 ) | ( n20408 & n20555 ) | ( ~n20546 & n20555 ) ;
  assign n20557 = ( n20408 & n20546 ) | ( n20408 & n20555 ) | ( n20546 & n20555 ) ;
  assign n20558 = ( n20546 & n20556 ) | ( n20546 & ~n20557 ) | ( n20556 & ~n20557 ) ;
  assign n20559 = n6584 & ~n19312 ;
  assign n20560 = n7022 & ~n19309 ;
  assign n20561 = n6588 & n18993 ;
  assign n20562 = n6587 & n19157 ;
  assign n20563 = n20561 | n20562 ;
  assign n20564 = ( ~n20559 & n20560 ) | ( ~n20559 & n20563 ) | ( n20560 & n20563 ) ;
  assign n20565 = ( ~x11 & n20559 ) | ( ~x11 & n20564 ) | ( n20559 & n20564 ) ;
  assign n20566 = ( n20559 & n20564 ) | ( n20559 & ~n20565 ) | ( n20564 & ~n20565 ) ;
  assign n20567 = ( x11 & n20565 ) | ( x11 & ~n20566 ) | ( n20565 & ~n20566 ) ;
  assign n20568 = ( n20420 & ~n20558 ) | ( n20420 & n20567 ) | ( ~n20558 & n20567 ) ;
  assign n20569 = ( n20420 & n20558 ) | ( n20420 & n20567 ) | ( n20558 & n20567 ) ;
  assign n20570 = ( n20558 & n20568 ) | ( n20558 & ~n20569 ) | ( n20568 & ~n20569 ) ;
  assign n20571 = ( x8 & n20432 ) | ( x8 & ~n20570 ) | ( n20432 & ~n20570 ) ;
  assign n20572 = ( x8 & n20432 ) | ( x8 & n20570 ) | ( n20432 & n20570 ) ;
  assign n20573 = ( n20570 & n20571 ) | ( n20570 & ~n20572 ) | ( n20571 & ~n20572 ) ;
  assign n20574 = ( n20439 & n20442 ) | ( n20439 & ~n20573 ) | ( n20442 & ~n20573 ) ;
  assign n20575 = ( n20439 & n20442 ) | ( n20439 & n20573 ) | ( n20442 & n20573 ) ;
  assign n20576 = ( n20573 & n20574 ) | ( n20573 & ~n20575 ) | ( n20574 & ~n20575 ) ;
  assign n20577 = n20445 & ~n20576 ;
  assign n20578 = n20445 & n20576 ;
  assign n20579 = ( n20576 & n20577 ) | ( n20576 & ~n20578 ) | ( n20577 & ~n20578 ) ;
  assign n20580 = n6584 & ~n19472 ;
  assign n20581 = n6588 & n19157 ;
  assign n20582 = n6587 & ~n19309 ;
  assign n20583 = n20581 | n20582 ;
  assign n20584 = ~n20580 & n20583 ;
  assign n20585 = ( ~x11 & n20580 ) | ( ~x11 & n20584 ) | ( n20580 & n20584 ) ;
  assign n20586 = ( n20580 & n20584 ) | ( n20580 & ~n20585 ) | ( n20584 & ~n20585 ) ;
  assign n20587 = ( x11 & n20585 ) | ( x11 & ~n20586 ) | ( n20585 & ~n20586 ) ;
  assign n20588 = n5508 & ~n18416 ;
  assign n20589 = n5507 & n16015 ;
  assign n20590 = n5504 & n16019 ;
  assign n20591 = n5666 & ~n16017 ;
  assign n20592 = n20590 | n20591 ;
  assign n20593 = ( ~n20588 & n20589 ) | ( ~n20588 & n20592 ) | ( n20589 & n20592 ) ;
  assign n20594 = ( ~x17 & n20588 ) | ( ~x17 & n20593 ) | ( n20588 & n20593 ) ;
  assign n20595 = ( n20588 & n20593 ) | ( n20588 & ~n20594 ) | ( n20593 & ~n20594 ) ;
  assign n20596 = ( x17 & n20594 ) | ( x17 & ~n20595 ) | ( n20594 & ~n20595 ) ;
  assign n20597 = n113 | n959 ;
  assign n20598 = n2167 | n20597 ;
  assign n20599 = n928 | n1528 ;
  assign n20600 = n577 | n990 ;
  assign n20601 = ( n10132 & ~n20599 ) | ( n10132 & n20600 ) | ( ~n20599 & n20600 ) ;
  assign n20602 = n20599 | n20601 ;
  assign n20603 = ( n1700 & ~n2457 ) | ( n1700 & n10590 ) | ( ~n2457 & n10590 ) ;
  assign n20604 = n2457 | n20603 ;
  assign n20605 = ( ~n20598 & n20602 ) | ( ~n20598 & n20604 ) | ( n20602 & n20604 ) ;
  assign n20606 = n20598 | n20605 ;
  assign n20607 = n1643 | n2940 ;
  assign n20608 = ( n3497 & n20606 ) | ( n3497 & ~n20607 ) | ( n20606 & ~n20607 ) ;
  assign n20609 = ~n20606 & n20608 ;
  assign n20610 = ( x8 & ~n20340 ) | ( x8 & n20609 ) | ( ~n20340 & n20609 ) ;
  assign n20611 = ( x8 & n20609 ) | ( x8 & ~n20610 ) | ( n20609 & ~n20610 ) ;
  assign n20612 = ( n20340 & n20610 ) | ( n20340 & ~n20611 ) | ( n20610 & ~n20611 ) ;
  assign n20613 = n607 & ~n16049 ;
  assign n20614 = n1250 & ~n16047 ;
  assign n20615 = n20613 | n20614 ;
  assign n20616 = n606 & n16045 ;
  assign n20617 = ( n606 & n20615 ) | ( n606 & ~n20616 ) | ( n20615 & ~n20616 ) ;
  assign n20618 = n1248 & n16876 ;
  assign n20619 = ( n1248 & n20617 ) | ( n1248 & ~n20618 ) | ( n20617 & ~n20618 ) ;
  assign n20620 = ( ~n20477 & n20612 ) | ( ~n20477 & n20619 ) | ( n20612 & n20619 ) ;
  assign n20621 = ( n20612 & n20619 ) | ( n20612 & ~n20620 ) | ( n20619 & ~n20620 ) ;
  assign n20622 = ( n20477 & n20620 ) | ( n20477 & ~n20621 ) | ( n20620 & ~n20621 ) ;
  assign n20623 = n3800 & ~n17051 ;
  assign n20624 = n3799 & n16039 ;
  assign n20625 = n3700 & ~n16043 ;
  assign n20626 = n3802 & n16041 ;
  assign n20627 = n20625 | n20626 ;
  assign n20628 = ( ~n20623 & n20624 ) | ( ~n20623 & n20627 ) | ( n20624 & n20627 ) ;
  assign n20629 = ( ~x29 & n20623 ) | ( ~x29 & n20628 ) | ( n20623 & n20628 ) ;
  assign n20630 = ( n20623 & n20628 ) | ( n20623 & ~n20629 ) | ( n20628 & ~n20629 ) ;
  assign n20631 = ( x29 & n20629 ) | ( x29 & ~n20630 ) | ( n20629 & ~n20630 ) ;
  assign n20632 = ( n20487 & ~n20622 ) | ( n20487 & n20631 ) | ( ~n20622 & n20631 ) ;
  assign n20633 = ( n20487 & n20622 ) | ( n20487 & n20631 ) | ( n20622 & n20631 ) ;
  assign n20634 = ( n20622 & n20632 ) | ( n20622 & ~n20633 ) | ( n20632 & ~n20633 ) ;
  assign n20635 = n4202 & ~n17412 ;
  assign n20636 = n4201 & ~n16033 ;
  assign n20637 = n4200 & ~n16037 ;
  assign n20638 = n4345 & n16035 ;
  assign n20639 = n20637 | n20638 ;
  assign n20640 = ( ~n20635 & n20636 ) | ( ~n20635 & n20639 ) | ( n20636 & n20639 ) ;
  assign n20641 = ( ~x26 & n20635 ) | ( ~x26 & n20640 ) | ( n20635 & n20640 ) ;
  assign n20642 = ( n20635 & n20640 ) | ( n20635 & ~n20641 ) | ( n20640 & ~n20641 ) ;
  assign n20643 = ( x26 & n20641 ) | ( x26 & ~n20642 ) | ( n20641 & ~n20642 ) ;
  assign n20644 = ( n20508 & ~n20634 ) | ( n20508 & n20643 ) | ( ~n20634 & n20643 ) ;
  assign n20645 = ( n20508 & n20634 ) | ( n20508 & n20643 ) | ( n20634 & n20643 ) ;
  assign n20646 = ( n20634 & n20644 ) | ( n20634 & ~n20645 ) | ( n20644 & ~n20645 ) ;
  assign n20647 = n4713 & n17634 ;
  assign n20648 = n4712 & ~n16027 ;
  assign n20649 = n4709 & n16031 ;
  assign n20650 = n4792 & ~n16029 ;
  assign n20651 = n20649 | n20650 ;
  assign n20652 = ( ~n20647 & n20648 ) | ( ~n20647 & n20651 ) | ( n20648 & n20651 ) ;
  assign n20653 = ( ~x23 & n20647 ) | ( ~x23 & n20652 ) | ( n20647 & n20652 ) ;
  assign n20654 = ( n20647 & n20652 ) | ( n20647 & ~n20653 ) | ( n20652 & ~n20653 ) ;
  assign n20655 = ( x23 & n20653 ) | ( x23 & ~n20654 ) | ( n20653 & ~n20654 ) ;
  assign n20656 = ( n20520 & ~n20646 ) | ( n20520 & n20655 ) | ( ~n20646 & n20655 ) ;
  assign n20657 = ( n20520 & n20646 ) | ( n20520 & n20655 ) | ( n20646 & n20655 ) ;
  assign n20658 = ( n20646 & n20656 ) | ( n20646 & ~n20657 ) | ( n20656 & ~n20657 ) ;
  assign n20659 = n4974 & ~n18091 ;
  assign n20660 = n5398 & n16021 ;
  assign n20661 = n4973 & ~n16025 ;
  assign n20662 = n4972 & n16023 ;
  assign n20663 = n20661 | n20662 ;
  assign n20664 = ( ~n20659 & n20660 ) | ( ~n20659 & n20663 ) | ( n20660 & n20663 ) ;
  assign n20665 = ( ~x20 & n20659 ) | ( ~x20 & n20664 ) | ( n20659 & n20664 ) ;
  assign n20666 = ( n20659 & n20664 ) | ( n20659 & ~n20665 ) | ( n20664 & ~n20665 ) ;
  assign n20667 = ( x20 & n20665 ) | ( x20 & ~n20666 ) | ( n20665 & ~n20666 ) ;
  assign n20668 = ( n20532 & ~n20658 ) | ( n20532 & n20667 ) | ( ~n20658 & n20667 ) ;
  assign n20669 = ( n20532 & n20658 ) | ( n20532 & n20667 ) | ( n20658 & n20667 ) ;
  assign n20670 = ( n20658 & n20668 ) | ( n20658 & ~n20669 ) | ( n20668 & ~n20669 ) ;
  assign n20671 = ( n20544 & n20596 ) | ( n20544 & ~n20670 ) | ( n20596 & ~n20670 ) ;
  assign n20672 = ( ~n20544 & n20596 ) | ( ~n20544 & n20670 ) | ( n20596 & n20670 ) ;
  assign n20673 = ( ~n20596 & n20671 ) | ( ~n20596 & n20672 ) | ( n20671 & n20672 ) ;
  assign n20674 = n5966 & n18996 ;
  assign n20675 = n6464 & n18993 ;
  assign n20676 = n5970 & ~n16013 ;
  assign n20677 = n5969 & n16138 ;
  assign n20678 = n20676 | n20677 ;
  assign n20679 = ( ~n20674 & n20675 ) | ( ~n20674 & n20678 ) | ( n20675 & n20678 ) ;
  assign n20680 = ( ~x14 & n20674 ) | ( ~x14 & n20679 ) | ( n20674 & n20679 ) ;
  assign n20681 = ( n20674 & n20679 ) | ( n20674 & ~n20680 ) | ( n20679 & ~n20680 ) ;
  assign n20682 = ( x14 & n20680 ) | ( x14 & ~n20681 ) | ( n20680 & ~n20681 ) ;
  assign n20683 = ( n20556 & ~n20673 ) | ( n20556 & n20682 ) | ( ~n20673 & n20682 ) ;
  assign n20684 = ( n20556 & n20673 ) | ( n20556 & n20682 ) | ( n20673 & n20682 ) ;
  assign n20685 = ( n20673 & n20683 ) | ( n20673 & ~n20684 ) | ( n20683 & ~n20684 ) ;
  assign n20686 = ( n20568 & n20587 ) | ( n20568 & ~n20685 ) | ( n20587 & ~n20685 ) ;
  assign n20687 = ( ~n20568 & n20587 ) | ( ~n20568 & n20685 ) | ( n20587 & n20685 ) ;
  assign n20688 = ( ~n20587 & n20686 ) | ( ~n20587 & n20687 ) | ( n20686 & n20687 ) ;
  assign n20689 = ( n20571 & n20574 ) | ( n20571 & ~n20688 ) | ( n20574 & ~n20688 ) ;
  assign n20690 = ( n20571 & n20574 ) | ( n20571 & n20688 ) | ( n20574 & n20688 ) ;
  assign n20691 = ( n20688 & n20689 ) | ( n20688 & ~n20690 ) | ( n20689 & ~n20690 ) ;
  assign n20692 = n20577 & ~n20691 ;
  assign n20693 = ~n20577 & n20691 ;
  assign n20694 = n20692 | n20693 ;
  assign n20695 = n3800 & ~n17138 ;
  assign n20696 = n3799 & ~n16037 ;
  assign n20697 = n3700 & n16041 ;
  assign n20698 = n3802 & n16039 ;
  assign n20699 = n20697 | n20698 ;
  assign n20700 = ( ~n20695 & n20696 ) | ( ~n20695 & n20699 ) | ( n20696 & n20699 ) ;
  assign n20701 = ( ~x29 & n20695 ) | ( ~x29 & n20700 ) | ( n20695 & n20700 ) ;
  assign n20702 = ( n20695 & n20700 ) | ( n20695 & ~n20701 ) | ( n20700 & ~n20701 ) ;
  assign n20703 = ( x29 & n20701 ) | ( x29 & ~n20702 ) | ( n20701 & ~n20702 ) ;
  assign n20704 = n444 | n549 ;
  assign n20705 = ( n505 & n2516 ) | ( n505 & ~n20704 ) | ( n2516 & ~n20704 ) ;
  assign n20706 = n20704 | n20705 ;
  assign n20707 = ( n731 & ~n4870 ) | ( n731 & n11976 ) | ( ~n4870 & n11976 ) ;
  assign n20708 = n4870 | n20707 ;
  assign n20709 = n118 | n3473 ;
  assign n20710 = ( n884 & n11535 ) | ( n884 & ~n20709 ) | ( n11535 & ~n20709 ) ;
  assign n20711 = n20709 | n20710 ;
  assign n20712 = ( ~n20706 & n20708 ) | ( ~n20706 & n20711 ) | ( n20708 & n20711 ) ;
  assign n20713 = n20706 | n20712 ;
  assign n20714 = ~n1362 & n2679 ;
  assign n20715 = ( ~n10976 & n20713 ) | ( ~n10976 & n20714 ) | ( n20713 & n20714 ) ;
  assign n20716 = ~n20713 & n20715 ;
  assign n20717 = n607 & ~n16047 ;
  assign n20718 = n1250 & ~n16045 ;
  assign n20719 = n20717 | n20718 ;
  assign n20720 = n606 & n16043 ;
  assign n20721 = ( n606 & n20719 ) | ( n606 & ~n20720 ) | ( n20719 & ~n20720 ) ;
  assign n20722 = n1248 & n16957 ;
  assign n20723 = ( n1248 & n20721 ) | ( n1248 & ~n20722 ) | ( n20721 & ~n20722 ) ;
  assign n20724 = ( ~n20610 & n20716 ) | ( ~n20610 & n20723 ) | ( n20716 & n20723 ) ;
  assign n20725 = ( n20716 & n20723 ) | ( n20716 & ~n20724 ) | ( n20723 & ~n20724 ) ;
  assign n20726 = ( n20610 & n20724 ) | ( n20610 & ~n20725 ) | ( n20724 & ~n20725 ) ;
  assign n20727 = ( n20620 & n20703 ) | ( n20620 & ~n20726 ) | ( n20703 & ~n20726 ) ;
  assign n20728 = ( ~n20620 & n20703 ) | ( ~n20620 & n20726 ) | ( n20703 & n20726 ) ;
  assign n20729 = ( ~n20703 & n20727 ) | ( ~n20703 & n20728 ) | ( n20727 & n20728 ) ;
  assign n20730 = n4202 & ~n17516 ;
  assign n20731 = n4201 & n16031 ;
  assign n20732 = n4200 & n16035 ;
  assign n20733 = n4345 & ~n16033 ;
  assign n20734 = n20732 | n20733 ;
  assign n20735 = ( ~n20730 & n20731 ) | ( ~n20730 & n20734 ) | ( n20731 & n20734 ) ;
  assign n20736 = ( ~x26 & n20730 ) | ( ~x26 & n20735 ) | ( n20730 & n20735 ) ;
  assign n20737 = ( n20730 & n20735 ) | ( n20730 & ~n20736 ) | ( n20735 & ~n20736 ) ;
  assign n20738 = ( x26 & n20736 ) | ( x26 & ~n20737 ) | ( n20736 & ~n20737 ) ;
  assign n20739 = ( n20632 & ~n20729 ) | ( n20632 & n20738 ) | ( ~n20729 & n20738 ) ;
  assign n20740 = ( n20632 & n20729 ) | ( n20632 & n20738 ) | ( n20729 & n20738 ) ;
  assign n20741 = ( n20729 & n20739 ) | ( n20729 & ~n20740 ) | ( n20739 & ~n20740 ) ;
  assign n20742 = n4713 & ~n17746 ;
  assign n20743 = n4712 & ~n16025 ;
  assign n20744 = n4709 & ~n16029 ;
  assign n20745 = n4792 & ~n16027 ;
  assign n20746 = n20744 | n20745 ;
  assign n20747 = ( ~n20742 & n20743 ) | ( ~n20742 & n20746 ) | ( n20743 & n20746 ) ;
  assign n20748 = ( ~x23 & n20742 ) | ( ~x23 & n20747 ) | ( n20742 & n20747 ) ;
  assign n20749 = ( n20742 & n20747 ) | ( n20742 & ~n20748 ) | ( n20747 & ~n20748 ) ;
  assign n20750 = ( x23 & n20748 ) | ( x23 & ~n20749 ) | ( n20748 & ~n20749 ) ;
  assign n20751 = ( n20644 & ~n20741 ) | ( n20644 & n20750 ) | ( ~n20741 & n20750 ) ;
  assign n20752 = ( n20644 & n20741 ) | ( n20644 & n20750 ) | ( n20741 & n20750 ) ;
  assign n20753 = ( n20741 & n20751 ) | ( n20741 & ~n20752 ) | ( n20751 & ~n20752 ) ;
  assign n20754 = n4974 & n18103 ;
  assign n20755 = n5398 & n16019 ;
  assign n20756 = n4973 & n16023 ;
  assign n20757 = n4972 & n16021 ;
  assign n20758 = n20756 | n20757 ;
  assign n20759 = ( ~n20754 & n20755 ) | ( ~n20754 & n20758 ) | ( n20755 & n20758 ) ;
  assign n20760 = ( ~x20 & n20754 ) | ( ~x20 & n20759 ) | ( n20754 & n20759 ) ;
  assign n20761 = ( n20754 & n20759 ) | ( n20754 & ~n20760 ) | ( n20759 & ~n20760 ) ;
  assign n20762 = ( x20 & n20760 ) | ( x20 & ~n20761 ) | ( n20760 & ~n20761 ) ;
  assign n20763 = ( n20656 & ~n20753 ) | ( n20656 & n20762 ) | ( ~n20753 & n20762 ) ;
  assign n20764 = ( n20656 & n20753 ) | ( n20656 & n20762 ) | ( n20753 & n20762 ) ;
  assign n20765 = ( n20753 & n20763 ) | ( n20753 & ~n20764 ) | ( n20763 & ~n20764 ) ;
  assign n20766 = n5508 & ~n18694 ;
  assign n20767 = n5507 & ~n16013 ;
  assign n20768 = n5504 & ~n16017 ;
  assign n20769 = n5666 & n16015 ;
  assign n20770 = n20768 | n20769 ;
  assign n20771 = ( ~n20766 & n20767 ) | ( ~n20766 & n20770 ) | ( n20767 & n20770 ) ;
  assign n20772 = ( ~x17 & n20766 ) | ( ~x17 & n20771 ) | ( n20766 & n20771 ) ;
  assign n20773 = ( n20766 & n20771 ) | ( n20766 & ~n20772 ) | ( n20771 & ~n20772 ) ;
  assign n20774 = ( x17 & n20772 ) | ( x17 & ~n20773 ) | ( n20772 & ~n20773 ) ;
  assign n20775 = ( n20668 & ~n20765 ) | ( n20668 & n20774 ) | ( ~n20765 & n20774 ) ;
  assign n20776 = ( n20668 & n20765 ) | ( n20668 & n20774 ) | ( n20765 & n20774 ) ;
  assign n20777 = ( n20765 & n20775 ) | ( n20765 & ~n20776 ) | ( n20775 & ~n20776 ) ;
  assign n20778 = n5966 & n19160 ;
  assign n20779 = n6464 & n19157 ;
  assign n20780 = n5970 & n16138 ;
  assign n20781 = n5969 & n18993 ;
  assign n20782 = n20780 | n20781 ;
  assign n20783 = ( ~n20778 & n20779 ) | ( ~n20778 & n20782 ) | ( n20779 & n20782 ) ;
  assign n20784 = ( ~x14 & n20778 ) | ( ~x14 & n20783 ) | ( n20778 & n20783 ) ;
  assign n20785 = ( n20778 & n20783 ) | ( n20778 & ~n20784 ) | ( n20783 & ~n20784 ) ;
  assign n20786 = ( x14 & n20784 ) | ( x14 & ~n20785 ) | ( n20784 & ~n20785 ) ;
  assign n20787 = ( n20671 & ~n20777 ) | ( n20671 & n20786 ) | ( ~n20777 & n20786 ) ;
  assign n20788 = ( n20671 & n20777 ) | ( n20671 & n20786 ) | ( n20777 & n20786 ) ;
  assign n20789 = ( n20777 & n20787 ) | ( n20777 & ~n20788 ) | ( n20787 & ~n20788 ) ;
  assign n20790 = n6588 & ~n19309 ;
  assign n20791 = ~x11 & n20790 ;
  assign n20792 = n20790 & ~n20791 ;
  assign n20793 = ( x11 & n20791 ) | ( x11 & ~n20792 ) | ( n20791 & ~n20792 ) ;
  assign n20794 = ( n20683 & ~n20789 ) | ( n20683 & n20793 ) | ( ~n20789 & n20793 ) ;
  assign n20795 = ( n20683 & n20789 ) | ( n20683 & n20793 ) | ( n20789 & n20793 ) ;
  assign n20796 = ( n20789 & n20794 ) | ( n20789 & ~n20795 ) | ( n20794 & ~n20795 ) ;
  assign n20797 = ( n20686 & n20689 ) | ( n20686 & ~n20796 ) | ( n20689 & ~n20796 ) ;
  assign n20798 = ( n20686 & n20689 ) | ( n20686 & n20796 ) | ( n20689 & n20796 ) ;
  assign n20799 = ( n20796 & n20797 ) | ( n20796 & ~n20798 ) | ( n20797 & ~n20798 ) ;
  assign n20800 = n20692 & ~n20799 ;
  assign n20801 = n20692 & n20799 ;
  assign n20802 = ( n20799 & n20800 ) | ( n20799 & ~n20801 ) | ( n20800 & ~n20801 ) ;
  assign n20803 = n773 | n2093 ;
  assign n20804 = ( n2362 & n3523 ) | ( n2362 & ~n20803 ) | ( n3523 & ~n20803 ) ;
  assign n20805 = n20803 | n20804 ;
  assign n20806 = n1005 | n1861 ;
  assign n20807 = ( n3564 & n10144 ) | ( n3564 & ~n20806 ) | ( n10144 & ~n20806 ) ;
  assign n20808 = n20806 | n20807 ;
  assign n20809 = ( n83 & n122 ) | ( n83 & n865 ) | ( n122 & n865 ) ;
  assign n20810 = ( n507 & n1496 ) | ( n507 & ~n20809 ) | ( n1496 & ~n20809 ) ;
  assign n20811 = n20809 | n20810 ;
  assign n20812 = ( ~n20805 & n20808 ) | ( ~n20805 & n20811 ) | ( n20808 & n20811 ) ;
  assign n20813 = n20805 | n20812 ;
  assign n20814 = ( n5220 & n10586 ) | ( n5220 & ~n11517 ) | ( n10586 & ~n11517 ) ;
  assign n20815 = n11517 | n20814 ;
  assign n20816 = ( n20332 & ~n20813 ) | ( n20332 & n20815 ) | ( ~n20813 & n20815 ) ;
  assign n20817 = n20813 | n20816 ;
  assign n20818 = ( n20716 & n20724 ) | ( n20716 & n20817 ) | ( n20724 & n20817 ) ;
  assign n20819 = ( n20716 & ~n20724 ) | ( n20716 & n20817 ) | ( ~n20724 & n20817 ) ;
  assign n20820 = ( n20724 & ~n20818 ) | ( n20724 & n20819 ) | ( ~n20818 & n20819 ) ;
  assign n20821 = n3800 & ~n17313 ;
  assign n20822 = n3799 & n16035 ;
  assign n20823 = n3700 & n16039 ;
  assign n20824 = n3802 & ~n16037 ;
  assign n20825 = n20823 | n20824 ;
  assign n20826 = ( ~n20821 & n20822 ) | ( ~n20821 & n20825 ) | ( n20822 & n20825 ) ;
  assign n20827 = ( ~x29 & n20821 ) | ( ~x29 & n20826 ) | ( n20821 & n20826 ) ;
  assign n20828 = ( n20821 & n20826 ) | ( n20821 & ~n20827 ) | ( n20826 & ~n20827 ) ;
  assign n20829 = ( x29 & n20827 ) | ( x29 & ~n20828 ) | ( n20827 & ~n20828 ) ;
  assign n20830 = n607 & ~n16045 ;
  assign n20831 = n1250 & ~n16043 ;
  assign n20832 = n20830 | n20831 ;
  assign n20833 = n606 & ~n16041 ;
  assign n20834 = ( n606 & n20832 ) | ( n606 & ~n20833 ) | ( n20832 & ~n20833 ) ;
  assign n20835 = n1248 & ~n16969 ;
  assign n20836 = ( n1248 & n20834 ) | ( n1248 & ~n20835 ) | ( n20834 & ~n20835 ) ;
  assign n20837 = ( n20820 & n20829 ) | ( n20820 & n20836 ) | ( n20829 & n20836 ) ;
  assign n20838 = ( ~n20820 & n20829 ) | ( ~n20820 & n20836 ) | ( n20829 & n20836 ) ;
  assign n20839 = ( n20820 & ~n20837 ) | ( n20820 & n20838 ) | ( ~n20837 & n20838 ) ;
  assign n20840 = n4202 & ~n17528 ;
  assign n20841 = n4201 & ~n16029 ;
  assign n20842 = n4200 & ~n16033 ;
  assign n20843 = n4345 & n16031 ;
  assign n20844 = n20842 | n20843 ;
  assign n20845 = ( ~n20840 & n20841 ) | ( ~n20840 & n20844 ) | ( n20841 & n20844 ) ;
  assign n20846 = ( ~x26 & n20840 ) | ( ~x26 & n20845 ) | ( n20840 & n20845 ) ;
  assign n20847 = ( n20840 & n20845 ) | ( n20840 & ~n20846 ) | ( n20845 & ~n20846 ) ;
  assign n20848 = ( x26 & n20846 ) | ( x26 & ~n20847 ) | ( n20846 & ~n20847 ) ;
  assign n20849 = ( n20727 & n20839 ) | ( n20727 & n20848 ) | ( n20839 & n20848 ) ;
  assign n20850 = ( n20727 & ~n20839 ) | ( n20727 & n20848 ) | ( ~n20839 & n20848 ) ;
  assign n20851 = ( n20839 & ~n20849 ) | ( n20839 & n20850 ) | ( ~n20849 & n20850 ) ;
  assign n20852 = n4713 & n17968 ;
  assign n20853 = n4712 & n16023 ;
  assign n20854 = n4709 & ~n16027 ;
  assign n20855 = n4792 & ~n16025 ;
  assign n20856 = n20854 | n20855 ;
  assign n20857 = ( ~n20852 & n20853 ) | ( ~n20852 & n20856 ) | ( n20853 & n20856 ) ;
  assign n20858 = ( ~x23 & n20852 ) | ( ~x23 & n20857 ) | ( n20852 & n20857 ) ;
  assign n20859 = ( n20852 & n20857 ) | ( n20852 & ~n20858 ) | ( n20857 & ~n20858 ) ;
  assign n20860 = ( x23 & n20858 ) | ( x23 & ~n20859 ) | ( n20858 & ~n20859 ) ;
  assign n20861 = ( n20739 & n20851 ) | ( n20739 & n20860 ) | ( n20851 & n20860 ) ;
  assign n20862 = ( n20739 & ~n20851 ) | ( n20739 & n20860 ) | ( ~n20851 & n20860 ) ;
  assign n20863 = ( n20851 & ~n20861 ) | ( n20851 & n20862 ) | ( ~n20861 & n20862 ) ;
  assign n20864 = n4974 & ~n18267 ;
  assign n20865 = n5398 & ~n16017 ;
  assign n20866 = n4973 & n16021 ;
  assign n20867 = n4972 & n16019 ;
  assign n20868 = n20866 | n20867 ;
  assign n20869 = ( ~n20864 & n20865 ) | ( ~n20864 & n20868 ) | ( n20865 & n20868 ) ;
  assign n20870 = ( ~x20 & n20864 ) | ( ~x20 & n20869 ) | ( n20864 & n20869 ) ;
  assign n20871 = ( n20864 & n20869 ) | ( n20864 & ~n20870 ) | ( n20869 & ~n20870 ) ;
  assign n20872 = ( x20 & n20870 ) | ( x20 & ~n20871 ) | ( n20870 & ~n20871 ) ;
  assign n20873 = ( n20751 & n20863 ) | ( n20751 & n20872 ) | ( n20863 & n20872 ) ;
  assign n20874 = ( n20751 & ~n20863 ) | ( n20751 & n20872 ) | ( ~n20863 & n20872 ) ;
  assign n20875 = ( n20863 & ~n20873 ) | ( n20863 & n20874 ) | ( ~n20873 & n20874 ) ;
  assign n20876 = n5508 & ~n16144 ;
  assign n20877 = n5507 & n16138 ;
  assign n20878 = n5504 & n16015 ;
  assign n20879 = n5666 & ~n16013 ;
  assign n20880 = n20878 | n20879 ;
  assign n20881 = ( ~n20876 & n20877 ) | ( ~n20876 & n20880 ) | ( n20877 & n20880 ) ;
  assign n20882 = ( ~x17 & n20876 ) | ( ~x17 & n20881 ) | ( n20876 & n20881 ) ;
  assign n20883 = ( n20876 & n20881 ) | ( n20876 & ~n20882 ) | ( n20881 & ~n20882 ) ;
  assign n20884 = ( x17 & n20882 ) | ( x17 & ~n20883 ) | ( n20882 & ~n20883 ) ;
  assign n20885 = ( n20763 & n20875 ) | ( n20763 & n20884 ) | ( n20875 & n20884 ) ;
  assign n20886 = ( n20763 & ~n20875 ) | ( n20763 & n20884 ) | ( ~n20875 & n20884 ) ;
  assign n20887 = ( n20875 & ~n20885 ) | ( n20875 & n20886 ) | ( ~n20885 & n20886 ) ;
  assign n20888 = n5966 & ~n19312 ;
  assign n20889 = n6464 & ~n19309 ;
  assign n20890 = n5970 & n18993 ;
  assign n20891 = n5969 & n19157 ;
  assign n20892 = n20890 | n20891 ;
  assign n20893 = ( ~n20888 & n20889 ) | ( ~n20888 & n20892 ) | ( n20889 & n20892 ) ;
  assign n20894 = ( ~x14 & n20888 ) | ( ~x14 & n20893 ) | ( n20888 & n20893 ) ;
  assign n20895 = ( n20888 & n20893 ) | ( n20888 & ~n20894 ) | ( n20893 & ~n20894 ) ;
  assign n20896 = ( x14 & n20894 ) | ( x14 & ~n20895 ) | ( n20894 & ~n20895 ) ;
  assign n20897 = ( n20775 & n20887 ) | ( n20775 & n20896 ) | ( n20887 & n20896 ) ;
  assign n20898 = ( n20775 & ~n20887 ) | ( n20775 & n20896 ) | ( ~n20887 & n20896 ) ;
  assign n20899 = ( n20887 & ~n20897 ) | ( n20887 & n20898 ) | ( ~n20897 & n20898 ) ;
  assign n20900 = ( x11 & n20787 ) | ( x11 & n20899 ) | ( n20787 & n20899 ) ;
  assign n20901 = ( ~x11 & n20787 ) | ( ~x11 & n20899 ) | ( n20787 & n20899 ) ;
  assign n20902 = ( x11 & ~n20900 ) | ( x11 & n20901 ) | ( ~n20900 & n20901 ) ;
  assign n20903 = ( n20794 & n20797 ) | ( n20794 & n20902 ) | ( n20797 & n20902 ) ;
  assign n20904 = ( n20794 & ~n20797 ) | ( n20794 & n20902 ) | ( ~n20797 & n20902 ) ;
  assign n20905 = ( n20797 & ~n20903 ) | ( n20797 & n20904 ) | ( ~n20903 & n20904 ) ;
  assign n20906 = n20800 & n20905 ;
  assign n20907 = n20800 | n20905 ;
  assign n20908 = ~n20906 & n20907 ;
  assign n20909 = n5966 & ~n19472 ;
  assign n20910 = n5970 & n19157 ;
  assign n20911 = n5969 & ~n19309 ;
  assign n20912 = n20910 | n20911 ;
  assign n20913 = ~n20909 & n20912 ;
  assign n20914 = ( ~x14 & n20909 ) | ( ~x14 & n20913 ) | ( n20909 & n20913 ) ;
  assign n20915 = ( n20909 & n20913 ) | ( n20909 & ~n20914 ) | ( n20913 & ~n20914 ) ;
  assign n20916 = ( x14 & n20914 ) | ( x14 & ~n20915 ) | ( n20914 & ~n20915 ) ;
  assign n20917 = n4974 & ~n18416 ;
  assign n20918 = n5398 & n16015 ;
  assign n20919 = n4973 & n16019 ;
  assign n20920 = n4972 & ~n16017 ;
  assign n20921 = n20919 | n20920 ;
  assign n20922 = ( ~n20917 & n20918 ) | ( ~n20917 & n20921 ) | ( n20918 & n20921 ) ;
  assign n20923 = ( ~x20 & n20917 ) | ( ~x20 & n20922 ) | ( n20917 & n20922 ) ;
  assign n20924 = ( n20917 & n20922 ) | ( n20917 & ~n20923 ) | ( n20922 & ~n20923 ) ;
  assign n20925 = ( x20 & n20923 ) | ( x20 & ~n20924 ) | ( n20923 & ~n20924 ) ;
  assign n20926 = n402 | n824 ;
  assign n20927 = n135 | n20926 ;
  assign n20928 = n287 | n1512 ;
  assign n20929 = ( ~n5019 & n10215 ) | ( ~n5019 & n20928 ) | ( n10215 & n20928 ) ;
  assign n20930 = ( n5019 & ~n20927 ) | ( n5019 & n20929 ) | ( ~n20927 & n20929 ) ;
  assign n20931 = n20927 | n20930 ;
  assign n20932 = n2422 | n4995 ;
  assign n20933 = n647 | n3420 ;
  assign n20934 = ( n3070 & n3571 ) | ( n3070 & ~n20933 ) | ( n3571 & ~n20933 ) ;
  assign n20935 = n20933 | n20934 ;
  assign n20936 = ( ~n20931 & n20932 ) | ( ~n20931 & n20935 ) | ( n20932 & n20935 ) ;
  assign n20937 = n20931 | n20936 ;
  assign n20938 = ( ~n1504 & n2451 ) | ( ~n1504 & n20937 ) | ( n2451 & n20937 ) ;
  assign n20939 = ~n20937 & n20938 ;
  assign n20940 = ( x11 & n20716 ) | ( x11 & n20939 ) | ( n20716 & n20939 ) ;
  assign n20941 = ( ~x11 & n20716 ) | ( ~x11 & n20939 ) | ( n20716 & n20939 ) ;
  assign n20942 = ( x11 & ~n20940 ) | ( x11 & n20941 ) | ( ~n20940 & n20941 ) ;
  assign n20943 = n607 & ~n16043 ;
  assign n20944 = n1250 & n16041 ;
  assign n20945 = n20943 | n20944 ;
  assign n20946 = n606 & ~n16039 ;
  assign n20947 = ( n606 & n20945 ) | ( n606 & ~n20946 ) | ( n20945 & ~n20946 ) ;
  assign n20948 = n1248 & ~n17051 ;
  assign n20949 = n20947 | n20948 ;
  assign n20950 = ( n20818 & ~n20942 ) | ( n20818 & n20949 ) | ( ~n20942 & n20949 ) ;
  assign n20951 = ( n20818 & n20942 ) | ( n20818 & n20949 ) | ( n20942 & n20949 ) ;
  assign n20952 = ( n20942 & n20950 ) | ( n20942 & ~n20951 ) | ( n20950 & ~n20951 ) ;
  assign n20953 = n3800 & ~n17412 ;
  assign n20954 = n3799 & ~n16033 ;
  assign n20955 = n3700 & ~n16037 ;
  assign n20956 = n3802 & n16035 ;
  assign n20957 = n20955 | n20956 ;
  assign n20958 = ( ~n20953 & n20954 ) | ( ~n20953 & n20957 ) | ( n20954 & n20957 ) ;
  assign n20959 = ( ~x29 & n20953 ) | ( ~x29 & n20958 ) | ( n20953 & n20958 ) ;
  assign n20960 = ( n20953 & n20958 ) | ( n20953 & ~n20959 ) | ( n20958 & ~n20959 ) ;
  assign n20961 = ( x29 & n20959 ) | ( x29 & ~n20960 ) | ( n20959 & ~n20960 ) ;
  assign n20962 = ( n20837 & ~n20952 ) | ( n20837 & n20961 ) | ( ~n20952 & n20961 ) ;
  assign n20963 = ( n20837 & n20952 ) | ( n20837 & n20961 ) | ( n20952 & n20961 ) ;
  assign n20964 = ( n20952 & n20962 ) | ( n20952 & ~n20963 ) | ( n20962 & ~n20963 ) ;
  assign n20965 = n4202 & n17634 ;
  assign n20966 = n4201 & ~n16027 ;
  assign n20967 = n4200 & n16031 ;
  assign n20968 = n4345 & ~n16029 ;
  assign n20969 = n20967 | n20968 ;
  assign n20970 = ( ~n20965 & n20966 ) | ( ~n20965 & n20969 ) | ( n20966 & n20969 ) ;
  assign n20971 = ( ~x26 & n20965 ) | ( ~x26 & n20970 ) | ( n20965 & n20970 ) ;
  assign n20972 = ( n20965 & n20970 ) | ( n20965 & ~n20971 ) | ( n20970 & ~n20971 ) ;
  assign n20973 = ( x26 & n20971 ) | ( x26 & ~n20972 ) | ( n20971 & ~n20972 ) ;
  assign n20974 = ( n20849 & ~n20964 ) | ( n20849 & n20973 ) | ( ~n20964 & n20973 ) ;
  assign n20975 = ( n20849 & n20964 ) | ( n20849 & n20973 ) | ( n20964 & n20973 ) ;
  assign n20976 = ( n20964 & n20974 ) | ( n20964 & ~n20975 ) | ( n20974 & ~n20975 ) ;
  assign n20977 = n4713 & ~n18091 ;
  assign n20978 = n4712 & n16021 ;
  assign n20979 = n4709 & ~n16025 ;
  assign n20980 = n4792 & n16023 ;
  assign n20981 = n20979 | n20980 ;
  assign n20982 = ( ~n20977 & n20978 ) | ( ~n20977 & n20981 ) | ( n20978 & n20981 ) ;
  assign n20983 = ( ~x23 & n20977 ) | ( ~x23 & n20982 ) | ( n20977 & n20982 ) ;
  assign n20984 = ( n20977 & n20982 ) | ( n20977 & ~n20983 ) | ( n20982 & ~n20983 ) ;
  assign n20985 = ( x23 & n20983 ) | ( x23 & ~n20984 ) | ( n20983 & ~n20984 ) ;
  assign n20986 = ( n20861 & ~n20976 ) | ( n20861 & n20985 ) | ( ~n20976 & n20985 ) ;
  assign n20987 = ( n20861 & n20976 ) | ( n20861 & n20985 ) | ( n20976 & n20985 ) ;
  assign n20988 = ( n20976 & n20986 ) | ( n20976 & ~n20987 ) | ( n20986 & ~n20987 ) ;
  assign n20989 = ( n20873 & n20925 ) | ( n20873 & ~n20988 ) | ( n20925 & ~n20988 ) ;
  assign n20990 = ( ~n20873 & n20925 ) | ( ~n20873 & n20988 ) | ( n20925 & n20988 ) ;
  assign n20991 = ( ~n20925 & n20989 ) | ( ~n20925 & n20990 ) | ( n20989 & n20990 ) ;
  assign n20992 = n5508 & n18996 ;
  assign n20993 = n5507 & n18993 ;
  assign n20994 = n5504 & ~n16013 ;
  assign n20995 = n5666 & n16138 ;
  assign n20996 = n20994 | n20995 ;
  assign n20997 = ( ~n20992 & n20993 ) | ( ~n20992 & n20996 ) | ( n20993 & n20996 ) ;
  assign n20998 = ( ~x17 & n20992 ) | ( ~x17 & n20997 ) | ( n20992 & n20997 ) ;
  assign n20999 = ( n20992 & n20997 ) | ( n20992 & ~n20998 ) | ( n20997 & ~n20998 ) ;
  assign n21000 = ( x17 & n20998 ) | ( x17 & ~n20999 ) | ( n20998 & ~n20999 ) ;
  assign n21001 = ( n20885 & ~n20991 ) | ( n20885 & n21000 ) | ( ~n20991 & n21000 ) ;
  assign n21002 = ( n20885 & n20991 ) | ( n20885 & n21000 ) | ( n20991 & n21000 ) ;
  assign n21003 = ( n20991 & n21001 ) | ( n20991 & ~n21002 ) | ( n21001 & ~n21002 ) ;
  assign n21004 = ( n20897 & n20916 ) | ( n20897 & ~n21003 ) | ( n20916 & ~n21003 ) ;
  assign n21005 = ( ~n20897 & n20916 ) | ( ~n20897 & n21003 ) | ( n20916 & n21003 ) ;
  assign n21006 = ( ~n20916 & n21004 ) | ( ~n20916 & n21005 ) | ( n21004 & n21005 ) ;
  assign n21007 = ( n20900 & n20903 ) | ( n20900 & ~n21006 ) | ( n20903 & ~n21006 ) ;
  assign n21008 = ( n20900 & n20903 ) | ( n20900 & n21006 ) | ( n20903 & n21006 ) ;
  assign n21009 = ( n21006 & n21007 ) | ( n21006 & ~n21008 ) | ( n21007 & ~n21008 ) ;
  assign n21010 = n20906 & ~n21009 ;
  assign n21011 = n20906 & n21009 ;
  assign n21012 = ( n21009 & n21010 ) | ( n21009 & ~n21011 ) | ( n21010 & ~n21011 ) ;
  assign n21013 = n607 & n16041 ;
  assign n21014 = n1250 & n16039 ;
  assign n21015 = n21013 | n21014 ;
  assign n21016 = n606 & n16037 ;
  assign n21017 = ( n606 & n21015 ) | ( n606 & ~n21016 ) | ( n21015 & ~n21016 ) ;
  assign n21018 = n1248 & n17138 ;
  assign n21019 = ( n1248 & n21017 ) | ( n1248 & ~n21018 ) | ( n21017 & ~n21018 ) ;
  assign n21020 = ( ~n10224 & n11529 ) | ( ~n10224 & n19338 ) | ( n11529 & n19338 ) ;
  assign n21021 = n595 | n1652 ;
  assign n21022 = ( n656 & n2443 ) | ( n656 & ~n21021 ) | ( n2443 & ~n21021 ) ;
  assign n21023 = n21021 | n21022 ;
  assign n21024 = ( n1278 & n2493 ) | ( n1278 & ~n10430 ) | ( n2493 & ~n10430 ) ;
  assign n21025 = n10430 | n21024 ;
  assign n21026 = ( n3030 & n3109 ) | ( n3030 & ~n3289 ) | ( n3109 & ~n3289 ) ;
  assign n21027 = n3289 | n21026 ;
  assign n21028 = ( ~n21023 & n21025 ) | ( ~n21023 & n21027 ) | ( n21025 & n21027 ) ;
  assign n21029 = n21023 | n21028 ;
  assign n21030 = ( ~n19338 & n19636 ) | ( ~n19338 & n21029 ) | ( n19636 & n21029 ) ;
  assign n21031 = ( ~n10224 & n21020 ) | ( ~n10224 & n21030 ) | ( n21020 & n21030 ) ;
  assign n21032 = n10224 | n21031 ;
  assign n21033 = ( n20940 & ~n21019 ) | ( n20940 & n21032 ) | ( ~n21019 & n21032 ) ;
  assign n21034 = ( n20940 & n21019 ) | ( n20940 & n21032 ) | ( n21019 & n21032 ) ;
  assign n21035 = ( n21019 & n21033 ) | ( n21019 & ~n21034 ) | ( n21033 & ~n21034 ) ;
  assign n21036 = n3800 & ~n17516 ;
  assign n21037 = n3799 & n16031 ;
  assign n21038 = n3700 & n16035 ;
  assign n21039 = n3802 & ~n16033 ;
  assign n21040 = n21038 | n21039 ;
  assign n21041 = ( ~n21036 & n21037 ) | ( ~n21036 & n21040 ) | ( n21037 & n21040 ) ;
  assign n21042 = ( ~x29 & n21036 ) | ( ~x29 & n21041 ) | ( n21036 & n21041 ) ;
  assign n21043 = ( n21036 & n21041 ) | ( n21036 & ~n21042 ) | ( n21041 & ~n21042 ) ;
  assign n21044 = ( x29 & n21042 ) | ( x29 & ~n21043 ) | ( n21042 & ~n21043 ) ;
  assign n21045 = ( n20950 & n21035 ) | ( n20950 & n21044 ) | ( n21035 & n21044 ) ;
  assign n21046 = ( ~n20950 & n21035 ) | ( ~n20950 & n21044 ) | ( n21035 & n21044 ) ;
  assign n21047 = ( n20950 & ~n21045 ) | ( n20950 & n21046 ) | ( ~n21045 & n21046 ) ;
  assign n21048 = n4202 & ~n17746 ;
  assign n21049 = n4201 & ~n16025 ;
  assign n21050 = n4200 & ~n16029 ;
  assign n21051 = n4345 & ~n16027 ;
  assign n21052 = n21050 | n21051 ;
  assign n21053 = ( ~n21048 & n21049 ) | ( ~n21048 & n21052 ) | ( n21049 & n21052 ) ;
  assign n21054 = ( ~x26 & n21048 ) | ( ~x26 & n21053 ) | ( n21048 & n21053 ) ;
  assign n21055 = ( n21048 & n21053 ) | ( n21048 & ~n21054 ) | ( n21053 & ~n21054 ) ;
  assign n21056 = ( x26 & n21054 ) | ( x26 & ~n21055 ) | ( n21054 & ~n21055 ) ;
  assign n21057 = ( n20962 & n21047 ) | ( n20962 & n21056 ) | ( n21047 & n21056 ) ;
  assign n21058 = ( n20962 & ~n21047 ) | ( n20962 & n21056 ) | ( ~n21047 & n21056 ) ;
  assign n21059 = ( n21047 & ~n21057 ) | ( n21047 & n21058 ) | ( ~n21057 & n21058 ) ;
  assign n21060 = n4713 & n18103 ;
  assign n21061 = n4712 & n16019 ;
  assign n21062 = n4709 & n16023 ;
  assign n21063 = n4792 & n16021 ;
  assign n21064 = n21062 | n21063 ;
  assign n21065 = ( ~n21060 & n21061 ) | ( ~n21060 & n21064 ) | ( n21061 & n21064 ) ;
  assign n21066 = ( ~x23 & n21060 ) | ( ~x23 & n21065 ) | ( n21060 & n21065 ) ;
  assign n21067 = ( n21060 & n21065 ) | ( n21060 & ~n21066 ) | ( n21065 & ~n21066 ) ;
  assign n21068 = ( x23 & n21066 ) | ( x23 & ~n21067 ) | ( n21066 & ~n21067 ) ;
  assign n21069 = ( n20974 & n21059 ) | ( n20974 & n21068 ) | ( n21059 & n21068 ) ;
  assign n21070 = ( n20974 & ~n21059 ) | ( n20974 & n21068 ) | ( ~n21059 & n21068 ) ;
  assign n21071 = ( n21059 & ~n21069 ) | ( n21059 & n21070 ) | ( ~n21069 & n21070 ) ;
  assign n21072 = n4974 & ~n18694 ;
  assign n21073 = n5398 & ~n16013 ;
  assign n21074 = n4973 & ~n16017 ;
  assign n21075 = n4972 & n16015 ;
  assign n21076 = n21074 | n21075 ;
  assign n21077 = ( ~n21072 & n21073 ) | ( ~n21072 & n21076 ) | ( n21073 & n21076 ) ;
  assign n21078 = ( ~x20 & n21072 ) | ( ~x20 & n21077 ) | ( n21072 & n21077 ) ;
  assign n21079 = ( n21072 & n21077 ) | ( n21072 & ~n21078 ) | ( n21077 & ~n21078 ) ;
  assign n21080 = ( x20 & n21078 ) | ( x20 & ~n21079 ) | ( n21078 & ~n21079 ) ;
  assign n21081 = ( n20986 & n21071 ) | ( n20986 & n21080 ) | ( n21071 & n21080 ) ;
  assign n21082 = ( n20986 & ~n21071 ) | ( n20986 & n21080 ) | ( ~n21071 & n21080 ) ;
  assign n21083 = ( n21071 & ~n21081 ) | ( n21071 & n21082 ) | ( ~n21081 & n21082 ) ;
  assign n21084 = n5508 & n19160 ;
  assign n21085 = n5507 & n19157 ;
  assign n21086 = n5504 & n16138 ;
  assign n21087 = n5666 & n18993 ;
  assign n21088 = n21086 | n21087 ;
  assign n21089 = ( ~n21084 & n21085 ) | ( ~n21084 & n21088 ) | ( n21085 & n21088 ) ;
  assign n21090 = ( ~x17 & n21084 ) | ( ~x17 & n21089 ) | ( n21084 & n21089 ) ;
  assign n21091 = ( n21084 & n21089 ) | ( n21084 & ~n21090 ) | ( n21089 & ~n21090 ) ;
  assign n21092 = ( x17 & n21090 ) | ( x17 & ~n21091 ) | ( n21090 & ~n21091 ) ;
  assign n21093 = ( n20989 & n21083 ) | ( n20989 & n21092 ) | ( n21083 & n21092 ) ;
  assign n21094 = ( n20989 & ~n21083 ) | ( n20989 & n21092 ) | ( ~n21083 & n21092 ) ;
  assign n21095 = ( n21083 & ~n21093 ) | ( n21083 & n21094 ) | ( ~n21093 & n21094 ) ;
  assign n21096 = n5970 & ~n19309 ;
  assign n21097 = ~x14 & n21096 ;
  assign n21098 = n21096 & ~n21097 ;
  assign n21099 = ( x14 & n21097 ) | ( x14 & ~n21098 ) | ( n21097 & ~n21098 ) ;
  assign n21100 = ( n21001 & n21095 ) | ( n21001 & n21099 ) | ( n21095 & n21099 ) ;
  assign n21101 = ( n21001 & ~n21095 ) | ( n21001 & n21099 ) | ( ~n21095 & n21099 ) ;
  assign n21102 = ( n21095 & ~n21100 ) | ( n21095 & n21101 ) | ( ~n21100 & n21101 ) ;
  assign n21103 = ( n21004 & n21007 ) | ( n21004 & n21102 ) | ( n21007 & n21102 ) ;
  assign n21104 = ( ~n21004 & n21007 ) | ( ~n21004 & n21102 ) | ( n21007 & n21102 ) ;
  assign n21105 = ( n21004 & ~n21103 ) | ( n21004 & n21104 ) | ( ~n21103 & n21104 ) ;
  assign n21106 = n21010 & n21105 ;
  assign n21107 = n21010 | n21105 ;
  assign n21108 = ~n21106 & n21107 ;
  assign n21109 = n607 & n16039 ;
  assign n21110 = n1250 & ~n16037 ;
  assign n21111 = n21109 | n21110 ;
  assign n21112 = n606 & ~n16035 ;
  assign n21113 = ( n606 & n21111 ) | ( n606 & ~n21112 ) | ( n21111 & ~n21112 ) ;
  assign n21114 = n1248 & n17313 ;
  assign n21115 = ( n1248 & n21113 ) | ( n1248 & ~n21114 ) | ( n21113 & ~n21114 ) ;
  assign n21116 = n562 | n760 ;
  assign n21117 = ( n489 & n1376 ) | ( n489 & ~n21116 ) | ( n1376 & ~n21116 ) ;
  assign n21118 = n21116 | n21117 ;
  assign n21119 = ( n346 & ~n923 ) | ( n346 & n1892 ) | ( ~n923 & n1892 ) ;
  assign n21120 = n923 | n21119 ;
  assign n21121 = n328 | n353 ;
  assign n21122 = ( n657 & n762 ) | ( n657 & ~n21121 ) | ( n762 & ~n21121 ) ;
  assign n21123 = n21121 | n21122 ;
  assign n21124 = ( ~n21118 & n21120 ) | ( ~n21118 & n21123 ) | ( n21120 & n21123 ) ;
  assign n21125 = n21118 | n21124 ;
  assign n21126 = n3072 | n3338 ;
  assign n21127 = ( n882 & ~n21125 ) | ( n882 & n21126 ) | ( ~n21125 & n21126 ) ;
  assign n21128 = n21125 | n21127 ;
  assign n21129 = ( n201 & ~n4024 ) | ( n201 & n21128 ) | ( ~n4024 & n21128 ) ;
  assign n21130 = ~n710 & n5129 ;
  assign n21131 = ( ~n4024 & n21129 ) | ( ~n4024 & n21130 ) | ( n21129 & n21130 ) ;
  assign n21132 = ~n21129 & n21131 ;
  assign n21133 = ( n21032 & ~n21115 ) | ( n21032 & n21132 ) | ( ~n21115 & n21132 ) ;
  assign n21134 = ( n21032 & n21115 ) | ( n21032 & n21132 ) | ( n21115 & n21132 ) ;
  assign n21135 = ( n21115 & n21133 ) | ( n21115 & ~n21134 ) | ( n21133 & ~n21134 ) ;
  assign n21136 = ( ~n21033 & n21045 ) | ( ~n21033 & n21135 ) | ( n21045 & n21135 ) ;
  assign n21137 = ( n21045 & n21135 ) | ( n21045 & ~n21136 ) | ( n21135 & ~n21136 ) ;
  assign n21138 = ( n21033 & n21136 ) | ( n21033 & ~n21137 ) | ( n21136 & ~n21137 ) ;
  assign n21139 = n4202 & n17968 ;
  assign n21140 = n4201 & n16023 ;
  assign n21141 = n4200 & ~n16027 ;
  assign n21142 = n4345 & ~n16025 ;
  assign n21143 = n21141 | n21142 ;
  assign n21144 = ( ~n21139 & n21140 ) | ( ~n21139 & n21143 ) | ( n21140 & n21143 ) ;
  assign n21145 = ( ~x26 & n21139 ) | ( ~x26 & n21144 ) | ( n21139 & n21144 ) ;
  assign n21146 = ( n21139 & n21144 ) | ( n21139 & ~n21145 ) | ( n21144 & ~n21145 ) ;
  assign n21147 = ( x26 & n21145 ) | ( x26 & ~n21146 ) | ( n21145 & ~n21146 ) ;
  assign n21148 = n3800 & ~n17528 ;
  assign n21149 = n3799 & ~n16029 ;
  assign n21150 = n3700 & ~n16033 ;
  assign n21151 = n3802 & n16031 ;
  assign n21152 = n21150 | n21151 ;
  assign n21153 = ( ~n21148 & n21149 ) | ( ~n21148 & n21152 ) | ( n21149 & n21152 ) ;
  assign n21154 = ( ~x29 & n21148 ) | ( ~x29 & n21153 ) | ( n21148 & n21153 ) ;
  assign n21155 = ( n21148 & n21153 ) | ( n21148 & ~n21154 ) | ( n21153 & ~n21154 ) ;
  assign n21156 = ( x29 & n21154 ) | ( x29 & ~n21155 ) | ( n21154 & ~n21155 ) ;
  assign n21157 = ( ~n21138 & n21147 ) | ( ~n21138 & n21156 ) | ( n21147 & n21156 ) ;
  assign n21158 = ( n21147 & n21156 ) | ( n21147 & ~n21157 ) | ( n21156 & ~n21157 ) ;
  assign n21159 = ( n21138 & n21157 ) | ( n21138 & ~n21158 ) | ( n21157 & ~n21158 ) ;
  assign n21160 = n4713 & ~n18267 ;
  assign n21161 = n4712 & ~n16017 ;
  assign n21162 = n4709 & n16021 ;
  assign n21163 = n4792 & n16019 ;
  assign n21164 = n21162 | n21163 ;
  assign n21165 = ( ~n21160 & n21161 ) | ( ~n21160 & n21164 ) | ( n21161 & n21164 ) ;
  assign n21166 = ( ~x23 & n21160 ) | ( ~x23 & n21165 ) | ( n21160 & n21165 ) ;
  assign n21167 = ( n21160 & n21165 ) | ( n21160 & ~n21166 ) | ( n21165 & ~n21166 ) ;
  assign n21168 = ( x23 & n21166 ) | ( x23 & ~n21167 ) | ( n21166 & ~n21167 ) ;
  assign n21169 = ( n21057 & ~n21159 ) | ( n21057 & n21168 ) | ( ~n21159 & n21168 ) ;
  assign n21170 = ( n21057 & n21159 ) | ( n21057 & n21168 ) | ( n21159 & n21168 ) ;
  assign n21171 = ( n21159 & n21169 ) | ( n21159 & ~n21170 ) | ( n21169 & ~n21170 ) ;
  assign n21172 = n4974 & ~n16144 ;
  assign n21173 = n5398 & n16138 ;
  assign n21174 = n4973 & n16015 ;
  assign n21175 = n4972 & ~n16013 ;
  assign n21176 = n21174 | n21175 ;
  assign n21177 = ( ~n21172 & n21173 ) | ( ~n21172 & n21176 ) | ( n21173 & n21176 ) ;
  assign n21178 = ( ~x20 & n21172 ) | ( ~x20 & n21177 ) | ( n21172 & n21177 ) ;
  assign n21179 = ( n21172 & n21177 ) | ( n21172 & ~n21178 ) | ( n21177 & ~n21178 ) ;
  assign n21180 = ( x20 & n21178 ) | ( x20 & ~n21179 ) | ( n21178 & ~n21179 ) ;
  assign n21181 = ( n21069 & ~n21171 ) | ( n21069 & n21180 ) | ( ~n21171 & n21180 ) ;
  assign n21182 = ( n21069 & n21171 ) | ( n21069 & n21180 ) | ( n21171 & n21180 ) ;
  assign n21183 = ( n21171 & n21181 ) | ( n21171 & ~n21182 ) | ( n21181 & ~n21182 ) ;
  assign n21184 = n5508 & ~n19312 ;
  assign n21185 = n5507 & ~n19309 ;
  assign n21186 = n5504 & n18993 ;
  assign n21187 = n5666 & n19157 ;
  assign n21188 = n21186 | n21187 ;
  assign n21189 = ( ~n21184 & n21185 ) | ( ~n21184 & n21188 ) | ( n21185 & n21188 ) ;
  assign n21190 = ( ~x17 & n21184 ) | ( ~x17 & n21189 ) | ( n21184 & n21189 ) ;
  assign n21191 = ( n21184 & n21189 ) | ( n21184 & ~n21190 ) | ( n21189 & ~n21190 ) ;
  assign n21192 = ( x17 & n21190 ) | ( x17 & ~n21191 ) | ( n21190 & ~n21191 ) ;
  assign n21193 = ( n21081 & ~n21183 ) | ( n21081 & n21192 ) | ( ~n21183 & n21192 ) ;
  assign n21194 = ( n21081 & n21183 ) | ( n21081 & n21192 ) | ( n21183 & n21192 ) ;
  assign n21195 = ( n21183 & n21193 ) | ( n21183 & ~n21194 ) | ( n21193 & ~n21194 ) ;
  assign n21196 = ( x14 & n21093 ) | ( x14 & ~n21195 ) | ( n21093 & ~n21195 ) ;
  assign n21197 = ( x14 & n21093 ) | ( x14 & n21195 ) | ( n21093 & n21195 ) ;
  assign n21198 = ( n21195 & n21196 ) | ( n21195 & ~n21197 ) | ( n21196 & ~n21197 ) ;
  assign n21199 = ( n21100 & n21103 ) | ( n21100 & ~n21198 ) | ( n21103 & ~n21198 ) ;
  assign n21200 = ( n21100 & n21103 ) | ( n21100 & n21198 ) | ( n21103 & n21198 ) ;
  assign n21201 = ( n21198 & n21199 ) | ( n21198 & ~n21200 ) | ( n21199 & ~n21200 ) ;
  assign n21202 = n21106 & ~n21201 ;
  assign n21203 = n21106 & n21201 ;
  assign n21204 = ( n21201 & n21202 ) | ( n21201 & ~n21203 ) | ( n21202 & ~n21203 ) ;
  assign n21205 = n5508 & ~n19472 ;
  assign n21206 = n5666 & ~n19309 ;
  assign n21207 = ~n5504 & n19157 ;
  assign n21208 = ( n19157 & n21206 ) | ( n19157 & ~n21207 ) | ( n21206 & ~n21207 ) ;
  assign n21209 = ( ~x17 & n21205 ) | ( ~x17 & n21208 ) | ( n21205 & n21208 ) ;
  assign n21210 = ( n21205 & n21208 ) | ( n21205 & ~n21209 ) | ( n21208 & ~n21209 ) ;
  assign n21211 = ( x17 & n21209 ) | ( x17 & ~n21210 ) | ( n21209 & ~n21210 ) ;
  assign n21212 = n4713 & ~n18416 ;
  assign n21213 = n4712 & n16015 ;
  assign n21214 = n4709 & n16019 ;
  assign n21215 = n4792 & ~n16017 ;
  assign n21216 = n21214 | n21215 ;
  assign n21217 = ( ~n21212 & n21213 ) | ( ~n21212 & n21216 ) | ( n21213 & n21216 ) ;
  assign n21218 = ( ~x23 & n21212 ) | ( ~x23 & n21217 ) | ( n21212 & n21217 ) ;
  assign n21219 = ( n21212 & n21217 ) | ( n21212 & ~n21218 ) | ( n21217 & ~n21218 ) ;
  assign n21220 = ( x23 & n21218 ) | ( x23 & ~n21219 ) | ( n21218 & ~n21219 ) ;
  assign n21221 = n3370 | n11406 ;
  assign n21222 = n148 | n298 ;
  assign n21223 = ( ~n1613 & n11103 ) | ( ~n1613 & n21222 ) | ( n11103 & n21222 ) ;
  assign n21224 = ( n1599 & n1613 ) | ( n1599 & ~n21223 ) | ( n1613 & ~n21223 ) ;
  assign n21225 = n21223 | n21224 ;
  assign n21226 = ( n3988 & ~n21221 ) | ( n3988 & n21225 ) | ( ~n21221 & n21225 ) ;
  assign n21227 = n21221 | n21226 ;
  assign n21228 = ( n2151 & n2373 ) | ( n2151 & n6036 ) | ( n2373 & n6036 ) ;
  assign n21229 = n6036 & ~n21228 ;
  assign n21230 = ( ~n10826 & n21227 ) | ( ~n10826 & n21229 ) | ( n21227 & n21229 ) ;
  assign n21231 = ~n21227 & n21230 ;
  assign n21232 = ( x14 & ~n21032 ) | ( x14 & n21231 ) | ( ~n21032 & n21231 ) ;
  assign n21233 = ( x14 & n21231 ) | ( x14 & ~n21232 ) | ( n21231 & ~n21232 ) ;
  assign n21234 = ( n21032 & n21232 ) | ( n21032 & ~n21233 ) | ( n21232 & ~n21233 ) ;
  assign n21235 = n607 & ~n16037 ;
  assign n21236 = n1250 & n16035 ;
  assign n21237 = n21235 | n21236 ;
  assign n21238 = n606 & n16033 ;
  assign n21239 = ( n606 & n21237 ) | ( n606 & ~n21238 ) | ( n21237 & ~n21238 ) ;
  assign n21240 = n1248 & n17412 ;
  assign n21241 = ( n1248 & n21239 ) | ( n1248 & ~n21240 ) | ( n21239 & ~n21240 ) ;
  assign n21242 = ( ~n21133 & n21234 ) | ( ~n21133 & n21241 ) | ( n21234 & n21241 ) ;
  assign n21243 = ( n21234 & n21241 ) | ( n21234 & ~n21242 ) | ( n21241 & ~n21242 ) ;
  assign n21244 = ( n21133 & n21242 ) | ( n21133 & ~n21243 ) | ( n21242 & ~n21243 ) ;
  assign n21245 = n3800 & n17634 ;
  assign n21246 = n3799 & ~n16027 ;
  assign n21247 = n3700 & n16031 ;
  assign n21248 = n3802 & ~n16029 ;
  assign n21249 = n21247 | n21248 ;
  assign n21250 = ( ~n21245 & n21246 ) | ( ~n21245 & n21249 ) | ( n21246 & n21249 ) ;
  assign n21251 = ( ~x29 & n21245 ) | ( ~x29 & n21250 ) | ( n21245 & n21250 ) ;
  assign n21252 = ( n21245 & n21250 ) | ( n21245 & ~n21251 ) | ( n21250 & ~n21251 ) ;
  assign n21253 = ( x29 & n21251 ) | ( x29 & ~n21252 ) | ( n21251 & ~n21252 ) ;
  assign n21254 = ( n21136 & ~n21244 ) | ( n21136 & n21253 ) | ( ~n21244 & n21253 ) ;
  assign n21255 = ( n21136 & n21244 ) | ( n21136 & n21253 ) | ( n21244 & n21253 ) ;
  assign n21256 = ( n21244 & n21254 ) | ( n21244 & ~n21255 ) | ( n21254 & ~n21255 ) ;
  assign n21257 = n4202 & ~n18091 ;
  assign n21258 = n4201 & n16021 ;
  assign n21259 = n4200 & ~n16025 ;
  assign n21260 = n4345 & n16023 ;
  assign n21261 = n21259 | n21260 ;
  assign n21262 = ( ~n21257 & n21258 ) | ( ~n21257 & n21261 ) | ( n21258 & n21261 ) ;
  assign n21263 = ( ~x26 & n21257 ) | ( ~x26 & n21262 ) | ( n21257 & n21262 ) ;
  assign n21264 = ( n21257 & n21262 ) | ( n21257 & ~n21263 ) | ( n21262 & ~n21263 ) ;
  assign n21265 = ( x26 & n21263 ) | ( x26 & ~n21264 ) | ( n21263 & ~n21264 ) ;
  assign n21266 = ( n21157 & ~n21256 ) | ( n21157 & n21265 ) | ( ~n21256 & n21265 ) ;
  assign n21267 = ( n21157 & n21256 ) | ( n21157 & n21265 ) | ( n21256 & n21265 ) ;
  assign n21268 = ( n21256 & n21266 ) | ( n21256 & ~n21267 ) | ( n21266 & ~n21267 ) ;
  assign n21269 = ( n21169 & n21220 ) | ( n21169 & ~n21268 ) | ( n21220 & ~n21268 ) ;
  assign n21270 = ( ~n21169 & n21220 ) | ( ~n21169 & n21268 ) | ( n21220 & n21268 ) ;
  assign n21271 = ( ~n21220 & n21269 ) | ( ~n21220 & n21270 ) | ( n21269 & n21270 ) ;
  assign n21272 = n4974 & n18996 ;
  assign n21273 = n5398 & n18993 ;
  assign n21274 = n4973 & ~n16013 ;
  assign n21275 = n4972 & n16138 ;
  assign n21276 = n21274 | n21275 ;
  assign n21277 = ( ~n21272 & n21273 ) | ( ~n21272 & n21276 ) | ( n21273 & n21276 ) ;
  assign n21278 = ( ~x20 & n21272 ) | ( ~x20 & n21277 ) | ( n21272 & n21277 ) ;
  assign n21279 = ( n21272 & n21277 ) | ( n21272 & ~n21278 ) | ( n21277 & ~n21278 ) ;
  assign n21280 = ( x20 & n21278 ) | ( x20 & ~n21279 ) | ( n21278 & ~n21279 ) ;
  assign n21281 = ( n21181 & ~n21271 ) | ( n21181 & n21280 ) | ( ~n21271 & n21280 ) ;
  assign n21282 = ( n21181 & n21271 ) | ( n21181 & n21280 ) | ( n21271 & n21280 ) ;
  assign n21283 = ( n21271 & n21281 ) | ( n21271 & ~n21282 ) | ( n21281 & ~n21282 ) ;
  assign n21284 = ( n21193 & n21211 ) | ( n21193 & ~n21283 ) | ( n21211 & ~n21283 ) ;
  assign n21285 = ( ~n21193 & n21211 ) | ( ~n21193 & n21283 ) | ( n21211 & n21283 ) ;
  assign n21286 = ( ~n21211 & n21284 ) | ( ~n21211 & n21285 ) | ( n21284 & n21285 ) ;
  assign n21287 = ( n21196 & n21199 ) | ( n21196 & ~n21286 ) | ( n21199 & ~n21286 ) ;
  assign n21288 = ( n21196 & n21199 ) | ( n21196 & n21286 ) | ( n21199 & n21286 ) ;
  assign n21289 = ( n21286 & n21287 ) | ( n21286 & ~n21288 ) | ( n21287 & ~n21288 ) ;
  assign n21290 = n21202 & ~n21289 ;
  assign n21291 = ~n21202 & n21289 ;
  assign n21292 = n21290 | n21291 ;
  assign n21293 = n3800 & ~n17746 ;
  assign n21294 = n3799 & ~n16025 ;
  assign n21295 = n3700 & ~n16029 ;
  assign n21296 = n3802 & ~n16027 ;
  assign n21297 = n21295 | n21296 ;
  assign n21298 = ( ~n21293 & n21294 ) | ( ~n21293 & n21297 ) | ( n21294 & n21297 ) ;
  assign n21299 = ( ~x29 & n21293 ) | ( ~x29 & n21298 ) | ( n21293 & n21298 ) ;
  assign n21300 = ( n21293 & n21298 ) | ( n21293 & ~n21299 ) | ( n21298 & ~n21299 ) ;
  assign n21301 = ( x29 & n21299 ) | ( x29 & ~n21300 ) | ( n21299 & ~n21300 ) ;
  assign n21302 = ( n3497 & n5000 ) | ( n3497 & n5521 ) | ( n5000 & n5521 ) ;
  assign n21303 = n648 | n2791 ;
  assign n21304 = n11810 | n21303 ;
  assign n21305 = n1315 | n2163 ;
  assign n21306 = n887 | n1032 ;
  assign n21307 = n138 | n291 ;
  assign n21308 = ( n806 & n2480 ) | ( n806 & ~n21307 ) | ( n2480 & ~n21307 ) ;
  assign n21309 = n21307 | n21308 ;
  assign n21310 = ( ~n21305 & n21306 ) | ( ~n21305 & n21309 ) | ( n21306 & n21309 ) ;
  assign n21311 = n21305 | n21310 ;
  assign n21312 = ( n210 & ~n21304 ) | ( n210 & n21311 ) | ( ~n21304 & n21311 ) ;
  assign n21313 = n21304 | n21312 ;
  assign n21314 = ( ~n5521 & n11008 ) | ( ~n5521 & n21313 ) | ( n11008 & n21313 ) ;
  assign n21315 = ( n3497 & n21302 ) | ( n3497 & n21314 ) | ( n21302 & n21314 ) ;
  assign n21316 = n3497 & ~n21315 ;
  assign n21317 = n607 & n16035 ;
  assign n21318 = n1250 & ~n16033 ;
  assign n21319 = n21317 | n21318 ;
  assign n21320 = n606 & ~n16031 ;
  assign n21321 = ( n606 & n21319 ) | ( n606 & ~n21320 ) | ( n21319 & ~n21320 ) ;
  assign n21322 = n1248 & n17516 ;
  assign n21323 = ( n1248 & n21321 ) | ( n1248 & ~n21322 ) | ( n21321 & ~n21322 ) ;
  assign n21324 = ( ~n21232 & n21316 ) | ( ~n21232 & n21323 ) | ( n21316 & n21323 ) ;
  assign n21325 = ( n21316 & n21323 ) | ( n21316 & ~n21324 ) | ( n21323 & ~n21324 ) ;
  assign n21326 = ( n21232 & n21324 ) | ( n21232 & ~n21325 ) | ( n21324 & ~n21325 ) ;
  assign n21327 = ( n21242 & n21301 ) | ( n21242 & ~n21326 ) | ( n21301 & ~n21326 ) ;
  assign n21328 = ( ~n21242 & n21301 ) | ( ~n21242 & n21326 ) | ( n21301 & n21326 ) ;
  assign n21329 = ( ~n21301 & n21327 ) | ( ~n21301 & n21328 ) | ( n21327 & n21328 ) ;
  assign n21330 = n4202 & n18103 ;
  assign n21331 = n4201 & n16019 ;
  assign n21332 = n4200 & n16023 ;
  assign n21333 = n4345 & n16021 ;
  assign n21334 = n21332 | n21333 ;
  assign n21335 = ( ~n21330 & n21331 ) | ( ~n21330 & n21334 ) | ( n21331 & n21334 ) ;
  assign n21336 = ( ~x26 & n21330 ) | ( ~x26 & n21335 ) | ( n21330 & n21335 ) ;
  assign n21337 = ( n21330 & n21335 ) | ( n21330 & ~n21336 ) | ( n21335 & ~n21336 ) ;
  assign n21338 = ( x26 & n21336 ) | ( x26 & ~n21337 ) | ( n21336 & ~n21337 ) ;
  assign n21339 = ( n21254 & ~n21329 ) | ( n21254 & n21338 ) | ( ~n21329 & n21338 ) ;
  assign n21340 = ( n21254 & n21329 ) | ( n21254 & n21338 ) | ( n21329 & n21338 ) ;
  assign n21341 = ( n21329 & n21339 ) | ( n21329 & ~n21340 ) | ( n21339 & ~n21340 ) ;
  assign n21342 = n4713 & ~n18694 ;
  assign n21343 = n4712 & ~n16013 ;
  assign n21344 = n4709 & ~n16017 ;
  assign n21345 = n4792 & n16015 ;
  assign n21346 = n21344 | n21345 ;
  assign n21347 = ( ~n21342 & n21343 ) | ( ~n21342 & n21346 ) | ( n21343 & n21346 ) ;
  assign n21348 = ( ~x23 & n21342 ) | ( ~x23 & n21347 ) | ( n21342 & n21347 ) ;
  assign n21349 = ( n21342 & n21347 ) | ( n21342 & ~n21348 ) | ( n21347 & ~n21348 ) ;
  assign n21350 = ( x23 & n21348 ) | ( x23 & ~n21349 ) | ( n21348 & ~n21349 ) ;
  assign n21351 = ( n21266 & ~n21341 ) | ( n21266 & n21350 ) | ( ~n21341 & n21350 ) ;
  assign n21352 = ( n21266 & n21341 ) | ( n21266 & n21350 ) | ( n21341 & n21350 ) ;
  assign n21353 = ( n21341 & n21351 ) | ( n21341 & ~n21352 ) | ( n21351 & ~n21352 ) ;
  assign n21354 = n4974 & n19160 ;
  assign n21355 = n5398 & n19157 ;
  assign n21356 = n4973 & n16138 ;
  assign n21357 = n4972 & n18993 ;
  assign n21358 = n21356 | n21357 ;
  assign n21359 = ( ~n21354 & n21355 ) | ( ~n21354 & n21358 ) | ( n21355 & n21358 ) ;
  assign n21360 = ( ~x20 & n21354 ) | ( ~x20 & n21359 ) | ( n21354 & n21359 ) ;
  assign n21361 = ( n21354 & n21359 ) | ( n21354 & ~n21360 ) | ( n21359 & ~n21360 ) ;
  assign n21362 = ( x20 & n21360 ) | ( x20 & ~n21361 ) | ( n21360 & ~n21361 ) ;
  assign n21363 = ( n21269 & ~n21353 ) | ( n21269 & n21362 ) | ( ~n21353 & n21362 ) ;
  assign n21364 = ( n21269 & n21353 ) | ( n21269 & n21362 ) | ( n21353 & n21362 ) ;
  assign n21365 = ( n21353 & n21363 ) | ( n21353 & ~n21364 ) | ( n21363 & ~n21364 ) ;
  assign n21366 = n5504 & ~n19309 ;
  assign n21367 = ~x17 & n21366 ;
  assign n21368 = n21366 & ~n21367 ;
  assign n21369 = ( x17 & n21367 ) | ( x17 & ~n21368 ) | ( n21367 & ~n21368 ) ;
  assign n21370 = ( n21281 & ~n21365 ) | ( n21281 & n21369 ) | ( ~n21365 & n21369 ) ;
  assign n21371 = ( n21281 & n21365 ) | ( n21281 & n21369 ) | ( n21365 & n21369 ) ;
  assign n21372 = ( n21365 & n21370 ) | ( n21365 & ~n21371 ) | ( n21370 & ~n21371 ) ;
  assign n21373 = ( n21284 & n21287 ) | ( n21284 & ~n21372 ) | ( n21287 & ~n21372 ) ;
  assign n21374 = ( n21284 & n21287 ) | ( n21284 & n21372 ) | ( n21287 & n21372 ) ;
  assign n21375 = ( n21372 & n21373 ) | ( n21372 & ~n21374 ) | ( n21373 & ~n21374 ) ;
  assign n21376 = n21290 & ~n21375 ;
  assign n21377 = n21290 & n21375 ;
  assign n21378 = ( n21375 & n21376 ) | ( n21375 & ~n21377 ) | ( n21376 & ~n21377 ) ;
  assign n21379 = n1652 | n2798 ;
  assign n21380 = n1736 | n1800 ;
  assign n21381 = ( n2443 & n2914 ) | ( n2443 & ~n21380 ) | ( n2914 & ~n21380 ) ;
  assign n21382 = n21380 | n21381 ;
  assign n21383 = n239 | n796 ;
  assign n21384 = ( n666 & n775 ) | ( n666 & ~n21383 ) | ( n775 & ~n21383 ) ;
  assign n21385 = n21383 | n21384 ;
  assign n21386 = ( ~n21379 & n21382 ) | ( ~n21379 & n21385 ) | ( n21382 & n21385 ) ;
  assign n21387 = n21379 | n21386 ;
  assign n21388 = ( n571 & ~n3319 ) | ( n571 & n21387 ) | ( ~n3319 & n21387 ) ;
  assign n21389 = n824 | n11921 ;
  assign n21390 = ( n3319 & ~n21388 ) | ( n3319 & n21389 ) | ( ~n21388 & n21389 ) ;
  assign n21391 = n21388 | n21390 ;
  assign n21392 = n1037 | n2230 ;
  assign n21393 = ( n5101 & ~n21391 ) | ( n5101 & n21392 ) | ( ~n21391 & n21392 ) ;
  assign n21394 = n21391 | n21393 ;
  assign n21395 = ( n21316 & ~n21324 ) | ( n21316 & n21394 ) | ( ~n21324 & n21394 ) ;
  assign n21396 = ( n21316 & n21394 ) | ( n21316 & ~n21395 ) | ( n21394 & ~n21395 ) ;
  assign n21397 = ( n21324 & n21395 ) | ( n21324 & ~n21396 ) | ( n21395 & ~n21396 ) ;
  assign n21398 = n3800 & n17968 ;
  assign n21399 = n3799 & n16023 ;
  assign n21400 = n3700 & ~n16027 ;
  assign n21401 = n3802 & ~n16025 ;
  assign n21402 = n21400 | n21401 ;
  assign n21403 = ( ~n21398 & n21399 ) | ( ~n21398 & n21402 ) | ( n21399 & n21402 ) ;
  assign n21404 = ( ~x29 & n21398 ) | ( ~x29 & n21403 ) | ( n21398 & n21403 ) ;
  assign n21405 = ( n21398 & n21403 ) | ( n21398 & ~n21404 ) | ( n21403 & ~n21404 ) ;
  assign n21406 = ( x29 & n21404 ) | ( x29 & ~n21405 ) | ( n21404 & ~n21405 ) ;
  assign n21407 = n607 & ~n16033 ;
  assign n21408 = n1250 & n16031 ;
  assign n21409 = n21407 | n21408 ;
  assign n21410 = n606 & n16029 ;
  assign n21411 = ( n606 & n21409 ) | ( n606 & ~n21410 ) | ( n21409 & ~n21410 ) ;
  assign n21412 = n1248 & n17528 ;
  assign n21413 = ( n1248 & n21411 ) | ( n1248 & ~n21412 ) | ( n21411 & ~n21412 ) ;
  assign n21414 = ( n21397 & n21406 ) | ( n21397 & n21413 ) | ( n21406 & n21413 ) ;
  assign n21415 = ( ~n21397 & n21406 ) | ( ~n21397 & n21413 ) | ( n21406 & n21413 ) ;
  assign n21416 = ( n21397 & ~n21414 ) | ( n21397 & n21415 ) | ( ~n21414 & n21415 ) ;
  assign n21417 = n4202 & ~n18267 ;
  assign n21418 = n4201 & ~n16017 ;
  assign n21419 = n4200 & n16021 ;
  assign n21420 = n4345 & n16019 ;
  assign n21421 = n21419 | n21420 ;
  assign n21422 = ( ~n21417 & n21418 ) | ( ~n21417 & n21421 ) | ( n21418 & n21421 ) ;
  assign n21423 = ( ~x26 & n21417 ) | ( ~x26 & n21422 ) | ( n21417 & n21422 ) ;
  assign n21424 = ( n21417 & n21422 ) | ( n21417 & ~n21423 ) | ( n21422 & ~n21423 ) ;
  assign n21425 = ( x26 & n21423 ) | ( x26 & ~n21424 ) | ( n21423 & ~n21424 ) ;
  assign n21426 = ( n21327 & n21416 ) | ( n21327 & n21425 ) | ( n21416 & n21425 ) ;
  assign n21427 = ( n21327 & ~n21416 ) | ( n21327 & n21425 ) | ( ~n21416 & n21425 ) ;
  assign n21428 = ( n21416 & ~n21426 ) | ( n21416 & n21427 ) | ( ~n21426 & n21427 ) ;
  assign n21429 = n4713 & ~n16144 ;
  assign n21430 = n4712 & n16138 ;
  assign n21431 = n4709 & n16015 ;
  assign n21432 = n4792 & ~n16013 ;
  assign n21433 = n21431 | n21432 ;
  assign n21434 = ( ~n21429 & n21430 ) | ( ~n21429 & n21433 ) | ( n21430 & n21433 ) ;
  assign n21435 = ( ~x23 & n21429 ) | ( ~x23 & n21434 ) | ( n21429 & n21434 ) ;
  assign n21436 = ( n21429 & n21434 ) | ( n21429 & ~n21435 ) | ( n21434 & ~n21435 ) ;
  assign n21437 = ( x23 & n21435 ) | ( x23 & ~n21436 ) | ( n21435 & ~n21436 ) ;
  assign n21438 = ( n21339 & n21428 ) | ( n21339 & n21437 ) | ( n21428 & n21437 ) ;
  assign n21439 = ( n21339 & ~n21428 ) | ( n21339 & n21437 ) | ( ~n21428 & n21437 ) ;
  assign n21440 = ( n21428 & ~n21438 ) | ( n21428 & n21439 ) | ( ~n21438 & n21439 ) ;
  assign n21441 = n4974 & ~n19312 ;
  assign n21442 = n5398 & ~n19309 ;
  assign n21443 = n4973 & n18993 ;
  assign n21444 = n4972 & n19157 ;
  assign n21445 = n21443 | n21444 ;
  assign n21446 = ( ~n21441 & n21442 ) | ( ~n21441 & n21445 ) | ( n21442 & n21445 ) ;
  assign n21447 = ( ~x20 & n21441 ) | ( ~x20 & n21446 ) | ( n21441 & n21446 ) ;
  assign n21448 = ( n21441 & n21446 ) | ( n21441 & ~n21447 ) | ( n21446 & ~n21447 ) ;
  assign n21449 = ( x20 & n21447 ) | ( x20 & ~n21448 ) | ( n21447 & ~n21448 ) ;
  assign n21450 = ( n21351 & n21440 ) | ( n21351 & n21449 ) | ( n21440 & n21449 ) ;
  assign n21451 = ( n21351 & ~n21440 ) | ( n21351 & n21449 ) | ( ~n21440 & n21449 ) ;
  assign n21452 = ( n21440 & ~n21450 ) | ( n21440 & n21451 ) | ( ~n21450 & n21451 ) ;
  assign n21453 = ( x17 & n21363 ) | ( x17 & n21452 ) | ( n21363 & n21452 ) ;
  assign n21454 = ( ~x17 & n21363 ) | ( ~x17 & n21452 ) | ( n21363 & n21452 ) ;
  assign n21455 = ( x17 & ~n21453 ) | ( x17 & n21454 ) | ( ~n21453 & n21454 ) ;
  assign n21456 = ( n21370 & n21373 ) | ( n21370 & n21455 ) | ( n21373 & n21455 ) ;
  assign n21457 = ( n21370 & ~n21373 ) | ( n21370 & n21455 ) | ( ~n21373 & n21455 ) ;
  assign n21458 = ( n21373 & ~n21456 ) | ( n21373 & n21457 ) | ( ~n21456 & n21457 ) ;
  assign n21459 = n21376 & n21458 ;
  assign n21460 = n21376 | n21458 ;
  assign n21461 = ~n21459 & n21460 ;
  assign n21462 = n4713 & n18996 ;
  assign n21463 = n4712 & n18993 ;
  assign n21464 = n4709 & ~n16013 ;
  assign n21465 = n4792 & n16138 ;
  assign n21466 = n21464 | n21465 ;
  assign n21467 = ( ~n21462 & n21463 ) | ( ~n21462 & n21466 ) | ( n21463 & n21466 ) ;
  assign n21468 = ( ~x23 & n21462 ) | ( ~x23 & n21467 ) | ( n21462 & n21467 ) ;
  assign n21469 = ( n21462 & n21467 ) | ( n21462 & ~n21468 ) | ( n21467 & ~n21468 ) ;
  assign n21470 = ( x23 & n21468 ) | ( x23 & ~n21469 ) | ( n21468 & ~n21469 ) ;
  assign n21471 = n3800 & ~n18091 ;
  assign n21472 = n3799 & n16021 ;
  assign n21473 = n3700 & ~n16025 ;
  assign n21474 = n3802 & n16023 ;
  assign n21475 = n21473 | n21474 ;
  assign n21476 = ( ~n21471 & n21472 ) | ( ~n21471 & n21475 ) | ( n21472 & n21475 ) ;
  assign n21477 = ( ~x29 & n21471 ) | ( ~x29 & n21476 ) | ( n21471 & n21476 ) ;
  assign n21478 = ( n21471 & n21476 ) | ( n21471 & ~n21477 ) | ( n21476 & ~n21477 ) ;
  assign n21479 = ( x29 & n21477 ) | ( x29 & ~n21478 ) | ( n21477 & ~n21478 ) ;
  assign n21480 = n607 & n16031 ;
  assign n21481 = n1250 & ~n16029 ;
  assign n21482 = n21480 | n21481 ;
  assign n21483 = n606 & n16027 ;
  assign n21484 = ( n606 & n21482 ) | ( n606 & ~n21483 ) | ( n21482 & ~n21483 ) ;
  assign n21485 = n1248 & ~n17634 ;
  assign n21486 = ( n1248 & n21484 ) | ( n1248 & ~n21485 ) | ( n21484 & ~n21485 ) ;
  assign n21487 = ( n963 & ~n1692 ) | ( n963 & n2046 ) | ( ~n1692 & n2046 ) ;
  assign n21488 = ( n1692 & ~n4221 ) | ( n1692 & n21487 ) | ( ~n4221 & n21487 ) ;
  assign n21489 = n4221 | n21488 ;
  assign n21490 = ( n1818 & ~n2190 ) | ( n1818 & n18476 ) | ( ~n2190 & n18476 ) ;
  assign n21491 = n2190 | n21490 ;
  assign n21492 = ( n2076 & n3507 ) | ( n2076 & ~n10085 ) | ( n3507 & ~n10085 ) ;
  assign n21493 = n10085 | n21492 ;
  assign n21494 = ( ~n21489 & n21491 ) | ( ~n21489 & n21493 ) | ( n21491 & n21493 ) ;
  assign n21495 = n21489 | n21494 ;
  assign n21496 = ( n4269 & n4843 ) | ( n4269 & ~n21495 ) | ( n4843 & ~n21495 ) ;
  assign n21497 = n21495 | n21496 ;
  assign n21498 = ( ~x17 & n21394 ) | ( ~x17 & n21497 ) | ( n21394 & n21497 ) ;
  assign n21499 = ( x17 & n21394 ) | ( x17 & n21497 ) | ( n21394 & n21497 ) ;
  assign n21500 = ( x17 & n21498 ) | ( x17 & ~n21499 ) | ( n21498 & ~n21499 ) ;
  assign n21501 = ( n21395 & ~n21486 ) | ( n21395 & n21500 ) | ( ~n21486 & n21500 ) ;
  assign n21502 = ( n21395 & n21486 ) | ( n21395 & n21500 ) | ( n21486 & n21500 ) ;
  assign n21503 = ( n21486 & n21501 ) | ( n21486 & ~n21502 ) | ( n21501 & ~n21502 ) ;
  assign n21504 = ( n21414 & n21479 ) | ( n21414 & n21503 ) | ( n21479 & n21503 ) ;
  assign n21505 = ( ~n21414 & n21479 ) | ( ~n21414 & n21503 ) | ( n21479 & n21503 ) ;
  assign n21506 = ( n21414 & ~n21504 ) | ( n21414 & n21505 ) | ( ~n21504 & n21505 ) ;
  assign n21507 = n4202 & ~n18416 ;
  assign n21508 = n4201 & n16015 ;
  assign n21509 = n4200 & n16019 ;
  assign n21510 = n4345 & ~n16017 ;
  assign n21511 = n21509 | n21510 ;
  assign n21512 = ( ~n21507 & n21508 ) | ( ~n21507 & n21511 ) | ( n21508 & n21511 ) ;
  assign n21513 = ( ~x26 & n21507 ) | ( ~x26 & n21512 ) | ( n21507 & n21512 ) ;
  assign n21514 = ( n21507 & n21512 ) | ( n21507 & ~n21513 ) | ( n21512 & ~n21513 ) ;
  assign n21515 = ( x26 & n21513 ) | ( x26 & ~n21514 ) | ( n21513 & ~n21514 ) ;
  assign n21516 = ( n21426 & n21506 ) | ( n21426 & n21515 ) | ( n21506 & n21515 ) ;
  assign n21517 = ( ~n21426 & n21506 ) | ( ~n21426 & n21515 ) | ( n21506 & n21515 ) ;
  assign n21518 = ( n21426 & ~n21516 ) | ( n21426 & n21517 ) | ( ~n21516 & n21517 ) ;
  assign n21519 = ( n21438 & n21470 ) | ( n21438 & n21518 ) | ( n21470 & n21518 ) ;
  assign n21520 = ( n21438 & ~n21470 ) | ( n21438 & n21518 ) | ( ~n21470 & n21518 ) ;
  assign n21521 = ( n21470 & ~n21519 ) | ( n21470 & n21520 ) | ( ~n21519 & n21520 ) ;
  assign n21522 = n4974 & ~n19472 ;
  assign n21523 = n4973 & n19157 ;
  assign n21524 = n4972 & ~n19309 ;
  assign n21525 = n21523 | n21524 ;
  assign n21526 = ~n21522 & n21525 ;
  assign n21527 = ( ~x20 & n21522 ) | ( ~x20 & n21526 ) | ( n21522 & n21526 ) ;
  assign n21528 = ( n21522 & n21526 ) | ( n21522 & ~n21527 ) | ( n21526 & ~n21527 ) ;
  assign n21529 = ( x20 & n21527 ) | ( x20 & ~n21528 ) | ( n21527 & ~n21528 ) ;
  assign n21530 = ( n21450 & n21521 ) | ( n21450 & n21529 ) | ( n21521 & n21529 ) ;
  assign n21531 = ( ~n21450 & n21521 ) | ( ~n21450 & n21529 ) | ( n21521 & n21529 ) ;
  assign n21532 = ( n21450 & ~n21530 ) | ( n21450 & n21531 ) | ( ~n21530 & n21531 ) ;
  assign n21533 = ( n21453 & n21456 ) | ( n21453 & n21532 ) | ( n21456 & n21532 ) ;
  assign n21534 = ( ~n21453 & n21456 ) | ( ~n21453 & n21532 ) | ( n21456 & n21532 ) ;
  assign n21535 = ( n21453 & ~n21533 ) | ( n21453 & n21534 ) | ( ~n21533 & n21534 ) ;
  assign n21536 = n21459 & n21535 ;
  assign n21537 = n21459 & ~n21535 ;
  assign n21538 = ( n21535 & ~n21536 ) | ( n21535 & n21537 ) | ( ~n21536 & n21537 ) ;
  assign n21539 = n1475 | n3374 ;
  assign n21540 = ( n6234 & n20458 ) | ( n6234 & ~n21539 ) | ( n20458 & ~n21539 ) ;
  assign n21541 = ( n1793 & n1915 ) | ( n1793 & ~n4397 ) | ( n1915 & ~n4397 ) ;
  assign n21542 = n4397 | n21541 ;
  assign n21543 = n3431 | n10250 ;
  assign n21544 = n197 | n295 ;
  assign n21545 = n361 | n1225 ;
  assign n21546 = ( n148 & n917 ) | ( n148 & ~n21545 ) | ( n917 & ~n21545 ) ;
  assign n21547 = n21545 | n21546 ;
  assign n21548 = ( n1024 & ~n21544 ) | ( n1024 & n21547 ) | ( ~n21544 & n21547 ) ;
  assign n21549 = n21544 | n21548 ;
  assign n21550 = ( ~n21542 & n21543 ) | ( ~n21542 & n21549 ) | ( n21543 & n21549 ) ;
  assign n21551 = n21542 | n21550 ;
  assign n21552 = ( n6234 & n21540 ) | ( n6234 & n21551 ) | ( n21540 & n21551 ) ;
  assign n21553 = n21540 & ~n21552 ;
  assign n21554 = n607 & ~n16029 ;
  assign n21555 = n1250 & ~n16027 ;
  assign n21556 = n21554 | n21555 ;
  assign n21557 = n606 & n16025 ;
  assign n21558 = ( n606 & n21556 ) | ( n606 & ~n21557 ) | ( n21556 & ~n21557 ) ;
  assign n21559 = n1248 & n17746 ;
  assign n21560 = ( n1248 & n21558 ) | ( n1248 & ~n21559 ) | ( n21558 & ~n21559 ) ;
  assign n21561 = ( n21498 & n21553 ) | ( n21498 & n21560 ) | ( n21553 & n21560 ) ;
  assign n21562 = ( n21498 & ~n21553 ) | ( n21498 & n21560 ) | ( ~n21553 & n21560 ) ;
  assign n21563 = ( n21553 & ~n21561 ) | ( n21553 & n21562 ) | ( ~n21561 & n21562 ) ;
  assign n21564 = n3800 & n18103 ;
  assign n21565 = n3799 & n16019 ;
  assign n21566 = n3700 & n16023 ;
  assign n21567 = n3802 & n16021 ;
  assign n21568 = n21566 | n21567 ;
  assign n21569 = ( ~n21564 & n21565 ) | ( ~n21564 & n21568 ) | ( n21565 & n21568 ) ;
  assign n21570 = ( ~x29 & n21564 ) | ( ~x29 & n21569 ) | ( n21564 & n21569 ) ;
  assign n21571 = ( n21564 & n21569 ) | ( n21564 & ~n21570 ) | ( n21569 & ~n21570 ) ;
  assign n21572 = ( x29 & n21570 ) | ( x29 & ~n21571 ) | ( n21570 & ~n21571 ) ;
  assign n21573 = ( ~n21501 & n21563 ) | ( ~n21501 & n21572 ) | ( n21563 & n21572 ) ;
  assign n21574 = ( n21563 & n21572 ) | ( n21563 & ~n21573 ) | ( n21572 & ~n21573 ) ;
  assign n21575 = ( n21501 & n21573 ) | ( n21501 & ~n21574 ) | ( n21573 & ~n21574 ) ;
  assign n21576 = n4202 & ~n18694 ;
  assign n21577 = n4201 & ~n16013 ;
  assign n21578 = n4200 & ~n16017 ;
  assign n21579 = n4345 & n16015 ;
  assign n21580 = n21578 | n21579 ;
  assign n21581 = ( ~n21576 & n21577 ) | ( ~n21576 & n21580 ) | ( n21577 & n21580 ) ;
  assign n21582 = ( ~x26 & n21576 ) | ( ~x26 & n21581 ) | ( n21576 & n21581 ) ;
  assign n21583 = ( n21576 & n21581 ) | ( n21576 & ~n21582 ) | ( n21581 & ~n21582 ) ;
  assign n21584 = ( x26 & n21582 ) | ( x26 & ~n21583 ) | ( n21582 & ~n21583 ) ;
  assign n21585 = ( n21504 & ~n21575 ) | ( n21504 & n21584 ) | ( ~n21575 & n21584 ) ;
  assign n21586 = ( n21504 & n21575 ) | ( n21504 & n21584 ) | ( n21575 & n21584 ) ;
  assign n21587 = ( n21575 & n21585 ) | ( n21575 & ~n21586 ) | ( n21585 & ~n21586 ) ;
  assign n21588 = n4713 & n19160 ;
  assign n21589 = n4712 & n19157 ;
  assign n21590 = n4709 & n16138 ;
  assign n21591 = n4792 & n18993 ;
  assign n21592 = n21590 | n21591 ;
  assign n21593 = ( ~n21588 & n21589 ) | ( ~n21588 & n21592 ) | ( n21589 & n21592 ) ;
  assign n21594 = ( ~x23 & n21588 ) | ( ~x23 & n21593 ) | ( n21588 & n21593 ) ;
  assign n21595 = ( n21588 & n21593 ) | ( n21588 & ~n21594 ) | ( n21593 & ~n21594 ) ;
  assign n21596 = ( x23 & n21594 ) | ( x23 & ~n21595 ) | ( n21594 & ~n21595 ) ;
  assign n21597 = ( n21516 & ~n21587 ) | ( n21516 & n21596 ) | ( ~n21587 & n21596 ) ;
  assign n21598 = ( n21516 & n21587 ) | ( n21516 & n21596 ) | ( n21587 & n21596 ) ;
  assign n21599 = ( n21587 & n21597 ) | ( n21587 & ~n21598 ) | ( n21597 & ~n21598 ) ;
  assign n21600 = n4973 & ~n19309 ;
  assign n21601 = ~x20 & n21600 ;
  assign n21602 = n21600 & ~n21601 ;
  assign n21603 = ( x20 & n21601 ) | ( x20 & ~n21602 ) | ( n21601 & ~n21602 ) ;
  assign n21604 = ( n21519 & ~n21599 ) | ( n21519 & n21603 ) | ( ~n21599 & n21603 ) ;
  assign n21605 = ( n21519 & n21599 ) | ( n21519 & n21603 ) | ( n21599 & n21603 ) ;
  assign n21606 = ( n21599 & n21604 ) | ( n21599 & ~n21605 ) | ( n21604 & ~n21605 ) ;
  assign n21607 = ( n21530 & n21533 ) | ( n21530 & ~n21606 ) | ( n21533 & ~n21606 ) ;
  assign n21608 = ( n21530 & n21533 ) | ( n21530 & n21606 ) | ( n21533 & n21606 ) ;
  assign n21609 = ( n21606 & n21607 ) | ( n21606 & ~n21608 ) | ( n21607 & ~n21608 ) ;
  assign n21610 = n21536 & ~n21609 ;
  assign n21611 = ~n21536 & n21609 ;
  assign n21612 = n21610 | n21611 ;
  assign n21613 = n1693 | n3484 ;
  assign n21614 = n878 | n960 ;
  assign n21615 = ( n1005 & n10189 ) | ( n1005 & ~n21614 ) | ( n10189 & ~n21614 ) ;
  assign n21616 = n21614 | n21615 ;
  assign n21617 = ( n21389 & ~n21613 ) | ( n21389 & n21616 ) | ( ~n21613 & n21616 ) ;
  assign n21618 = ( n10599 & n21613 ) | ( n10599 & ~n21617 ) | ( n21613 & ~n21617 ) ;
  assign n21619 = n21617 | n21618 ;
  assign n21620 = ( n4260 & n19919 ) | ( n4260 & ~n21619 ) | ( n19919 & ~n21619 ) ;
  assign n21621 = n21619 | n21620 ;
  assign n21622 = ( n1822 & n4605 ) | ( n1822 & n21621 ) | ( n4605 & n21621 ) ;
  assign n21623 = ( n4605 & ~n6191 ) | ( n4605 & n21622 ) | ( ~n6191 & n21622 ) ;
  assign n21624 = ~n21622 & n21623 ;
  assign n21625 = n607 & ~n16027 ;
  assign n21626 = n1250 & ~n16025 ;
  assign n21627 = n21625 | n21626 ;
  assign n21628 = n606 & ~n16023 ;
  assign n21629 = ( n606 & n21627 ) | ( n606 & ~n21628 ) | ( n21627 & ~n21628 ) ;
  assign n21630 = n1248 & ~n17968 ;
  assign n21631 = ( n1248 & n21629 ) | ( n1248 & ~n21630 ) | ( n21629 & ~n21630 ) ;
  assign n21632 = ( n21553 & ~n21624 ) | ( n21553 & n21631 ) | ( ~n21624 & n21631 ) ;
  assign n21633 = ( n21553 & n21624 ) | ( n21553 & n21631 ) | ( n21624 & n21631 ) ;
  assign n21634 = ( n21624 & n21632 ) | ( n21624 & ~n21633 ) | ( n21632 & ~n21633 ) ;
  assign n21635 = ( n21561 & n21573 ) | ( n21561 & ~n21634 ) | ( n21573 & ~n21634 ) ;
  assign n21636 = ( n21561 & ~n21573 ) | ( n21561 & n21634 ) | ( ~n21573 & n21634 ) ;
  assign n21637 = ( ~n21561 & n21635 ) | ( ~n21561 & n21636 ) | ( n21635 & n21636 ) ;
  assign n21638 = n4202 & ~n16144 ;
  assign n21639 = n4201 & n16138 ;
  assign n21640 = n4200 & n16015 ;
  assign n21641 = n4345 & ~n16013 ;
  assign n21642 = n21640 | n21641 ;
  assign n21643 = ( ~n21638 & n21639 ) | ( ~n21638 & n21642 ) | ( n21639 & n21642 ) ;
  assign n21644 = ( ~x26 & n21638 ) | ( ~x26 & n21643 ) | ( n21638 & n21643 ) ;
  assign n21645 = ( n21638 & n21643 ) | ( n21638 & ~n21644 ) | ( n21643 & ~n21644 ) ;
  assign n21646 = ( x26 & n21644 ) | ( x26 & ~n21645 ) | ( n21644 & ~n21645 ) ;
  assign n21647 = n3800 & ~n18267 ;
  assign n21648 = n3799 & ~n16017 ;
  assign n21649 = n3700 & n16021 ;
  assign n21650 = n3802 & n16019 ;
  assign n21651 = n21649 | n21650 ;
  assign n21652 = ( ~n21647 & n21648 ) | ( ~n21647 & n21651 ) | ( n21648 & n21651 ) ;
  assign n21653 = ( ~x29 & n21647 ) | ( ~x29 & n21652 ) | ( n21647 & n21652 ) ;
  assign n21654 = ( n21647 & n21652 ) | ( n21647 & ~n21653 ) | ( n21652 & ~n21653 ) ;
  assign n21655 = ( x29 & n21653 ) | ( x29 & ~n21654 ) | ( n21653 & ~n21654 ) ;
  assign n21656 = ( ~n21637 & n21646 ) | ( ~n21637 & n21655 ) | ( n21646 & n21655 ) ;
  assign n21657 = ( n21646 & n21655 ) | ( n21646 & ~n21656 ) | ( n21655 & ~n21656 ) ;
  assign n21658 = ( n21637 & n21656 ) | ( n21637 & ~n21657 ) | ( n21656 & ~n21657 ) ;
  assign n21659 = n4713 & ~n19312 ;
  assign n21660 = n4712 & ~n19309 ;
  assign n21661 = n4709 & n18993 ;
  assign n21662 = n4792 & n19157 ;
  assign n21663 = n21661 | n21662 ;
  assign n21664 = ( ~n21659 & n21660 ) | ( ~n21659 & n21663 ) | ( n21660 & n21663 ) ;
  assign n21665 = ( ~x23 & n21659 ) | ( ~x23 & n21664 ) | ( n21659 & n21664 ) ;
  assign n21666 = ( n21659 & n21664 ) | ( n21659 & ~n21665 ) | ( n21664 & ~n21665 ) ;
  assign n21667 = ( x23 & n21665 ) | ( x23 & ~n21666 ) | ( n21665 & ~n21666 ) ;
  assign n21668 = ( n21585 & ~n21658 ) | ( n21585 & n21667 ) | ( ~n21658 & n21667 ) ;
  assign n21669 = ( n21585 & n21658 ) | ( n21585 & n21667 ) | ( n21658 & n21667 ) ;
  assign n21670 = ( n21658 & n21668 ) | ( n21658 & ~n21669 ) | ( n21668 & ~n21669 ) ;
  assign n21671 = ( x20 & n21597 ) | ( x20 & ~n21670 ) | ( n21597 & ~n21670 ) ;
  assign n21672 = ( x20 & n21597 ) | ( x20 & n21670 ) | ( n21597 & n21670 ) ;
  assign n21673 = ( n21670 & n21671 ) | ( n21670 & ~n21672 ) | ( n21671 & ~n21672 ) ;
  assign n21674 = ( n21604 & n21607 ) | ( n21604 & ~n21673 ) | ( n21607 & ~n21673 ) ;
  assign n21675 = ( n21604 & n21607 ) | ( n21604 & n21673 ) | ( n21607 & n21673 ) ;
  assign n21676 = ( n21673 & n21674 ) | ( n21673 & ~n21675 ) | ( n21674 & ~n21675 ) ;
  assign n21677 = n21610 & ~n21676 ;
  assign n21678 = n21610 & n21676 ;
  assign n21679 = ( n21676 & n21677 ) | ( n21676 & ~n21678 ) | ( n21677 & ~n21678 ) ;
  assign n21680 = n4713 & ~n19472 ;
  assign n21681 = n4709 & n19157 ;
  assign n21682 = n4792 & ~n19309 ;
  assign n21683 = n21681 | n21682 ;
  assign n21684 = ~n21680 & n21683 ;
  assign n21685 = ( ~x23 & n21680 ) | ( ~x23 & n21684 ) | ( n21680 & n21684 ) ;
  assign n21686 = ( n21680 & n21684 ) | ( n21680 & ~n21685 ) | ( n21684 & ~n21685 ) ;
  assign n21687 = ( x23 & n21685 ) | ( x23 & ~n21686 ) | ( n21685 & ~n21686 ) ;
  assign n21688 = n3800 & ~n18416 ;
  assign n21689 = n3799 & n16015 ;
  assign n21690 = n3700 & n16019 ;
  assign n21691 = n3802 & ~n16017 ;
  assign n21692 = n21690 | n21691 ;
  assign n21693 = ( ~n21688 & n21689 ) | ( ~n21688 & n21692 ) | ( n21689 & n21692 ) ;
  assign n21694 = ( ~x29 & n21688 ) | ( ~x29 & n21693 ) | ( n21688 & n21693 ) ;
  assign n21695 = ( n21688 & n21693 ) | ( n21688 & ~n21694 ) | ( n21693 & ~n21694 ) ;
  assign n21696 = ( x29 & n21694 ) | ( x29 & ~n21695 ) | ( n21694 & ~n21695 ) ;
  assign n21697 = n3319 | n11375 ;
  assign n21698 = n2142 | n21697 ;
  assign n21699 = n1300 | n1835 ;
  assign n21700 = ( ~n1003 & n11899 ) | ( ~n1003 & n21699 ) | ( n11899 & n21699 ) ;
  assign n21701 = ~n21699 & n21700 ;
  assign n21702 = n1356 | n1515 ;
  assign n21703 = ( n1113 & n1564 ) | ( n1113 & ~n10517 ) | ( n1564 & ~n10517 ) ;
  assign n21704 = n10517 | n21703 ;
  assign n21705 = n241 | n562 ;
  assign n21706 = ( n298 & n783 ) | ( n298 & ~n21705 ) | ( n783 & ~n21705 ) ;
  assign n21707 = n21705 | n21706 ;
  assign n21708 = ( ~n21702 & n21704 ) | ( ~n21702 & n21707 ) | ( n21704 & n21707 ) ;
  assign n21709 = n21702 | n21708 ;
  assign n21710 = ( n21697 & n21701 ) | ( n21697 & ~n21709 ) | ( n21701 & ~n21709 ) ;
  assign n21711 = ( n4486 & ~n21698 ) | ( n4486 & n21710 ) | ( ~n21698 & n21710 ) ;
  assign n21712 = ~n4486 & n21711 ;
  assign n21713 = ( x20 & n21553 ) | ( x20 & n21712 ) | ( n21553 & n21712 ) ;
  assign n21714 = ( ~x20 & n21553 ) | ( ~x20 & n21712 ) | ( n21553 & n21712 ) ;
  assign n21715 = ( x20 & ~n21713 ) | ( x20 & n21714 ) | ( ~n21713 & n21714 ) ;
  assign n21716 = n607 & ~n16025 ;
  assign n21717 = n1250 & n16023 ;
  assign n21718 = n21716 | n21717 ;
  assign n21719 = n606 & ~n16021 ;
  assign n21720 = ( n606 & n21718 ) | ( n606 & ~n21719 ) | ( n21718 & ~n21719 ) ;
  assign n21721 = n1248 & ~n18091 ;
  assign n21722 = n21720 | n21721 ;
  assign n21723 = ( n21632 & ~n21715 ) | ( n21632 & n21722 ) | ( ~n21715 & n21722 ) ;
  assign n21724 = ( n21632 & n21715 ) | ( n21632 & n21722 ) | ( n21715 & n21722 ) ;
  assign n21725 = ( n21715 & n21723 ) | ( n21715 & ~n21724 ) | ( n21723 & ~n21724 ) ;
  assign n21726 = ( n21635 & n21696 ) | ( n21635 & ~n21725 ) | ( n21696 & ~n21725 ) ;
  assign n21727 = ( ~n21635 & n21696 ) | ( ~n21635 & n21725 ) | ( n21696 & n21725 ) ;
  assign n21728 = ( ~n21696 & n21726 ) | ( ~n21696 & n21727 ) | ( n21726 & n21727 ) ;
  assign n21729 = n4202 & n18996 ;
  assign n21730 = n4201 & n18993 ;
  assign n21731 = n4200 & ~n16013 ;
  assign n21732 = n4345 & n16138 ;
  assign n21733 = n21731 | n21732 ;
  assign n21734 = ( ~n21729 & n21730 ) | ( ~n21729 & n21733 ) | ( n21730 & n21733 ) ;
  assign n21735 = ( ~x26 & n21729 ) | ( ~x26 & n21734 ) | ( n21729 & n21734 ) ;
  assign n21736 = ( n21729 & n21734 ) | ( n21729 & ~n21735 ) | ( n21734 & ~n21735 ) ;
  assign n21737 = ( x26 & n21735 ) | ( x26 & ~n21736 ) | ( n21735 & ~n21736 ) ;
  assign n21738 = ( n21656 & ~n21728 ) | ( n21656 & n21737 ) | ( ~n21728 & n21737 ) ;
  assign n21739 = ( n21656 & n21728 ) | ( n21656 & n21737 ) | ( n21728 & n21737 ) ;
  assign n21740 = ( n21728 & n21738 ) | ( n21728 & ~n21739 ) | ( n21738 & ~n21739 ) ;
  assign n21741 = ( n21668 & n21687 ) | ( n21668 & ~n21740 ) | ( n21687 & ~n21740 ) ;
  assign n21742 = ( ~n21668 & n21687 ) | ( ~n21668 & n21740 ) | ( n21687 & n21740 ) ;
  assign n21743 = ( ~n21687 & n21741 ) | ( ~n21687 & n21742 ) | ( n21741 & n21742 ) ;
  assign n21744 = ( n21671 & n21674 ) | ( n21671 & ~n21743 ) | ( n21674 & ~n21743 ) ;
  assign n21745 = ( n21671 & n21674 ) | ( n21671 & n21743 ) | ( n21674 & n21743 ) ;
  assign n21746 = ( n21743 & n21744 ) | ( n21743 & ~n21745 ) | ( n21744 & ~n21745 ) ;
  assign n21747 = n21677 & ~n21746 ;
  assign n21748 = ~n21677 & n21746 ;
  assign n21749 = n21747 | n21748 ;
  assign n21750 = n607 & n16023 ;
  assign n21751 = n1250 & n16021 ;
  assign n21752 = n21750 | n21751 ;
  assign n21753 = n606 & ~n16019 ;
  assign n21754 = ( n606 & n21752 ) | ( n606 & ~n21753 ) | ( n21752 & ~n21753 ) ;
  assign n21755 = n1248 & ~n18103 ;
  assign n21756 = ( n1248 & n21754 ) | ( n1248 & ~n21755 ) | ( n21754 & ~n21755 ) ;
  assign n21757 = ( n112 & n952 ) | ( n112 & ~n1556 ) | ( n952 & ~n1556 ) ;
  assign n21758 = n1556 | n21757 ;
  assign n21759 = ( n686 & ~n2558 ) | ( n686 & n21758 ) | ( ~n2558 & n21758 ) ;
  assign n21760 = ( n1560 & n2558 ) | ( n1560 & ~n21759 ) | ( n2558 & ~n21759 ) ;
  assign n21761 = n21759 | n21760 ;
  assign n21762 = ( n3986 & ~n11815 ) | ( n3986 & n21761 ) | ( ~n11815 & n21761 ) ;
  assign n21763 = n2683 | n4872 ;
  assign n21764 = ( n2610 & n11939 ) | ( n2610 & ~n21763 ) | ( n11939 & ~n21763 ) ;
  assign n21765 = n21763 | n21764 ;
  assign n21766 = ( n11815 & ~n21762 ) | ( n11815 & n21765 ) | ( ~n21762 & n21765 ) ;
  assign n21767 = n21762 | n21766 ;
  assign n21768 = n2659 | n4269 ;
  assign n21769 = ( n10118 & ~n21767 ) | ( n10118 & n21768 ) | ( ~n21767 & n21768 ) ;
  assign n21770 = n21767 | n21769 ;
  assign n21771 = ( n21713 & n21756 ) | ( n21713 & n21770 ) | ( n21756 & n21770 ) ;
  assign n21772 = ( n21713 & ~n21756 ) | ( n21713 & n21770 ) | ( ~n21756 & n21770 ) ;
  assign n21773 = ( n21756 & ~n21771 ) | ( n21756 & n21772 ) | ( ~n21771 & n21772 ) ;
  assign n21774 = n3800 & ~n18694 ;
  assign n21775 = n3799 & ~n16013 ;
  assign n21776 = n3700 & ~n16017 ;
  assign n21777 = n3802 & n16015 ;
  assign n21778 = n21776 | n21777 ;
  assign n21779 = ( ~n21774 & n21775 ) | ( ~n21774 & n21778 ) | ( n21775 & n21778 ) ;
  assign n21780 = ( ~x29 & n21774 ) | ( ~x29 & n21779 ) | ( n21774 & n21779 ) ;
  assign n21781 = ( n21774 & n21779 ) | ( n21774 & ~n21780 ) | ( n21779 & ~n21780 ) ;
  assign n21782 = ( x29 & n21780 ) | ( x29 & ~n21781 ) | ( n21780 & ~n21781 ) ;
  assign n21783 = ( n21723 & n21773 ) | ( n21723 & n21782 ) | ( n21773 & n21782 ) ;
  assign n21784 = ( ~n21723 & n21773 ) | ( ~n21723 & n21782 ) | ( n21773 & n21782 ) ;
  assign n21785 = ( n21723 & ~n21783 ) | ( n21723 & n21784 ) | ( ~n21783 & n21784 ) ;
  assign n21786 = n4202 & n19160 ;
  assign n21787 = n4201 & n19157 ;
  assign n21788 = n4200 & n16138 ;
  assign n21789 = n4345 & n18993 ;
  assign n21790 = n21788 | n21789 ;
  assign n21791 = ( ~n21786 & n21787 ) | ( ~n21786 & n21790 ) | ( n21787 & n21790 ) ;
  assign n21792 = ( ~x26 & n21786 ) | ( ~x26 & n21791 ) | ( n21786 & n21791 ) ;
  assign n21793 = ( n21786 & n21791 ) | ( n21786 & ~n21792 ) | ( n21791 & ~n21792 ) ;
  assign n21794 = ( x26 & n21792 ) | ( x26 & ~n21793 ) | ( n21792 & ~n21793 ) ;
  assign n21795 = ( n21726 & n21785 ) | ( n21726 & n21794 ) | ( n21785 & n21794 ) ;
  assign n21796 = ( n21726 & ~n21785 ) | ( n21726 & n21794 ) | ( ~n21785 & n21794 ) ;
  assign n21797 = ( n21785 & ~n21795 ) | ( n21785 & n21796 ) | ( ~n21795 & n21796 ) ;
  assign n21798 = n4709 & ~n19309 ;
  assign n21799 = ~x23 & n21798 ;
  assign n21800 = n21798 & ~n21799 ;
  assign n21801 = ( x23 & n21799 ) | ( x23 & ~n21800 ) | ( n21799 & ~n21800 ) ;
  assign n21802 = ( n21738 & n21797 ) | ( n21738 & n21801 ) | ( n21797 & n21801 ) ;
  assign n21803 = ( ~n21738 & n21797 ) | ( ~n21738 & n21801 ) | ( n21797 & n21801 ) ;
  assign n21804 = ( n21738 & ~n21802 ) | ( n21738 & n21803 ) | ( ~n21802 & n21803 ) ;
  assign n21805 = ( n21741 & n21744 ) | ( n21741 & n21804 ) | ( n21744 & n21804 ) ;
  assign n21806 = ( ~n21741 & n21744 ) | ( ~n21741 & n21804 ) | ( n21744 & n21804 ) ;
  assign n21807 = ( n21741 & ~n21805 ) | ( n21741 & n21806 ) | ( ~n21805 & n21806 ) ;
  assign n21808 = n21747 & n21807 ;
  assign n21809 = n21747 & ~n21807 ;
  assign n21810 = ( n21807 & ~n21808 ) | ( n21807 & n21809 ) | ( ~n21808 & n21809 ) ;
  assign n21811 = n309 | n1155 ;
  assign n21812 = n686 | n2207 ;
  assign n21813 = n172 | n1005 ;
  assign n21814 = ( n913 & n1085 ) | ( n913 & ~n21813 ) | ( n1085 & ~n21813 ) ;
  assign n21815 = n21813 | n21814 ;
  assign n21816 = n356 | n885 ;
  assign n21817 = ( n713 & n1341 ) | ( n713 & ~n21816 ) | ( n1341 & ~n21816 ) ;
  assign n21818 = n21816 | n21817 ;
  assign n21819 = ( ~n21812 & n21815 ) | ( ~n21812 & n21818 ) | ( n21815 & n21818 ) ;
  assign n21820 = n21812 | n21819 ;
  assign n21821 = ( n10259 & n12006 ) | ( n10259 & ~n21820 ) | ( n12006 & ~n21820 ) ;
  assign n21822 = n21820 | n21821 ;
  assign n21823 = ( ~n309 & n20464 ) | ( ~n309 & n21822 ) | ( n20464 & n21822 ) ;
  assign n21824 = ( n18165 & n21811 ) | ( n18165 & n21823 ) | ( n21811 & n21823 ) ;
  assign n21825 = n18165 & ~n21824 ;
  assign n21826 = ( n21770 & ~n21772 ) | ( n21770 & n21825 ) | ( ~n21772 & n21825 ) ;
  assign n21827 = ( n21713 & ~n21771 ) | ( n21713 & n21825 ) | ( ~n21771 & n21825 ) ;
  assign n21828 = ( ~n21825 & n21826 ) | ( ~n21825 & n21827 ) | ( n21826 & n21827 ) ;
  assign n21829 = n607 & n16021 ;
  assign n21830 = n1250 & n16019 ;
  assign n21831 = n21829 | n21830 ;
  assign n21832 = n606 & n16017 ;
  assign n21833 = ( n606 & n21831 ) | ( n606 & ~n21832 ) | ( n21831 & ~n21832 ) ;
  assign n21834 = n1248 & n18267 ;
  assign n21835 = ( n1248 & n21833 ) | ( n1248 & ~n21834 ) | ( n21833 & ~n21834 ) ;
  assign n21836 = ( n21783 & ~n21828 ) | ( n21783 & n21835 ) | ( ~n21828 & n21835 ) ;
  assign n21837 = ( n21783 & n21828 ) | ( n21783 & n21835 ) | ( n21828 & n21835 ) ;
  assign n21838 = ( n21828 & n21836 ) | ( n21828 & ~n21837 ) | ( n21836 & ~n21837 ) ;
  assign n21839 = n4202 & ~n19312 ;
  assign n21840 = n4201 & ~n19309 ;
  assign n21841 = n4200 & n18993 ;
  assign n21842 = n4345 & n19157 ;
  assign n21843 = n21841 | n21842 ;
  assign n21844 = ( ~n21839 & n21840 ) | ( ~n21839 & n21843 ) | ( n21840 & n21843 ) ;
  assign n21845 = ( ~x26 & n21839 ) | ( ~x26 & n21844 ) | ( n21839 & n21844 ) ;
  assign n21846 = ( n21839 & n21844 ) | ( n21839 & ~n21845 ) | ( n21844 & ~n21845 ) ;
  assign n21847 = ( x26 & n21845 ) | ( x26 & ~n21846 ) | ( n21845 & ~n21846 ) ;
  assign n21848 = n3800 & ~n16144 ;
  assign n21849 = n3799 & n16138 ;
  assign n21850 = n3700 & n16015 ;
  assign n21851 = n3802 & ~n16013 ;
  assign n21852 = n21850 | n21851 ;
  assign n21853 = ( ~n21848 & n21849 ) | ( ~n21848 & n21852 ) | ( n21849 & n21852 ) ;
  assign n21854 = ( ~x29 & n21848 ) | ( ~x29 & n21853 ) | ( n21848 & n21853 ) ;
  assign n21855 = ( n21848 & n21853 ) | ( n21848 & ~n21854 ) | ( n21853 & ~n21854 ) ;
  assign n21856 = ( x29 & n21854 ) | ( x29 & ~n21855 ) | ( n21854 & ~n21855 ) ;
  assign n21857 = ( ~n21838 & n21847 ) | ( ~n21838 & n21856 ) | ( n21847 & n21856 ) ;
  assign n21858 = ( n21847 & n21856 ) | ( n21847 & ~n21857 ) | ( n21856 & ~n21857 ) ;
  assign n21859 = ( n21838 & n21857 ) | ( n21838 & ~n21858 ) | ( n21857 & ~n21858 ) ;
  assign n21860 = ( x23 & n21795 ) | ( x23 & ~n21859 ) | ( n21795 & ~n21859 ) ;
  assign n21861 = ( x23 & n21795 ) | ( x23 & n21859 ) | ( n21795 & n21859 ) ;
  assign n21862 = ( n21859 & n21860 ) | ( n21859 & ~n21861 ) | ( n21860 & ~n21861 ) ;
  assign n21863 = ( n21802 & n21805 ) | ( n21802 & ~n21862 ) | ( n21805 & ~n21862 ) ;
  assign n21864 = ( n21802 & n21805 ) | ( n21802 & n21862 ) | ( n21805 & n21862 ) ;
  assign n21865 = ( n21862 & n21863 ) | ( n21862 & ~n21864 ) | ( n21863 & ~n21864 ) ;
  assign n21866 = n21808 & ~n21865 ;
  assign n21867 = ~n21808 & n21865 ;
  assign n21868 = n21866 | n21867 ;
  assign n21869 = n4202 & ~n19472 ;
  assign n21870 = n4200 & n19157 ;
  assign n21871 = n4345 & ~n19309 ;
  assign n21872 = n21870 | n21871 ;
  assign n21873 = ~n21869 & n21872 ;
  assign n21874 = ( ~x26 & n21869 ) | ( ~x26 & n21873 ) | ( n21869 & n21873 ) ;
  assign n21875 = ( n21869 & n21873 ) | ( n21869 & ~n21874 ) | ( n21873 & ~n21874 ) ;
  assign n21876 = ( x26 & n21874 ) | ( x26 & ~n21875 ) | ( n21874 & ~n21875 ) ;
  assign n21877 = n344 & ~n400 ;
  assign n21878 = ( n66 & n83 ) | ( n66 & n97 ) | ( n83 & n97 ) ;
  assign n21879 = ( n51 & n500 ) | ( n51 & ~n21878 ) | ( n500 & ~n21878 ) ;
  assign n21880 = n21878 | n21879 ;
  assign n21881 = n1056 | n4847 ;
  assign n21882 = n21880 | n21881 ;
  assign n21883 = ( n48 & n75 ) | ( n48 & n145 ) | ( n75 & n145 ) ;
  assign n21884 = n630 | n21883 ;
  assign n21885 = ( ~n69 & n11993 ) | ( ~n69 & n21884 ) | ( n11993 & n21884 ) ;
  assign n21886 = n69 | n21885 ;
  assign n21887 = ( ~n400 & n21882 ) | ( ~n400 & n21886 ) | ( n21882 & n21886 ) ;
  assign n21888 = ( n9887 & n21877 ) | ( n9887 & ~n21887 ) | ( n21877 & ~n21887 ) ;
  assign n21889 = ~n9887 & n21888 ;
  assign n21890 = ( x23 & n21825 ) | ( x23 & n21889 ) | ( n21825 & n21889 ) ;
  assign n21891 = ( ~x23 & n21825 ) | ( ~x23 & n21889 ) | ( n21825 & n21889 ) ;
  assign n21892 = ( x23 & ~n21890 ) | ( x23 & n21891 ) | ( ~n21890 & n21891 ) ;
  assign n21893 = n607 & n16019 ;
  assign n21894 = n1250 & ~n16017 ;
  assign n21895 = n21893 | n21894 ;
  assign n21896 = n606 & ~n16015 ;
  assign n21897 = ( n606 & n21895 ) | ( n606 & ~n21896 ) | ( n21895 & ~n21896 ) ;
  assign n21898 = n1248 & n18416 ;
  assign n21899 = ( n1248 & n21897 ) | ( n1248 & ~n21898 ) | ( n21897 & ~n21898 ) ;
  assign n21900 = ( n21826 & ~n21892 ) | ( n21826 & n21899 ) | ( ~n21892 & n21899 ) ;
  assign n21901 = ( n21826 & n21892 ) | ( n21826 & n21899 ) | ( n21892 & n21899 ) ;
  assign n21902 = ( n21892 & n21900 ) | ( n21892 & ~n21901 ) | ( n21900 & ~n21901 ) ;
  assign n21903 = n3800 & n18996 ;
  assign n21904 = n3799 & n18993 ;
  assign n21905 = n3700 & ~n16013 ;
  assign n21906 = n3802 & n16138 ;
  assign n21907 = n21905 | n21906 ;
  assign n21908 = ( ~n21903 & n21904 ) | ( ~n21903 & n21907 ) | ( n21904 & n21907 ) ;
  assign n21909 = ( ~x29 & n21903 ) | ( ~x29 & n21908 ) | ( n21903 & n21908 ) ;
  assign n21910 = ( n21903 & n21908 ) | ( n21903 & ~n21909 ) | ( n21908 & ~n21909 ) ;
  assign n21911 = ( x29 & n21909 ) | ( x29 & ~n21910 ) | ( n21909 & ~n21910 ) ;
  assign n21912 = ( n21836 & ~n21902 ) | ( n21836 & n21911 ) | ( ~n21902 & n21911 ) ;
  assign n21913 = ( n21836 & n21902 ) | ( n21836 & n21911 ) | ( n21902 & n21911 ) ;
  assign n21914 = ( n21902 & n21912 ) | ( n21902 & ~n21913 ) | ( n21912 & ~n21913 ) ;
  assign n21915 = ( n21857 & n21876 ) | ( n21857 & ~n21914 ) | ( n21876 & ~n21914 ) ;
  assign n21916 = ( ~n21857 & n21876 ) | ( ~n21857 & n21914 ) | ( n21876 & n21914 ) ;
  assign n21917 = ( ~n21876 & n21915 ) | ( ~n21876 & n21916 ) | ( n21915 & n21916 ) ;
  assign n21918 = ( n21860 & n21863 ) | ( n21860 & ~n21917 ) | ( n21863 & ~n21917 ) ;
  assign n21919 = ( n21860 & n21863 ) | ( n21860 & n21917 ) | ( n21863 & n21917 ) ;
  assign n21920 = ( n21917 & n21918 ) | ( n21917 & ~n21919 ) | ( n21918 & ~n21919 ) ;
  assign n21921 = n21866 & ~n21920 ;
  assign n21922 = n21866 & n21920 ;
  assign n21923 = ( n21920 & n21921 ) | ( n21920 & ~n21922 ) | ( n21921 & ~n21922 ) ;
  assign n21924 = n241 | n313 ;
  assign n21925 = n112 | n21924 ;
  assign n21926 = n782 | n1323 ;
  assign n21927 = ( n648 & n836 ) | ( n648 & ~n21926 ) | ( n836 & ~n21926 ) ;
  assign n21928 = n21926 | n21927 ;
  assign n21929 = ( ~n325 & n21925 ) | ( ~n325 & n21928 ) | ( n21925 & n21928 ) ;
  assign n21930 = n690 | n2680 ;
  assign n21931 = n4114 | n21930 ;
  assign n21932 = n6116 | n11407 ;
  assign n21933 = n21931 | n21932 ;
  assign n21934 = ( n325 & ~n21929 ) | ( n325 & n21933 ) | ( ~n21929 & n21933 ) ;
  assign n21935 = n21929 | n21934 ;
  assign n21936 = n414 | n1229 ;
  assign n21937 = ( n12003 & ~n21935 ) | ( n12003 & n21936 ) | ( ~n21935 & n21936 ) ;
  assign n21938 = n21935 | n21937 ;
  assign n21939 = n1248 & n18694 ;
  assign n21940 = n607 & ~n16017 ;
  assign n21941 = ( n606 & ~n16013 ) | ( n606 & n21940 ) | ( ~n16013 & n21940 ) ;
  assign n21942 = n1250 & ~n16015 ;
  assign n21943 = ( n1250 & n21941 ) | ( n1250 & ~n21942 ) | ( n21941 & ~n21942 ) ;
  assign n21944 = ( n1248 & ~n21939 ) | ( n1248 & n21943 ) | ( ~n21939 & n21943 ) ;
  assign n21945 = ( n21890 & n21938 ) | ( n21890 & ~n21944 ) | ( n21938 & ~n21944 ) ;
  assign n21946 = ( ~n21890 & n21938 ) | ( ~n21890 & n21944 ) | ( n21938 & n21944 ) ;
  assign n21947 = ( ~n21938 & n21945 ) | ( ~n21938 & n21946 ) | ( n21945 & n21946 ) ;
  assign n21948 = n3800 & n19160 ;
  assign n21949 = n3799 & n19157 ;
  assign n21950 = n3700 & n16138 ;
  assign n21951 = ( n3802 & n18993 ) | ( n3802 & n21950 ) | ( n18993 & n21950 ) ;
  assign n21952 = ( ~n21948 & n21949 ) | ( ~n21948 & n21951 ) | ( n21949 & n21951 ) ;
  assign n21953 = ( ~x29 & n21948 ) | ( ~x29 & n21952 ) | ( n21948 & n21952 ) ;
  assign n21954 = ( n21948 & n21952 ) | ( n21948 & ~n21953 ) | ( n21952 & ~n21953 ) ;
  assign n21955 = ( x29 & n21953 ) | ( x29 & ~n21954 ) | ( n21953 & ~n21954 ) ;
  assign n21956 = ( n21900 & n21947 ) | ( n21900 & n21955 ) | ( n21947 & n21955 ) ;
  assign n21957 = ( ~n21900 & n21947 ) | ( ~n21900 & n21955 ) | ( n21947 & n21955 ) ;
  assign n21958 = ( n21900 & ~n21956 ) | ( n21900 & n21957 ) | ( ~n21956 & n21957 ) ;
  assign n21959 = n4200 & ~n19309 ;
  assign n21960 = ~x26 & n21959 ;
  assign n21961 = n21959 & ~n21960 ;
  assign n21962 = ( x26 & n21960 ) | ( x26 & ~n21961 ) | ( n21960 & ~n21961 ) ;
  assign n21963 = ( n21912 & n21958 ) | ( n21912 & n21962 ) | ( n21958 & n21962 ) ;
  assign n21964 = ( n21912 & ~n21958 ) | ( n21912 & n21962 ) | ( ~n21958 & n21962 ) ;
  assign n21965 = ( n21958 & ~n21963 ) | ( n21958 & n21964 ) | ( ~n21963 & n21964 ) ;
  assign n21966 = ( n21915 & n21918 ) | ( n21915 & n21965 ) | ( n21918 & n21965 ) ;
  assign n21967 = ( ~n21915 & n21918 ) | ( ~n21915 & n21965 ) | ( n21918 & n21965 ) ;
  assign n21968 = ( n21915 & ~n21966 ) | ( n21915 & n21967 ) | ( ~n21966 & n21967 ) ;
  assign n21969 = n21921 & n21968 ;
  assign n21970 = n21921 | n21968 ;
  assign n21971 = ~n21969 & n21970 ;
  assign n21972 = n1273 | n3086 ;
  assign n21973 = ( n366 & ~n3651 ) | ( n366 & n10293 ) | ( ~n3651 & n10293 ) ;
  assign n21974 = n3651 | n21973 ;
  assign n21975 = ( n3641 & n21972 ) | ( n3641 & ~n21974 ) | ( n21972 & ~n21974 ) ;
  assign n21976 = ( n414 & n21972 ) | ( n414 & n21975 ) | ( n21972 & n21975 ) ;
  assign n21977 = n21975 & ~n21976 ;
  assign n21978 = ( n21938 & n21945 ) | ( n21938 & n21977 ) | ( n21945 & n21977 ) ;
  assign n21979 = ( ~n21938 & n21945 ) | ( ~n21938 & n21977 ) | ( n21945 & n21977 ) ;
  assign n21980 = ( n21938 & ~n21978 ) | ( n21938 & n21979 ) | ( ~n21978 & n21979 ) ;
  assign n21981 = n607 & n16015 ;
  assign n21982 = n1250 & ~n16013 ;
  assign n21983 = n21981 | n21982 ;
  assign n21984 = n606 & ~n16138 ;
  assign n21985 = ( n606 & n21983 ) | ( n606 & ~n21984 ) | ( n21983 & ~n21984 ) ;
  assign n21986 = n1248 & n16144 ;
  assign n21987 = ( n1248 & n21985 ) | ( n1248 & ~n21986 ) | ( n21985 & ~n21986 ) ;
  assign n21988 = ( n21956 & ~n21980 ) | ( n21956 & n21987 ) | ( ~n21980 & n21987 ) ;
  assign n21989 = ( n21956 & n21980 ) | ( n21956 & n21987 ) | ( n21980 & n21987 ) ;
  assign n21990 = ( n21980 & n21988 ) | ( n21980 & ~n21989 ) | ( n21988 & ~n21989 ) ;
  assign n21991 = n3800 & ~n19312 ;
  assign n21992 = n3799 & ~n19309 ;
  assign n21993 = n3700 & n18993 ;
  assign n21994 = n3802 & n19157 ;
  assign n21995 = n21993 | n21994 ;
  assign n21996 = ( ~n21991 & n21992 ) | ( ~n21991 & n21995 ) | ( n21992 & n21995 ) ;
  assign n21997 = ( ~x29 & n21991 ) | ( ~x29 & n21996 ) | ( n21991 & n21996 ) ;
  assign n21998 = ( n21991 & n21996 ) | ( n21991 & ~n21997 ) | ( n21996 & ~n21997 ) ;
  assign n21999 = ( x29 & n21997 ) | ( x29 & ~n21998 ) | ( n21997 & ~n21998 ) ;
  assign n22000 = x26 & n21999 ;
  assign n22001 = x26 | n21999 ;
  assign n22002 = ~n22000 & n22001 ;
  assign n22003 = ~n21990 & n22002 ;
  assign n22004 = ( n21990 & n22000 ) | ( n21990 & ~n22001 ) | ( n22000 & ~n22001 ) ;
  assign n22005 = n22003 | n22004 ;
  assign n22006 = ( n21963 & n21966 ) | ( n21963 & ~n22005 ) | ( n21966 & ~n22005 ) ;
  assign n22007 = ( n21963 & n21966 ) | ( n21963 & n22005 ) | ( n21966 & n22005 ) ;
  assign n22008 = ( n22005 & n22006 ) | ( n22005 & ~n22007 ) | ( n22006 & ~n22007 ) ;
  assign n22009 = n21969 & ~n22008 ;
  assign n22010 = n21969 & n22008 ;
  assign n22011 = ( n22008 & n22009 ) | ( n22008 & ~n22010 ) | ( n22009 & ~n22010 ) ;
  assign n22012 = ( ~n22000 & n22003 ) | ( ~n22000 & n22006 ) | ( n22003 & n22006 ) ;
  assign n22013 = ( n22003 & n22006 ) | ( n22003 & ~n22012 ) | ( n22006 & ~n22012 ) ;
  assign n22014 = ( n22000 & n22012 ) | ( n22000 & ~n22013 ) | ( n22012 & ~n22013 ) ;
  assign n22015 = n3656 | n3688 ;
  assign n22016 = n3700 & n19157 ;
  assign n22017 = n3800 & ~n19472 ;
  assign n22018 = n22016 | n22017 ;
  assign n22019 = n607 & ~n16013 ;
  assign n22020 = n1250 & n16138 ;
  assign n22021 = n22019 | n22020 ;
  assign n22022 = n606 & ~n18993 ;
  assign n22023 = ( n606 & n22021 ) | ( n606 & ~n22022 ) | ( n22021 & ~n22022 ) ;
  assign n22024 = n1248 & ~n18996 ;
  assign n22025 = ( n1248 & n22023 ) | ( n1248 & ~n22024 ) | ( n22023 & ~n22024 ) ;
  assign n22026 = ( ~x29 & n22018 ) | ( ~x29 & n22025 ) | ( n22018 & n22025 ) ;
  assign n22027 = ( n22018 & n22025 ) | ( n22018 & ~n22026 ) | ( n22025 & ~n22026 ) ;
  assign n22028 = ( x29 & n22026 ) | ( x29 & ~n22027 ) | ( n22026 & ~n22027 ) ;
  assign n22029 = ( ~n21978 & n21988 ) | ( ~n21978 & n22028 ) | ( n21988 & n22028 ) ;
  assign n22030 = ( n21988 & n22028 ) | ( n21988 & ~n22029 ) | ( n22028 & ~n22029 ) ;
  assign n22031 = ( n21978 & n22029 ) | ( n21978 & ~n22030 ) | ( n22029 & ~n22030 ) ;
  assign n22032 = ( ~x26 & n22015 ) | ( ~x26 & n22031 ) | ( n22015 & n22031 ) ;
  assign n22033 = ( n22015 & n22031 ) | ( n22015 & ~n22032 ) | ( n22031 & ~n22032 ) ;
  assign n22034 = ( x26 & n22032 ) | ( x26 & ~n22033 ) | ( n22032 & ~n22033 ) ;
  assign n22035 = ( ~n21938 & n22014 ) | ( ~n21938 & n22034 ) | ( n22014 & n22034 ) ;
  assign n22036 = ( n22014 & n22034 ) | ( n22014 & ~n22035 ) | ( n22034 & ~n22035 ) ;
  assign n22037 = ( n21938 & n22035 ) | ( n21938 & ~n22036 ) | ( n22035 & ~n22036 ) ;
  assign n22038 = ~n22009 & n22037 ;
  assign n22039 = n22037 & ~n22038 ;
  assign n22040 = ( n22009 & n22038 ) | ( n22009 & ~n22039 ) | ( n22038 & ~n22039 ) ;
  assign y0 = n18843 ;
  assign y1 = n19011 ;
  assign y2 = ~n19175 ;
  assign y3 = ~n19327 ;
  assign y4 = ~n19485 ;
  assign y5 = ~n19628 ;
  assign y6 = ~n19775 ;
  assign y7 = ~n19914 ;
  assign y8 = n20055 ;
  assign y9 = n20185 ;
  assign y10 = n20313 ;
  assign y11 = n20447 ;
  assign y12 = ~n20579 ;
  assign y13 = ~n20694 ;
  assign y14 = ~n20802 ;
  assign y15 = n20908 ;
  assign y16 = ~n21012 ;
  assign y17 = n21108 ;
  assign y18 = ~n21204 ;
  assign y19 = ~n21292 ;
  assign y20 = ~n21378 ;
  assign y21 = n21461 ;
  assign y22 = n21538 ;
  assign y23 = ~n21612 ;
  assign y24 = ~n21679 ;
  assign y25 = ~n21749 ;
  assign y26 = n21810 ;
  assign y27 = ~n21868 ;
  assign y28 = ~n21923 ;
  assign y29 = n21971 ;
  assign y30 = ~n22011 ;
  assign y31 = n22040 ;
endmodule
