module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n8 = ( x2 & ~x3 ) | ( x2 & x4 ) | ( ~x3 & x4 ) ;
  assign n9 = ~x4 & n8 ;
  assign n10 = x1 & n9 ;
  assign n11 = x0 | x1 ;
  assign n12 = x2 | n11 ;
  assign n13 = x3 & x4 ;
  assign n14 = ( n10 & n12 ) | ( n10 & n13 ) | ( n12 & n13 ) ;
  assign n15 = x0 & ~x1 ;
  assign n16 = ~x3 & x4 ;
  assign n17 = ~x2 & n16 ;
  assign n18 = ~x0 & n17 ;
  assign n19 = ~x2 & x4 ;
  assign n20 = ( ~x2 & x3 ) | ( ~x2 & x4 ) | ( x3 & x4 ) ;
  assign n21 = x0 & x1 ;
  assign n22 = n13 & ~n21 ;
  assign n23 = x2 & n22 ;
  assign n24 = ( n20 & ~n22 ) | ( n20 & n23 ) | ( ~n22 & n23 ) ;
  assign n25 = ( x1 & x4 ) | ( x1 & n24 ) | ( x4 & n24 ) ;
  assign n26 = ( ~x4 & n8 ) | ( ~x4 & n13 ) | ( n8 & n13 ) ;
  assign n27 = ( x1 & n18 ) | ( x1 & n26 ) | ( n18 & n26 ) ;
  assign n28 = ( n19 & ~n25 ) | ( n19 & n27 ) | ( ~n25 & n27 ) ;
  assign n29 = ( n17 & ~n18 ) | ( n17 & n28 ) | ( ~n18 & n28 ) ;
  assign n30 = ( n10 & ~n15 ) | ( n10 & n29 ) | ( ~n15 & n29 ) ;
  assign n31 = x3 & ~x4 ;
  assign n32 = x1 & n31 ;
  assign n33 = ~x2 & x3 ;
  assign n34 = ( ~n14 & n16 ) | ( ~n14 & n33 ) | ( n16 & n33 ) ;
  assign n35 = ( n28 & n32 ) | ( n28 & n34 ) | ( n32 & n34 ) ;
  assign n36 = ~n32 & n34 ;
  assign n37 = x0 & x2 ;
  assign n38 = n16 & n37 ;
  assign n39 = ( x1 & n16 ) | ( x1 & n33 ) | ( n16 & n33 ) ;
  assign n40 = ( ~x6 & n17 ) | ( ~x6 & n19 ) | ( n17 & n19 ) ;
  assign n41 = n39 & ~n40 ;
  assign n42 = x0 & n41 ;
  assign n43 = x5 & n39 ;
  assign n44 = ( ~x4 & n33 ) | ( ~x4 & n43 ) | ( n33 & n43 ) ;
  assign n45 = ( n22 & n42 ) | ( n22 & n44 ) | ( n42 & n44 ) ;
  assign n46 = n38 | n45 ;
  assign n47 = ( ~n12 & n13 ) | ( ~n12 & n37 ) | ( n13 & n37 ) ;
  assign n48 = n10 | n47 ;
  assign n49 = ( n16 & ~n28 ) | ( n16 & n33 ) | ( ~n28 & n33 ) ;
  assign n50 = x3 | x4 ;
  assign n51 = n12 | n50 ;
  assign n52 = ( x4 & n10 ) | ( x4 & n12 ) | ( n10 & n12 ) ;
  assign n53 = n33 | n52 ;
  assign n54 = n37 & ~n50 ;
  assign n55 = ~x0 & n9 ;
  assign n56 = x2 & n31 ;
  assign n57 = ~n11 & n56 ;
  assign n58 = n15 & n56 ;
  assign n59 = n32 & n37 ;
  assign n60 = ~x0 & x2 ;
  assign n61 = n32 & n60 ;
  assign n62 = x0 & n44 ;
  assign n63 = n23 | n62 ;
  assign n64 = ~n41 & n62 ;
  assign n65 = n63 & ~n64 ;
  assign n66 = ( ~n11 & n17 ) | ( ~n11 & n21 ) | ( n17 & n21 ) ;
  assign n67 = n15 & n17 ;
  assign y0 = n14 ;
  assign y1 = n30 ;
  assign y2 = n35 ;
  assign y3 = n36 ;
  assign y4 = n46 ;
  assign y5 = n41 ;
  assign y6 = n24 ;
  assign y7 = n48 ;
  assign y8 = n27 ;
  assign y9 = n28 ;
  assign y10 = n49 ;
  assign y11 = ~n51 ;
  assign y12 = n53 ;
  assign y13 = n54 ;
  assign y14 = n55 ;
  assign y15 = n57 ;
  assign y16 = n58 ;
  assign y17 = n59 ;
  assign y18 = n61 ;
  assign y19 = n9 ;
  assign y20 = n63 ;
  assign y21 = n64 ;
  assign y22 = n65 ;
  assign y23 = ~1'b0 ;
  assign y24 = n66 ;
  assign y25 = n67 ;
endmodule
