module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 ;
  assign n129 = ~x1 & x64 ;
  assign n130 = ~x59 & x64 ;
  assign n131 = ~x61 & x64 ;
  assign n132 = x126 | x127 ;
  assign n133 = x125 | n132 ;
  assign n134 = x124 | n133 ;
  assign n135 = x123 | n134 ;
  assign n136 = x122 | n135 ;
  assign n137 = x121 | n136 ;
  assign n138 = x120 | n137 ;
  assign n139 = x119 | n138 ;
  assign n140 = x118 | n139 ;
  assign n141 = x117 | n140 ;
  assign n142 = x116 | n141 ;
  assign n143 = x115 | n142 ;
  assign n144 = x114 | n143 ;
  assign n145 = x113 | n144 ;
  assign n146 = x112 | n145 ;
  assign n147 = x111 | n146 ;
  assign n148 = x110 | n147 ;
  assign n149 = x109 | n148 ;
  assign n150 = x108 | n149 ;
  assign n151 = x107 | n150 ;
  assign n152 = x106 | n151 ;
  assign n153 = x105 | n152 ;
  assign n154 = x104 | n153 ;
  assign n155 = x103 | n154 ;
  assign n156 = x101 | x102 ;
  assign n157 = n155 | n156 ;
  assign n158 = x100 | n157 ;
  assign n159 = x99 | n158 ;
  assign n160 = x97 | x98 ;
  assign n161 = n159 | n160 ;
  assign n162 = x96 | n161 ;
  assign n163 = x95 | n162 ;
  assign n164 = x94 | n163 ;
  assign n165 = x93 | n164 ;
  assign n166 = x92 | n165 ;
  assign n167 = x91 | n166 ;
  assign n168 = x90 | n167 ;
  assign n169 = x89 | n168 ;
  assign n170 = x88 | n169 ;
  assign n171 = x86 | x87 ;
  assign n172 = n170 | n171 ;
  assign n173 = x84 | x85 ;
  assign n174 = n172 | n173 ;
  assign n175 = x82 | x83 ;
  assign n176 = n174 | n175 ;
  assign n177 = x80 | x81 ;
  assign n178 = n176 | n177 ;
  assign n179 = x78 | x79 ;
  assign n180 = n178 | n179 ;
  assign n181 = x73 | x74 ;
  assign n182 = x75 | n181 ;
  assign n183 = x72 | n182 ;
  assign n184 = x76 | x77 ;
  assign n185 = n183 | n184 ;
  assign n186 = n180 | n185 ;
  assign n187 = x70 | x71 ;
  assign n188 = x69 | n187 ;
  assign n189 = x68 | n188 ;
  assign n190 = n186 | n189 ;
  assign n191 = x67 | n190 ;
  assign n192 = ~x62 & x64 ;
  assign n193 = x65 | x66 ;
  assign n194 = ( x66 & n192 ) | ( x66 & n193 ) | ( n192 & n193 ) ;
  assign n195 = n191 | n194 ;
  assign n196 = x63 & ~x64 ;
  assign n197 = n191 | n193 ;
  assign n198 = ( x63 & n196 ) | ( x63 & n197 ) | ( n196 & n197 ) ;
  assign n199 = ( x65 & n192 ) | ( x65 & ~n198 ) | ( n192 & ~n198 ) ;
  assign n200 = n195 | n199 ;
  assign n201 = n180 | n184 ;
  assign n202 = n182 | n201 ;
  assign n203 = x64 & ~n202 ;
  assign n204 = x62 & ~n203 ;
  assign n205 = ( x62 & n200 ) | ( x62 & n204 ) | ( n200 & n204 ) ;
  assign n206 = ( x65 & n131 ) | ( x65 & ~n205 ) | ( n131 & ~n205 ) ;
  assign n207 = x65 & ~n195 ;
  assign n208 = n198 & ~n207 ;
  assign n209 = ( x66 & n206 ) | ( x66 & ~n208 ) | ( n206 & ~n208 ) ;
  assign n210 = n191 | n209 ;
  assign n211 = ( x61 & ~x64 ) | ( x61 & n210 ) | ( ~x64 & n210 ) ;
  assign n212 = ~x61 & n210 ;
  assign n213 = ( n131 & n211 ) | ( n131 & ~n212 ) | ( n211 & ~n212 ) ;
  assign n214 = ~x60 & x64 ;
  assign n215 = ( x65 & ~n213 ) | ( x65 & n214 ) | ( ~n213 & n214 ) ;
  assign n216 = ( x65 & n131 ) | ( x65 & ~n210 ) | ( n131 & ~n210 ) ;
  assign n217 = x65 & n131 ;
  assign n218 = ( ~n205 & n216 ) | ( ~n205 & n217 ) | ( n216 & n217 ) ;
  assign n219 = ( n205 & n216 ) | ( n205 & n217 ) | ( n216 & n217 ) ;
  assign n220 = ( n205 & n218 ) | ( n205 & ~n219 ) | ( n218 & ~n219 ) ;
  assign n221 = ( x66 & n215 ) | ( x66 & ~n220 ) | ( n215 & ~n220 ) ;
  assign n222 = x66 & n206 ;
  assign n223 = ( x66 & ~n191 ) | ( x66 & n206 ) | ( ~n191 & n206 ) ;
  assign n224 = ( n208 & n222 ) | ( n208 & ~n223 ) | ( n222 & ~n223 ) ;
  assign n225 = ( x67 & n221 ) | ( x67 & ~n224 ) | ( n221 & ~n224 ) ;
  assign n226 = x72 | n189 ;
  assign n227 = n203 & ~n226 ;
  assign n228 = ( x60 & ~n225 ) | ( x60 & n227 ) | ( ~n225 & n227 ) ;
  assign n229 = x60 & ~n227 ;
  assign n230 = x60 & ~n225 ;
  assign n231 = ( n228 & n229 ) | ( n228 & ~n230 ) | ( n229 & ~n230 ) ;
  assign n232 = ( x65 & n130 ) | ( x65 & ~n231 ) | ( n130 & ~n231 ) ;
  assign n233 = n190 | n225 ;
  assign n234 = ( x65 & n214 ) | ( x65 & n233 ) | ( n214 & n233 ) ;
  assign n235 = x65 | n214 ;
  assign n236 = ( n213 & ~n234 ) | ( n213 & n235 ) | ( ~n234 & n235 ) ;
  assign n237 = ( n213 & n234 ) | ( n213 & n235 ) | ( n234 & n235 ) ;
  assign n238 = ( n234 & n236 ) | ( n234 & ~n237 ) | ( n236 & ~n237 ) ;
  assign n239 = ( x66 & n232 ) | ( x66 & ~n238 ) | ( n232 & ~n238 ) ;
  assign n240 = ( x66 & n215 ) | ( x66 & ~n233 ) | ( n215 & ~n233 ) ;
  assign n241 = x66 & n215 ;
  assign n242 = ( ~n220 & n240 ) | ( ~n220 & n241 ) | ( n240 & n241 ) ;
  assign n243 = ( n220 & n240 ) | ( n220 & n241 ) | ( n240 & n241 ) ;
  assign n244 = ( n220 & n242 ) | ( n220 & ~n243 ) | ( n242 & ~n243 ) ;
  assign n245 = ( x67 & n239 ) | ( x67 & ~n244 ) | ( n239 & ~n244 ) ;
  assign n246 = x67 & n221 ;
  assign n247 = ( x67 & ~n190 ) | ( x67 & n221 ) | ( ~n190 & n221 ) ;
  assign n248 = ( n224 & n246 ) | ( n224 & ~n247 ) | ( n246 & ~n247 ) ;
  assign n249 = ( x68 & n245 ) | ( x68 & ~n248 ) | ( n245 & ~n248 ) ;
  assign n250 = n183 | n188 ;
  assign n251 = n201 | n250 ;
  assign n252 = n249 | n251 ;
  assign n253 = ( x59 & ~x64 ) | ( x59 & n252 ) | ( ~x64 & n252 ) ;
  assign n254 = ~x59 & n252 ;
  assign n255 = ( n130 & n253 ) | ( n130 & ~n254 ) | ( n253 & ~n254 ) ;
  assign n256 = ~x58 & x64 ;
  assign n257 = ( x65 & ~n255 ) | ( x65 & n256 ) | ( ~n255 & n256 ) ;
  assign n258 = ( x65 & n130 ) | ( x65 & ~n252 ) | ( n130 & ~n252 ) ;
  assign n259 = x65 & n130 ;
  assign n260 = ( n231 & n258 ) | ( n231 & n259 ) | ( n258 & n259 ) ;
  assign n261 = ( ~n231 & n258 ) | ( ~n231 & n259 ) | ( n258 & n259 ) ;
  assign n262 = ( n231 & ~n260 ) | ( n231 & n261 ) | ( ~n260 & n261 ) ;
  assign n263 = ( x66 & n257 ) | ( x66 & ~n262 ) | ( n257 & ~n262 ) ;
  assign n264 = ( x66 & n232 ) | ( x66 & ~n252 ) | ( n232 & ~n252 ) ;
  assign n265 = x66 & n232 ;
  assign n266 = ( n238 & n264 ) | ( n238 & n265 ) | ( n264 & n265 ) ;
  assign n267 = ( ~n238 & n264 ) | ( ~n238 & n265 ) | ( n264 & n265 ) ;
  assign n268 = ( n238 & ~n266 ) | ( n238 & n267 ) | ( ~n266 & n267 ) ;
  assign n269 = ( x67 & n263 ) | ( x67 & ~n268 ) | ( n263 & ~n268 ) ;
  assign n270 = ( x67 & n239 ) | ( x67 & ~n252 ) | ( n239 & ~n252 ) ;
  assign n271 = x67 & n239 ;
  assign n272 = ( n244 & n270 ) | ( n244 & n271 ) | ( n270 & n271 ) ;
  assign n273 = ( ~n244 & n270 ) | ( ~n244 & n271 ) | ( n270 & n271 ) ;
  assign n274 = ( n244 & ~n272 ) | ( n244 & n273 ) | ( ~n272 & n273 ) ;
  assign n275 = ( x68 & n269 ) | ( x68 & ~n274 ) | ( n269 & ~n274 ) ;
  assign n276 = x68 & n245 ;
  assign n277 = ( x68 & n245 ) | ( x68 & ~n251 ) | ( n245 & ~n251 ) ;
  assign n278 = ( n248 & n276 ) | ( n248 & ~n277 ) | ( n276 & ~n277 ) ;
  assign n279 = ~n251 & n278 ;
  assign n280 = ~n275 & n279 ;
  assign n281 = ( x69 & n186 ) | ( x69 & ~n278 ) | ( n186 & ~n278 ) ;
  assign n282 = ~n279 & n281 ;
  assign n283 = ( ~x69 & n187 ) | ( ~x69 & n278 ) | ( n187 & n278 ) ;
  assign n284 = n275 | n283 ;
  assign n285 = ( ~n279 & n282 ) | ( ~n279 & n284 ) | ( n282 & n284 ) ;
  assign n286 = ( n278 & n280 ) | ( n278 & n285 ) | ( n280 & n285 ) ;
  assign n287 = ( x58 & x64 ) | ( x58 & ~n285 ) | ( x64 & ~n285 ) ;
  assign n288 = x58 & n285 ;
  assign n289 = x58 & x64 ;
  assign n290 = ( n287 & n288 ) | ( n287 & ~n289 ) | ( n288 & ~n289 ) ;
  assign n291 = ~x57 & x64 ;
  assign n292 = ( x65 & ~n290 ) | ( x65 & n291 ) | ( ~n290 & n291 ) ;
  assign n293 = ( x65 & n256 ) | ( x65 & n285 ) | ( n256 & n285 ) ;
  assign n294 = x65 | n256 ;
  assign n295 = ( ~n255 & n293 ) | ( ~n255 & n294 ) | ( n293 & n294 ) ;
  assign n296 = ( n255 & n293 ) | ( n255 & n294 ) | ( n293 & n294 ) ;
  assign n297 = ( n255 & n295 ) | ( n255 & ~n296 ) | ( n295 & ~n296 ) ;
  assign n298 = ( x66 & n292 ) | ( x66 & ~n297 ) | ( n292 & ~n297 ) ;
  assign n299 = ( x66 & n257 ) | ( x66 & ~n285 ) | ( n257 & ~n285 ) ;
  assign n300 = x66 & n257 ;
  assign n301 = ( ~n262 & n299 ) | ( ~n262 & n300 ) | ( n299 & n300 ) ;
  assign n302 = ( n262 & n299 ) | ( n262 & n300 ) | ( n299 & n300 ) ;
  assign n303 = ( n262 & n301 ) | ( n262 & ~n302 ) | ( n301 & ~n302 ) ;
  assign n304 = ( x67 & n298 ) | ( x67 & ~n303 ) | ( n298 & ~n303 ) ;
  assign n305 = ( x67 & n263 ) | ( x67 & ~n285 ) | ( n263 & ~n285 ) ;
  assign n306 = x67 & n263 ;
  assign n307 = ( n268 & n305 ) | ( n268 & n306 ) | ( n305 & n306 ) ;
  assign n308 = ( ~n268 & n305 ) | ( ~n268 & n306 ) | ( n305 & n306 ) ;
  assign n309 = ( n268 & ~n307 ) | ( n268 & n308 ) | ( ~n307 & n308 ) ;
  assign n310 = ( x68 & n304 ) | ( x68 & ~n309 ) | ( n304 & ~n309 ) ;
  assign n311 = ( x68 & n269 ) | ( x68 & ~n285 ) | ( n269 & ~n285 ) ;
  assign n312 = x68 & n269 ;
  assign n313 = ( n274 & n311 ) | ( n274 & n312 ) | ( n311 & n312 ) ;
  assign n314 = ( ~n274 & n311 ) | ( ~n274 & n312 ) | ( n311 & n312 ) ;
  assign n315 = ( n274 & ~n313 ) | ( n274 & n314 ) | ( ~n313 & n314 ) ;
  assign n316 = ( x69 & n310 ) | ( x69 & ~n315 ) | ( n310 & ~n315 ) ;
  assign n317 = x70 | n316 ;
  assign n318 = x71 | n186 ;
  assign n319 = ( x70 & n316 ) | ( x70 & n318 ) | ( n316 & n318 ) ;
  assign n320 = ( n286 & ~n317 ) | ( n286 & n319 ) | ( ~n317 & n319 ) ;
  assign n321 = ( x70 & ~n286 ) | ( x70 & n316 ) | ( ~n286 & n316 ) ;
  assign n322 = x64 & ~x71 ;
  assign n323 = ~n186 & n322 ;
  assign n324 = ( x57 & ~n321 ) | ( x57 & n323 ) | ( ~n321 & n323 ) ;
  assign n325 = x57 & ~n323 ;
  assign n326 = x57 & ~n321 ;
  assign n327 = ( n324 & n325 ) | ( n324 & ~n326 ) | ( n325 & ~n326 ) ;
  assign n328 = ~x56 & x64 ;
  assign n329 = ( x65 & ~n327 ) | ( x65 & n328 ) | ( ~n327 & n328 ) ;
  assign n330 = n318 | n321 ;
  assign n331 = ( x65 & n291 ) | ( x65 & n330 ) | ( n291 & n330 ) ;
  assign n332 = x65 | n291 ;
  assign n333 = ( n290 & ~n331 ) | ( n290 & n332 ) | ( ~n331 & n332 ) ;
  assign n334 = ( n290 & n331 ) | ( n290 & n332 ) | ( n331 & n332 ) ;
  assign n335 = ( n331 & n333 ) | ( n331 & ~n334 ) | ( n333 & ~n334 ) ;
  assign n336 = ( x66 & n329 ) | ( x66 & ~n335 ) | ( n329 & ~n335 ) ;
  assign n337 = ( x66 & n292 ) | ( x66 & n330 ) | ( n292 & n330 ) ;
  assign n338 = x66 | n292 ;
  assign n339 = ( ~n297 & n337 ) | ( ~n297 & n338 ) | ( n337 & n338 ) ;
  assign n340 = ( n297 & n337 ) | ( n297 & n338 ) | ( n337 & n338 ) ;
  assign n341 = ( n297 & n339 ) | ( n297 & ~n340 ) | ( n339 & ~n340 ) ;
  assign n342 = ( x67 & n336 ) | ( x67 & ~n341 ) | ( n336 & ~n341 ) ;
  assign n343 = ( x67 & n298 ) | ( x67 & ~n330 ) | ( n298 & ~n330 ) ;
  assign n344 = x67 & n298 ;
  assign n345 = ( ~n303 & n343 ) | ( ~n303 & n344 ) | ( n343 & n344 ) ;
  assign n346 = ( n303 & n343 ) | ( n303 & n344 ) | ( n343 & n344 ) ;
  assign n347 = ( n303 & n345 ) | ( n303 & ~n346 ) | ( n345 & ~n346 ) ;
  assign n348 = ( x68 & n342 ) | ( x68 & ~n347 ) | ( n342 & ~n347 ) ;
  assign n349 = ( x68 & n304 ) | ( x68 & ~n330 ) | ( n304 & ~n330 ) ;
  assign n350 = x68 & n304 ;
  assign n351 = ( n309 & n349 ) | ( n309 & n350 ) | ( n349 & n350 ) ;
  assign n352 = ( ~n309 & n349 ) | ( ~n309 & n350 ) | ( n349 & n350 ) ;
  assign n353 = ( n309 & ~n351 ) | ( n309 & n352 ) | ( ~n351 & n352 ) ;
  assign n354 = ( x69 & n348 ) | ( x69 & ~n353 ) | ( n348 & ~n353 ) ;
  assign n355 = ( x69 & n310 ) | ( x69 & ~n330 ) | ( n310 & ~n330 ) ;
  assign n356 = x69 & n310 ;
  assign n357 = ( n315 & n355 ) | ( n315 & n356 ) | ( n355 & n356 ) ;
  assign n358 = ( ~n315 & n355 ) | ( ~n315 & n356 ) | ( n355 & n356 ) ;
  assign n359 = ( n315 & ~n357 ) | ( n315 & n358 ) | ( ~n357 & n358 ) ;
  assign n360 = ( x70 & n354 ) | ( x70 & ~n359 ) | ( n354 & ~n359 ) ;
  assign n361 = ( x71 & ~n320 ) | ( x71 & n360 ) | ( ~n320 & n360 ) ;
  assign n362 = ~x72 & n203 ;
  assign n363 = ( x56 & ~n361 ) | ( x56 & n362 ) | ( ~n361 & n362 ) ;
  assign n364 = x56 & ~n362 ;
  assign n365 = x56 & ~n361 ;
  assign n366 = ( n363 & n364 ) | ( n363 & ~n365 ) | ( n364 & ~n365 ) ;
  assign n367 = ~x55 & x64 ;
  assign n368 = ( x65 & ~n366 ) | ( x65 & n367 ) | ( ~n366 & n367 ) ;
  assign n369 = n186 | n361 ;
  assign n370 = ( x65 & n328 ) | ( x65 & n369 ) | ( n328 & n369 ) ;
  assign n371 = x65 | n328 ;
  assign n372 = ( n327 & ~n370 ) | ( n327 & n371 ) | ( ~n370 & n371 ) ;
  assign n373 = ( n327 & n370 ) | ( n327 & n371 ) | ( n370 & n371 ) ;
  assign n374 = ( n370 & n372 ) | ( n370 & ~n373 ) | ( n372 & ~n373 ) ;
  assign n375 = ( x66 & n368 ) | ( x66 & ~n374 ) | ( n368 & ~n374 ) ;
  assign n376 = ( x66 & n329 ) | ( x66 & n369 ) | ( n329 & n369 ) ;
  assign n377 = x66 | n329 ;
  assign n378 = ( ~n335 & n376 ) | ( ~n335 & n377 ) | ( n376 & n377 ) ;
  assign n379 = ( n335 & n376 ) | ( n335 & n377 ) | ( n376 & n377 ) ;
  assign n380 = ( n335 & n378 ) | ( n335 & ~n379 ) | ( n378 & ~n379 ) ;
  assign n381 = ( x67 & n375 ) | ( x67 & ~n380 ) | ( n375 & ~n380 ) ;
  assign n382 = ( x67 & n336 ) | ( x67 & ~n369 ) | ( n336 & ~n369 ) ;
  assign n383 = x67 & n336 ;
  assign n384 = ( ~n341 & n382 ) | ( ~n341 & n383 ) | ( n382 & n383 ) ;
  assign n385 = ( n341 & n382 ) | ( n341 & n383 ) | ( n382 & n383 ) ;
  assign n386 = ( n341 & n384 ) | ( n341 & ~n385 ) | ( n384 & ~n385 ) ;
  assign n387 = ( x68 & n381 ) | ( x68 & ~n386 ) | ( n381 & ~n386 ) ;
  assign n388 = ( x68 & n342 ) | ( x68 & ~n369 ) | ( n342 & ~n369 ) ;
  assign n389 = x68 & n342 ;
  assign n390 = ( n347 & n388 ) | ( n347 & n389 ) | ( n388 & n389 ) ;
  assign n391 = ( ~n347 & n388 ) | ( ~n347 & n389 ) | ( n388 & n389 ) ;
  assign n392 = ( n347 & ~n390 ) | ( n347 & n391 ) | ( ~n390 & n391 ) ;
  assign n393 = ( x69 & n387 ) | ( x69 & ~n392 ) | ( n387 & ~n392 ) ;
  assign n394 = ( x69 & n348 ) | ( x69 & ~n369 ) | ( n348 & ~n369 ) ;
  assign n395 = x69 & n348 ;
  assign n396 = ( ~n353 & n394 ) | ( ~n353 & n395 ) | ( n394 & n395 ) ;
  assign n397 = ( n353 & n394 ) | ( n353 & n395 ) | ( n394 & n395 ) ;
  assign n398 = ( n353 & n396 ) | ( n353 & ~n397 ) | ( n396 & ~n397 ) ;
  assign n399 = ( x70 & n393 ) | ( x70 & ~n398 ) | ( n393 & ~n398 ) ;
  assign n400 = ( x70 & n354 ) | ( x70 & ~n369 ) | ( n354 & ~n369 ) ;
  assign n401 = x70 & n354 ;
  assign n402 = ( ~n359 & n400 ) | ( ~n359 & n401 ) | ( n400 & n401 ) ;
  assign n403 = ( n359 & n400 ) | ( n359 & n401 ) | ( n400 & n401 ) ;
  assign n404 = ( n359 & n402 ) | ( n359 & ~n403 ) | ( n402 & ~n403 ) ;
  assign n405 = ( x71 & n399 ) | ( x71 & ~n404 ) | ( n399 & ~n404 ) ;
  assign n406 = ( n186 & n202 ) | ( n186 & ~n286 ) | ( n202 & ~n286 ) ;
  assign n407 = n405 | n406 ;
  assign n408 = n320 & n369 ;
  assign n409 = ~n186 & n408 ;
  assign n410 = ( n280 & n408 ) | ( n280 & ~n409 ) | ( n408 & ~n409 ) ;
  assign n411 = ( n280 & n407 ) | ( n280 & n410 ) | ( n407 & n410 ) ;
  assign n412 = n407 & ~n409 ;
  assign n413 = ( x55 & x64 ) | ( x55 & ~n412 ) | ( x64 & ~n412 ) ;
  assign n414 = x55 & n412 ;
  assign n415 = x55 & x64 ;
  assign n416 = ( n413 & n414 ) | ( n413 & ~n415 ) | ( n414 & ~n415 ) ;
  assign n417 = ~x54 & x64 ;
  assign n418 = ( x65 & ~n416 ) | ( x65 & n417 ) | ( ~n416 & n417 ) ;
  assign n419 = ( x65 & n367 ) | ( x65 & n412 ) | ( n367 & n412 ) ;
  assign n420 = x65 | n367 ;
  assign n421 = ( ~n366 & n419 ) | ( ~n366 & n420 ) | ( n419 & n420 ) ;
  assign n422 = ( n366 & n419 ) | ( n366 & n420 ) | ( n419 & n420 ) ;
  assign n423 = ( n366 & n421 ) | ( n366 & ~n422 ) | ( n421 & ~n422 ) ;
  assign n424 = ( x66 & n418 ) | ( x66 & ~n423 ) | ( n418 & ~n423 ) ;
  assign n425 = ( x66 & n368 ) | ( x66 & n412 ) | ( n368 & n412 ) ;
  assign n426 = x66 | n368 ;
  assign n427 = ( n374 & n425 ) | ( n374 & n426 ) | ( n425 & n426 ) ;
  assign n428 = ( ~n374 & n425 ) | ( ~n374 & n426 ) | ( n425 & n426 ) ;
  assign n429 = ( n374 & ~n427 ) | ( n374 & n428 ) | ( ~n427 & n428 ) ;
  assign n430 = ( x67 & n424 ) | ( x67 & ~n429 ) | ( n424 & ~n429 ) ;
  assign n431 = ( x67 & n375 ) | ( x67 & ~n412 ) | ( n375 & ~n412 ) ;
  assign n432 = x67 & n375 ;
  assign n433 = ( n380 & n431 ) | ( n380 & n432 ) | ( n431 & n432 ) ;
  assign n434 = ( ~n380 & n431 ) | ( ~n380 & n432 ) | ( n431 & n432 ) ;
  assign n435 = ( n380 & ~n433 ) | ( n380 & n434 ) | ( ~n433 & n434 ) ;
  assign n436 = ( x68 & n430 ) | ( x68 & ~n435 ) | ( n430 & ~n435 ) ;
  assign n437 = ( x68 & n381 ) | ( x68 & ~n412 ) | ( n381 & ~n412 ) ;
  assign n438 = x68 & n381 ;
  assign n439 = ( ~n386 & n437 ) | ( ~n386 & n438 ) | ( n437 & n438 ) ;
  assign n440 = ( n386 & n437 ) | ( n386 & n438 ) | ( n437 & n438 ) ;
  assign n441 = ( n386 & n439 ) | ( n386 & ~n440 ) | ( n439 & ~n440 ) ;
  assign n442 = ( x69 & n436 ) | ( x69 & ~n441 ) | ( n436 & ~n441 ) ;
  assign n443 = ( x69 & n387 ) | ( x69 & ~n412 ) | ( n387 & ~n412 ) ;
  assign n444 = x69 & n387 ;
  assign n445 = ( n392 & n443 ) | ( n392 & n444 ) | ( n443 & n444 ) ;
  assign n446 = ( ~n392 & n443 ) | ( ~n392 & n444 ) | ( n443 & n444 ) ;
  assign n447 = ( n392 & ~n445 ) | ( n392 & n446 ) | ( ~n445 & n446 ) ;
  assign n448 = ( x70 & n442 ) | ( x70 & ~n447 ) | ( n442 & ~n447 ) ;
  assign n449 = ( x70 & n393 ) | ( x70 & ~n412 ) | ( n393 & ~n412 ) ;
  assign n450 = x70 & n393 ;
  assign n451 = ( ~n398 & n449 ) | ( ~n398 & n450 ) | ( n449 & n450 ) ;
  assign n452 = ( n398 & n449 ) | ( n398 & n450 ) | ( n449 & n450 ) ;
  assign n453 = ( n398 & n451 ) | ( n398 & ~n452 ) | ( n451 & ~n452 ) ;
  assign n454 = ( x71 & n448 ) | ( x71 & ~n453 ) | ( n448 & ~n453 ) ;
  assign n455 = ( x71 & n399 ) | ( x71 & n404 ) | ( n399 & n404 ) ;
  assign n456 = n412 | n455 ;
  assign n457 = ( n404 & n407 ) | ( n404 & ~n456 ) | ( n407 & ~n456 ) ;
  assign n458 = ( x72 & n454 ) | ( x72 & ~n457 ) | ( n454 & ~n457 ) ;
  assign n459 = x73 | n458 ;
  assign n460 = x74 | x75 ;
  assign n461 = n201 | n460 ;
  assign n462 = ( x73 & n458 ) | ( x73 & n461 ) | ( n458 & n461 ) ;
  assign n463 = ( n411 & ~n459 ) | ( n411 & n462 ) | ( ~n459 & n462 ) ;
  assign n464 = ( x73 & ~n411 ) | ( x73 & n458 ) | ( ~n411 & n458 ) ;
  assign n465 = n461 | n464 ;
  assign n466 = ( x54 & ~x64 ) | ( x54 & n465 ) | ( ~x64 & n465 ) ;
  assign n467 = ~x54 & n465 ;
  assign n468 = ( n417 & n466 ) | ( n417 & ~n467 ) | ( n466 & ~n467 ) ;
  assign n469 = ~x53 & x64 ;
  assign n470 = ( x65 & ~n468 ) | ( x65 & n469 ) | ( ~n468 & n469 ) ;
  assign n471 = ( x65 & n417 ) | ( x65 & ~n465 ) | ( n417 & ~n465 ) ;
  assign n472 = x65 & n417 ;
  assign n473 = ( n416 & n471 ) | ( n416 & n472 ) | ( n471 & n472 ) ;
  assign n474 = ( ~n416 & n471 ) | ( ~n416 & n472 ) | ( n471 & n472 ) ;
  assign n475 = ( n416 & ~n473 ) | ( n416 & n474 ) | ( ~n473 & n474 ) ;
  assign n476 = ( x66 & n470 ) | ( x66 & ~n475 ) | ( n470 & ~n475 ) ;
  assign n477 = ( x66 & n418 ) | ( x66 & n465 ) | ( n418 & n465 ) ;
  assign n478 = x66 | n418 ;
  assign n479 = ( ~n423 & n477 ) | ( ~n423 & n478 ) | ( n477 & n478 ) ;
  assign n480 = ( n423 & n477 ) | ( n423 & n478 ) | ( n477 & n478 ) ;
  assign n481 = ( n423 & n479 ) | ( n423 & ~n480 ) | ( n479 & ~n480 ) ;
  assign n482 = ( x67 & n476 ) | ( x67 & ~n481 ) | ( n476 & ~n481 ) ;
  assign n483 = ( x67 & n424 ) | ( x67 & ~n465 ) | ( n424 & ~n465 ) ;
  assign n484 = x67 & n424 ;
  assign n485 = ( ~n429 & n483 ) | ( ~n429 & n484 ) | ( n483 & n484 ) ;
  assign n486 = ( n429 & n483 ) | ( n429 & n484 ) | ( n483 & n484 ) ;
  assign n487 = ( n429 & n485 ) | ( n429 & ~n486 ) | ( n485 & ~n486 ) ;
  assign n488 = ( x68 & n482 ) | ( x68 & ~n487 ) | ( n482 & ~n487 ) ;
  assign n489 = ( x68 & n430 ) | ( x68 & ~n465 ) | ( n430 & ~n465 ) ;
  assign n490 = x68 & n430 ;
  assign n491 = ( n435 & n489 ) | ( n435 & n490 ) | ( n489 & n490 ) ;
  assign n492 = ( ~n435 & n489 ) | ( ~n435 & n490 ) | ( n489 & n490 ) ;
  assign n493 = ( n435 & ~n491 ) | ( n435 & n492 ) | ( ~n491 & n492 ) ;
  assign n494 = ( x69 & n488 ) | ( x69 & ~n493 ) | ( n488 & ~n493 ) ;
  assign n495 = ( x69 & n436 ) | ( x69 & ~n465 ) | ( n436 & ~n465 ) ;
  assign n496 = x69 & n436 ;
  assign n497 = ( ~n441 & n495 ) | ( ~n441 & n496 ) | ( n495 & n496 ) ;
  assign n498 = ( n441 & n495 ) | ( n441 & n496 ) | ( n495 & n496 ) ;
  assign n499 = ( n441 & n497 ) | ( n441 & ~n498 ) | ( n497 & ~n498 ) ;
  assign n500 = ( x70 & n494 ) | ( x70 & ~n499 ) | ( n494 & ~n499 ) ;
  assign n501 = ( x70 & n442 ) | ( x70 & ~n465 ) | ( n442 & ~n465 ) ;
  assign n502 = x70 & n442 ;
  assign n503 = ( n447 & n501 ) | ( n447 & n502 ) | ( n501 & n502 ) ;
  assign n504 = ( ~n447 & n501 ) | ( ~n447 & n502 ) | ( n501 & n502 ) ;
  assign n505 = ( n447 & ~n503 ) | ( n447 & n504 ) | ( ~n503 & n504 ) ;
  assign n506 = ( x71 & n500 ) | ( x71 & ~n505 ) | ( n500 & ~n505 ) ;
  assign n507 = ( x71 & n448 ) | ( x71 & ~n465 ) | ( n448 & ~n465 ) ;
  assign n508 = x71 & n448 ;
  assign n509 = ( ~n453 & n507 ) | ( ~n453 & n508 ) | ( n507 & n508 ) ;
  assign n510 = ( n453 & n507 ) | ( n453 & n508 ) | ( n507 & n508 ) ;
  assign n511 = ( n453 & n509 ) | ( n453 & ~n510 ) | ( n509 & ~n510 ) ;
  assign n512 = ( x72 & n506 ) | ( x72 & ~n511 ) | ( n506 & ~n511 ) ;
  assign n513 = ( x72 & n454 ) | ( x72 & ~n465 ) | ( n454 & ~n465 ) ;
  assign n514 = x72 & n454 ;
  assign n515 = ( ~n457 & n513 ) | ( ~n457 & n514 ) | ( n513 & n514 ) ;
  assign n516 = ( n457 & n513 ) | ( n457 & n514 ) | ( n513 & n514 ) ;
  assign n517 = ( n457 & n515 ) | ( n457 & ~n516 ) | ( n515 & ~n516 ) ;
  assign n518 = ( x73 & n512 ) | ( x73 & ~n517 ) | ( n512 & ~n517 ) ;
  assign n519 = x74 | n518 ;
  assign n520 = x75 | n201 ;
  assign n521 = ( x74 & n518 ) | ( x74 & n520 ) | ( n518 & n520 ) ;
  assign n522 = ( n463 & ~n519 ) | ( n463 & n521 ) | ( ~n519 & n521 ) ;
  assign n523 = ( x74 & ~n463 ) | ( x74 & n518 ) | ( ~n463 & n518 ) ;
  assign n524 = n520 | n523 ;
  assign n525 = ( x53 & ~x64 ) | ( x53 & n524 ) | ( ~x64 & n524 ) ;
  assign n526 = ~x53 & n524 ;
  assign n527 = ( n469 & n525 ) | ( n469 & ~n526 ) | ( n525 & ~n526 ) ;
  assign n528 = ~x52 & x64 ;
  assign n529 = ( x65 & ~n527 ) | ( x65 & n528 ) | ( ~n527 & n528 ) ;
  assign n530 = ( x65 & n469 ) | ( x65 & ~n524 ) | ( n469 & ~n524 ) ;
  assign n531 = x65 & n469 ;
  assign n532 = ( n468 & n530 ) | ( n468 & n531 ) | ( n530 & n531 ) ;
  assign n533 = ( ~n468 & n530 ) | ( ~n468 & n531 ) | ( n530 & n531 ) ;
  assign n534 = ( n468 & ~n532 ) | ( n468 & n533 ) | ( ~n532 & n533 ) ;
  assign n535 = ( x66 & n529 ) | ( x66 & ~n534 ) | ( n529 & ~n534 ) ;
  assign n536 = ( x66 & n470 ) | ( x66 & n524 ) | ( n470 & n524 ) ;
  assign n537 = x66 | n470 ;
  assign n538 = ( ~n475 & n536 ) | ( ~n475 & n537 ) | ( n536 & n537 ) ;
  assign n539 = ( n475 & n536 ) | ( n475 & n537 ) | ( n536 & n537 ) ;
  assign n540 = ( n475 & n538 ) | ( n475 & ~n539 ) | ( n538 & ~n539 ) ;
  assign n541 = ( x67 & n535 ) | ( x67 & ~n540 ) | ( n535 & ~n540 ) ;
  assign n542 = ( x67 & n476 ) | ( x67 & ~n524 ) | ( n476 & ~n524 ) ;
  assign n543 = x67 & n476 ;
  assign n544 = ( ~n481 & n542 ) | ( ~n481 & n543 ) | ( n542 & n543 ) ;
  assign n545 = ( n481 & n542 ) | ( n481 & n543 ) | ( n542 & n543 ) ;
  assign n546 = ( n481 & n544 ) | ( n481 & ~n545 ) | ( n544 & ~n545 ) ;
  assign n547 = ( x68 & n541 ) | ( x68 & ~n546 ) | ( n541 & ~n546 ) ;
  assign n548 = ( x68 & n482 ) | ( x68 & ~n524 ) | ( n482 & ~n524 ) ;
  assign n549 = x68 & n482 ;
  assign n550 = ( n487 & n548 ) | ( n487 & n549 ) | ( n548 & n549 ) ;
  assign n551 = ( ~n487 & n548 ) | ( ~n487 & n549 ) | ( n548 & n549 ) ;
  assign n552 = ( n487 & ~n550 ) | ( n487 & n551 ) | ( ~n550 & n551 ) ;
  assign n553 = ( x69 & n547 ) | ( x69 & ~n552 ) | ( n547 & ~n552 ) ;
  assign n554 = ( x69 & n488 ) | ( x69 & ~n524 ) | ( n488 & ~n524 ) ;
  assign n555 = x69 & n488 ;
  assign n556 = ( ~n493 & n554 ) | ( ~n493 & n555 ) | ( n554 & n555 ) ;
  assign n557 = ( n493 & n554 ) | ( n493 & n555 ) | ( n554 & n555 ) ;
  assign n558 = ( n493 & n556 ) | ( n493 & ~n557 ) | ( n556 & ~n557 ) ;
  assign n559 = ( x70 & n553 ) | ( x70 & ~n558 ) | ( n553 & ~n558 ) ;
  assign n560 = ( x70 & n494 ) | ( x70 & ~n524 ) | ( n494 & ~n524 ) ;
  assign n561 = x70 & n494 ;
  assign n562 = ( n499 & n560 ) | ( n499 & n561 ) | ( n560 & n561 ) ;
  assign n563 = ( ~n499 & n560 ) | ( ~n499 & n561 ) | ( n560 & n561 ) ;
  assign n564 = ( n499 & ~n562 ) | ( n499 & n563 ) | ( ~n562 & n563 ) ;
  assign n565 = ( x71 & n559 ) | ( x71 & ~n564 ) | ( n559 & ~n564 ) ;
  assign n566 = ( x71 & n500 ) | ( x71 & ~n524 ) | ( n500 & ~n524 ) ;
  assign n567 = x71 & n500 ;
  assign n568 = ( ~n505 & n566 ) | ( ~n505 & n567 ) | ( n566 & n567 ) ;
  assign n569 = ( n505 & n566 ) | ( n505 & n567 ) | ( n566 & n567 ) ;
  assign n570 = ( n505 & n568 ) | ( n505 & ~n569 ) | ( n568 & ~n569 ) ;
  assign n571 = ( x72 & n565 ) | ( x72 & ~n570 ) | ( n565 & ~n570 ) ;
  assign n572 = ( x72 & n506 ) | ( x72 & ~n524 ) | ( n506 & ~n524 ) ;
  assign n573 = x72 & n506 ;
  assign n574 = ( n511 & n572 ) | ( n511 & n573 ) | ( n572 & n573 ) ;
  assign n575 = ( ~n511 & n572 ) | ( ~n511 & n573 ) | ( n572 & n573 ) ;
  assign n576 = ( n511 & ~n574 ) | ( n511 & n575 ) | ( ~n574 & n575 ) ;
  assign n577 = ( x73 & n571 ) | ( x73 & ~n576 ) | ( n571 & ~n576 ) ;
  assign n578 = ( x73 & n512 ) | ( x73 & ~n524 ) | ( n512 & ~n524 ) ;
  assign n579 = x73 & n512 ;
  assign n580 = ( n517 & n578 ) | ( n517 & n579 ) | ( n578 & n579 ) ;
  assign n581 = ( ~n517 & n578 ) | ( ~n517 & n579 ) | ( n578 & n579 ) ;
  assign n582 = ( n517 & ~n580 ) | ( n517 & n581 ) | ( ~n580 & n581 ) ;
  assign n583 = ( x74 & n577 ) | ( x74 & ~n582 ) | ( n577 & ~n582 ) ;
  assign n584 = ( x75 & ~n522 ) | ( x75 & n583 ) | ( ~n522 & n583 ) ;
  assign n585 = n201 | n584 ;
  assign n586 = n522 & n585 ;
  assign n587 = n280 | n586 ;
  assign n588 = ( x52 & ~x64 ) | ( x52 & n585 ) | ( ~x64 & n585 ) ;
  assign n589 = ~x52 & n585 ;
  assign n590 = ( n528 & n588 ) | ( n528 & ~n589 ) | ( n588 & ~n589 ) ;
  assign n591 = ~x51 & x64 ;
  assign n592 = ( x65 & ~n590 ) | ( x65 & n591 ) | ( ~n590 & n591 ) ;
  assign n593 = ( x65 & n528 ) | ( x65 & ~n585 ) | ( n528 & ~n585 ) ;
  assign n594 = x65 & n528 ;
  assign n595 = ( n527 & n593 ) | ( n527 & n594 ) | ( n593 & n594 ) ;
  assign n596 = ( ~n527 & n593 ) | ( ~n527 & n594 ) | ( n593 & n594 ) ;
  assign n597 = ( n527 & ~n595 ) | ( n527 & n596 ) | ( ~n595 & n596 ) ;
  assign n598 = ( x66 & n592 ) | ( x66 & ~n597 ) | ( n592 & ~n597 ) ;
  assign n599 = ( x66 & n529 ) | ( x66 & ~n585 ) | ( n529 & ~n585 ) ;
  assign n600 = x66 & n529 ;
  assign n601 = ( n534 & n599 ) | ( n534 & n600 ) | ( n599 & n600 ) ;
  assign n602 = ( ~n534 & n599 ) | ( ~n534 & n600 ) | ( n599 & n600 ) ;
  assign n603 = ( n534 & ~n601 ) | ( n534 & n602 ) | ( ~n601 & n602 ) ;
  assign n604 = ( x67 & n598 ) | ( x67 & ~n603 ) | ( n598 & ~n603 ) ;
  assign n605 = ( x67 & n535 ) | ( x67 & ~n585 ) | ( n535 & ~n585 ) ;
  assign n606 = x67 & n535 ;
  assign n607 = ( ~n540 & n605 ) | ( ~n540 & n606 ) | ( n605 & n606 ) ;
  assign n608 = ( n540 & n605 ) | ( n540 & n606 ) | ( n605 & n606 ) ;
  assign n609 = ( n540 & n607 ) | ( n540 & ~n608 ) | ( n607 & ~n608 ) ;
  assign n610 = ( x68 & n604 ) | ( x68 & ~n609 ) | ( n604 & ~n609 ) ;
  assign n611 = ( x68 & n541 ) | ( x68 & ~n585 ) | ( n541 & ~n585 ) ;
  assign n612 = x68 & n541 ;
  assign n613 = ( n546 & n611 ) | ( n546 & n612 ) | ( n611 & n612 ) ;
  assign n614 = ( ~n546 & n611 ) | ( ~n546 & n612 ) | ( n611 & n612 ) ;
  assign n615 = ( n546 & ~n613 ) | ( n546 & n614 ) | ( ~n613 & n614 ) ;
  assign n616 = ( x69 & n610 ) | ( x69 & ~n615 ) | ( n610 & ~n615 ) ;
  assign n617 = ( x69 & n547 ) | ( x69 & ~n585 ) | ( n547 & ~n585 ) ;
  assign n618 = x69 & n547 ;
  assign n619 = ( ~n552 & n617 ) | ( ~n552 & n618 ) | ( n617 & n618 ) ;
  assign n620 = ( n552 & n617 ) | ( n552 & n618 ) | ( n617 & n618 ) ;
  assign n621 = ( n552 & n619 ) | ( n552 & ~n620 ) | ( n619 & ~n620 ) ;
  assign n622 = ( x70 & n616 ) | ( x70 & ~n621 ) | ( n616 & ~n621 ) ;
  assign n623 = ( x70 & n553 ) | ( x70 & ~n585 ) | ( n553 & ~n585 ) ;
  assign n624 = x70 & n553 ;
  assign n625 = ( n558 & n623 ) | ( n558 & n624 ) | ( n623 & n624 ) ;
  assign n626 = ( ~n558 & n623 ) | ( ~n558 & n624 ) | ( n623 & n624 ) ;
  assign n627 = ( n558 & ~n625 ) | ( n558 & n626 ) | ( ~n625 & n626 ) ;
  assign n628 = ( x71 & n622 ) | ( x71 & ~n627 ) | ( n622 & ~n627 ) ;
  assign n629 = ( x71 & n559 ) | ( x71 & ~n585 ) | ( n559 & ~n585 ) ;
  assign n630 = x71 & n559 ;
  assign n631 = ( ~n564 & n629 ) | ( ~n564 & n630 ) | ( n629 & n630 ) ;
  assign n632 = ( n564 & n629 ) | ( n564 & n630 ) | ( n629 & n630 ) ;
  assign n633 = ( n564 & n631 ) | ( n564 & ~n632 ) | ( n631 & ~n632 ) ;
  assign n634 = ( x72 & n628 ) | ( x72 & ~n633 ) | ( n628 & ~n633 ) ;
  assign n635 = ( x72 & n565 ) | ( x72 & ~n585 ) | ( n565 & ~n585 ) ;
  assign n636 = x72 & n565 ;
  assign n637 = ( n570 & n635 ) | ( n570 & n636 ) | ( n635 & n636 ) ;
  assign n638 = ( ~n570 & n635 ) | ( ~n570 & n636 ) | ( n635 & n636 ) ;
  assign n639 = ( n570 & ~n637 ) | ( n570 & n638 ) | ( ~n637 & n638 ) ;
  assign n640 = ( x73 & n634 ) | ( x73 & ~n639 ) | ( n634 & ~n639 ) ;
  assign n641 = ( x73 & n571 ) | ( x73 & ~n585 ) | ( n571 & ~n585 ) ;
  assign n642 = x73 & n571 ;
  assign n643 = ( ~n576 & n641 ) | ( ~n576 & n642 ) | ( n641 & n642 ) ;
  assign n644 = ( n576 & n641 ) | ( n576 & n642 ) | ( n641 & n642 ) ;
  assign n645 = ( n576 & n643 ) | ( n576 & ~n644 ) | ( n643 & ~n644 ) ;
  assign n646 = ( x74 & n640 ) | ( x74 & ~n645 ) | ( n640 & ~n645 ) ;
  assign n647 = ( x74 & n577 ) | ( x74 & ~n585 ) | ( n577 & ~n585 ) ;
  assign n648 = x74 & n577 ;
  assign n649 = ( ~n582 & n647 ) | ( ~n582 & n648 ) | ( n647 & n648 ) ;
  assign n650 = ( n582 & n647 ) | ( n582 & n648 ) | ( n647 & n648 ) ;
  assign n651 = ( n582 & n649 ) | ( n582 & ~n650 ) | ( n649 & ~n650 ) ;
  assign n652 = ( x75 & n646 ) | ( x75 & ~n651 ) | ( n646 & ~n651 ) ;
  assign n653 = x76 | n652 ;
  assign n654 = x77 | n180 ;
  assign n655 = ( x76 & n652 ) | ( x76 & n654 ) | ( n652 & n654 ) ;
  assign n656 = ( n587 & ~n653 ) | ( n587 & n655 ) | ( ~n653 & n655 ) ;
  assign n657 = ( x76 & ~n587 ) | ( x76 & n652 ) | ( ~n587 & n652 ) ;
  assign n658 = n654 | n657 ;
  assign n659 = ( x51 & ~x64 ) | ( x51 & n658 ) | ( ~x64 & n658 ) ;
  assign n660 = ~x51 & n658 ;
  assign n661 = ( n591 & n659 ) | ( n591 & ~n660 ) | ( n659 & ~n660 ) ;
  assign n662 = ~x50 & x64 ;
  assign n663 = ( x65 & ~n661 ) | ( x65 & n662 ) | ( ~n661 & n662 ) ;
  assign n664 = ( x65 & n591 ) | ( x65 & ~n658 ) | ( n591 & ~n658 ) ;
  assign n665 = x65 & n591 ;
  assign n666 = ( n590 & n664 ) | ( n590 & n665 ) | ( n664 & n665 ) ;
  assign n667 = ( ~n590 & n664 ) | ( ~n590 & n665 ) | ( n664 & n665 ) ;
  assign n668 = ( n590 & ~n666 ) | ( n590 & n667 ) | ( ~n666 & n667 ) ;
  assign n669 = ( x66 & n663 ) | ( x66 & ~n668 ) | ( n663 & ~n668 ) ;
  assign n670 = ( x66 & n592 ) | ( x66 & ~n658 ) | ( n592 & ~n658 ) ;
  assign n671 = x66 & n592 ;
  assign n672 = ( n597 & n670 ) | ( n597 & n671 ) | ( n670 & n671 ) ;
  assign n673 = ( ~n597 & n670 ) | ( ~n597 & n671 ) | ( n670 & n671 ) ;
  assign n674 = ( n597 & ~n672 ) | ( n597 & n673 ) | ( ~n672 & n673 ) ;
  assign n675 = ( x67 & n669 ) | ( x67 & ~n674 ) | ( n669 & ~n674 ) ;
  assign n676 = ( x67 & n598 ) | ( x67 & ~n658 ) | ( n598 & ~n658 ) ;
  assign n677 = x67 & n598 ;
  assign n678 = ( ~n603 & n676 ) | ( ~n603 & n677 ) | ( n676 & n677 ) ;
  assign n679 = ( n603 & n676 ) | ( n603 & n677 ) | ( n676 & n677 ) ;
  assign n680 = ( n603 & n678 ) | ( n603 & ~n679 ) | ( n678 & ~n679 ) ;
  assign n681 = ( x68 & n675 ) | ( x68 & ~n680 ) | ( n675 & ~n680 ) ;
  assign n682 = ( x68 & n604 ) | ( x68 & ~n658 ) | ( n604 & ~n658 ) ;
  assign n683 = x68 & n604 ;
  assign n684 = ( n609 & n682 ) | ( n609 & n683 ) | ( n682 & n683 ) ;
  assign n685 = ( ~n609 & n682 ) | ( ~n609 & n683 ) | ( n682 & n683 ) ;
  assign n686 = ( n609 & ~n684 ) | ( n609 & n685 ) | ( ~n684 & n685 ) ;
  assign n687 = ( x69 & n681 ) | ( x69 & ~n686 ) | ( n681 & ~n686 ) ;
  assign n688 = ( x69 & n610 ) | ( x69 & ~n658 ) | ( n610 & ~n658 ) ;
  assign n689 = x69 & n610 ;
  assign n690 = ( ~n615 & n688 ) | ( ~n615 & n689 ) | ( n688 & n689 ) ;
  assign n691 = ( n615 & n688 ) | ( n615 & n689 ) | ( n688 & n689 ) ;
  assign n692 = ( n615 & n690 ) | ( n615 & ~n691 ) | ( n690 & ~n691 ) ;
  assign n693 = ( x70 & n687 ) | ( x70 & ~n692 ) | ( n687 & ~n692 ) ;
  assign n694 = ( x70 & n616 ) | ( x70 & ~n658 ) | ( n616 & ~n658 ) ;
  assign n695 = x70 & n616 ;
  assign n696 = ( n621 & n694 ) | ( n621 & n695 ) | ( n694 & n695 ) ;
  assign n697 = ( ~n621 & n694 ) | ( ~n621 & n695 ) | ( n694 & n695 ) ;
  assign n698 = ( n621 & ~n696 ) | ( n621 & n697 ) | ( ~n696 & n697 ) ;
  assign n699 = ( x71 & n693 ) | ( x71 & ~n698 ) | ( n693 & ~n698 ) ;
  assign n700 = ( x71 & n622 ) | ( x71 & ~n658 ) | ( n622 & ~n658 ) ;
  assign n701 = x71 & n622 ;
  assign n702 = ( ~n627 & n700 ) | ( ~n627 & n701 ) | ( n700 & n701 ) ;
  assign n703 = ( n627 & n700 ) | ( n627 & n701 ) | ( n700 & n701 ) ;
  assign n704 = ( n627 & n702 ) | ( n627 & ~n703 ) | ( n702 & ~n703 ) ;
  assign n705 = ( x72 & n699 ) | ( x72 & ~n704 ) | ( n699 & ~n704 ) ;
  assign n706 = ( x72 & n628 ) | ( x72 & ~n658 ) | ( n628 & ~n658 ) ;
  assign n707 = x72 & n628 ;
  assign n708 = ( n633 & n706 ) | ( n633 & n707 ) | ( n706 & n707 ) ;
  assign n709 = ( ~n633 & n706 ) | ( ~n633 & n707 ) | ( n706 & n707 ) ;
  assign n710 = ( n633 & ~n708 ) | ( n633 & n709 ) | ( ~n708 & n709 ) ;
  assign n711 = ( x73 & n705 ) | ( x73 & ~n710 ) | ( n705 & ~n710 ) ;
  assign n712 = ( x73 & n634 ) | ( x73 & ~n658 ) | ( n634 & ~n658 ) ;
  assign n713 = x73 & n634 ;
  assign n714 = ( ~n639 & n712 ) | ( ~n639 & n713 ) | ( n712 & n713 ) ;
  assign n715 = ( n639 & n712 ) | ( n639 & n713 ) | ( n712 & n713 ) ;
  assign n716 = ( n639 & n714 ) | ( n639 & ~n715 ) | ( n714 & ~n715 ) ;
  assign n717 = ( x74 & n711 ) | ( x74 & ~n716 ) | ( n711 & ~n716 ) ;
  assign n718 = ( x74 & n640 ) | ( x74 & ~n658 ) | ( n640 & ~n658 ) ;
  assign n719 = x74 & n640 ;
  assign n720 = ( n645 & n718 ) | ( n645 & n719 ) | ( n718 & n719 ) ;
  assign n721 = ( ~n645 & n718 ) | ( ~n645 & n719 ) | ( n718 & n719 ) ;
  assign n722 = ( n645 & ~n720 ) | ( n645 & n721 ) | ( ~n720 & n721 ) ;
  assign n723 = ( x75 & n717 ) | ( x75 & ~n722 ) | ( n717 & ~n722 ) ;
  assign n724 = ( x75 & n646 ) | ( x75 & ~n658 ) | ( n646 & ~n658 ) ;
  assign n725 = x75 & n646 ;
  assign n726 = ( n651 & n724 ) | ( n651 & n725 ) | ( n724 & n725 ) ;
  assign n727 = ( ~n651 & n724 ) | ( ~n651 & n725 ) | ( n724 & n725 ) ;
  assign n728 = ( n651 & ~n726 ) | ( n651 & n727 ) | ( ~n726 & n727 ) ;
  assign n729 = ( x76 & n723 ) | ( x76 & ~n728 ) | ( n723 & ~n728 ) ;
  assign n730 = x77 | n729 ;
  assign n731 = ( x77 & n180 ) | ( x77 & n729 ) | ( n180 & n729 ) ;
  assign n732 = ( n656 & ~n730 ) | ( n656 & n731 ) | ( ~n730 & n731 ) ;
  assign n733 = ( x77 & ~n656 ) | ( x77 & n729 ) | ( ~n656 & n729 ) ;
  assign n734 = n180 | n733 ;
  assign n735 = ( x50 & ~x64 ) | ( x50 & n734 ) | ( ~x64 & n734 ) ;
  assign n736 = ~x50 & n734 ;
  assign n737 = ( n662 & n735 ) | ( n662 & ~n736 ) | ( n735 & ~n736 ) ;
  assign n738 = ~x49 & x64 ;
  assign n739 = ( x65 & ~n737 ) | ( x65 & n738 ) | ( ~n737 & n738 ) ;
  assign n740 = ( x65 & n662 ) | ( x65 & ~n734 ) | ( n662 & ~n734 ) ;
  assign n741 = x65 & n662 ;
  assign n742 = ( n661 & n740 ) | ( n661 & n741 ) | ( n740 & n741 ) ;
  assign n743 = ( ~n661 & n740 ) | ( ~n661 & n741 ) | ( n740 & n741 ) ;
  assign n744 = ( n661 & ~n742 ) | ( n661 & n743 ) | ( ~n742 & n743 ) ;
  assign n745 = ( x66 & n739 ) | ( x66 & ~n744 ) | ( n739 & ~n744 ) ;
  assign n746 = ( x66 & n663 ) | ( x66 & n734 ) | ( n663 & n734 ) ;
  assign n747 = x66 | n663 ;
  assign n748 = ( ~n668 & n746 ) | ( ~n668 & n747 ) | ( n746 & n747 ) ;
  assign n749 = ( n668 & n746 ) | ( n668 & n747 ) | ( n746 & n747 ) ;
  assign n750 = ( n668 & n748 ) | ( n668 & ~n749 ) | ( n748 & ~n749 ) ;
  assign n751 = ( x67 & n745 ) | ( x67 & ~n750 ) | ( n745 & ~n750 ) ;
  assign n752 = ( x67 & n669 ) | ( x67 & ~n734 ) | ( n669 & ~n734 ) ;
  assign n753 = x67 & n669 ;
  assign n754 = ( ~n674 & n752 ) | ( ~n674 & n753 ) | ( n752 & n753 ) ;
  assign n755 = ( n674 & n752 ) | ( n674 & n753 ) | ( n752 & n753 ) ;
  assign n756 = ( n674 & n754 ) | ( n674 & ~n755 ) | ( n754 & ~n755 ) ;
  assign n757 = ( x68 & n751 ) | ( x68 & ~n756 ) | ( n751 & ~n756 ) ;
  assign n758 = ( x68 & n675 ) | ( x68 & ~n734 ) | ( n675 & ~n734 ) ;
  assign n759 = x68 & n675 ;
  assign n760 = ( n680 & n758 ) | ( n680 & n759 ) | ( n758 & n759 ) ;
  assign n761 = ( ~n680 & n758 ) | ( ~n680 & n759 ) | ( n758 & n759 ) ;
  assign n762 = ( n680 & ~n760 ) | ( n680 & n761 ) | ( ~n760 & n761 ) ;
  assign n763 = ( x69 & n757 ) | ( x69 & ~n762 ) | ( n757 & ~n762 ) ;
  assign n764 = ( x69 & n681 ) | ( x69 & ~n734 ) | ( n681 & ~n734 ) ;
  assign n765 = x69 & n681 ;
  assign n766 = ( ~n686 & n764 ) | ( ~n686 & n765 ) | ( n764 & n765 ) ;
  assign n767 = ( n686 & n764 ) | ( n686 & n765 ) | ( n764 & n765 ) ;
  assign n768 = ( n686 & n766 ) | ( n686 & ~n767 ) | ( n766 & ~n767 ) ;
  assign n769 = ( x70 & n763 ) | ( x70 & ~n768 ) | ( n763 & ~n768 ) ;
  assign n770 = ( x70 & n687 ) | ( x70 & ~n734 ) | ( n687 & ~n734 ) ;
  assign n771 = x70 & n687 ;
  assign n772 = ( n692 & n770 ) | ( n692 & n771 ) | ( n770 & n771 ) ;
  assign n773 = ( ~n692 & n770 ) | ( ~n692 & n771 ) | ( n770 & n771 ) ;
  assign n774 = ( n692 & ~n772 ) | ( n692 & n773 ) | ( ~n772 & n773 ) ;
  assign n775 = ( x71 & n769 ) | ( x71 & ~n774 ) | ( n769 & ~n774 ) ;
  assign n776 = ( x71 & n693 ) | ( x71 & ~n734 ) | ( n693 & ~n734 ) ;
  assign n777 = x71 & n693 ;
  assign n778 = ( ~n698 & n776 ) | ( ~n698 & n777 ) | ( n776 & n777 ) ;
  assign n779 = ( n698 & n776 ) | ( n698 & n777 ) | ( n776 & n777 ) ;
  assign n780 = ( n698 & n778 ) | ( n698 & ~n779 ) | ( n778 & ~n779 ) ;
  assign n781 = ( x72 & n775 ) | ( x72 & ~n780 ) | ( n775 & ~n780 ) ;
  assign n782 = ( x72 & n699 ) | ( x72 & ~n734 ) | ( n699 & ~n734 ) ;
  assign n783 = x72 & n699 ;
  assign n784 = ( n704 & n782 ) | ( n704 & n783 ) | ( n782 & n783 ) ;
  assign n785 = ( ~n704 & n782 ) | ( ~n704 & n783 ) | ( n782 & n783 ) ;
  assign n786 = ( n704 & ~n784 ) | ( n704 & n785 ) | ( ~n784 & n785 ) ;
  assign n787 = ( x73 & n781 ) | ( x73 & ~n786 ) | ( n781 & ~n786 ) ;
  assign n788 = ( x73 & n705 ) | ( x73 & ~n734 ) | ( n705 & ~n734 ) ;
  assign n789 = x73 & n705 ;
  assign n790 = ( ~n710 & n788 ) | ( ~n710 & n789 ) | ( n788 & n789 ) ;
  assign n791 = ( n710 & n788 ) | ( n710 & n789 ) | ( n788 & n789 ) ;
  assign n792 = ( n710 & n790 ) | ( n710 & ~n791 ) | ( n790 & ~n791 ) ;
  assign n793 = ( x74 & n787 ) | ( x74 & ~n792 ) | ( n787 & ~n792 ) ;
  assign n794 = ( x74 & n711 ) | ( x74 & ~n734 ) | ( n711 & ~n734 ) ;
  assign n795 = x74 & n711 ;
  assign n796 = ( n716 & n794 ) | ( n716 & n795 ) | ( n794 & n795 ) ;
  assign n797 = ( ~n716 & n794 ) | ( ~n716 & n795 ) | ( n794 & n795 ) ;
  assign n798 = ( n716 & ~n796 ) | ( n716 & n797 ) | ( ~n796 & n797 ) ;
  assign n799 = ( x75 & n793 ) | ( x75 & ~n798 ) | ( n793 & ~n798 ) ;
  assign n800 = ( x75 & n717 ) | ( x75 & ~n734 ) | ( n717 & ~n734 ) ;
  assign n801 = x75 & n717 ;
  assign n802 = ( ~n722 & n800 ) | ( ~n722 & n801 ) | ( n800 & n801 ) ;
  assign n803 = ( n722 & n800 ) | ( n722 & n801 ) | ( n800 & n801 ) ;
  assign n804 = ( n722 & n802 ) | ( n722 & ~n803 ) | ( n802 & ~n803 ) ;
  assign n805 = ( x76 & n799 ) | ( x76 & ~n804 ) | ( n799 & ~n804 ) ;
  assign n806 = ( x76 & n723 ) | ( x76 & ~n734 ) | ( n723 & ~n734 ) ;
  assign n807 = x76 & n723 ;
  assign n808 = ( ~n728 & n806 ) | ( ~n728 & n807 ) | ( n806 & n807 ) ;
  assign n809 = ( n728 & n806 ) | ( n728 & n807 ) | ( n806 & n807 ) ;
  assign n810 = ( n728 & n808 ) | ( n728 & ~n809 ) | ( n808 & ~n809 ) ;
  assign n811 = ( x77 & n805 ) | ( x77 & ~n810 ) | ( n805 & ~n810 ) ;
  assign n812 = x78 | n811 ;
  assign n813 = x79 | n178 ;
  assign n814 = ( x78 & n811 ) | ( x78 & n813 ) | ( n811 & n813 ) ;
  assign n815 = ( n732 & ~n812 ) | ( n732 & n814 ) | ( ~n812 & n814 ) ;
  assign n816 = ( x78 & ~n732 ) | ( x78 & n811 ) | ( ~n732 & n811 ) ;
  assign n817 = n813 | n816 ;
  assign n818 = ( x49 & ~x64 ) | ( x49 & n817 ) | ( ~x64 & n817 ) ;
  assign n819 = ~x49 & n817 ;
  assign n820 = ( n738 & n818 ) | ( n738 & ~n819 ) | ( n818 & ~n819 ) ;
  assign n821 = ~x48 & x64 ;
  assign n822 = ( x65 & ~n820 ) | ( x65 & n821 ) | ( ~n820 & n821 ) ;
  assign n823 = ( x65 & n738 ) | ( x65 & ~n817 ) | ( n738 & ~n817 ) ;
  assign n824 = x65 & n738 ;
  assign n825 = ( n737 & n823 ) | ( n737 & n824 ) | ( n823 & n824 ) ;
  assign n826 = ( ~n737 & n823 ) | ( ~n737 & n824 ) | ( n823 & n824 ) ;
  assign n827 = ( n737 & ~n825 ) | ( n737 & n826 ) | ( ~n825 & n826 ) ;
  assign n828 = ( x66 & n822 ) | ( x66 & ~n827 ) | ( n822 & ~n827 ) ;
  assign n829 = ( x66 & n739 ) | ( x66 & n817 ) | ( n739 & n817 ) ;
  assign n830 = x66 | n739 ;
  assign n831 = ( ~n744 & n829 ) | ( ~n744 & n830 ) | ( n829 & n830 ) ;
  assign n832 = ( n744 & n829 ) | ( n744 & n830 ) | ( n829 & n830 ) ;
  assign n833 = ( n744 & n831 ) | ( n744 & ~n832 ) | ( n831 & ~n832 ) ;
  assign n834 = ( x67 & n828 ) | ( x67 & ~n833 ) | ( n828 & ~n833 ) ;
  assign n835 = ( x67 & n745 ) | ( x67 & ~n817 ) | ( n745 & ~n817 ) ;
  assign n836 = x67 & n745 ;
  assign n837 = ( ~n750 & n835 ) | ( ~n750 & n836 ) | ( n835 & n836 ) ;
  assign n838 = ( n750 & n835 ) | ( n750 & n836 ) | ( n835 & n836 ) ;
  assign n839 = ( n750 & n837 ) | ( n750 & ~n838 ) | ( n837 & ~n838 ) ;
  assign n840 = ( x68 & n834 ) | ( x68 & ~n839 ) | ( n834 & ~n839 ) ;
  assign n841 = ( x68 & n751 ) | ( x68 & ~n817 ) | ( n751 & ~n817 ) ;
  assign n842 = x68 & n751 ;
  assign n843 = ( n756 & n841 ) | ( n756 & n842 ) | ( n841 & n842 ) ;
  assign n844 = ( ~n756 & n841 ) | ( ~n756 & n842 ) | ( n841 & n842 ) ;
  assign n845 = ( n756 & ~n843 ) | ( n756 & n844 ) | ( ~n843 & n844 ) ;
  assign n846 = ( x69 & n840 ) | ( x69 & ~n845 ) | ( n840 & ~n845 ) ;
  assign n847 = ( x69 & n757 ) | ( x69 & ~n817 ) | ( n757 & ~n817 ) ;
  assign n848 = x69 & n757 ;
  assign n849 = ( ~n762 & n847 ) | ( ~n762 & n848 ) | ( n847 & n848 ) ;
  assign n850 = ( n762 & n847 ) | ( n762 & n848 ) | ( n847 & n848 ) ;
  assign n851 = ( n762 & n849 ) | ( n762 & ~n850 ) | ( n849 & ~n850 ) ;
  assign n852 = ( x70 & n846 ) | ( x70 & ~n851 ) | ( n846 & ~n851 ) ;
  assign n853 = ( x70 & n763 ) | ( x70 & ~n817 ) | ( n763 & ~n817 ) ;
  assign n854 = x70 & n763 ;
  assign n855 = ( n768 & n853 ) | ( n768 & n854 ) | ( n853 & n854 ) ;
  assign n856 = ( ~n768 & n853 ) | ( ~n768 & n854 ) | ( n853 & n854 ) ;
  assign n857 = ( n768 & ~n855 ) | ( n768 & n856 ) | ( ~n855 & n856 ) ;
  assign n858 = ( x71 & n852 ) | ( x71 & ~n857 ) | ( n852 & ~n857 ) ;
  assign n859 = ( x71 & n769 ) | ( x71 & ~n817 ) | ( n769 & ~n817 ) ;
  assign n860 = x71 & n769 ;
  assign n861 = ( ~n774 & n859 ) | ( ~n774 & n860 ) | ( n859 & n860 ) ;
  assign n862 = ( n774 & n859 ) | ( n774 & n860 ) | ( n859 & n860 ) ;
  assign n863 = ( n774 & n861 ) | ( n774 & ~n862 ) | ( n861 & ~n862 ) ;
  assign n864 = ( x72 & n858 ) | ( x72 & ~n863 ) | ( n858 & ~n863 ) ;
  assign n865 = ( x72 & n775 ) | ( x72 & ~n817 ) | ( n775 & ~n817 ) ;
  assign n866 = x72 & n775 ;
  assign n867 = ( n780 & n865 ) | ( n780 & n866 ) | ( n865 & n866 ) ;
  assign n868 = ( ~n780 & n865 ) | ( ~n780 & n866 ) | ( n865 & n866 ) ;
  assign n869 = ( n780 & ~n867 ) | ( n780 & n868 ) | ( ~n867 & n868 ) ;
  assign n870 = ( x73 & n864 ) | ( x73 & ~n869 ) | ( n864 & ~n869 ) ;
  assign n871 = ( x73 & n781 ) | ( x73 & ~n817 ) | ( n781 & ~n817 ) ;
  assign n872 = x73 & n781 ;
  assign n873 = ( ~n786 & n871 ) | ( ~n786 & n872 ) | ( n871 & n872 ) ;
  assign n874 = ( n786 & n871 ) | ( n786 & n872 ) | ( n871 & n872 ) ;
  assign n875 = ( n786 & n873 ) | ( n786 & ~n874 ) | ( n873 & ~n874 ) ;
  assign n876 = ( x74 & n870 ) | ( x74 & ~n875 ) | ( n870 & ~n875 ) ;
  assign n877 = ( x74 & n787 ) | ( x74 & ~n817 ) | ( n787 & ~n817 ) ;
  assign n878 = x74 & n787 ;
  assign n879 = ( n792 & n877 ) | ( n792 & n878 ) | ( n877 & n878 ) ;
  assign n880 = ( ~n792 & n877 ) | ( ~n792 & n878 ) | ( n877 & n878 ) ;
  assign n881 = ( n792 & ~n879 ) | ( n792 & n880 ) | ( ~n879 & n880 ) ;
  assign n882 = ( x75 & n876 ) | ( x75 & ~n881 ) | ( n876 & ~n881 ) ;
  assign n883 = ( x75 & n793 ) | ( x75 & ~n817 ) | ( n793 & ~n817 ) ;
  assign n884 = x75 & n793 ;
  assign n885 = ( ~n798 & n883 ) | ( ~n798 & n884 ) | ( n883 & n884 ) ;
  assign n886 = ( n798 & n883 ) | ( n798 & n884 ) | ( n883 & n884 ) ;
  assign n887 = ( n798 & n885 ) | ( n798 & ~n886 ) | ( n885 & ~n886 ) ;
  assign n888 = ( x76 & n882 ) | ( x76 & ~n887 ) | ( n882 & ~n887 ) ;
  assign n889 = ( x76 & n799 ) | ( x76 & ~n817 ) | ( n799 & ~n817 ) ;
  assign n890 = x76 & n799 ;
  assign n891 = ( n804 & n889 ) | ( n804 & n890 ) | ( n889 & n890 ) ;
  assign n892 = ( ~n804 & n889 ) | ( ~n804 & n890 ) | ( n889 & n890 ) ;
  assign n893 = ( n804 & ~n891 ) | ( n804 & n892 ) | ( ~n891 & n892 ) ;
  assign n894 = ( x77 & n888 ) | ( x77 & ~n893 ) | ( n888 & ~n893 ) ;
  assign n895 = ( x77 & n805 ) | ( x77 & ~n817 ) | ( n805 & ~n817 ) ;
  assign n896 = x77 & n805 ;
  assign n897 = ( n810 & n895 ) | ( n810 & n896 ) | ( n895 & n896 ) ;
  assign n898 = ( ~n810 & n895 ) | ( ~n810 & n896 ) | ( n895 & n896 ) ;
  assign n899 = ( n810 & ~n897 ) | ( n810 & n898 ) | ( ~n897 & n898 ) ;
  assign n900 = ( x78 & n894 ) | ( x78 & ~n899 ) | ( n894 & ~n899 ) ;
  assign n901 = x79 | n900 ;
  assign n902 = ( x79 & n178 ) | ( x79 & n900 ) | ( n178 & n900 ) ;
  assign n903 = ( n815 & ~n901 ) | ( n815 & n902 ) | ( ~n901 & n902 ) ;
  assign n904 = ( x79 & ~n815 ) | ( x79 & n900 ) | ( ~n815 & n900 ) ;
  assign n905 = n178 | n904 ;
  assign n906 = ( x48 & ~x64 ) | ( x48 & n905 ) | ( ~x64 & n905 ) ;
  assign n907 = ~x48 & n905 ;
  assign n908 = ( n821 & n906 ) | ( n821 & ~n907 ) | ( n906 & ~n907 ) ;
  assign n909 = ~x47 & x64 ;
  assign n910 = ( x65 & ~n908 ) | ( x65 & n909 ) | ( ~n908 & n909 ) ;
  assign n911 = ( x65 & n821 ) | ( x65 & ~n905 ) | ( n821 & ~n905 ) ;
  assign n912 = x65 & n821 ;
  assign n913 = ( n820 & n911 ) | ( n820 & n912 ) | ( n911 & n912 ) ;
  assign n914 = ( ~n820 & n911 ) | ( ~n820 & n912 ) | ( n911 & n912 ) ;
  assign n915 = ( n820 & ~n913 ) | ( n820 & n914 ) | ( ~n913 & n914 ) ;
  assign n916 = ( x66 & n910 ) | ( x66 & ~n915 ) | ( n910 & ~n915 ) ;
  assign n917 = ( x66 & n822 ) | ( x66 & ~n905 ) | ( n822 & ~n905 ) ;
  assign n918 = x66 & n822 ;
  assign n919 = ( n827 & n917 ) | ( n827 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ( ~n827 & n917 ) | ( ~n827 & n918 ) | ( n917 & n918 ) ;
  assign n921 = ( n827 & ~n919 ) | ( n827 & n920 ) | ( ~n919 & n920 ) ;
  assign n922 = ( x67 & n916 ) | ( x67 & ~n921 ) | ( n916 & ~n921 ) ;
  assign n923 = ( x67 & n828 ) | ( x67 & ~n905 ) | ( n828 & ~n905 ) ;
  assign n924 = x67 & n828 ;
  assign n925 = ( ~n833 & n923 ) | ( ~n833 & n924 ) | ( n923 & n924 ) ;
  assign n926 = ( n833 & n923 ) | ( n833 & n924 ) | ( n923 & n924 ) ;
  assign n927 = ( n833 & n925 ) | ( n833 & ~n926 ) | ( n925 & ~n926 ) ;
  assign n928 = ( x68 & n922 ) | ( x68 & ~n927 ) | ( n922 & ~n927 ) ;
  assign n929 = ( x68 & n834 ) | ( x68 & ~n905 ) | ( n834 & ~n905 ) ;
  assign n930 = x68 & n834 ;
  assign n931 = ( n839 & n929 ) | ( n839 & n930 ) | ( n929 & n930 ) ;
  assign n932 = ( ~n839 & n929 ) | ( ~n839 & n930 ) | ( n929 & n930 ) ;
  assign n933 = ( n839 & ~n931 ) | ( n839 & n932 ) | ( ~n931 & n932 ) ;
  assign n934 = ( x69 & n928 ) | ( x69 & ~n933 ) | ( n928 & ~n933 ) ;
  assign n935 = ( x69 & n840 ) | ( x69 & ~n905 ) | ( n840 & ~n905 ) ;
  assign n936 = x69 & n840 ;
  assign n937 = ( ~n845 & n935 ) | ( ~n845 & n936 ) | ( n935 & n936 ) ;
  assign n938 = ( n845 & n935 ) | ( n845 & n936 ) | ( n935 & n936 ) ;
  assign n939 = ( n845 & n937 ) | ( n845 & ~n938 ) | ( n937 & ~n938 ) ;
  assign n940 = ( x70 & n934 ) | ( x70 & ~n939 ) | ( n934 & ~n939 ) ;
  assign n941 = ( x70 & n846 ) | ( x70 & ~n905 ) | ( n846 & ~n905 ) ;
  assign n942 = x70 & n846 ;
  assign n943 = ( n851 & n941 ) | ( n851 & n942 ) | ( n941 & n942 ) ;
  assign n944 = ( ~n851 & n941 ) | ( ~n851 & n942 ) | ( n941 & n942 ) ;
  assign n945 = ( n851 & ~n943 ) | ( n851 & n944 ) | ( ~n943 & n944 ) ;
  assign n946 = ( x71 & n940 ) | ( x71 & ~n945 ) | ( n940 & ~n945 ) ;
  assign n947 = ( x71 & n852 ) | ( x71 & ~n905 ) | ( n852 & ~n905 ) ;
  assign n948 = x71 & n852 ;
  assign n949 = ( ~n857 & n947 ) | ( ~n857 & n948 ) | ( n947 & n948 ) ;
  assign n950 = ( n857 & n947 ) | ( n857 & n948 ) | ( n947 & n948 ) ;
  assign n951 = ( n857 & n949 ) | ( n857 & ~n950 ) | ( n949 & ~n950 ) ;
  assign n952 = ( x72 & n946 ) | ( x72 & ~n951 ) | ( n946 & ~n951 ) ;
  assign n953 = ( x72 & n858 ) | ( x72 & ~n905 ) | ( n858 & ~n905 ) ;
  assign n954 = x72 & n858 ;
  assign n955 = ( n863 & n953 ) | ( n863 & n954 ) | ( n953 & n954 ) ;
  assign n956 = ( ~n863 & n953 ) | ( ~n863 & n954 ) | ( n953 & n954 ) ;
  assign n957 = ( n863 & ~n955 ) | ( n863 & n956 ) | ( ~n955 & n956 ) ;
  assign n958 = ( x73 & n952 ) | ( x73 & ~n957 ) | ( n952 & ~n957 ) ;
  assign n959 = ( x73 & n864 ) | ( x73 & ~n905 ) | ( n864 & ~n905 ) ;
  assign n960 = x73 & n864 ;
  assign n961 = ( ~n869 & n959 ) | ( ~n869 & n960 ) | ( n959 & n960 ) ;
  assign n962 = ( n869 & n959 ) | ( n869 & n960 ) | ( n959 & n960 ) ;
  assign n963 = ( n869 & n961 ) | ( n869 & ~n962 ) | ( n961 & ~n962 ) ;
  assign n964 = ( x74 & n958 ) | ( x74 & ~n963 ) | ( n958 & ~n963 ) ;
  assign n965 = ( x74 & n870 ) | ( x74 & ~n905 ) | ( n870 & ~n905 ) ;
  assign n966 = x74 & n870 ;
  assign n967 = ( n875 & n965 ) | ( n875 & n966 ) | ( n965 & n966 ) ;
  assign n968 = ( ~n875 & n965 ) | ( ~n875 & n966 ) | ( n965 & n966 ) ;
  assign n969 = ( n875 & ~n967 ) | ( n875 & n968 ) | ( ~n967 & n968 ) ;
  assign n970 = ( x75 & n964 ) | ( x75 & ~n969 ) | ( n964 & ~n969 ) ;
  assign n971 = ( x75 & n876 ) | ( x75 & ~n905 ) | ( n876 & ~n905 ) ;
  assign n972 = x75 & n876 ;
  assign n973 = ( ~n881 & n971 ) | ( ~n881 & n972 ) | ( n971 & n972 ) ;
  assign n974 = ( n881 & n971 ) | ( n881 & n972 ) | ( n971 & n972 ) ;
  assign n975 = ( n881 & n973 ) | ( n881 & ~n974 ) | ( n973 & ~n974 ) ;
  assign n976 = ( x76 & n970 ) | ( x76 & ~n975 ) | ( n970 & ~n975 ) ;
  assign n977 = ( x76 & n882 ) | ( x76 & ~n905 ) | ( n882 & ~n905 ) ;
  assign n978 = x76 & n882 ;
  assign n979 = ( n887 & n977 ) | ( n887 & n978 ) | ( n977 & n978 ) ;
  assign n980 = ( ~n887 & n977 ) | ( ~n887 & n978 ) | ( n977 & n978 ) ;
  assign n981 = ( n887 & ~n979 ) | ( n887 & n980 ) | ( ~n979 & n980 ) ;
  assign n982 = ( x77 & n976 ) | ( x77 & ~n981 ) | ( n976 & ~n981 ) ;
  assign n983 = ( x77 & n888 ) | ( x77 & ~n905 ) | ( n888 & ~n905 ) ;
  assign n984 = x77 & n888 ;
  assign n985 = ( ~n893 & n983 ) | ( ~n893 & n984 ) | ( n983 & n984 ) ;
  assign n986 = ( n893 & n983 ) | ( n893 & n984 ) | ( n983 & n984 ) ;
  assign n987 = ( n893 & n985 ) | ( n893 & ~n986 ) | ( n985 & ~n986 ) ;
  assign n988 = ( x78 & n982 ) | ( x78 & ~n987 ) | ( n982 & ~n987 ) ;
  assign n989 = ( x78 & n894 ) | ( x78 & ~n905 ) | ( n894 & ~n905 ) ;
  assign n990 = x78 & n894 ;
  assign n991 = ( ~n899 & n989 ) | ( ~n899 & n990 ) | ( n989 & n990 ) ;
  assign n992 = ( n899 & n989 ) | ( n899 & n990 ) | ( n989 & n990 ) ;
  assign n993 = ( n899 & n991 ) | ( n899 & ~n992 ) | ( n991 & ~n992 ) ;
  assign n994 = ( x79 & n988 ) | ( x79 & ~n993 ) | ( n988 & ~n993 ) ;
  assign n995 = x80 | n994 ;
  assign n996 = x81 | x82 ;
  assign n997 = x83 | n174 ;
  assign n998 = n996 | n997 ;
  assign n999 = ( x80 & n994 ) | ( x80 & n998 ) | ( n994 & n998 ) ;
  assign n1000 = ( n903 & ~n995 ) | ( n903 & n999 ) | ( ~n995 & n999 ) ;
  assign n1001 = ( x80 & ~n903 ) | ( x80 & n994 ) | ( ~n903 & n994 ) ;
  assign n1002 = n998 | n1001 ;
  assign n1003 = ( x47 & ~x64 ) | ( x47 & n1002 ) | ( ~x64 & n1002 ) ;
  assign n1004 = ~x47 & n1002 ;
  assign n1005 = ( n909 & n1003 ) | ( n909 & ~n1004 ) | ( n1003 & ~n1004 ) ;
  assign n1006 = ~x46 & x64 ;
  assign n1007 = ( x65 & ~n1005 ) | ( x65 & n1006 ) | ( ~n1005 & n1006 ) ;
  assign n1008 = ( x65 & n909 ) | ( x65 & ~n1002 ) | ( n909 & ~n1002 ) ;
  assign n1009 = x65 & n909 ;
  assign n1010 = ( n908 & n1008 ) | ( n908 & n1009 ) | ( n1008 & n1009 ) ;
  assign n1011 = ( ~n908 & n1008 ) | ( ~n908 & n1009 ) | ( n1008 & n1009 ) ;
  assign n1012 = ( n908 & ~n1010 ) | ( n908 & n1011 ) | ( ~n1010 & n1011 ) ;
  assign n1013 = ( x66 & n1007 ) | ( x66 & ~n1012 ) | ( n1007 & ~n1012 ) ;
  assign n1014 = ( x66 & n910 ) | ( x66 & n1002 ) | ( n910 & n1002 ) ;
  assign n1015 = x66 | n910 ;
  assign n1016 = ( ~n915 & n1014 ) | ( ~n915 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1017 = ( n915 & n1014 ) | ( n915 & n1015 ) | ( n1014 & n1015 ) ;
  assign n1018 = ( n915 & n1016 ) | ( n915 & ~n1017 ) | ( n1016 & ~n1017 ) ;
  assign n1019 = ( x67 & n1013 ) | ( x67 & ~n1018 ) | ( n1013 & ~n1018 ) ;
  assign n1020 = ( x67 & n916 ) | ( x67 & ~n1002 ) | ( n916 & ~n1002 ) ;
  assign n1021 = x67 & n916 ;
  assign n1022 = ( ~n921 & n1020 ) | ( ~n921 & n1021 ) | ( n1020 & n1021 ) ;
  assign n1023 = ( n921 & n1020 ) | ( n921 & n1021 ) | ( n1020 & n1021 ) ;
  assign n1024 = ( n921 & n1022 ) | ( n921 & ~n1023 ) | ( n1022 & ~n1023 ) ;
  assign n1025 = ( x68 & n1019 ) | ( x68 & ~n1024 ) | ( n1019 & ~n1024 ) ;
  assign n1026 = ( x68 & n922 ) | ( x68 & ~n1002 ) | ( n922 & ~n1002 ) ;
  assign n1027 = x68 & n922 ;
  assign n1028 = ( n927 & n1026 ) | ( n927 & n1027 ) | ( n1026 & n1027 ) ;
  assign n1029 = ( ~n927 & n1026 ) | ( ~n927 & n1027 ) | ( n1026 & n1027 ) ;
  assign n1030 = ( n927 & ~n1028 ) | ( n927 & n1029 ) | ( ~n1028 & n1029 ) ;
  assign n1031 = ( x69 & n1025 ) | ( x69 & ~n1030 ) | ( n1025 & ~n1030 ) ;
  assign n1032 = ( x69 & n928 ) | ( x69 & ~n1002 ) | ( n928 & ~n1002 ) ;
  assign n1033 = x69 & n928 ;
  assign n1034 = ( ~n933 & n1032 ) | ( ~n933 & n1033 ) | ( n1032 & n1033 ) ;
  assign n1035 = ( n933 & n1032 ) | ( n933 & n1033 ) | ( n1032 & n1033 ) ;
  assign n1036 = ( n933 & n1034 ) | ( n933 & ~n1035 ) | ( n1034 & ~n1035 ) ;
  assign n1037 = ( x70 & n1031 ) | ( x70 & ~n1036 ) | ( n1031 & ~n1036 ) ;
  assign n1038 = ( x70 & n934 ) | ( x70 & ~n1002 ) | ( n934 & ~n1002 ) ;
  assign n1039 = x70 & n934 ;
  assign n1040 = ( n939 & n1038 ) | ( n939 & n1039 ) | ( n1038 & n1039 ) ;
  assign n1041 = ( ~n939 & n1038 ) | ( ~n939 & n1039 ) | ( n1038 & n1039 ) ;
  assign n1042 = ( n939 & ~n1040 ) | ( n939 & n1041 ) | ( ~n1040 & n1041 ) ;
  assign n1043 = ( x71 & n1037 ) | ( x71 & ~n1042 ) | ( n1037 & ~n1042 ) ;
  assign n1044 = ( x71 & n940 ) | ( x71 & ~n1002 ) | ( n940 & ~n1002 ) ;
  assign n1045 = x71 & n940 ;
  assign n1046 = ( ~n945 & n1044 ) | ( ~n945 & n1045 ) | ( n1044 & n1045 ) ;
  assign n1047 = ( n945 & n1044 ) | ( n945 & n1045 ) | ( n1044 & n1045 ) ;
  assign n1048 = ( n945 & n1046 ) | ( n945 & ~n1047 ) | ( n1046 & ~n1047 ) ;
  assign n1049 = ( x72 & n1043 ) | ( x72 & ~n1048 ) | ( n1043 & ~n1048 ) ;
  assign n1050 = ( x72 & n946 ) | ( x72 & ~n1002 ) | ( n946 & ~n1002 ) ;
  assign n1051 = x72 & n946 ;
  assign n1052 = ( n951 & n1050 ) | ( n951 & n1051 ) | ( n1050 & n1051 ) ;
  assign n1053 = ( ~n951 & n1050 ) | ( ~n951 & n1051 ) | ( n1050 & n1051 ) ;
  assign n1054 = ( n951 & ~n1052 ) | ( n951 & n1053 ) | ( ~n1052 & n1053 ) ;
  assign n1055 = ( x73 & n1049 ) | ( x73 & ~n1054 ) | ( n1049 & ~n1054 ) ;
  assign n1056 = ( x73 & n952 ) | ( x73 & ~n1002 ) | ( n952 & ~n1002 ) ;
  assign n1057 = x73 & n952 ;
  assign n1058 = ( ~n957 & n1056 ) | ( ~n957 & n1057 ) | ( n1056 & n1057 ) ;
  assign n1059 = ( n957 & n1056 ) | ( n957 & n1057 ) | ( n1056 & n1057 ) ;
  assign n1060 = ( n957 & n1058 ) | ( n957 & ~n1059 ) | ( n1058 & ~n1059 ) ;
  assign n1061 = ( x74 & n1055 ) | ( x74 & ~n1060 ) | ( n1055 & ~n1060 ) ;
  assign n1062 = ( x74 & n958 ) | ( x74 & ~n1002 ) | ( n958 & ~n1002 ) ;
  assign n1063 = x74 & n958 ;
  assign n1064 = ( n963 & n1062 ) | ( n963 & n1063 ) | ( n1062 & n1063 ) ;
  assign n1065 = ( ~n963 & n1062 ) | ( ~n963 & n1063 ) | ( n1062 & n1063 ) ;
  assign n1066 = ( n963 & ~n1064 ) | ( n963 & n1065 ) | ( ~n1064 & n1065 ) ;
  assign n1067 = ( x75 & n1061 ) | ( x75 & ~n1066 ) | ( n1061 & ~n1066 ) ;
  assign n1068 = ( x75 & n964 ) | ( x75 & ~n1002 ) | ( n964 & ~n1002 ) ;
  assign n1069 = x75 & n964 ;
  assign n1070 = ( ~n969 & n1068 ) | ( ~n969 & n1069 ) | ( n1068 & n1069 ) ;
  assign n1071 = ( n969 & n1068 ) | ( n969 & n1069 ) | ( n1068 & n1069 ) ;
  assign n1072 = ( n969 & n1070 ) | ( n969 & ~n1071 ) | ( n1070 & ~n1071 ) ;
  assign n1073 = ( x76 & n1067 ) | ( x76 & ~n1072 ) | ( n1067 & ~n1072 ) ;
  assign n1074 = ( x76 & n970 ) | ( x76 & ~n1002 ) | ( n970 & ~n1002 ) ;
  assign n1075 = x76 & n970 ;
  assign n1076 = ( n975 & n1074 ) | ( n975 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1077 = ( ~n975 & n1074 ) | ( ~n975 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1078 = ( n975 & ~n1076 ) | ( n975 & n1077 ) | ( ~n1076 & n1077 ) ;
  assign n1079 = ( x77 & n1073 ) | ( x77 & ~n1078 ) | ( n1073 & ~n1078 ) ;
  assign n1080 = ( x77 & n976 ) | ( x77 & ~n1002 ) | ( n976 & ~n1002 ) ;
  assign n1081 = x77 & n976 ;
  assign n1082 = ( ~n981 & n1080 ) | ( ~n981 & n1081 ) | ( n1080 & n1081 ) ;
  assign n1083 = ( n981 & n1080 ) | ( n981 & n1081 ) | ( n1080 & n1081 ) ;
  assign n1084 = ( n981 & n1082 ) | ( n981 & ~n1083 ) | ( n1082 & ~n1083 ) ;
  assign n1085 = ( x78 & n1079 ) | ( x78 & ~n1084 ) | ( n1079 & ~n1084 ) ;
  assign n1086 = ( x78 & n982 ) | ( x78 & ~n1002 ) | ( n982 & ~n1002 ) ;
  assign n1087 = x78 & n982 ;
  assign n1088 = ( n987 & n1086 ) | ( n987 & n1087 ) | ( n1086 & n1087 ) ;
  assign n1089 = ( ~n987 & n1086 ) | ( ~n987 & n1087 ) | ( n1086 & n1087 ) ;
  assign n1090 = ( n987 & ~n1088 ) | ( n987 & n1089 ) | ( ~n1088 & n1089 ) ;
  assign n1091 = ( x79 & n1085 ) | ( x79 & ~n1090 ) | ( n1085 & ~n1090 ) ;
  assign n1092 = ( x79 & n988 ) | ( x79 & ~n1002 ) | ( n988 & ~n1002 ) ;
  assign n1093 = x79 & n988 ;
  assign n1094 = ( n993 & n1092 ) | ( n993 & n1093 ) | ( n1092 & n1093 ) ;
  assign n1095 = ( ~n993 & n1092 ) | ( ~n993 & n1093 ) | ( n1092 & n1093 ) ;
  assign n1096 = ( n993 & ~n1094 ) | ( n993 & n1095 ) | ( ~n1094 & n1095 ) ;
  assign n1097 = ( x80 & n1091 ) | ( x80 & ~n1096 ) | ( n1091 & ~n1096 ) ;
  assign n1098 = ( n998 & ~n1000 ) | ( n998 & n1097 ) | ( ~n1000 & n1097 ) ;
  assign n1099 = n176 | n1098 ;
  assign n1100 = n1000 & n1099 ;
  assign n1101 = n280 | n1100 ;
  assign n1102 = ( x46 & ~x64 ) | ( x46 & n1099 ) | ( ~x64 & n1099 ) ;
  assign n1103 = ~x46 & n1099 ;
  assign n1104 = ( n1006 & n1102 ) | ( n1006 & ~n1103 ) | ( n1102 & ~n1103 ) ;
  assign n1105 = ~x45 & x64 ;
  assign n1106 = ( x65 & ~n1104 ) | ( x65 & n1105 ) | ( ~n1104 & n1105 ) ;
  assign n1107 = ( x65 & n1006 ) | ( x65 & ~n1099 ) | ( n1006 & ~n1099 ) ;
  assign n1108 = x65 & n1006 ;
  assign n1109 = ( n1005 & n1107 ) | ( n1005 & n1108 ) | ( n1107 & n1108 ) ;
  assign n1110 = ( ~n1005 & n1107 ) | ( ~n1005 & n1108 ) | ( n1107 & n1108 ) ;
  assign n1111 = ( n1005 & ~n1109 ) | ( n1005 & n1110 ) | ( ~n1109 & n1110 ) ;
  assign n1112 = ( x66 & n1106 ) | ( x66 & ~n1111 ) | ( n1106 & ~n1111 ) ;
  assign n1113 = ( x66 & n1007 ) | ( x66 & ~n1099 ) | ( n1007 & ~n1099 ) ;
  assign n1114 = x66 & n1007 ;
  assign n1115 = ( n1012 & n1113 ) | ( n1012 & n1114 ) | ( n1113 & n1114 ) ;
  assign n1116 = ( ~n1012 & n1113 ) | ( ~n1012 & n1114 ) | ( n1113 & n1114 ) ;
  assign n1117 = ( n1012 & ~n1115 ) | ( n1012 & n1116 ) | ( ~n1115 & n1116 ) ;
  assign n1118 = ( x67 & n1112 ) | ( x67 & ~n1117 ) | ( n1112 & ~n1117 ) ;
  assign n1119 = ( x67 & n1013 ) | ( x67 & ~n1099 ) | ( n1013 & ~n1099 ) ;
  assign n1120 = x67 & n1013 ;
  assign n1121 = ( ~n1018 & n1119 ) | ( ~n1018 & n1120 ) | ( n1119 & n1120 ) ;
  assign n1122 = ( n1018 & n1119 ) | ( n1018 & n1120 ) | ( n1119 & n1120 ) ;
  assign n1123 = ( n1018 & n1121 ) | ( n1018 & ~n1122 ) | ( n1121 & ~n1122 ) ;
  assign n1124 = ( x68 & n1118 ) | ( x68 & ~n1123 ) | ( n1118 & ~n1123 ) ;
  assign n1125 = ( x68 & n1019 ) | ( x68 & ~n1099 ) | ( n1019 & ~n1099 ) ;
  assign n1126 = x68 & n1019 ;
  assign n1127 = ( n1024 & n1125 ) | ( n1024 & n1126 ) | ( n1125 & n1126 ) ;
  assign n1128 = ( ~n1024 & n1125 ) | ( ~n1024 & n1126 ) | ( n1125 & n1126 ) ;
  assign n1129 = ( n1024 & ~n1127 ) | ( n1024 & n1128 ) | ( ~n1127 & n1128 ) ;
  assign n1130 = ( x69 & n1124 ) | ( x69 & ~n1129 ) | ( n1124 & ~n1129 ) ;
  assign n1131 = ( x69 & n1025 ) | ( x69 & ~n1099 ) | ( n1025 & ~n1099 ) ;
  assign n1132 = x69 & n1025 ;
  assign n1133 = ( ~n1030 & n1131 ) | ( ~n1030 & n1132 ) | ( n1131 & n1132 ) ;
  assign n1134 = ( n1030 & n1131 ) | ( n1030 & n1132 ) | ( n1131 & n1132 ) ;
  assign n1135 = ( n1030 & n1133 ) | ( n1030 & ~n1134 ) | ( n1133 & ~n1134 ) ;
  assign n1136 = ( x70 & n1130 ) | ( x70 & ~n1135 ) | ( n1130 & ~n1135 ) ;
  assign n1137 = ( x70 & n1031 ) | ( x70 & ~n1099 ) | ( n1031 & ~n1099 ) ;
  assign n1138 = x70 & n1031 ;
  assign n1139 = ( n1036 & n1137 ) | ( n1036 & n1138 ) | ( n1137 & n1138 ) ;
  assign n1140 = ( ~n1036 & n1137 ) | ( ~n1036 & n1138 ) | ( n1137 & n1138 ) ;
  assign n1141 = ( n1036 & ~n1139 ) | ( n1036 & n1140 ) | ( ~n1139 & n1140 ) ;
  assign n1142 = ( x71 & n1136 ) | ( x71 & ~n1141 ) | ( n1136 & ~n1141 ) ;
  assign n1143 = ( x71 & n1037 ) | ( x71 & ~n1099 ) | ( n1037 & ~n1099 ) ;
  assign n1144 = x71 & n1037 ;
  assign n1145 = ( ~n1042 & n1143 ) | ( ~n1042 & n1144 ) | ( n1143 & n1144 ) ;
  assign n1146 = ( n1042 & n1143 ) | ( n1042 & n1144 ) | ( n1143 & n1144 ) ;
  assign n1147 = ( n1042 & n1145 ) | ( n1042 & ~n1146 ) | ( n1145 & ~n1146 ) ;
  assign n1148 = ( x72 & n1142 ) | ( x72 & ~n1147 ) | ( n1142 & ~n1147 ) ;
  assign n1149 = ( x72 & n1043 ) | ( x72 & ~n1099 ) | ( n1043 & ~n1099 ) ;
  assign n1150 = x72 & n1043 ;
  assign n1151 = ( n1048 & n1149 ) | ( n1048 & n1150 ) | ( n1149 & n1150 ) ;
  assign n1152 = ( ~n1048 & n1149 ) | ( ~n1048 & n1150 ) | ( n1149 & n1150 ) ;
  assign n1153 = ( n1048 & ~n1151 ) | ( n1048 & n1152 ) | ( ~n1151 & n1152 ) ;
  assign n1154 = ( x73 & n1148 ) | ( x73 & ~n1153 ) | ( n1148 & ~n1153 ) ;
  assign n1155 = ( x73 & n1049 ) | ( x73 & ~n1099 ) | ( n1049 & ~n1099 ) ;
  assign n1156 = x73 & n1049 ;
  assign n1157 = ( ~n1054 & n1155 ) | ( ~n1054 & n1156 ) | ( n1155 & n1156 ) ;
  assign n1158 = ( n1054 & n1155 ) | ( n1054 & n1156 ) | ( n1155 & n1156 ) ;
  assign n1159 = ( n1054 & n1157 ) | ( n1054 & ~n1158 ) | ( n1157 & ~n1158 ) ;
  assign n1160 = ( x74 & n1154 ) | ( x74 & ~n1159 ) | ( n1154 & ~n1159 ) ;
  assign n1161 = ( x74 & n1055 ) | ( x74 & ~n1099 ) | ( n1055 & ~n1099 ) ;
  assign n1162 = x74 & n1055 ;
  assign n1163 = ( n1060 & n1161 ) | ( n1060 & n1162 ) | ( n1161 & n1162 ) ;
  assign n1164 = ( ~n1060 & n1161 ) | ( ~n1060 & n1162 ) | ( n1161 & n1162 ) ;
  assign n1165 = ( n1060 & ~n1163 ) | ( n1060 & n1164 ) | ( ~n1163 & n1164 ) ;
  assign n1166 = ( x75 & n1160 ) | ( x75 & ~n1165 ) | ( n1160 & ~n1165 ) ;
  assign n1167 = ( x75 & n1061 ) | ( x75 & ~n1099 ) | ( n1061 & ~n1099 ) ;
  assign n1168 = x75 & n1061 ;
  assign n1169 = ( ~n1066 & n1167 ) | ( ~n1066 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1170 = ( n1066 & n1167 ) | ( n1066 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1171 = ( n1066 & n1169 ) | ( n1066 & ~n1170 ) | ( n1169 & ~n1170 ) ;
  assign n1172 = ( x76 & n1166 ) | ( x76 & ~n1171 ) | ( n1166 & ~n1171 ) ;
  assign n1173 = ( x76 & n1067 ) | ( x76 & ~n1099 ) | ( n1067 & ~n1099 ) ;
  assign n1174 = x76 & n1067 ;
  assign n1175 = ( n1072 & n1173 ) | ( n1072 & n1174 ) | ( n1173 & n1174 ) ;
  assign n1176 = ( ~n1072 & n1173 ) | ( ~n1072 & n1174 ) | ( n1173 & n1174 ) ;
  assign n1177 = ( n1072 & ~n1175 ) | ( n1072 & n1176 ) | ( ~n1175 & n1176 ) ;
  assign n1178 = ( x77 & n1172 ) | ( x77 & ~n1177 ) | ( n1172 & ~n1177 ) ;
  assign n1179 = ( x77 & n1073 ) | ( x77 & ~n1099 ) | ( n1073 & ~n1099 ) ;
  assign n1180 = x77 & n1073 ;
  assign n1181 = ( ~n1078 & n1179 ) | ( ~n1078 & n1180 ) | ( n1179 & n1180 ) ;
  assign n1182 = ( n1078 & n1179 ) | ( n1078 & n1180 ) | ( n1179 & n1180 ) ;
  assign n1183 = ( n1078 & n1181 ) | ( n1078 & ~n1182 ) | ( n1181 & ~n1182 ) ;
  assign n1184 = ( x78 & n1178 ) | ( x78 & ~n1183 ) | ( n1178 & ~n1183 ) ;
  assign n1185 = ( x78 & n1079 ) | ( x78 & ~n1099 ) | ( n1079 & ~n1099 ) ;
  assign n1186 = x78 & n1079 ;
  assign n1187 = ( n1084 & n1185 ) | ( n1084 & n1186 ) | ( n1185 & n1186 ) ;
  assign n1188 = ( ~n1084 & n1185 ) | ( ~n1084 & n1186 ) | ( n1185 & n1186 ) ;
  assign n1189 = ( n1084 & ~n1187 ) | ( n1084 & n1188 ) | ( ~n1187 & n1188 ) ;
  assign n1190 = ( x79 & n1184 ) | ( x79 & ~n1189 ) | ( n1184 & ~n1189 ) ;
  assign n1191 = ( x79 & n1085 ) | ( x79 & ~n1099 ) | ( n1085 & ~n1099 ) ;
  assign n1192 = x79 & n1085 ;
  assign n1193 = ( ~n1090 & n1191 ) | ( ~n1090 & n1192 ) | ( n1191 & n1192 ) ;
  assign n1194 = ( n1090 & n1191 ) | ( n1090 & n1192 ) | ( n1191 & n1192 ) ;
  assign n1195 = ( n1090 & n1193 ) | ( n1090 & ~n1194 ) | ( n1193 & ~n1194 ) ;
  assign n1196 = ( x80 & n1190 ) | ( x80 & ~n1195 ) | ( n1190 & ~n1195 ) ;
  assign n1197 = ( x80 & n1091 ) | ( x80 & ~n1099 ) | ( n1091 & ~n1099 ) ;
  assign n1198 = x80 & n1091 ;
  assign n1199 = ( ~n1096 & n1197 ) | ( ~n1096 & n1198 ) | ( n1197 & n1198 ) ;
  assign n1200 = ( n1096 & n1197 ) | ( n1096 & n1198 ) | ( n1197 & n1198 ) ;
  assign n1201 = ( n1096 & n1199 ) | ( n1096 & ~n1200 ) | ( n1199 & ~n1200 ) ;
  assign n1202 = ( x81 & n1196 ) | ( x81 & ~n1201 ) | ( n1196 & ~n1201 ) ;
  assign n1203 = x82 | n1202 ;
  assign n1204 = ( x82 & n997 ) | ( x82 & n1202 ) | ( n997 & n1202 ) ;
  assign n1205 = ( n1101 & ~n1203 ) | ( n1101 & n1204 ) | ( ~n1203 & n1204 ) ;
  assign n1206 = ( x82 & ~n1101 ) | ( x82 & n1202 ) | ( ~n1101 & n1202 ) ;
  assign n1207 = n997 | n1206 ;
  assign n1208 = ( x45 & ~x64 ) | ( x45 & n1207 ) | ( ~x64 & n1207 ) ;
  assign n1209 = ~x45 & n1207 ;
  assign n1210 = ( n1105 & n1208 ) | ( n1105 & ~n1209 ) | ( n1208 & ~n1209 ) ;
  assign n1211 = ~x44 & x64 ;
  assign n1212 = ( x65 & ~n1210 ) | ( x65 & n1211 ) | ( ~n1210 & n1211 ) ;
  assign n1213 = ( x65 & n1105 ) | ( x65 & ~n1207 ) | ( n1105 & ~n1207 ) ;
  assign n1214 = x65 & n1105 ;
  assign n1215 = ( n1104 & n1213 ) | ( n1104 & n1214 ) | ( n1213 & n1214 ) ;
  assign n1216 = ( ~n1104 & n1213 ) | ( ~n1104 & n1214 ) | ( n1213 & n1214 ) ;
  assign n1217 = ( n1104 & ~n1215 ) | ( n1104 & n1216 ) | ( ~n1215 & n1216 ) ;
  assign n1218 = ( x66 & n1212 ) | ( x66 & ~n1217 ) | ( n1212 & ~n1217 ) ;
  assign n1219 = ( x66 & n1106 ) | ( x66 & ~n1207 ) | ( n1106 & ~n1207 ) ;
  assign n1220 = x66 & n1106 ;
  assign n1221 = ( n1111 & n1219 ) | ( n1111 & n1220 ) | ( n1219 & n1220 ) ;
  assign n1222 = ( ~n1111 & n1219 ) | ( ~n1111 & n1220 ) | ( n1219 & n1220 ) ;
  assign n1223 = ( n1111 & ~n1221 ) | ( n1111 & n1222 ) | ( ~n1221 & n1222 ) ;
  assign n1224 = ( x67 & n1218 ) | ( x67 & ~n1223 ) | ( n1218 & ~n1223 ) ;
  assign n1225 = ( x67 & n1112 ) | ( x67 & ~n1207 ) | ( n1112 & ~n1207 ) ;
  assign n1226 = x67 & n1112 ;
  assign n1227 = ( ~n1117 & n1225 ) | ( ~n1117 & n1226 ) | ( n1225 & n1226 ) ;
  assign n1228 = ( n1117 & n1225 ) | ( n1117 & n1226 ) | ( n1225 & n1226 ) ;
  assign n1229 = ( n1117 & n1227 ) | ( n1117 & ~n1228 ) | ( n1227 & ~n1228 ) ;
  assign n1230 = ( x68 & n1224 ) | ( x68 & ~n1229 ) | ( n1224 & ~n1229 ) ;
  assign n1231 = ( x68 & n1118 ) | ( x68 & ~n1207 ) | ( n1118 & ~n1207 ) ;
  assign n1232 = x68 & n1118 ;
  assign n1233 = ( n1123 & n1231 ) | ( n1123 & n1232 ) | ( n1231 & n1232 ) ;
  assign n1234 = ( ~n1123 & n1231 ) | ( ~n1123 & n1232 ) | ( n1231 & n1232 ) ;
  assign n1235 = ( n1123 & ~n1233 ) | ( n1123 & n1234 ) | ( ~n1233 & n1234 ) ;
  assign n1236 = ( x69 & n1230 ) | ( x69 & ~n1235 ) | ( n1230 & ~n1235 ) ;
  assign n1237 = ( x69 & n1124 ) | ( x69 & ~n1207 ) | ( n1124 & ~n1207 ) ;
  assign n1238 = x69 & n1124 ;
  assign n1239 = ( ~n1129 & n1237 ) | ( ~n1129 & n1238 ) | ( n1237 & n1238 ) ;
  assign n1240 = ( n1129 & n1237 ) | ( n1129 & n1238 ) | ( n1237 & n1238 ) ;
  assign n1241 = ( n1129 & n1239 ) | ( n1129 & ~n1240 ) | ( n1239 & ~n1240 ) ;
  assign n1242 = ( x70 & n1236 ) | ( x70 & ~n1241 ) | ( n1236 & ~n1241 ) ;
  assign n1243 = ( x70 & n1130 ) | ( x70 & ~n1207 ) | ( n1130 & ~n1207 ) ;
  assign n1244 = x70 & n1130 ;
  assign n1245 = ( n1135 & n1243 ) | ( n1135 & n1244 ) | ( n1243 & n1244 ) ;
  assign n1246 = ( ~n1135 & n1243 ) | ( ~n1135 & n1244 ) | ( n1243 & n1244 ) ;
  assign n1247 = ( n1135 & ~n1245 ) | ( n1135 & n1246 ) | ( ~n1245 & n1246 ) ;
  assign n1248 = ( x71 & n1242 ) | ( x71 & ~n1247 ) | ( n1242 & ~n1247 ) ;
  assign n1249 = ( x71 & n1136 ) | ( x71 & ~n1207 ) | ( n1136 & ~n1207 ) ;
  assign n1250 = x71 & n1136 ;
  assign n1251 = ( ~n1141 & n1249 ) | ( ~n1141 & n1250 ) | ( n1249 & n1250 ) ;
  assign n1252 = ( n1141 & n1249 ) | ( n1141 & n1250 ) | ( n1249 & n1250 ) ;
  assign n1253 = ( n1141 & n1251 ) | ( n1141 & ~n1252 ) | ( n1251 & ~n1252 ) ;
  assign n1254 = ( x72 & n1248 ) | ( x72 & ~n1253 ) | ( n1248 & ~n1253 ) ;
  assign n1255 = ( x72 & n1142 ) | ( x72 & ~n1207 ) | ( n1142 & ~n1207 ) ;
  assign n1256 = x72 & n1142 ;
  assign n1257 = ( n1147 & n1255 ) | ( n1147 & n1256 ) | ( n1255 & n1256 ) ;
  assign n1258 = ( ~n1147 & n1255 ) | ( ~n1147 & n1256 ) | ( n1255 & n1256 ) ;
  assign n1259 = ( n1147 & ~n1257 ) | ( n1147 & n1258 ) | ( ~n1257 & n1258 ) ;
  assign n1260 = ( x73 & n1254 ) | ( x73 & ~n1259 ) | ( n1254 & ~n1259 ) ;
  assign n1261 = ( x73 & n1148 ) | ( x73 & ~n1207 ) | ( n1148 & ~n1207 ) ;
  assign n1262 = x73 & n1148 ;
  assign n1263 = ( ~n1153 & n1261 ) | ( ~n1153 & n1262 ) | ( n1261 & n1262 ) ;
  assign n1264 = ( n1153 & n1261 ) | ( n1153 & n1262 ) | ( n1261 & n1262 ) ;
  assign n1265 = ( n1153 & n1263 ) | ( n1153 & ~n1264 ) | ( n1263 & ~n1264 ) ;
  assign n1266 = ( x74 & n1260 ) | ( x74 & ~n1265 ) | ( n1260 & ~n1265 ) ;
  assign n1267 = ( x74 & n1154 ) | ( x74 & ~n1207 ) | ( n1154 & ~n1207 ) ;
  assign n1268 = x74 & n1154 ;
  assign n1269 = ( n1159 & n1267 ) | ( n1159 & n1268 ) | ( n1267 & n1268 ) ;
  assign n1270 = ( ~n1159 & n1267 ) | ( ~n1159 & n1268 ) | ( n1267 & n1268 ) ;
  assign n1271 = ( n1159 & ~n1269 ) | ( n1159 & n1270 ) | ( ~n1269 & n1270 ) ;
  assign n1272 = ( x75 & n1266 ) | ( x75 & ~n1271 ) | ( n1266 & ~n1271 ) ;
  assign n1273 = ( x75 & n1160 ) | ( x75 & ~n1207 ) | ( n1160 & ~n1207 ) ;
  assign n1274 = x75 & n1160 ;
  assign n1275 = ( ~n1165 & n1273 ) | ( ~n1165 & n1274 ) | ( n1273 & n1274 ) ;
  assign n1276 = ( n1165 & n1273 ) | ( n1165 & n1274 ) | ( n1273 & n1274 ) ;
  assign n1277 = ( n1165 & n1275 ) | ( n1165 & ~n1276 ) | ( n1275 & ~n1276 ) ;
  assign n1278 = ( x76 & n1272 ) | ( x76 & ~n1277 ) | ( n1272 & ~n1277 ) ;
  assign n1279 = ( x76 & n1166 ) | ( x76 & ~n1207 ) | ( n1166 & ~n1207 ) ;
  assign n1280 = x76 & n1166 ;
  assign n1281 = ( n1171 & n1279 ) | ( n1171 & n1280 ) | ( n1279 & n1280 ) ;
  assign n1282 = ( ~n1171 & n1279 ) | ( ~n1171 & n1280 ) | ( n1279 & n1280 ) ;
  assign n1283 = ( n1171 & ~n1281 ) | ( n1171 & n1282 ) | ( ~n1281 & n1282 ) ;
  assign n1284 = ( x77 & n1278 ) | ( x77 & ~n1283 ) | ( n1278 & ~n1283 ) ;
  assign n1285 = ( x77 & n1172 ) | ( x77 & ~n1207 ) | ( n1172 & ~n1207 ) ;
  assign n1286 = x77 & n1172 ;
  assign n1287 = ( ~n1177 & n1285 ) | ( ~n1177 & n1286 ) | ( n1285 & n1286 ) ;
  assign n1288 = ( n1177 & n1285 ) | ( n1177 & n1286 ) | ( n1285 & n1286 ) ;
  assign n1289 = ( n1177 & n1287 ) | ( n1177 & ~n1288 ) | ( n1287 & ~n1288 ) ;
  assign n1290 = ( x78 & n1284 ) | ( x78 & ~n1289 ) | ( n1284 & ~n1289 ) ;
  assign n1291 = ( x78 & n1178 ) | ( x78 & ~n1207 ) | ( n1178 & ~n1207 ) ;
  assign n1292 = x78 & n1178 ;
  assign n1293 = ( n1183 & n1291 ) | ( n1183 & n1292 ) | ( n1291 & n1292 ) ;
  assign n1294 = ( ~n1183 & n1291 ) | ( ~n1183 & n1292 ) | ( n1291 & n1292 ) ;
  assign n1295 = ( n1183 & ~n1293 ) | ( n1183 & n1294 ) | ( ~n1293 & n1294 ) ;
  assign n1296 = ( x79 & n1290 ) | ( x79 & ~n1295 ) | ( n1290 & ~n1295 ) ;
  assign n1297 = ( x79 & n1184 ) | ( x79 & ~n1207 ) | ( n1184 & ~n1207 ) ;
  assign n1298 = x79 & n1184 ;
  assign n1299 = ( ~n1189 & n1297 ) | ( ~n1189 & n1298 ) | ( n1297 & n1298 ) ;
  assign n1300 = ( n1189 & n1297 ) | ( n1189 & n1298 ) | ( n1297 & n1298 ) ;
  assign n1301 = ( n1189 & n1299 ) | ( n1189 & ~n1300 ) | ( n1299 & ~n1300 ) ;
  assign n1302 = ( x80 & n1296 ) | ( x80 & ~n1301 ) | ( n1296 & ~n1301 ) ;
  assign n1303 = ( x80 & n1190 ) | ( x80 & ~n1207 ) | ( n1190 & ~n1207 ) ;
  assign n1304 = x80 & n1190 ;
  assign n1305 = ( n1195 & n1303 ) | ( n1195 & n1304 ) | ( n1303 & n1304 ) ;
  assign n1306 = ( ~n1195 & n1303 ) | ( ~n1195 & n1304 ) | ( n1303 & n1304 ) ;
  assign n1307 = ( n1195 & ~n1305 ) | ( n1195 & n1306 ) | ( ~n1305 & n1306 ) ;
  assign n1308 = ( x81 & n1302 ) | ( x81 & ~n1307 ) | ( n1302 & ~n1307 ) ;
  assign n1309 = ( x81 & n1196 ) | ( x81 & ~n1207 ) | ( n1196 & ~n1207 ) ;
  assign n1310 = x81 & n1196 ;
  assign n1311 = ( n1201 & n1309 ) | ( n1201 & n1310 ) | ( n1309 & n1310 ) ;
  assign n1312 = ( ~n1201 & n1309 ) | ( ~n1201 & n1310 ) | ( n1309 & n1310 ) ;
  assign n1313 = ( n1201 & ~n1311 ) | ( n1201 & n1312 ) | ( ~n1311 & n1312 ) ;
  assign n1314 = ( x82 & n1308 ) | ( x82 & ~n1313 ) | ( n1308 & ~n1313 ) ;
  assign n1315 = x83 & n1314 ;
  assign n1316 = ( x83 & ~n174 ) | ( x83 & n1314 ) | ( ~n174 & n1314 ) ;
  assign n1317 = ( n1205 & n1315 ) | ( n1205 & ~n1316 ) | ( n1315 & ~n1316 ) ;
  assign n1318 = ( x83 & ~n1205 ) | ( x83 & n1314 ) | ( ~n1205 & n1314 ) ;
  assign n1319 = n174 | n1318 ;
  assign n1320 = ( x44 & ~x64 ) | ( x44 & n1319 ) | ( ~x64 & n1319 ) ;
  assign n1321 = ~x44 & n1319 ;
  assign n1322 = ( n1211 & n1320 ) | ( n1211 & ~n1321 ) | ( n1320 & ~n1321 ) ;
  assign n1323 = ~x43 & x64 ;
  assign n1324 = ( x65 & ~n1322 ) | ( x65 & n1323 ) | ( ~n1322 & n1323 ) ;
  assign n1325 = ( x65 & n1211 ) | ( x65 & ~n1319 ) | ( n1211 & ~n1319 ) ;
  assign n1326 = x65 & n1211 ;
  assign n1327 = ( n1210 & n1325 ) | ( n1210 & n1326 ) | ( n1325 & n1326 ) ;
  assign n1328 = ( ~n1210 & n1325 ) | ( ~n1210 & n1326 ) | ( n1325 & n1326 ) ;
  assign n1329 = ( n1210 & ~n1327 ) | ( n1210 & n1328 ) | ( ~n1327 & n1328 ) ;
  assign n1330 = ( x66 & n1324 ) | ( x66 & ~n1329 ) | ( n1324 & ~n1329 ) ;
  assign n1331 = ( x66 & n1212 ) | ( x66 & ~n1319 ) | ( n1212 & ~n1319 ) ;
  assign n1332 = x66 & n1212 ;
  assign n1333 = ( n1217 & n1331 ) | ( n1217 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1334 = ( ~n1217 & n1331 ) | ( ~n1217 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1335 = ( n1217 & ~n1333 ) | ( n1217 & n1334 ) | ( ~n1333 & n1334 ) ;
  assign n1336 = ( x67 & n1330 ) | ( x67 & ~n1335 ) | ( n1330 & ~n1335 ) ;
  assign n1337 = ( x67 & n1218 ) | ( x67 & ~n1319 ) | ( n1218 & ~n1319 ) ;
  assign n1338 = x67 & n1218 ;
  assign n1339 = ( ~n1223 & n1337 ) | ( ~n1223 & n1338 ) | ( n1337 & n1338 ) ;
  assign n1340 = ( n1223 & n1337 ) | ( n1223 & n1338 ) | ( n1337 & n1338 ) ;
  assign n1341 = ( n1223 & n1339 ) | ( n1223 & ~n1340 ) | ( n1339 & ~n1340 ) ;
  assign n1342 = ( x68 & n1336 ) | ( x68 & ~n1341 ) | ( n1336 & ~n1341 ) ;
  assign n1343 = ( x68 & n1224 ) | ( x68 & ~n1319 ) | ( n1224 & ~n1319 ) ;
  assign n1344 = x68 & n1224 ;
  assign n1345 = ( n1229 & n1343 ) | ( n1229 & n1344 ) | ( n1343 & n1344 ) ;
  assign n1346 = ( ~n1229 & n1343 ) | ( ~n1229 & n1344 ) | ( n1343 & n1344 ) ;
  assign n1347 = ( n1229 & ~n1345 ) | ( n1229 & n1346 ) | ( ~n1345 & n1346 ) ;
  assign n1348 = ( x69 & n1342 ) | ( x69 & ~n1347 ) | ( n1342 & ~n1347 ) ;
  assign n1349 = ( x69 & n1230 ) | ( x69 & ~n1319 ) | ( n1230 & ~n1319 ) ;
  assign n1350 = x69 & n1230 ;
  assign n1351 = ( ~n1235 & n1349 ) | ( ~n1235 & n1350 ) | ( n1349 & n1350 ) ;
  assign n1352 = ( n1235 & n1349 ) | ( n1235 & n1350 ) | ( n1349 & n1350 ) ;
  assign n1353 = ( n1235 & n1351 ) | ( n1235 & ~n1352 ) | ( n1351 & ~n1352 ) ;
  assign n1354 = ( x70 & n1348 ) | ( x70 & ~n1353 ) | ( n1348 & ~n1353 ) ;
  assign n1355 = ( x70 & n1236 ) | ( x70 & ~n1319 ) | ( n1236 & ~n1319 ) ;
  assign n1356 = x70 & n1236 ;
  assign n1357 = ( n1241 & n1355 ) | ( n1241 & n1356 ) | ( n1355 & n1356 ) ;
  assign n1358 = ( ~n1241 & n1355 ) | ( ~n1241 & n1356 ) | ( n1355 & n1356 ) ;
  assign n1359 = ( n1241 & ~n1357 ) | ( n1241 & n1358 ) | ( ~n1357 & n1358 ) ;
  assign n1360 = ( x71 & n1354 ) | ( x71 & ~n1359 ) | ( n1354 & ~n1359 ) ;
  assign n1361 = ( x71 & n1242 ) | ( x71 & ~n1319 ) | ( n1242 & ~n1319 ) ;
  assign n1362 = x71 & n1242 ;
  assign n1363 = ( ~n1247 & n1361 ) | ( ~n1247 & n1362 ) | ( n1361 & n1362 ) ;
  assign n1364 = ( n1247 & n1361 ) | ( n1247 & n1362 ) | ( n1361 & n1362 ) ;
  assign n1365 = ( n1247 & n1363 ) | ( n1247 & ~n1364 ) | ( n1363 & ~n1364 ) ;
  assign n1366 = ( x72 & n1360 ) | ( x72 & ~n1365 ) | ( n1360 & ~n1365 ) ;
  assign n1367 = ( x72 & n1248 ) | ( x72 & ~n1319 ) | ( n1248 & ~n1319 ) ;
  assign n1368 = x72 & n1248 ;
  assign n1369 = ( n1253 & n1367 ) | ( n1253 & n1368 ) | ( n1367 & n1368 ) ;
  assign n1370 = ( ~n1253 & n1367 ) | ( ~n1253 & n1368 ) | ( n1367 & n1368 ) ;
  assign n1371 = ( n1253 & ~n1369 ) | ( n1253 & n1370 ) | ( ~n1369 & n1370 ) ;
  assign n1372 = ( x73 & n1366 ) | ( x73 & ~n1371 ) | ( n1366 & ~n1371 ) ;
  assign n1373 = ( x73 & n1254 ) | ( x73 & ~n1319 ) | ( n1254 & ~n1319 ) ;
  assign n1374 = x73 & n1254 ;
  assign n1375 = ( ~n1259 & n1373 ) | ( ~n1259 & n1374 ) | ( n1373 & n1374 ) ;
  assign n1376 = ( n1259 & n1373 ) | ( n1259 & n1374 ) | ( n1373 & n1374 ) ;
  assign n1377 = ( n1259 & n1375 ) | ( n1259 & ~n1376 ) | ( n1375 & ~n1376 ) ;
  assign n1378 = ( x74 & n1372 ) | ( x74 & ~n1377 ) | ( n1372 & ~n1377 ) ;
  assign n1379 = ( x74 & n1260 ) | ( x74 & ~n1319 ) | ( n1260 & ~n1319 ) ;
  assign n1380 = x74 & n1260 ;
  assign n1381 = ( n1265 & n1379 ) | ( n1265 & n1380 ) | ( n1379 & n1380 ) ;
  assign n1382 = ( ~n1265 & n1379 ) | ( ~n1265 & n1380 ) | ( n1379 & n1380 ) ;
  assign n1383 = ( n1265 & ~n1381 ) | ( n1265 & n1382 ) | ( ~n1381 & n1382 ) ;
  assign n1384 = ( x75 & n1378 ) | ( x75 & ~n1383 ) | ( n1378 & ~n1383 ) ;
  assign n1385 = ( x75 & n1266 ) | ( x75 & ~n1319 ) | ( n1266 & ~n1319 ) ;
  assign n1386 = x75 & n1266 ;
  assign n1387 = ( ~n1271 & n1385 ) | ( ~n1271 & n1386 ) | ( n1385 & n1386 ) ;
  assign n1388 = ( n1271 & n1385 ) | ( n1271 & n1386 ) | ( n1385 & n1386 ) ;
  assign n1389 = ( n1271 & n1387 ) | ( n1271 & ~n1388 ) | ( n1387 & ~n1388 ) ;
  assign n1390 = ( x76 & n1384 ) | ( x76 & ~n1389 ) | ( n1384 & ~n1389 ) ;
  assign n1391 = ( x76 & n1272 ) | ( x76 & ~n1319 ) | ( n1272 & ~n1319 ) ;
  assign n1392 = x76 & n1272 ;
  assign n1393 = ( n1277 & n1391 ) | ( n1277 & n1392 ) | ( n1391 & n1392 ) ;
  assign n1394 = ( ~n1277 & n1391 ) | ( ~n1277 & n1392 ) | ( n1391 & n1392 ) ;
  assign n1395 = ( n1277 & ~n1393 ) | ( n1277 & n1394 ) | ( ~n1393 & n1394 ) ;
  assign n1396 = ( x77 & n1390 ) | ( x77 & ~n1395 ) | ( n1390 & ~n1395 ) ;
  assign n1397 = ( x77 & n1278 ) | ( x77 & ~n1319 ) | ( n1278 & ~n1319 ) ;
  assign n1398 = x77 & n1278 ;
  assign n1399 = ( ~n1283 & n1397 ) | ( ~n1283 & n1398 ) | ( n1397 & n1398 ) ;
  assign n1400 = ( n1283 & n1397 ) | ( n1283 & n1398 ) | ( n1397 & n1398 ) ;
  assign n1401 = ( n1283 & n1399 ) | ( n1283 & ~n1400 ) | ( n1399 & ~n1400 ) ;
  assign n1402 = ( x78 & n1396 ) | ( x78 & ~n1401 ) | ( n1396 & ~n1401 ) ;
  assign n1403 = ( x78 & n1284 ) | ( x78 & ~n1319 ) | ( n1284 & ~n1319 ) ;
  assign n1404 = x78 & n1284 ;
  assign n1405 = ( n1289 & n1403 ) | ( n1289 & n1404 ) | ( n1403 & n1404 ) ;
  assign n1406 = ( ~n1289 & n1403 ) | ( ~n1289 & n1404 ) | ( n1403 & n1404 ) ;
  assign n1407 = ( n1289 & ~n1405 ) | ( n1289 & n1406 ) | ( ~n1405 & n1406 ) ;
  assign n1408 = ( x79 & n1402 ) | ( x79 & ~n1407 ) | ( n1402 & ~n1407 ) ;
  assign n1409 = ( x79 & n1290 ) | ( x79 & ~n1319 ) | ( n1290 & ~n1319 ) ;
  assign n1410 = x79 & n1290 ;
  assign n1411 = ( ~n1295 & n1409 ) | ( ~n1295 & n1410 ) | ( n1409 & n1410 ) ;
  assign n1412 = ( n1295 & n1409 ) | ( n1295 & n1410 ) | ( n1409 & n1410 ) ;
  assign n1413 = ( n1295 & n1411 ) | ( n1295 & ~n1412 ) | ( n1411 & ~n1412 ) ;
  assign n1414 = ( x80 & n1408 ) | ( x80 & ~n1413 ) | ( n1408 & ~n1413 ) ;
  assign n1415 = ( x80 & n1296 ) | ( x80 & ~n1319 ) | ( n1296 & ~n1319 ) ;
  assign n1416 = x80 & n1296 ;
  assign n1417 = ( n1301 & n1415 ) | ( n1301 & n1416 ) | ( n1415 & n1416 ) ;
  assign n1418 = ( ~n1301 & n1415 ) | ( ~n1301 & n1416 ) | ( n1415 & n1416 ) ;
  assign n1419 = ( n1301 & ~n1417 ) | ( n1301 & n1418 ) | ( ~n1417 & n1418 ) ;
  assign n1420 = ( x81 & n1414 ) | ( x81 & ~n1419 ) | ( n1414 & ~n1419 ) ;
  assign n1421 = ( x81 & n1302 ) | ( x81 & ~n1319 ) | ( n1302 & ~n1319 ) ;
  assign n1422 = x81 & n1302 ;
  assign n1423 = ( ~n1307 & n1421 ) | ( ~n1307 & n1422 ) | ( n1421 & n1422 ) ;
  assign n1424 = ( n1307 & n1421 ) | ( n1307 & n1422 ) | ( n1421 & n1422 ) ;
  assign n1425 = ( n1307 & n1423 ) | ( n1307 & ~n1424 ) | ( n1423 & ~n1424 ) ;
  assign n1426 = ( x82 & n1420 ) | ( x82 & ~n1425 ) | ( n1420 & ~n1425 ) ;
  assign n1427 = ( x82 & n1308 ) | ( x82 & ~n1319 ) | ( n1308 & ~n1319 ) ;
  assign n1428 = x82 & n1308 ;
  assign n1429 = ( ~n1313 & n1427 ) | ( ~n1313 & n1428 ) | ( n1427 & n1428 ) ;
  assign n1430 = ( n1313 & n1427 ) | ( n1313 & n1428 ) | ( n1427 & n1428 ) ;
  assign n1431 = ( n1313 & n1429 ) | ( n1313 & ~n1430 ) | ( n1429 & ~n1430 ) ;
  assign n1432 = ( x83 & n1426 ) | ( x83 & ~n1431 ) | ( n1426 & ~n1431 ) ;
  assign n1433 = ( n174 & ~n1317 ) | ( n174 & n1432 ) | ( ~n1317 & n1432 ) ;
  assign n1434 = x85 | n172 ;
  assign n1435 = n1433 | n1434 ;
  assign n1436 = n1317 & n1435 ;
  assign n1437 = n280 | n1436 ;
  assign n1438 = ( x43 & ~x64 ) | ( x43 & n1435 ) | ( ~x64 & n1435 ) ;
  assign n1439 = ~x43 & n1435 ;
  assign n1440 = ( n1323 & n1438 ) | ( n1323 & ~n1439 ) | ( n1438 & ~n1439 ) ;
  assign n1441 = ~x42 & x64 ;
  assign n1442 = ( x65 & ~n1440 ) | ( x65 & n1441 ) | ( ~n1440 & n1441 ) ;
  assign n1443 = ( x65 & n1323 ) | ( x65 & ~n1435 ) | ( n1323 & ~n1435 ) ;
  assign n1444 = x65 & n1323 ;
  assign n1445 = ( n1322 & n1443 ) | ( n1322 & n1444 ) | ( n1443 & n1444 ) ;
  assign n1446 = ( ~n1322 & n1443 ) | ( ~n1322 & n1444 ) | ( n1443 & n1444 ) ;
  assign n1447 = ( n1322 & ~n1445 ) | ( n1322 & n1446 ) | ( ~n1445 & n1446 ) ;
  assign n1448 = ( x66 & n1442 ) | ( x66 & ~n1447 ) | ( n1442 & ~n1447 ) ;
  assign n1449 = ( x66 & n1324 ) | ( x66 & ~n1435 ) | ( n1324 & ~n1435 ) ;
  assign n1450 = x66 & n1324 ;
  assign n1451 = ( n1329 & n1449 ) | ( n1329 & n1450 ) | ( n1449 & n1450 ) ;
  assign n1452 = ( ~n1329 & n1449 ) | ( ~n1329 & n1450 ) | ( n1449 & n1450 ) ;
  assign n1453 = ( n1329 & ~n1451 ) | ( n1329 & n1452 ) | ( ~n1451 & n1452 ) ;
  assign n1454 = ( x67 & n1448 ) | ( x67 & ~n1453 ) | ( n1448 & ~n1453 ) ;
  assign n1455 = ( x67 & n1330 ) | ( x67 & ~n1435 ) | ( n1330 & ~n1435 ) ;
  assign n1456 = x67 & n1330 ;
  assign n1457 = ( ~n1335 & n1455 ) | ( ~n1335 & n1456 ) | ( n1455 & n1456 ) ;
  assign n1458 = ( n1335 & n1455 ) | ( n1335 & n1456 ) | ( n1455 & n1456 ) ;
  assign n1459 = ( n1335 & n1457 ) | ( n1335 & ~n1458 ) | ( n1457 & ~n1458 ) ;
  assign n1460 = ( x68 & n1454 ) | ( x68 & ~n1459 ) | ( n1454 & ~n1459 ) ;
  assign n1461 = ( x68 & n1336 ) | ( x68 & ~n1435 ) | ( n1336 & ~n1435 ) ;
  assign n1462 = x68 & n1336 ;
  assign n1463 = ( n1341 & n1461 ) | ( n1341 & n1462 ) | ( n1461 & n1462 ) ;
  assign n1464 = ( ~n1341 & n1461 ) | ( ~n1341 & n1462 ) | ( n1461 & n1462 ) ;
  assign n1465 = ( n1341 & ~n1463 ) | ( n1341 & n1464 ) | ( ~n1463 & n1464 ) ;
  assign n1466 = ( x69 & n1460 ) | ( x69 & ~n1465 ) | ( n1460 & ~n1465 ) ;
  assign n1467 = ( x69 & n1342 ) | ( x69 & ~n1435 ) | ( n1342 & ~n1435 ) ;
  assign n1468 = x69 & n1342 ;
  assign n1469 = ( ~n1347 & n1467 ) | ( ~n1347 & n1468 ) | ( n1467 & n1468 ) ;
  assign n1470 = ( n1347 & n1467 ) | ( n1347 & n1468 ) | ( n1467 & n1468 ) ;
  assign n1471 = ( n1347 & n1469 ) | ( n1347 & ~n1470 ) | ( n1469 & ~n1470 ) ;
  assign n1472 = ( x70 & n1466 ) | ( x70 & ~n1471 ) | ( n1466 & ~n1471 ) ;
  assign n1473 = ( x70 & n1348 ) | ( x70 & ~n1435 ) | ( n1348 & ~n1435 ) ;
  assign n1474 = x70 & n1348 ;
  assign n1475 = ( n1353 & n1473 ) | ( n1353 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1476 = ( ~n1353 & n1473 ) | ( ~n1353 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1477 = ( n1353 & ~n1475 ) | ( n1353 & n1476 ) | ( ~n1475 & n1476 ) ;
  assign n1478 = ( x71 & n1472 ) | ( x71 & ~n1477 ) | ( n1472 & ~n1477 ) ;
  assign n1479 = ( x71 & n1354 ) | ( x71 & ~n1435 ) | ( n1354 & ~n1435 ) ;
  assign n1480 = x71 & n1354 ;
  assign n1481 = ( ~n1359 & n1479 ) | ( ~n1359 & n1480 ) | ( n1479 & n1480 ) ;
  assign n1482 = ( n1359 & n1479 ) | ( n1359 & n1480 ) | ( n1479 & n1480 ) ;
  assign n1483 = ( n1359 & n1481 ) | ( n1359 & ~n1482 ) | ( n1481 & ~n1482 ) ;
  assign n1484 = ( x72 & n1478 ) | ( x72 & ~n1483 ) | ( n1478 & ~n1483 ) ;
  assign n1485 = ( x72 & n1360 ) | ( x72 & ~n1435 ) | ( n1360 & ~n1435 ) ;
  assign n1486 = x72 & n1360 ;
  assign n1487 = ( n1365 & n1485 ) | ( n1365 & n1486 ) | ( n1485 & n1486 ) ;
  assign n1488 = ( ~n1365 & n1485 ) | ( ~n1365 & n1486 ) | ( n1485 & n1486 ) ;
  assign n1489 = ( n1365 & ~n1487 ) | ( n1365 & n1488 ) | ( ~n1487 & n1488 ) ;
  assign n1490 = ( x73 & n1484 ) | ( x73 & ~n1489 ) | ( n1484 & ~n1489 ) ;
  assign n1491 = ( x73 & n1366 ) | ( x73 & ~n1435 ) | ( n1366 & ~n1435 ) ;
  assign n1492 = x73 & n1366 ;
  assign n1493 = ( ~n1371 & n1491 ) | ( ~n1371 & n1492 ) | ( n1491 & n1492 ) ;
  assign n1494 = ( n1371 & n1491 ) | ( n1371 & n1492 ) | ( n1491 & n1492 ) ;
  assign n1495 = ( n1371 & n1493 ) | ( n1371 & ~n1494 ) | ( n1493 & ~n1494 ) ;
  assign n1496 = ( x74 & n1490 ) | ( x74 & ~n1495 ) | ( n1490 & ~n1495 ) ;
  assign n1497 = ( x74 & n1372 ) | ( x74 & ~n1435 ) | ( n1372 & ~n1435 ) ;
  assign n1498 = x74 & n1372 ;
  assign n1499 = ( n1377 & n1497 ) | ( n1377 & n1498 ) | ( n1497 & n1498 ) ;
  assign n1500 = ( ~n1377 & n1497 ) | ( ~n1377 & n1498 ) | ( n1497 & n1498 ) ;
  assign n1501 = ( n1377 & ~n1499 ) | ( n1377 & n1500 ) | ( ~n1499 & n1500 ) ;
  assign n1502 = ( x75 & n1496 ) | ( x75 & ~n1501 ) | ( n1496 & ~n1501 ) ;
  assign n1503 = ( x75 & n1378 ) | ( x75 & ~n1435 ) | ( n1378 & ~n1435 ) ;
  assign n1504 = x75 & n1378 ;
  assign n1505 = ( ~n1383 & n1503 ) | ( ~n1383 & n1504 ) | ( n1503 & n1504 ) ;
  assign n1506 = ( n1383 & n1503 ) | ( n1383 & n1504 ) | ( n1503 & n1504 ) ;
  assign n1507 = ( n1383 & n1505 ) | ( n1383 & ~n1506 ) | ( n1505 & ~n1506 ) ;
  assign n1508 = ( x76 & n1502 ) | ( x76 & ~n1507 ) | ( n1502 & ~n1507 ) ;
  assign n1509 = ( x76 & n1384 ) | ( x76 & ~n1435 ) | ( n1384 & ~n1435 ) ;
  assign n1510 = x76 & n1384 ;
  assign n1511 = ( n1389 & n1509 ) | ( n1389 & n1510 ) | ( n1509 & n1510 ) ;
  assign n1512 = ( ~n1389 & n1509 ) | ( ~n1389 & n1510 ) | ( n1509 & n1510 ) ;
  assign n1513 = ( n1389 & ~n1511 ) | ( n1389 & n1512 ) | ( ~n1511 & n1512 ) ;
  assign n1514 = ( x77 & n1508 ) | ( x77 & ~n1513 ) | ( n1508 & ~n1513 ) ;
  assign n1515 = ( x77 & n1390 ) | ( x77 & ~n1435 ) | ( n1390 & ~n1435 ) ;
  assign n1516 = x77 & n1390 ;
  assign n1517 = ( ~n1395 & n1515 ) | ( ~n1395 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1518 = ( n1395 & n1515 ) | ( n1395 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1519 = ( n1395 & n1517 ) | ( n1395 & ~n1518 ) | ( n1517 & ~n1518 ) ;
  assign n1520 = ( x78 & n1514 ) | ( x78 & ~n1519 ) | ( n1514 & ~n1519 ) ;
  assign n1521 = ( x78 & n1396 ) | ( x78 & ~n1435 ) | ( n1396 & ~n1435 ) ;
  assign n1522 = x78 & n1396 ;
  assign n1523 = ( n1401 & n1521 ) | ( n1401 & n1522 ) | ( n1521 & n1522 ) ;
  assign n1524 = ( ~n1401 & n1521 ) | ( ~n1401 & n1522 ) | ( n1521 & n1522 ) ;
  assign n1525 = ( n1401 & ~n1523 ) | ( n1401 & n1524 ) | ( ~n1523 & n1524 ) ;
  assign n1526 = ( x79 & n1520 ) | ( x79 & ~n1525 ) | ( n1520 & ~n1525 ) ;
  assign n1527 = ( x79 & n1402 ) | ( x79 & ~n1435 ) | ( n1402 & ~n1435 ) ;
  assign n1528 = x79 & n1402 ;
  assign n1529 = ( ~n1407 & n1527 ) | ( ~n1407 & n1528 ) | ( n1527 & n1528 ) ;
  assign n1530 = ( n1407 & n1527 ) | ( n1407 & n1528 ) | ( n1527 & n1528 ) ;
  assign n1531 = ( n1407 & n1529 ) | ( n1407 & ~n1530 ) | ( n1529 & ~n1530 ) ;
  assign n1532 = ( x80 & n1526 ) | ( x80 & ~n1531 ) | ( n1526 & ~n1531 ) ;
  assign n1533 = ( x80 & n1408 ) | ( x80 & ~n1435 ) | ( n1408 & ~n1435 ) ;
  assign n1534 = x80 & n1408 ;
  assign n1535 = ( n1413 & n1533 ) | ( n1413 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1536 = ( ~n1413 & n1533 ) | ( ~n1413 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1537 = ( n1413 & ~n1535 ) | ( n1413 & n1536 ) | ( ~n1535 & n1536 ) ;
  assign n1538 = ( x81 & n1532 ) | ( x81 & ~n1537 ) | ( n1532 & ~n1537 ) ;
  assign n1539 = ( x81 & n1414 ) | ( x81 & ~n1435 ) | ( n1414 & ~n1435 ) ;
  assign n1540 = x81 & n1414 ;
  assign n1541 = ( ~n1419 & n1539 ) | ( ~n1419 & n1540 ) | ( n1539 & n1540 ) ;
  assign n1542 = ( n1419 & n1539 ) | ( n1419 & n1540 ) | ( n1539 & n1540 ) ;
  assign n1543 = ( n1419 & n1541 ) | ( n1419 & ~n1542 ) | ( n1541 & ~n1542 ) ;
  assign n1544 = ( x82 & n1538 ) | ( x82 & ~n1543 ) | ( n1538 & ~n1543 ) ;
  assign n1545 = ( x82 & n1420 ) | ( x82 & ~n1435 ) | ( n1420 & ~n1435 ) ;
  assign n1546 = x82 & n1420 ;
  assign n1547 = ( n1425 & n1545 ) | ( n1425 & n1546 ) | ( n1545 & n1546 ) ;
  assign n1548 = ( ~n1425 & n1545 ) | ( ~n1425 & n1546 ) | ( n1545 & n1546 ) ;
  assign n1549 = ( n1425 & ~n1547 ) | ( n1425 & n1548 ) | ( ~n1547 & n1548 ) ;
  assign n1550 = ( x83 & n1544 ) | ( x83 & ~n1549 ) | ( n1544 & ~n1549 ) ;
  assign n1551 = ( x83 & n1426 ) | ( x83 & ~n1435 ) | ( n1426 & ~n1435 ) ;
  assign n1552 = x83 & n1426 ;
  assign n1553 = ( n1431 & n1551 ) | ( n1431 & n1552 ) | ( n1551 & n1552 ) ;
  assign n1554 = ( ~n1431 & n1551 ) | ( ~n1431 & n1552 ) | ( n1551 & n1552 ) ;
  assign n1555 = ( n1431 & ~n1553 ) | ( n1431 & n1554 ) | ( ~n1553 & n1554 ) ;
  assign n1556 = ( x84 & n1550 ) | ( x84 & ~n1555 ) | ( n1550 & ~n1555 ) ;
  assign n1557 = x85 | n1556 ;
  assign n1558 = ( x85 & n172 ) | ( x85 & n1556 ) | ( n172 & n1556 ) ;
  assign n1559 = ( n1437 & ~n1557 ) | ( n1437 & n1558 ) | ( ~n1557 & n1558 ) ;
  assign n1560 = ( x85 & ~n1437 ) | ( x85 & n1556 ) | ( ~n1437 & n1556 ) ;
  assign n1561 = n172 | n1560 ;
  assign n1562 = ( x42 & ~x64 ) | ( x42 & n1561 ) | ( ~x64 & n1561 ) ;
  assign n1563 = ~x42 & n1561 ;
  assign n1564 = ( n1441 & n1562 ) | ( n1441 & ~n1563 ) | ( n1562 & ~n1563 ) ;
  assign n1565 = ~x41 & x64 ;
  assign n1566 = ( x65 & ~n1564 ) | ( x65 & n1565 ) | ( ~n1564 & n1565 ) ;
  assign n1567 = ( x65 & n1441 ) | ( x65 & ~n1561 ) | ( n1441 & ~n1561 ) ;
  assign n1568 = x65 & n1441 ;
  assign n1569 = ( n1440 & n1567 ) | ( n1440 & n1568 ) | ( n1567 & n1568 ) ;
  assign n1570 = ( ~n1440 & n1567 ) | ( ~n1440 & n1568 ) | ( n1567 & n1568 ) ;
  assign n1571 = ( n1440 & ~n1569 ) | ( n1440 & n1570 ) | ( ~n1569 & n1570 ) ;
  assign n1572 = ( x66 & n1566 ) | ( x66 & ~n1571 ) | ( n1566 & ~n1571 ) ;
  assign n1573 = ( x66 & n1442 ) | ( x66 & ~n1561 ) | ( n1442 & ~n1561 ) ;
  assign n1574 = x66 & n1442 ;
  assign n1575 = ( n1447 & n1573 ) | ( n1447 & n1574 ) | ( n1573 & n1574 ) ;
  assign n1576 = ( ~n1447 & n1573 ) | ( ~n1447 & n1574 ) | ( n1573 & n1574 ) ;
  assign n1577 = ( n1447 & ~n1575 ) | ( n1447 & n1576 ) | ( ~n1575 & n1576 ) ;
  assign n1578 = ( x67 & n1572 ) | ( x67 & ~n1577 ) | ( n1572 & ~n1577 ) ;
  assign n1579 = ( x67 & n1448 ) | ( x67 & ~n1561 ) | ( n1448 & ~n1561 ) ;
  assign n1580 = x67 & n1448 ;
  assign n1581 = ( ~n1453 & n1579 ) | ( ~n1453 & n1580 ) | ( n1579 & n1580 ) ;
  assign n1582 = ( n1453 & n1579 ) | ( n1453 & n1580 ) | ( n1579 & n1580 ) ;
  assign n1583 = ( n1453 & n1581 ) | ( n1453 & ~n1582 ) | ( n1581 & ~n1582 ) ;
  assign n1584 = ( x68 & n1578 ) | ( x68 & ~n1583 ) | ( n1578 & ~n1583 ) ;
  assign n1585 = ( x68 & n1454 ) | ( x68 & ~n1561 ) | ( n1454 & ~n1561 ) ;
  assign n1586 = x68 & n1454 ;
  assign n1587 = ( n1459 & n1585 ) | ( n1459 & n1586 ) | ( n1585 & n1586 ) ;
  assign n1588 = ( ~n1459 & n1585 ) | ( ~n1459 & n1586 ) | ( n1585 & n1586 ) ;
  assign n1589 = ( n1459 & ~n1587 ) | ( n1459 & n1588 ) | ( ~n1587 & n1588 ) ;
  assign n1590 = ( x69 & n1584 ) | ( x69 & ~n1589 ) | ( n1584 & ~n1589 ) ;
  assign n1591 = ( x69 & n1460 ) | ( x69 & ~n1561 ) | ( n1460 & ~n1561 ) ;
  assign n1592 = x69 & n1460 ;
  assign n1593 = ( ~n1465 & n1591 ) | ( ~n1465 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = ( n1465 & n1591 ) | ( n1465 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1595 = ( n1465 & n1593 ) | ( n1465 & ~n1594 ) | ( n1593 & ~n1594 ) ;
  assign n1596 = ( x70 & n1590 ) | ( x70 & ~n1595 ) | ( n1590 & ~n1595 ) ;
  assign n1597 = ( x70 & n1466 ) | ( x70 & ~n1561 ) | ( n1466 & ~n1561 ) ;
  assign n1598 = x70 & n1466 ;
  assign n1599 = ( n1471 & n1597 ) | ( n1471 & n1598 ) | ( n1597 & n1598 ) ;
  assign n1600 = ( ~n1471 & n1597 ) | ( ~n1471 & n1598 ) | ( n1597 & n1598 ) ;
  assign n1601 = ( n1471 & ~n1599 ) | ( n1471 & n1600 ) | ( ~n1599 & n1600 ) ;
  assign n1602 = ( x71 & n1596 ) | ( x71 & ~n1601 ) | ( n1596 & ~n1601 ) ;
  assign n1603 = ( x71 & n1472 ) | ( x71 & ~n1561 ) | ( n1472 & ~n1561 ) ;
  assign n1604 = x71 & n1472 ;
  assign n1605 = ( ~n1477 & n1603 ) | ( ~n1477 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1606 = ( n1477 & n1603 ) | ( n1477 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1607 = ( n1477 & n1605 ) | ( n1477 & ~n1606 ) | ( n1605 & ~n1606 ) ;
  assign n1608 = ( x72 & n1602 ) | ( x72 & ~n1607 ) | ( n1602 & ~n1607 ) ;
  assign n1609 = ( x72 & n1478 ) | ( x72 & ~n1561 ) | ( n1478 & ~n1561 ) ;
  assign n1610 = x72 & n1478 ;
  assign n1611 = ( n1483 & n1609 ) | ( n1483 & n1610 ) | ( n1609 & n1610 ) ;
  assign n1612 = ( ~n1483 & n1609 ) | ( ~n1483 & n1610 ) | ( n1609 & n1610 ) ;
  assign n1613 = ( n1483 & ~n1611 ) | ( n1483 & n1612 ) | ( ~n1611 & n1612 ) ;
  assign n1614 = ( x73 & n1608 ) | ( x73 & ~n1613 ) | ( n1608 & ~n1613 ) ;
  assign n1615 = ( x73 & n1484 ) | ( x73 & ~n1561 ) | ( n1484 & ~n1561 ) ;
  assign n1616 = x73 & n1484 ;
  assign n1617 = ( ~n1489 & n1615 ) | ( ~n1489 & n1616 ) | ( n1615 & n1616 ) ;
  assign n1618 = ( n1489 & n1615 ) | ( n1489 & n1616 ) | ( n1615 & n1616 ) ;
  assign n1619 = ( n1489 & n1617 ) | ( n1489 & ~n1618 ) | ( n1617 & ~n1618 ) ;
  assign n1620 = ( x74 & n1614 ) | ( x74 & ~n1619 ) | ( n1614 & ~n1619 ) ;
  assign n1621 = ( x74 & n1490 ) | ( x74 & ~n1561 ) | ( n1490 & ~n1561 ) ;
  assign n1622 = x74 & n1490 ;
  assign n1623 = ( n1495 & n1621 ) | ( n1495 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1624 = ( ~n1495 & n1621 ) | ( ~n1495 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1625 = ( n1495 & ~n1623 ) | ( n1495 & n1624 ) | ( ~n1623 & n1624 ) ;
  assign n1626 = ( x75 & n1620 ) | ( x75 & ~n1625 ) | ( n1620 & ~n1625 ) ;
  assign n1627 = ( x75 & n1496 ) | ( x75 & ~n1561 ) | ( n1496 & ~n1561 ) ;
  assign n1628 = x75 & n1496 ;
  assign n1629 = ( ~n1501 & n1627 ) | ( ~n1501 & n1628 ) | ( n1627 & n1628 ) ;
  assign n1630 = ( n1501 & n1627 ) | ( n1501 & n1628 ) | ( n1627 & n1628 ) ;
  assign n1631 = ( n1501 & n1629 ) | ( n1501 & ~n1630 ) | ( n1629 & ~n1630 ) ;
  assign n1632 = ( x76 & n1626 ) | ( x76 & ~n1631 ) | ( n1626 & ~n1631 ) ;
  assign n1633 = ( x76 & n1502 ) | ( x76 & ~n1561 ) | ( n1502 & ~n1561 ) ;
  assign n1634 = x76 & n1502 ;
  assign n1635 = ( n1507 & n1633 ) | ( n1507 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1636 = ( ~n1507 & n1633 ) | ( ~n1507 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1637 = ( n1507 & ~n1635 ) | ( n1507 & n1636 ) | ( ~n1635 & n1636 ) ;
  assign n1638 = ( x77 & n1632 ) | ( x77 & ~n1637 ) | ( n1632 & ~n1637 ) ;
  assign n1639 = ( x77 & n1508 ) | ( x77 & ~n1561 ) | ( n1508 & ~n1561 ) ;
  assign n1640 = x77 & n1508 ;
  assign n1641 = ( ~n1513 & n1639 ) | ( ~n1513 & n1640 ) | ( n1639 & n1640 ) ;
  assign n1642 = ( n1513 & n1639 ) | ( n1513 & n1640 ) | ( n1639 & n1640 ) ;
  assign n1643 = ( n1513 & n1641 ) | ( n1513 & ~n1642 ) | ( n1641 & ~n1642 ) ;
  assign n1644 = ( x78 & n1638 ) | ( x78 & ~n1643 ) | ( n1638 & ~n1643 ) ;
  assign n1645 = ( x78 & n1514 ) | ( x78 & ~n1561 ) | ( n1514 & ~n1561 ) ;
  assign n1646 = x78 & n1514 ;
  assign n1647 = ( n1519 & n1645 ) | ( n1519 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1648 = ( ~n1519 & n1645 ) | ( ~n1519 & n1646 ) | ( n1645 & n1646 ) ;
  assign n1649 = ( n1519 & ~n1647 ) | ( n1519 & n1648 ) | ( ~n1647 & n1648 ) ;
  assign n1650 = ( x79 & n1644 ) | ( x79 & ~n1649 ) | ( n1644 & ~n1649 ) ;
  assign n1651 = ( x79 & n1520 ) | ( x79 & ~n1561 ) | ( n1520 & ~n1561 ) ;
  assign n1652 = x79 & n1520 ;
  assign n1653 = ( ~n1525 & n1651 ) | ( ~n1525 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1654 = ( n1525 & n1651 ) | ( n1525 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1655 = ( n1525 & n1653 ) | ( n1525 & ~n1654 ) | ( n1653 & ~n1654 ) ;
  assign n1656 = ( x80 & n1650 ) | ( x80 & ~n1655 ) | ( n1650 & ~n1655 ) ;
  assign n1657 = ( x80 & n1526 ) | ( x80 & ~n1561 ) | ( n1526 & ~n1561 ) ;
  assign n1658 = x80 & n1526 ;
  assign n1659 = ( n1531 & n1657 ) | ( n1531 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1660 = ( ~n1531 & n1657 ) | ( ~n1531 & n1658 ) | ( n1657 & n1658 ) ;
  assign n1661 = ( n1531 & ~n1659 ) | ( n1531 & n1660 ) | ( ~n1659 & n1660 ) ;
  assign n1662 = ( x81 & n1656 ) | ( x81 & ~n1661 ) | ( n1656 & ~n1661 ) ;
  assign n1663 = ( x81 & n1532 ) | ( x81 & ~n1561 ) | ( n1532 & ~n1561 ) ;
  assign n1664 = x81 & n1532 ;
  assign n1665 = ( ~n1537 & n1663 ) | ( ~n1537 & n1664 ) | ( n1663 & n1664 ) ;
  assign n1666 = ( n1537 & n1663 ) | ( n1537 & n1664 ) | ( n1663 & n1664 ) ;
  assign n1667 = ( n1537 & n1665 ) | ( n1537 & ~n1666 ) | ( n1665 & ~n1666 ) ;
  assign n1668 = ( x82 & n1662 ) | ( x82 & ~n1667 ) | ( n1662 & ~n1667 ) ;
  assign n1669 = ( x82 & n1538 ) | ( x82 & ~n1561 ) | ( n1538 & ~n1561 ) ;
  assign n1670 = x82 & n1538 ;
  assign n1671 = ( n1543 & n1669 ) | ( n1543 & n1670 ) | ( n1669 & n1670 ) ;
  assign n1672 = ( ~n1543 & n1669 ) | ( ~n1543 & n1670 ) | ( n1669 & n1670 ) ;
  assign n1673 = ( n1543 & ~n1671 ) | ( n1543 & n1672 ) | ( ~n1671 & n1672 ) ;
  assign n1674 = ( x83 & n1668 ) | ( x83 & ~n1673 ) | ( n1668 & ~n1673 ) ;
  assign n1675 = ( x83 & n1544 ) | ( x83 & ~n1561 ) | ( n1544 & ~n1561 ) ;
  assign n1676 = x83 & n1544 ;
  assign n1677 = ( ~n1549 & n1675 ) | ( ~n1549 & n1676 ) | ( n1675 & n1676 ) ;
  assign n1678 = ( n1549 & n1675 ) | ( n1549 & n1676 ) | ( n1675 & n1676 ) ;
  assign n1679 = ( n1549 & n1677 ) | ( n1549 & ~n1678 ) | ( n1677 & ~n1678 ) ;
  assign n1680 = ( x84 & n1674 ) | ( x84 & ~n1679 ) | ( n1674 & ~n1679 ) ;
  assign n1681 = ( x84 & n1550 ) | ( x84 & ~n1561 ) | ( n1550 & ~n1561 ) ;
  assign n1682 = x84 & n1550 ;
  assign n1683 = ( ~n1555 & n1681 ) | ( ~n1555 & n1682 ) | ( n1681 & n1682 ) ;
  assign n1684 = ( n1555 & n1681 ) | ( n1555 & n1682 ) | ( n1681 & n1682 ) ;
  assign n1685 = ( n1555 & n1683 ) | ( n1555 & ~n1684 ) | ( n1683 & ~n1684 ) ;
  assign n1686 = ( x85 & n1680 ) | ( x85 & ~n1685 ) | ( n1680 & ~n1685 ) ;
  assign n1687 = x86 | n1686 ;
  assign n1688 = x87 | n170 ;
  assign n1689 = ( x86 & n1686 ) | ( x86 & n1688 ) | ( n1686 & n1688 ) ;
  assign n1690 = ( n1559 & ~n1687 ) | ( n1559 & n1689 ) | ( ~n1687 & n1689 ) ;
  assign n1691 = ( x86 & ~n1559 ) | ( x86 & n1686 ) | ( ~n1559 & n1686 ) ;
  assign n1692 = n1688 | n1691 ;
  assign n1693 = ( x41 & ~x64 ) | ( x41 & n1692 ) | ( ~x64 & n1692 ) ;
  assign n1694 = ~x41 & n1692 ;
  assign n1695 = ( n1565 & n1693 ) | ( n1565 & ~n1694 ) | ( n1693 & ~n1694 ) ;
  assign n1696 = ~x40 & x64 ;
  assign n1697 = ( x65 & ~n1695 ) | ( x65 & n1696 ) | ( ~n1695 & n1696 ) ;
  assign n1698 = ( x65 & n1565 ) | ( x65 & ~n1692 ) | ( n1565 & ~n1692 ) ;
  assign n1699 = x65 & n1565 ;
  assign n1700 = ( n1564 & n1698 ) | ( n1564 & n1699 ) | ( n1698 & n1699 ) ;
  assign n1701 = ( ~n1564 & n1698 ) | ( ~n1564 & n1699 ) | ( n1698 & n1699 ) ;
  assign n1702 = ( n1564 & ~n1700 ) | ( n1564 & n1701 ) | ( ~n1700 & n1701 ) ;
  assign n1703 = ( x66 & n1697 ) | ( x66 & ~n1702 ) | ( n1697 & ~n1702 ) ;
  assign n1704 = ( x66 & n1566 ) | ( x66 & n1692 ) | ( n1566 & n1692 ) ;
  assign n1705 = x66 | n1566 ;
  assign n1706 = ( ~n1571 & n1704 ) | ( ~n1571 & n1705 ) | ( n1704 & n1705 ) ;
  assign n1707 = ( n1571 & n1704 ) | ( n1571 & n1705 ) | ( n1704 & n1705 ) ;
  assign n1708 = ( n1571 & n1706 ) | ( n1571 & ~n1707 ) | ( n1706 & ~n1707 ) ;
  assign n1709 = ( x67 & n1703 ) | ( x67 & ~n1708 ) | ( n1703 & ~n1708 ) ;
  assign n1710 = ( x67 & n1572 ) | ( x67 & ~n1692 ) | ( n1572 & ~n1692 ) ;
  assign n1711 = x67 & n1572 ;
  assign n1712 = ( ~n1577 & n1710 ) | ( ~n1577 & n1711 ) | ( n1710 & n1711 ) ;
  assign n1713 = ( n1577 & n1710 ) | ( n1577 & n1711 ) | ( n1710 & n1711 ) ;
  assign n1714 = ( n1577 & n1712 ) | ( n1577 & ~n1713 ) | ( n1712 & ~n1713 ) ;
  assign n1715 = ( x68 & n1709 ) | ( x68 & ~n1714 ) | ( n1709 & ~n1714 ) ;
  assign n1716 = ( x68 & n1578 ) | ( x68 & ~n1692 ) | ( n1578 & ~n1692 ) ;
  assign n1717 = x68 & n1578 ;
  assign n1718 = ( n1583 & n1716 ) | ( n1583 & n1717 ) | ( n1716 & n1717 ) ;
  assign n1719 = ( ~n1583 & n1716 ) | ( ~n1583 & n1717 ) | ( n1716 & n1717 ) ;
  assign n1720 = ( n1583 & ~n1718 ) | ( n1583 & n1719 ) | ( ~n1718 & n1719 ) ;
  assign n1721 = ( x69 & n1715 ) | ( x69 & ~n1720 ) | ( n1715 & ~n1720 ) ;
  assign n1722 = ( x69 & n1584 ) | ( x69 & ~n1692 ) | ( n1584 & ~n1692 ) ;
  assign n1723 = x69 & n1584 ;
  assign n1724 = ( ~n1589 & n1722 ) | ( ~n1589 & n1723 ) | ( n1722 & n1723 ) ;
  assign n1725 = ( n1589 & n1722 ) | ( n1589 & n1723 ) | ( n1722 & n1723 ) ;
  assign n1726 = ( n1589 & n1724 ) | ( n1589 & ~n1725 ) | ( n1724 & ~n1725 ) ;
  assign n1727 = ( x70 & n1721 ) | ( x70 & ~n1726 ) | ( n1721 & ~n1726 ) ;
  assign n1728 = ( x70 & n1590 ) | ( x70 & ~n1692 ) | ( n1590 & ~n1692 ) ;
  assign n1729 = x70 & n1590 ;
  assign n1730 = ( n1595 & n1728 ) | ( n1595 & n1729 ) | ( n1728 & n1729 ) ;
  assign n1731 = ( ~n1595 & n1728 ) | ( ~n1595 & n1729 ) | ( n1728 & n1729 ) ;
  assign n1732 = ( n1595 & ~n1730 ) | ( n1595 & n1731 ) | ( ~n1730 & n1731 ) ;
  assign n1733 = ( x71 & n1727 ) | ( x71 & ~n1732 ) | ( n1727 & ~n1732 ) ;
  assign n1734 = ( x71 & n1596 ) | ( x71 & ~n1692 ) | ( n1596 & ~n1692 ) ;
  assign n1735 = x71 & n1596 ;
  assign n1736 = ( ~n1601 & n1734 ) | ( ~n1601 & n1735 ) | ( n1734 & n1735 ) ;
  assign n1737 = ( n1601 & n1734 ) | ( n1601 & n1735 ) | ( n1734 & n1735 ) ;
  assign n1738 = ( n1601 & n1736 ) | ( n1601 & ~n1737 ) | ( n1736 & ~n1737 ) ;
  assign n1739 = ( x72 & n1733 ) | ( x72 & ~n1738 ) | ( n1733 & ~n1738 ) ;
  assign n1740 = ( x72 & n1602 ) | ( x72 & ~n1692 ) | ( n1602 & ~n1692 ) ;
  assign n1741 = x72 & n1602 ;
  assign n1742 = ( n1607 & n1740 ) | ( n1607 & n1741 ) | ( n1740 & n1741 ) ;
  assign n1743 = ( ~n1607 & n1740 ) | ( ~n1607 & n1741 ) | ( n1740 & n1741 ) ;
  assign n1744 = ( n1607 & ~n1742 ) | ( n1607 & n1743 ) | ( ~n1742 & n1743 ) ;
  assign n1745 = ( x73 & n1739 ) | ( x73 & ~n1744 ) | ( n1739 & ~n1744 ) ;
  assign n1746 = ( x73 & n1608 ) | ( x73 & ~n1692 ) | ( n1608 & ~n1692 ) ;
  assign n1747 = x73 & n1608 ;
  assign n1748 = ( ~n1613 & n1746 ) | ( ~n1613 & n1747 ) | ( n1746 & n1747 ) ;
  assign n1749 = ( n1613 & n1746 ) | ( n1613 & n1747 ) | ( n1746 & n1747 ) ;
  assign n1750 = ( n1613 & n1748 ) | ( n1613 & ~n1749 ) | ( n1748 & ~n1749 ) ;
  assign n1751 = ( x74 & n1745 ) | ( x74 & ~n1750 ) | ( n1745 & ~n1750 ) ;
  assign n1752 = ( x74 & n1614 ) | ( x74 & ~n1692 ) | ( n1614 & ~n1692 ) ;
  assign n1753 = x74 & n1614 ;
  assign n1754 = ( n1619 & n1752 ) | ( n1619 & n1753 ) | ( n1752 & n1753 ) ;
  assign n1755 = ( ~n1619 & n1752 ) | ( ~n1619 & n1753 ) | ( n1752 & n1753 ) ;
  assign n1756 = ( n1619 & ~n1754 ) | ( n1619 & n1755 ) | ( ~n1754 & n1755 ) ;
  assign n1757 = ( x75 & n1751 ) | ( x75 & ~n1756 ) | ( n1751 & ~n1756 ) ;
  assign n1758 = ( x75 & n1620 ) | ( x75 & ~n1692 ) | ( n1620 & ~n1692 ) ;
  assign n1759 = x75 & n1620 ;
  assign n1760 = ( ~n1625 & n1758 ) | ( ~n1625 & n1759 ) | ( n1758 & n1759 ) ;
  assign n1761 = ( n1625 & n1758 ) | ( n1625 & n1759 ) | ( n1758 & n1759 ) ;
  assign n1762 = ( n1625 & n1760 ) | ( n1625 & ~n1761 ) | ( n1760 & ~n1761 ) ;
  assign n1763 = ( x76 & n1757 ) | ( x76 & ~n1762 ) | ( n1757 & ~n1762 ) ;
  assign n1764 = ( x76 & n1626 ) | ( x76 & ~n1692 ) | ( n1626 & ~n1692 ) ;
  assign n1765 = x76 & n1626 ;
  assign n1766 = ( n1631 & n1764 ) | ( n1631 & n1765 ) | ( n1764 & n1765 ) ;
  assign n1767 = ( ~n1631 & n1764 ) | ( ~n1631 & n1765 ) | ( n1764 & n1765 ) ;
  assign n1768 = ( n1631 & ~n1766 ) | ( n1631 & n1767 ) | ( ~n1766 & n1767 ) ;
  assign n1769 = ( x77 & n1763 ) | ( x77 & ~n1768 ) | ( n1763 & ~n1768 ) ;
  assign n1770 = ( x77 & n1632 ) | ( x77 & ~n1692 ) | ( n1632 & ~n1692 ) ;
  assign n1771 = x77 & n1632 ;
  assign n1772 = ( ~n1637 & n1770 ) | ( ~n1637 & n1771 ) | ( n1770 & n1771 ) ;
  assign n1773 = ( n1637 & n1770 ) | ( n1637 & n1771 ) | ( n1770 & n1771 ) ;
  assign n1774 = ( n1637 & n1772 ) | ( n1637 & ~n1773 ) | ( n1772 & ~n1773 ) ;
  assign n1775 = ( x78 & n1769 ) | ( x78 & ~n1774 ) | ( n1769 & ~n1774 ) ;
  assign n1776 = ( x78 & n1638 ) | ( x78 & ~n1692 ) | ( n1638 & ~n1692 ) ;
  assign n1777 = x78 & n1638 ;
  assign n1778 = ( n1643 & n1776 ) | ( n1643 & n1777 ) | ( n1776 & n1777 ) ;
  assign n1779 = ( ~n1643 & n1776 ) | ( ~n1643 & n1777 ) | ( n1776 & n1777 ) ;
  assign n1780 = ( n1643 & ~n1778 ) | ( n1643 & n1779 ) | ( ~n1778 & n1779 ) ;
  assign n1781 = ( x79 & n1775 ) | ( x79 & ~n1780 ) | ( n1775 & ~n1780 ) ;
  assign n1782 = ( x79 & n1644 ) | ( x79 & ~n1692 ) | ( n1644 & ~n1692 ) ;
  assign n1783 = x79 & n1644 ;
  assign n1784 = ( ~n1649 & n1782 ) | ( ~n1649 & n1783 ) | ( n1782 & n1783 ) ;
  assign n1785 = ( n1649 & n1782 ) | ( n1649 & n1783 ) | ( n1782 & n1783 ) ;
  assign n1786 = ( n1649 & n1784 ) | ( n1649 & ~n1785 ) | ( n1784 & ~n1785 ) ;
  assign n1787 = ( x80 & n1781 ) | ( x80 & ~n1786 ) | ( n1781 & ~n1786 ) ;
  assign n1788 = ( x80 & n1650 ) | ( x80 & ~n1692 ) | ( n1650 & ~n1692 ) ;
  assign n1789 = x80 & n1650 ;
  assign n1790 = ( n1655 & n1788 ) | ( n1655 & n1789 ) | ( n1788 & n1789 ) ;
  assign n1791 = ( ~n1655 & n1788 ) | ( ~n1655 & n1789 ) | ( n1788 & n1789 ) ;
  assign n1792 = ( n1655 & ~n1790 ) | ( n1655 & n1791 ) | ( ~n1790 & n1791 ) ;
  assign n1793 = ( x81 & n1787 ) | ( x81 & ~n1792 ) | ( n1787 & ~n1792 ) ;
  assign n1794 = ( x81 & n1656 ) | ( x81 & ~n1692 ) | ( n1656 & ~n1692 ) ;
  assign n1795 = x81 & n1656 ;
  assign n1796 = ( ~n1661 & n1794 ) | ( ~n1661 & n1795 ) | ( n1794 & n1795 ) ;
  assign n1797 = ( n1661 & n1794 ) | ( n1661 & n1795 ) | ( n1794 & n1795 ) ;
  assign n1798 = ( n1661 & n1796 ) | ( n1661 & ~n1797 ) | ( n1796 & ~n1797 ) ;
  assign n1799 = ( x82 & n1793 ) | ( x82 & ~n1798 ) | ( n1793 & ~n1798 ) ;
  assign n1800 = ( x82 & n1662 ) | ( x82 & ~n1692 ) | ( n1662 & ~n1692 ) ;
  assign n1801 = x82 & n1662 ;
  assign n1802 = ( n1667 & n1800 ) | ( n1667 & n1801 ) | ( n1800 & n1801 ) ;
  assign n1803 = ( ~n1667 & n1800 ) | ( ~n1667 & n1801 ) | ( n1800 & n1801 ) ;
  assign n1804 = ( n1667 & ~n1802 ) | ( n1667 & n1803 ) | ( ~n1802 & n1803 ) ;
  assign n1805 = ( x83 & n1799 ) | ( x83 & ~n1804 ) | ( n1799 & ~n1804 ) ;
  assign n1806 = ( x83 & n1668 ) | ( x83 & ~n1692 ) | ( n1668 & ~n1692 ) ;
  assign n1807 = x83 & n1668 ;
  assign n1808 = ( ~n1673 & n1806 ) | ( ~n1673 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1809 = ( n1673 & n1806 ) | ( n1673 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1810 = ( n1673 & n1808 ) | ( n1673 & ~n1809 ) | ( n1808 & ~n1809 ) ;
  assign n1811 = ( x84 & n1805 ) | ( x84 & ~n1810 ) | ( n1805 & ~n1810 ) ;
  assign n1812 = ( x84 & n1674 ) | ( x84 & ~n1692 ) | ( n1674 & ~n1692 ) ;
  assign n1813 = x84 & n1674 ;
  assign n1814 = ( n1679 & n1812 ) | ( n1679 & n1813 ) | ( n1812 & n1813 ) ;
  assign n1815 = ( ~n1679 & n1812 ) | ( ~n1679 & n1813 ) | ( n1812 & n1813 ) ;
  assign n1816 = ( n1679 & ~n1814 ) | ( n1679 & n1815 ) | ( ~n1814 & n1815 ) ;
  assign n1817 = ( x85 & n1811 ) | ( x85 & ~n1816 ) | ( n1811 & ~n1816 ) ;
  assign n1818 = ( x85 & n1680 ) | ( x85 & ~n1692 ) | ( n1680 & ~n1692 ) ;
  assign n1819 = x85 & n1680 ;
  assign n1820 = ( n1685 & n1818 ) | ( n1685 & n1819 ) | ( n1818 & n1819 ) ;
  assign n1821 = ( ~n1685 & n1818 ) | ( ~n1685 & n1819 ) | ( n1818 & n1819 ) ;
  assign n1822 = ( n1685 & ~n1820 ) | ( n1685 & n1821 ) | ( ~n1820 & n1821 ) ;
  assign n1823 = ( x86 & n1817 ) | ( x86 & ~n1822 ) | ( n1817 & ~n1822 ) ;
  assign n1824 = ( x87 & ~n1690 ) | ( x87 & n1823 ) | ( ~n1690 & n1823 ) ;
  assign n1825 = n170 | n1824 ;
  assign n1826 = n1690 & n1825 ;
  assign n1827 = n280 | n1826 ;
  assign n1828 = ( x40 & ~x64 ) | ( x40 & n1825 ) | ( ~x64 & n1825 ) ;
  assign n1829 = ~x40 & n1825 ;
  assign n1830 = ( n1696 & n1828 ) | ( n1696 & ~n1829 ) | ( n1828 & ~n1829 ) ;
  assign n1831 = ~x39 & x64 ;
  assign n1832 = ( x65 & ~n1830 ) | ( x65 & n1831 ) | ( ~n1830 & n1831 ) ;
  assign n1833 = ( x65 & n1696 ) | ( x65 & ~n1825 ) | ( n1696 & ~n1825 ) ;
  assign n1834 = x65 & n1696 ;
  assign n1835 = ( n1695 & n1833 ) | ( n1695 & n1834 ) | ( n1833 & n1834 ) ;
  assign n1836 = ( ~n1695 & n1833 ) | ( ~n1695 & n1834 ) | ( n1833 & n1834 ) ;
  assign n1837 = ( n1695 & ~n1835 ) | ( n1695 & n1836 ) | ( ~n1835 & n1836 ) ;
  assign n1838 = ( x66 & n1832 ) | ( x66 & ~n1837 ) | ( n1832 & ~n1837 ) ;
  assign n1839 = ( x66 & n1697 ) | ( x66 & ~n1825 ) | ( n1697 & ~n1825 ) ;
  assign n1840 = x66 & n1697 ;
  assign n1841 = ( n1702 & n1839 ) | ( n1702 & n1840 ) | ( n1839 & n1840 ) ;
  assign n1842 = ( ~n1702 & n1839 ) | ( ~n1702 & n1840 ) | ( n1839 & n1840 ) ;
  assign n1843 = ( n1702 & ~n1841 ) | ( n1702 & n1842 ) | ( ~n1841 & n1842 ) ;
  assign n1844 = ( x67 & n1838 ) | ( x67 & ~n1843 ) | ( n1838 & ~n1843 ) ;
  assign n1845 = ( x67 & n1703 ) | ( x67 & ~n1825 ) | ( n1703 & ~n1825 ) ;
  assign n1846 = x67 & n1703 ;
  assign n1847 = ( ~n1708 & n1845 ) | ( ~n1708 & n1846 ) | ( n1845 & n1846 ) ;
  assign n1848 = ( n1708 & n1845 ) | ( n1708 & n1846 ) | ( n1845 & n1846 ) ;
  assign n1849 = ( n1708 & n1847 ) | ( n1708 & ~n1848 ) | ( n1847 & ~n1848 ) ;
  assign n1850 = ( x68 & n1844 ) | ( x68 & ~n1849 ) | ( n1844 & ~n1849 ) ;
  assign n1851 = ( x68 & n1709 ) | ( x68 & ~n1825 ) | ( n1709 & ~n1825 ) ;
  assign n1852 = x68 & n1709 ;
  assign n1853 = ( n1714 & n1851 ) | ( n1714 & n1852 ) | ( n1851 & n1852 ) ;
  assign n1854 = ( ~n1714 & n1851 ) | ( ~n1714 & n1852 ) | ( n1851 & n1852 ) ;
  assign n1855 = ( n1714 & ~n1853 ) | ( n1714 & n1854 ) | ( ~n1853 & n1854 ) ;
  assign n1856 = ( x69 & n1850 ) | ( x69 & ~n1855 ) | ( n1850 & ~n1855 ) ;
  assign n1857 = ( x69 & n1715 ) | ( x69 & ~n1825 ) | ( n1715 & ~n1825 ) ;
  assign n1858 = x69 & n1715 ;
  assign n1859 = ( ~n1720 & n1857 ) | ( ~n1720 & n1858 ) | ( n1857 & n1858 ) ;
  assign n1860 = ( n1720 & n1857 ) | ( n1720 & n1858 ) | ( n1857 & n1858 ) ;
  assign n1861 = ( n1720 & n1859 ) | ( n1720 & ~n1860 ) | ( n1859 & ~n1860 ) ;
  assign n1862 = ( x70 & n1856 ) | ( x70 & ~n1861 ) | ( n1856 & ~n1861 ) ;
  assign n1863 = ( x70 & n1721 ) | ( x70 & ~n1825 ) | ( n1721 & ~n1825 ) ;
  assign n1864 = x70 & n1721 ;
  assign n1865 = ( n1726 & n1863 ) | ( n1726 & n1864 ) | ( n1863 & n1864 ) ;
  assign n1866 = ( ~n1726 & n1863 ) | ( ~n1726 & n1864 ) | ( n1863 & n1864 ) ;
  assign n1867 = ( n1726 & ~n1865 ) | ( n1726 & n1866 ) | ( ~n1865 & n1866 ) ;
  assign n1868 = ( x71 & n1862 ) | ( x71 & ~n1867 ) | ( n1862 & ~n1867 ) ;
  assign n1869 = ( x71 & n1727 ) | ( x71 & ~n1825 ) | ( n1727 & ~n1825 ) ;
  assign n1870 = x71 & n1727 ;
  assign n1871 = ( ~n1732 & n1869 ) | ( ~n1732 & n1870 ) | ( n1869 & n1870 ) ;
  assign n1872 = ( n1732 & n1869 ) | ( n1732 & n1870 ) | ( n1869 & n1870 ) ;
  assign n1873 = ( n1732 & n1871 ) | ( n1732 & ~n1872 ) | ( n1871 & ~n1872 ) ;
  assign n1874 = ( x72 & n1868 ) | ( x72 & ~n1873 ) | ( n1868 & ~n1873 ) ;
  assign n1875 = ( x72 & n1733 ) | ( x72 & ~n1825 ) | ( n1733 & ~n1825 ) ;
  assign n1876 = x72 & n1733 ;
  assign n1877 = ( n1738 & n1875 ) | ( n1738 & n1876 ) | ( n1875 & n1876 ) ;
  assign n1878 = ( ~n1738 & n1875 ) | ( ~n1738 & n1876 ) | ( n1875 & n1876 ) ;
  assign n1879 = ( n1738 & ~n1877 ) | ( n1738 & n1878 ) | ( ~n1877 & n1878 ) ;
  assign n1880 = ( x73 & n1874 ) | ( x73 & ~n1879 ) | ( n1874 & ~n1879 ) ;
  assign n1881 = ( x73 & n1739 ) | ( x73 & ~n1825 ) | ( n1739 & ~n1825 ) ;
  assign n1882 = x73 & n1739 ;
  assign n1883 = ( ~n1744 & n1881 ) | ( ~n1744 & n1882 ) | ( n1881 & n1882 ) ;
  assign n1884 = ( n1744 & n1881 ) | ( n1744 & n1882 ) | ( n1881 & n1882 ) ;
  assign n1885 = ( n1744 & n1883 ) | ( n1744 & ~n1884 ) | ( n1883 & ~n1884 ) ;
  assign n1886 = ( x74 & n1880 ) | ( x74 & ~n1885 ) | ( n1880 & ~n1885 ) ;
  assign n1887 = ( x74 & n1745 ) | ( x74 & ~n1825 ) | ( n1745 & ~n1825 ) ;
  assign n1888 = x74 & n1745 ;
  assign n1889 = ( n1750 & n1887 ) | ( n1750 & n1888 ) | ( n1887 & n1888 ) ;
  assign n1890 = ( ~n1750 & n1887 ) | ( ~n1750 & n1888 ) | ( n1887 & n1888 ) ;
  assign n1891 = ( n1750 & ~n1889 ) | ( n1750 & n1890 ) | ( ~n1889 & n1890 ) ;
  assign n1892 = ( x75 & n1886 ) | ( x75 & ~n1891 ) | ( n1886 & ~n1891 ) ;
  assign n1893 = ( x75 & n1751 ) | ( x75 & ~n1825 ) | ( n1751 & ~n1825 ) ;
  assign n1894 = x75 & n1751 ;
  assign n1895 = ( ~n1756 & n1893 ) | ( ~n1756 & n1894 ) | ( n1893 & n1894 ) ;
  assign n1896 = ( n1756 & n1893 ) | ( n1756 & n1894 ) | ( n1893 & n1894 ) ;
  assign n1897 = ( n1756 & n1895 ) | ( n1756 & ~n1896 ) | ( n1895 & ~n1896 ) ;
  assign n1898 = ( x76 & n1892 ) | ( x76 & ~n1897 ) | ( n1892 & ~n1897 ) ;
  assign n1899 = ( x76 & n1757 ) | ( x76 & ~n1825 ) | ( n1757 & ~n1825 ) ;
  assign n1900 = x76 & n1757 ;
  assign n1901 = ( n1762 & n1899 ) | ( n1762 & n1900 ) | ( n1899 & n1900 ) ;
  assign n1902 = ( ~n1762 & n1899 ) | ( ~n1762 & n1900 ) | ( n1899 & n1900 ) ;
  assign n1903 = ( n1762 & ~n1901 ) | ( n1762 & n1902 ) | ( ~n1901 & n1902 ) ;
  assign n1904 = ( x77 & n1898 ) | ( x77 & ~n1903 ) | ( n1898 & ~n1903 ) ;
  assign n1905 = ( x77 & n1763 ) | ( x77 & ~n1825 ) | ( n1763 & ~n1825 ) ;
  assign n1906 = x77 & n1763 ;
  assign n1907 = ( ~n1768 & n1905 ) | ( ~n1768 & n1906 ) | ( n1905 & n1906 ) ;
  assign n1908 = ( n1768 & n1905 ) | ( n1768 & n1906 ) | ( n1905 & n1906 ) ;
  assign n1909 = ( n1768 & n1907 ) | ( n1768 & ~n1908 ) | ( n1907 & ~n1908 ) ;
  assign n1910 = ( x78 & n1904 ) | ( x78 & ~n1909 ) | ( n1904 & ~n1909 ) ;
  assign n1911 = ( x78 & n1769 ) | ( x78 & ~n1825 ) | ( n1769 & ~n1825 ) ;
  assign n1912 = x78 & n1769 ;
  assign n1913 = ( n1774 & n1911 ) | ( n1774 & n1912 ) | ( n1911 & n1912 ) ;
  assign n1914 = ( ~n1774 & n1911 ) | ( ~n1774 & n1912 ) | ( n1911 & n1912 ) ;
  assign n1915 = ( n1774 & ~n1913 ) | ( n1774 & n1914 ) | ( ~n1913 & n1914 ) ;
  assign n1916 = ( x79 & n1910 ) | ( x79 & ~n1915 ) | ( n1910 & ~n1915 ) ;
  assign n1917 = ( x79 & n1775 ) | ( x79 & ~n1825 ) | ( n1775 & ~n1825 ) ;
  assign n1918 = x79 & n1775 ;
  assign n1919 = ( ~n1780 & n1917 ) | ( ~n1780 & n1918 ) | ( n1917 & n1918 ) ;
  assign n1920 = ( n1780 & n1917 ) | ( n1780 & n1918 ) | ( n1917 & n1918 ) ;
  assign n1921 = ( n1780 & n1919 ) | ( n1780 & ~n1920 ) | ( n1919 & ~n1920 ) ;
  assign n1922 = ( x80 & n1916 ) | ( x80 & ~n1921 ) | ( n1916 & ~n1921 ) ;
  assign n1923 = ( x80 & n1781 ) | ( x80 & ~n1825 ) | ( n1781 & ~n1825 ) ;
  assign n1924 = x80 & n1781 ;
  assign n1925 = ( n1786 & n1923 ) | ( n1786 & n1924 ) | ( n1923 & n1924 ) ;
  assign n1926 = ( ~n1786 & n1923 ) | ( ~n1786 & n1924 ) | ( n1923 & n1924 ) ;
  assign n1927 = ( n1786 & ~n1925 ) | ( n1786 & n1926 ) | ( ~n1925 & n1926 ) ;
  assign n1928 = ( x81 & n1922 ) | ( x81 & ~n1927 ) | ( n1922 & ~n1927 ) ;
  assign n1929 = ( x81 & n1787 ) | ( x81 & ~n1825 ) | ( n1787 & ~n1825 ) ;
  assign n1930 = x81 & n1787 ;
  assign n1931 = ( ~n1792 & n1929 ) | ( ~n1792 & n1930 ) | ( n1929 & n1930 ) ;
  assign n1932 = ( n1792 & n1929 ) | ( n1792 & n1930 ) | ( n1929 & n1930 ) ;
  assign n1933 = ( n1792 & n1931 ) | ( n1792 & ~n1932 ) | ( n1931 & ~n1932 ) ;
  assign n1934 = ( x82 & n1928 ) | ( x82 & ~n1933 ) | ( n1928 & ~n1933 ) ;
  assign n1935 = ( x82 & n1793 ) | ( x82 & ~n1825 ) | ( n1793 & ~n1825 ) ;
  assign n1936 = x82 & n1793 ;
  assign n1937 = ( n1798 & n1935 ) | ( n1798 & n1936 ) | ( n1935 & n1936 ) ;
  assign n1938 = ( ~n1798 & n1935 ) | ( ~n1798 & n1936 ) | ( n1935 & n1936 ) ;
  assign n1939 = ( n1798 & ~n1937 ) | ( n1798 & n1938 ) | ( ~n1937 & n1938 ) ;
  assign n1940 = ( x83 & n1934 ) | ( x83 & ~n1939 ) | ( n1934 & ~n1939 ) ;
  assign n1941 = ( x83 & n1799 ) | ( x83 & ~n1825 ) | ( n1799 & ~n1825 ) ;
  assign n1942 = x83 & n1799 ;
  assign n1943 = ( ~n1804 & n1941 ) | ( ~n1804 & n1942 ) | ( n1941 & n1942 ) ;
  assign n1944 = ( n1804 & n1941 ) | ( n1804 & n1942 ) | ( n1941 & n1942 ) ;
  assign n1945 = ( n1804 & n1943 ) | ( n1804 & ~n1944 ) | ( n1943 & ~n1944 ) ;
  assign n1946 = ( x84 & n1940 ) | ( x84 & ~n1945 ) | ( n1940 & ~n1945 ) ;
  assign n1947 = ( x84 & n1805 ) | ( x84 & ~n1825 ) | ( n1805 & ~n1825 ) ;
  assign n1948 = x84 & n1805 ;
  assign n1949 = ( n1810 & n1947 ) | ( n1810 & n1948 ) | ( n1947 & n1948 ) ;
  assign n1950 = ( ~n1810 & n1947 ) | ( ~n1810 & n1948 ) | ( n1947 & n1948 ) ;
  assign n1951 = ( n1810 & ~n1949 ) | ( n1810 & n1950 ) | ( ~n1949 & n1950 ) ;
  assign n1952 = ( x85 & n1946 ) | ( x85 & ~n1951 ) | ( n1946 & ~n1951 ) ;
  assign n1953 = ( x85 & n1811 ) | ( x85 & ~n1825 ) | ( n1811 & ~n1825 ) ;
  assign n1954 = x85 & n1811 ;
  assign n1955 = ( ~n1816 & n1953 ) | ( ~n1816 & n1954 ) | ( n1953 & n1954 ) ;
  assign n1956 = ( n1816 & n1953 ) | ( n1816 & n1954 ) | ( n1953 & n1954 ) ;
  assign n1957 = ( n1816 & n1955 ) | ( n1816 & ~n1956 ) | ( n1955 & ~n1956 ) ;
  assign n1958 = ( x86 & n1952 ) | ( x86 & ~n1957 ) | ( n1952 & ~n1957 ) ;
  assign n1959 = ( x86 & n1817 ) | ( x86 & ~n1825 ) | ( n1817 & ~n1825 ) ;
  assign n1960 = x86 & n1817 ;
  assign n1961 = ( ~n1822 & n1959 ) | ( ~n1822 & n1960 ) | ( n1959 & n1960 ) ;
  assign n1962 = ( n1822 & n1959 ) | ( n1822 & n1960 ) | ( n1959 & n1960 ) ;
  assign n1963 = ( n1822 & n1961 ) | ( n1822 & ~n1962 ) | ( n1961 & ~n1962 ) ;
  assign n1964 = ( x87 & n1958 ) | ( x87 & ~n1963 ) | ( n1958 & ~n1963 ) ;
  assign n1965 = x88 | n1964 ;
  assign n1966 = ( x88 & n169 ) | ( x88 & n1964 ) | ( n169 & n1964 ) ;
  assign n1967 = ( n1827 & ~n1965 ) | ( n1827 & n1966 ) | ( ~n1965 & n1966 ) ;
  assign n1968 = ( x88 & ~n1827 ) | ( x88 & n1964 ) | ( ~n1827 & n1964 ) ;
  assign n1969 = n169 | n1968 ;
  assign n1970 = ( x39 & ~x64 ) | ( x39 & n1969 ) | ( ~x64 & n1969 ) ;
  assign n1971 = ~x39 & n1969 ;
  assign n1972 = ( n1831 & n1970 ) | ( n1831 & ~n1971 ) | ( n1970 & ~n1971 ) ;
  assign n1973 = ~x38 & x64 ;
  assign n1974 = ( x65 & ~n1972 ) | ( x65 & n1973 ) | ( ~n1972 & n1973 ) ;
  assign n1975 = ( x65 & n1831 ) | ( x65 & ~n1969 ) | ( n1831 & ~n1969 ) ;
  assign n1976 = x65 & n1831 ;
  assign n1977 = ( n1830 & n1975 ) | ( n1830 & n1976 ) | ( n1975 & n1976 ) ;
  assign n1978 = ( ~n1830 & n1975 ) | ( ~n1830 & n1976 ) | ( n1975 & n1976 ) ;
  assign n1979 = ( n1830 & ~n1977 ) | ( n1830 & n1978 ) | ( ~n1977 & n1978 ) ;
  assign n1980 = ( x66 & n1974 ) | ( x66 & ~n1979 ) | ( n1974 & ~n1979 ) ;
  assign n1981 = ( x66 & n1832 ) | ( x66 & ~n1969 ) | ( n1832 & ~n1969 ) ;
  assign n1982 = x66 & n1832 ;
  assign n1983 = ( n1837 & n1981 ) | ( n1837 & n1982 ) | ( n1981 & n1982 ) ;
  assign n1984 = ( ~n1837 & n1981 ) | ( ~n1837 & n1982 ) | ( n1981 & n1982 ) ;
  assign n1985 = ( n1837 & ~n1983 ) | ( n1837 & n1984 ) | ( ~n1983 & n1984 ) ;
  assign n1986 = ( x67 & n1980 ) | ( x67 & ~n1985 ) | ( n1980 & ~n1985 ) ;
  assign n1987 = ( x67 & n1838 ) | ( x67 & ~n1969 ) | ( n1838 & ~n1969 ) ;
  assign n1988 = x67 & n1838 ;
  assign n1989 = ( ~n1843 & n1987 ) | ( ~n1843 & n1988 ) | ( n1987 & n1988 ) ;
  assign n1990 = ( n1843 & n1987 ) | ( n1843 & n1988 ) | ( n1987 & n1988 ) ;
  assign n1991 = ( n1843 & n1989 ) | ( n1843 & ~n1990 ) | ( n1989 & ~n1990 ) ;
  assign n1992 = ( x68 & n1986 ) | ( x68 & ~n1991 ) | ( n1986 & ~n1991 ) ;
  assign n1993 = ( x68 & n1844 ) | ( x68 & ~n1969 ) | ( n1844 & ~n1969 ) ;
  assign n1994 = x68 & n1844 ;
  assign n1995 = ( n1849 & n1993 ) | ( n1849 & n1994 ) | ( n1993 & n1994 ) ;
  assign n1996 = ( ~n1849 & n1993 ) | ( ~n1849 & n1994 ) | ( n1993 & n1994 ) ;
  assign n1997 = ( n1849 & ~n1995 ) | ( n1849 & n1996 ) | ( ~n1995 & n1996 ) ;
  assign n1998 = ( x69 & n1992 ) | ( x69 & ~n1997 ) | ( n1992 & ~n1997 ) ;
  assign n1999 = ( x69 & n1850 ) | ( x69 & ~n1969 ) | ( n1850 & ~n1969 ) ;
  assign n2000 = x69 & n1850 ;
  assign n2001 = ( ~n1855 & n1999 ) | ( ~n1855 & n2000 ) | ( n1999 & n2000 ) ;
  assign n2002 = ( n1855 & n1999 ) | ( n1855 & n2000 ) | ( n1999 & n2000 ) ;
  assign n2003 = ( n1855 & n2001 ) | ( n1855 & ~n2002 ) | ( n2001 & ~n2002 ) ;
  assign n2004 = ( x70 & n1998 ) | ( x70 & ~n2003 ) | ( n1998 & ~n2003 ) ;
  assign n2005 = ( x70 & n1856 ) | ( x70 & ~n1969 ) | ( n1856 & ~n1969 ) ;
  assign n2006 = x70 & n1856 ;
  assign n2007 = ( n1861 & n2005 ) | ( n1861 & n2006 ) | ( n2005 & n2006 ) ;
  assign n2008 = ( ~n1861 & n2005 ) | ( ~n1861 & n2006 ) | ( n2005 & n2006 ) ;
  assign n2009 = ( n1861 & ~n2007 ) | ( n1861 & n2008 ) | ( ~n2007 & n2008 ) ;
  assign n2010 = ( x71 & n2004 ) | ( x71 & ~n2009 ) | ( n2004 & ~n2009 ) ;
  assign n2011 = ( x71 & n1862 ) | ( x71 & ~n1969 ) | ( n1862 & ~n1969 ) ;
  assign n2012 = x71 & n1862 ;
  assign n2013 = ( ~n1867 & n2011 ) | ( ~n1867 & n2012 ) | ( n2011 & n2012 ) ;
  assign n2014 = ( n1867 & n2011 ) | ( n1867 & n2012 ) | ( n2011 & n2012 ) ;
  assign n2015 = ( n1867 & n2013 ) | ( n1867 & ~n2014 ) | ( n2013 & ~n2014 ) ;
  assign n2016 = ( x72 & n2010 ) | ( x72 & ~n2015 ) | ( n2010 & ~n2015 ) ;
  assign n2017 = ( x72 & n1868 ) | ( x72 & ~n1969 ) | ( n1868 & ~n1969 ) ;
  assign n2018 = x72 & n1868 ;
  assign n2019 = ( n1873 & n2017 ) | ( n1873 & n2018 ) | ( n2017 & n2018 ) ;
  assign n2020 = ( ~n1873 & n2017 ) | ( ~n1873 & n2018 ) | ( n2017 & n2018 ) ;
  assign n2021 = ( n1873 & ~n2019 ) | ( n1873 & n2020 ) | ( ~n2019 & n2020 ) ;
  assign n2022 = ( x73 & n2016 ) | ( x73 & ~n2021 ) | ( n2016 & ~n2021 ) ;
  assign n2023 = ( x73 & n1874 ) | ( x73 & ~n1969 ) | ( n1874 & ~n1969 ) ;
  assign n2024 = x73 & n1874 ;
  assign n2025 = ( ~n1879 & n2023 ) | ( ~n1879 & n2024 ) | ( n2023 & n2024 ) ;
  assign n2026 = ( n1879 & n2023 ) | ( n1879 & n2024 ) | ( n2023 & n2024 ) ;
  assign n2027 = ( n1879 & n2025 ) | ( n1879 & ~n2026 ) | ( n2025 & ~n2026 ) ;
  assign n2028 = ( x74 & n2022 ) | ( x74 & ~n2027 ) | ( n2022 & ~n2027 ) ;
  assign n2029 = ( x74 & n1880 ) | ( x74 & ~n1969 ) | ( n1880 & ~n1969 ) ;
  assign n2030 = x74 & n1880 ;
  assign n2031 = ( n1885 & n2029 ) | ( n1885 & n2030 ) | ( n2029 & n2030 ) ;
  assign n2032 = ( ~n1885 & n2029 ) | ( ~n1885 & n2030 ) | ( n2029 & n2030 ) ;
  assign n2033 = ( n1885 & ~n2031 ) | ( n1885 & n2032 ) | ( ~n2031 & n2032 ) ;
  assign n2034 = ( x75 & n2028 ) | ( x75 & ~n2033 ) | ( n2028 & ~n2033 ) ;
  assign n2035 = ( x75 & n1886 ) | ( x75 & ~n1969 ) | ( n1886 & ~n1969 ) ;
  assign n2036 = x75 & n1886 ;
  assign n2037 = ( ~n1891 & n2035 ) | ( ~n1891 & n2036 ) | ( n2035 & n2036 ) ;
  assign n2038 = ( n1891 & n2035 ) | ( n1891 & n2036 ) | ( n2035 & n2036 ) ;
  assign n2039 = ( n1891 & n2037 ) | ( n1891 & ~n2038 ) | ( n2037 & ~n2038 ) ;
  assign n2040 = ( x76 & n2034 ) | ( x76 & ~n2039 ) | ( n2034 & ~n2039 ) ;
  assign n2041 = ( x76 & n1892 ) | ( x76 & ~n1969 ) | ( n1892 & ~n1969 ) ;
  assign n2042 = x76 & n1892 ;
  assign n2043 = ( n1897 & n2041 ) | ( n1897 & n2042 ) | ( n2041 & n2042 ) ;
  assign n2044 = ( ~n1897 & n2041 ) | ( ~n1897 & n2042 ) | ( n2041 & n2042 ) ;
  assign n2045 = ( n1897 & ~n2043 ) | ( n1897 & n2044 ) | ( ~n2043 & n2044 ) ;
  assign n2046 = ( x77 & n2040 ) | ( x77 & ~n2045 ) | ( n2040 & ~n2045 ) ;
  assign n2047 = ( x77 & n1898 ) | ( x77 & ~n1969 ) | ( n1898 & ~n1969 ) ;
  assign n2048 = x77 & n1898 ;
  assign n2049 = ( ~n1903 & n2047 ) | ( ~n1903 & n2048 ) | ( n2047 & n2048 ) ;
  assign n2050 = ( n1903 & n2047 ) | ( n1903 & n2048 ) | ( n2047 & n2048 ) ;
  assign n2051 = ( n1903 & n2049 ) | ( n1903 & ~n2050 ) | ( n2049 & ~n2050 ) ;
  assign n2052 = ( x78 & n2046 ) | ( x78 & ~n2051 ) | ( n2046 & ~n2051 ) ;
  assign n2053 = ( x78 & n1904 ) | ( x78 & ~n1969 ) | ( n1904 & ~n1969 ) ;
  assign n2054 = x78 & n1904 ;
  assign n2055 = ( n1909 & n2053 ) | ( n1909 & n2054 ) | ( n2053 & n2054 ) ;
  assign n2056 = ( ~n1909 & n2053 ) | ( ~n1909 & n2054 ) | ( n2053 & n2054 ) ;
  assign n2057 = ( n1909 & ~n2055 ) | ( n1909 & n2056 ) | ( ~n2055 & n2056 ) ;
  assign n2058 = ( x79 & n2052 ) | ( x79 & ~n2057 ) | ( n2052 & ~n2057 ) ;
  assign n2059 = ( x79 & n1910 ) | ( x79 & ~n1969 ) | ( n1910 & ~n1969 ) ;
  assign n2060 = x79 & n1910 ;
  assign n2061 = ( ~n1915 & n2059 ) | ( ~n1915 & n2060 ) | ( n2059 & n2060 ) ;
  assign n2062 = ( n1915 & n2059 ) | ( n1915 & n2060 ) | ( n2059 & n2060 ) ;
  assign n2063 = ( n1915 & n2061 ) | ( n1915 & ~n2062 ) | ( n2061 & ~n2062 ) ;
  assign n2064 = ( x80 & n2058 ) | ( x80 & ~n2063 ) | ( n2058 & ~n2063 ) ;
  assign n2065 = ( x80 & n1916 ) | ( x80 & ~n1969 ) | ( n1916 & ~n1969 ) ;
  assign n2066 = x80 & n1916 ;
  assign n2067 = ( n1921 & n2065 ) | ( n1921 & n2066 ) | ( n2065 & n2066 ) ;
  assign n2068 = ( ~n1921 & n2065 ) | ( ~n1921 & n2066 ) | ( n2065 & n2066 ) ;
  assign n2069 = ( n1921 & ~n2067 ) | ( n1921 & n2068 ) | ( ~n2067 & n2068 ) ;
  assign n2070 = ( x81 & n2064 ) | ( x81 & ~n2069 ) | ( n2064 & ~n2069 ) ;
  assign n2071 = ( x81 & n1922 ) | ( x81 & ~n1969 ) | ( n1922 & ~n1969 ) ;
  assign n2072 = x81 & n1922 ;
  assign n2073 = ( ~n1927 & n2071 ) | ( ~n1927 & n2072 ) | ( n2071 & n2072 ) ;
  assign n2074 = ( n1927 & n2071 ) | ( n1927 & n2072 ) | ( n2071 & n2072 ) ;
  assign n2075 = ( n1927 & n2073 ) | ( n1927 & ~n2074 ) | ( n2073 & ~n2074 ) ;
  assign n2076 = ( x82 & n2070 ) | ( x82 & ~n2075 ) | ( n2070 & ~n2075 ) ;
  assign n2077 = ( x82 & n1928 ) | ( x82 & ~n1969 ) | ( n1928 & ~n1969 ) ;
  assign n2078 = x82 & n1928 ;
  assign n2079 = ( n1933 & n2077 ) | ( n1933 & n2078 ) | ( n2077 & n2078 ) ;
  assign n2080 = ( ~n1933 & n2077 ) | ( ~n1933 & n2078 ) | ( n2077 & n2078 ) ;
  assign n2081 = ( n1933 & ~n2079 ) | ( n1933 & n2080 ) | ( ~n2079 & n2080 ) ;
  assign n2082 = ( x83 & n2076 ) | ( x83 & ~n2081 ) | ( n2076 & ~n2081 ) ;
  assign n2083 = ( x83 & n1934 ) | ( x83 & ~n1969 ) | ( n1934 & ~n1969 ) ;
  assign n2084 = x83 & n1934 ;
  assign n2085 = ( ~n1939 & n2083 ) | ( ~n1939 & n2084 ) | ( n2083 & n2084 ) ;
  assign n2086 = ( n1939 & n2083 ) | ( n1939 & n2084 ) | ( n2083 & n2084 ) ;
  assign n2087 = ( n1939 & n2085 ) | ( n1939 & ~n2086 ) | ( n2085 & ~n2086 ) ;
  assign n2088 = ( x84 & n2082 ) | ( x84 & ~n2087 ) | ( n2082 & ~n2087 ) ;
  assign n2089 = ( x84 & n1940 ) | ( x84 & ~n1969 ) | ( n1940 & ~n1969 ) ;
  assign n2090 = x84 & n1940 ;
  assign n2091 = ( n1945 & n2089 ) | ( n1945 & n2090 ) | ( n2089 & n2090 ) ;
  assign n2092 = ( ~n1945 & n2089 ) | ( ~n1945 & n2090 ) | ( n2089 & n2090 ) ;
  assign n2093 = ( n1945 & ~n2091 ) | ( n1945 & n2092 ) | ( ~n2091 & n2092 ) ;
  assign n2094 = ( x85 & n2088 ) | ( x85 & ~n2093 ) | ( n2088 & ~n2093 ) ;
  assign n2095 = ( x85 & n1946 ) | ( x85 & ~n1969 ) | ( n1946 & ~n1969 ) ;
  assign n2096 = x85 & n1946 ;
  assign n2097 = ( ~n1951 & n2095 ) | ( ~n1951 & n2096 ) | ( n2095 & n2096 ) ;
  assign n2098 = ( n1951 & n2095 ) | ( n1951 & n2096 ) | ( n2095 & n2096 ) ;
  assign n2099 = ( n1951 & n2097 ) | ( n1951 & ~n2098 ) | ( n2097 & ~n2098 ) ;
  assign n2100 = ( x86 & n2094 ) | ( x86 & ~n2099 ) | ( n2094 & ~n2099 ) ;
  assign n2101 = ( x86 & n1952 ) | ( x86 & ~n1969 ) | ( n1952 & ~n1969 ) ;
  assign n2102 = x86 & n1952 ;
  assign n2103 = ( n1957 & n2101 ) | ( n1957 & n2102 ) | ( n2101 & n2102 ) ;
  assign n2104 = ( ~n1957 & n2101 ) | ( ~n1957 & n2102 ) | ( n2101 & n2102 ) ;
  assign n2105 = ( n1957 & ~n2103 ) | ( n1957 & n2104 ) | ( ~n2103 & n2104 ) ;
  assign n2106 = ( x87 & n2100 ) | ( x87 & ~n2105 ) | ( n2100 & ~n2105 ) ;
  assign n2107 = ( x87 & n1958 ) | ( x87 & ~n1969 ) | ( n1958 & ~n1969 ) ;
  assign n2108 = x87 & n1958 ;
  assign n2109 = ( n1963 & n2107 ) | ( n1963 & n2108 ) | ( n2107 & n2108 ) ;
  assign n2110 = ( ~n1963 & n2107 ) | ( ~n1963 & n2108 ) | ( n2107 & n2108 ) ;
  assign n2111 = ( n1963 & ~n2109 ) | ( n1963 & n2110 ) | ( ~n2109 & n2110 ) ;
  assign n2112 = ( x88 & n2106 ) | ( x88 & ~n2111 ) | ( n2106 & ~n2111 ) ;
  assign n2113 = x89 & n2112 ;
  assign n2114 = ( x89 & ~n168 ) | ( x89 & n2112 ) | ( ~n168 & n2112 ) ;
  assign n2115 = ( n1967 & n2113 ) | ( n1967 & ~n2114 ) | ( n2113 & ~n2114 ) ;
  assign n2116 = ( x89 & ~n1967 ) | ( x89 & n2112 ) | ( ~n1967 & n2112 ) ;
  assign n2117 = n168 | n2116 ;
  assign n2118 = ( x38 & ~x64 ) | ( x38 & n2117 ) | ( ~x64 & n2117 ) ;
  assign n2119 = ~x38 & n2117 ;
  assign n2120 = ( n1973 & n2118 ) | ( n1973 & ~n2119 ) | ( n2118 & ~n2119 ) ;
  assign n2121 = ~x37 & x64 ;
  assign n2122 = ( x65 & ~n2120 ) | ( x65 & n2121 ) | ( ~n2120 & n2121 ) ;
  assign n2123 = ( x65 & n1973 ) | ( x65 & ~n2117 ) | ( n1973 & ~n2117 ) ;
  assign n2124 = x65 & n1973 ;
  assign n2125 = ( n1972 & n2123 ) | ( n1972 & n2124 ) | ( n2123 & n2124 ) ;
  assign n2126 = ( ~n1972 & n2123 ) | ( ~n1972 & n2124 ) | ( n2123 & n2124 ) ;
  assign n2127 = ( n1972 & ~n2125 ) | ( n1972 & n2126 ) | ( ~n2125 & n2126 ) ;
  assign n2128 = ( x66 & n2122 ) | ( x66 & ~n2127 ) | ( n2122 & ~n2127 ) ;
  assign n2129 = ( x66 & n1974 ) | ( x66 & ~n2117 ) | ( n1974 & ~n2117 ) ;
  assign n2130 = x66 & n1974 ;
  assign n2131 = ( n1979 & n2129 ) | ( n1979 & n2130 ) | ( n2129 & n2130 ) ;
  assign n2132 = ( ~n1979 & n2129 ) | ( ~n1979 & n2130 ) | ( n2129 & n2130 ) ;
  assign n2133 = ( n1979 & ~n2131 ) | ( n1979 & n2132 ) | ( ~n2131 & n2132 ) ;
  assign n2134 = ( x67 & n2128 ) | ( x67 & ~n2133 ) | ( n2128 & ~n2133 ) ;
  assign n2135 = ( x67 & n1980 ) | ( x67 & ~n2117 ) | ( n1980 & ~n2117 ) ;
  assign n2136 = x67 & n1980 ;
  assign n2137 = ( ~n1985 & n2135 ) | ( ~n1985 & n2136 ) | ( n2135 & n2136 ) ;
  assign n2138 = ( n1985 & n2135 ) | ( n1985 & n2136 ) | ( n2135 & n2136 ) ;
  assign n2139 = ( n1985 & n2137 ) | ( n1985 & ~n2138 ) | ( n2137 & ~n2138 ) ;
  assign n2140 = ( x68 & n2134 ) | ( x68 & ~n2139 ) | ( n2134 & ~n2139 ) ;
  assign n2141 = ( x68 & n1986 ) | ( x68 & ~n2117 ) | ( n1986 & ~n2117 ) ;
  assign n2142 = x68 & n1986 ;
  assign n2143 = ( n1991 & n2141 ) | ( n1991 & n2142 ) | ( n2141 & n2142 ) ;
  assign n2144 = ( ~n1991 & n2141 ) | ( ~n1991 & n2142 ) | ( n2141 & n2142 ) ;
  assign n2145 = ( n1991 & ~n2143 ) | ( n1991 & n2144 ) | ( ~n2143 & n2144 ) ;
  assign n2146 = ( x69 & n2140 ) | ( x69 & ~n2145 ) | ( n2140 & ~n2145 ) ;
  assign n2147 = ( x69 & n1992 ) | ( x69 & ~n2117 ) | ( n1992 & ~n2117 ) ;
  assign n2148 = x69 & n1992 ;
  assign n2149 = ( ~n1997 & n2147 ) | ( ~n1997 & n2148 ) | ( n2147 & n2148 ) ;
  assign n2150 = ( n1997 & n2147 ) | ( n1997 & n2148 ) | ( n2147 & n2148 ) ;
  assign n2151 = ( n1997 & n2149 ) | ( n1997 & ~n2150 ) | ( n2149 & ~n2150 ) ;
  assign n2152 = ( x70 & n2146 ) | ( x70 & ~n2151 ) | ( n2146 & ~n2151 ) ;
  assign n2153 = ( x70 & n1998 ) | ( x70 & ~n2117 ) | ( n1998 & ~n2117 ) ;
  assign n2154 = x70 & n1998 ;
  assign n2155 = ( n2003 & n2153 ) | ( n2003 & n2154 ) | ( n2153 & n2154 ) ;
  assign n2156 = ( ~n2003 & n2153 ) | ( ~n2003 & n2154 ) | ( n2153 & n2154 ) ;
  assign n2157 = ( n2003 & ~n2155 ) | ( n2003 & n2156 ) | ( ~n2155 & n2156 ) ;
  assign n2158 = ( x71 & n2152 ) | ( x71 & ~n2157 ) | ( n2152 & ~n2157 ) ;
  assign n2159 = ( x71 & n2004 ) | ( x71 & ~n2117 ) | ( n2004 & ~n2117 ) ;
  assign n2160 = x71 & n2004 ;
  assign n2161 = ( ~n2009 & n2159 ) | ( ~n2009 & n2160 ) | ( n2159 & n2160 ) ;
  assign n2162 = ( n2009 & n2159 ) | ( n2009 & n2160 ) | ( n2159 & n2160 ) ;
  assign n2163 = ( n2009 & n2161 ) | ( n2009 & ~n2162 ) | ( n2161 & ~n2162 ) ;
  assign n2164 = ( x72 & n2158 ) | ( x72 & ~n2163 ) | ( n2158 & ~n2163 ) ;
  assign n2165 = ( x72 & n2010 ) | ( x72 & ~n2117 ) | ( n2010 & ~n2117 ) ;
  assign n2166 = x72 & n2010 ;
  assign n2167 = ( n2015 & n2165 ) | ( n2015 & n2166 ) | ( n2165 & n2166 ) ;
  assign n2168 = ( ~n2015 & n2165 ) | ( ~n2015 & n2166 ) | ( n2165 & n2166 ) ;
  assign n2169 = ( n2015 & ~n2167 ) | ( n2015 & n2168 ) | ( ~n2167 & n2168 ) ;
  assign n2170 = ( x73 & n2164 ) | ( x73 & ~n2169 ) | ( n2164 & ~n2169 ) ;
  assign n2171 = ( x73 & n2016 ) | ( x73 & ~n2117 ) | ( n2016 & ~n2117 ) ;
  assign n2172 = x73 & n2016 ;
  assign n2173 = ( ~n2021 & n2171 ) | ( ~n2021 & n2172 ) | ( n2171 & n2172 ) ;
  assign n2174 = ( n2021 & n2171 ) | ( n2021 & n2172 ) | ( n2171 & n2172 ) ;
  assign n2175 = ( n2021 & n2173 ) | ( n2021 & ~n2174 ) | ( n2173 & ~n2174 ) ;
  assign n2176 = ( x74 & n2170 ) | ( x74 & ~n2175 ) | ( n2170 & ~n2175 ) ;
  assign n2177 = ( x74 & n2022 ) | ( x74 & ~n2117 ) | ( n2022 & ~n2117 ) ;
  assign n2178 = x74 & n2022 ;
  assign n2179 = ( n2027 & n2177 ) | ( n2027 & n2178 ) | ( n2177 & n2178 ) ;
  assign n2180 = ( ~n2027 & n2177 ) | ( ~n2027 & n2178 ) | ( n2177 & n2178 ) ;
  assign n2181 = ( n2027 & ~n2179 ) | ( n2027 & n2180 ) | ( ~n2179 & n2180 ) ;
  assign n2182 = ( x75 & n2176 ) | ( x75 & ~n2181 ) | ( n2176 & ~n2181 ) ;
  assign n2183 = ( x75 & n2028 ) | ( x75 & ~n2117 ) | ( n2028 & ~n2117 ) ;
  assign n2184 = x75 & n2028 ;
  assign n2185 = ( ~n2033 & n2183 ) | ( ~n2033 & n2184 ) | ( n2183 & n2184 ) ;
  assign n2186 = ( n2033 & n2183 ) | ( n2033 & n2184 ) | ( n2183 & n2184 ) ;
  assign n2187 = ( n2033 & n2185 ) | ( n2033 & ~n2186 ) | ( n2185 & ~n2186 ) ;
  assign n2188 = ( x76 & n2182 ) | ( x76 & ~n2187 ) | ( n2182 & ~n2187 ) ;
  assign n2189 = ( x76 & n2034 ) | ( x76 & ~n2117 ) | ( n2034 & ~n2117 ) ;
  assign n2190 = x76 & n2034 ;
  assign n2191 = ( n2039 & n2189 ) | ( n2039 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2192 = ( ~n2039 & n2189 ) | ( ~n2039 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2193 = ( n2039 & ~n2191 ) | ( n2039 & n2192 ) | ( ~n2191 & n2192 ) ;
  assign n2194 = ( x77 & n2188 ) | ( x77 & ~n2193 ) | ( n2188 & ~n2193 ) ;
  assign n2195 = ( x77 & n2040 ) | ( x77 & ~n2117 ) | ( n2040 & ~n2117 ) ;
  assign n2196 = x77 & n2040 ;
  assign n2197 = ( ~n2045 & n2195 ) | ( ~n2045 & n2196 ) | ( n2195 & n2196 ) ;
  assign n2198 = ( n2045 & n2195 ) | ( n2045 & n2196 ) | ( n2195 & n2196 ) ;
  assign n2199 = ( n2045 & n2197 ) | ( n2045 & ~n2198 ) | ( n2197 & ~n2198 ) ;
  assign n2200 = ( x78 & n2194 ) | ( x78 & ~n2199 ) | ( n2194 & ~n2199 ) ;
  assign n2201 = ( x78 & n2046 ) | ( x78 & ~n2117 ) | ( n2046 & ~n2117 ) ;
  assign n2202 = x78 & n2046 ;
  assign n2203 = ( n2051 & n2201 ) | ( n2051 & n2202 ) | ( n2201 & n2202 ) ;
  assign n2204 = ( ~n2051 & n2201 ) | ( ~n2051 & n2202 ) | ( n2201 & n2202 ) ;
  assign n2205 = ( n2051 & ~n2203 ) | ( n2051 & n2204 ) | ( ~n2203 & n2204 ) ;
  assign n2206 = ( x79 & n2200 ) | ( x79 & ~n2205 ) | ( n2200 & ~n2205 ) ;
  assign n2207 = ( x79 & n2052 ) | ( x79 & ~n2117 ) | ( n2052 & ~n2117 ) ;
  assign n2208 = x79 & n2052 ;
  assign n2209 = ( ~n2057 & n2207 ) | ( ~n2057 & n2208 ) | ( n2207 & n2208 ) ;
  assign n2210 = ( n2057 & n2207 ) | ( n2057 & n2208 ) | ( n2207 & n2208 ) ;
  assign n2211 = ( n2057 & n2209 ) | ( n2057 & ~n2210 ) | ( n2209 & ~n2210 ) ;
  assign n2212 = ( x80 & n2206 ) | ( x80 & ~n2211 ) | ( n2206 & ~n2211 ) ;
  assign n2213 = ( x80 & n2058 ) | ( x80 & ~n2117 ) | ( n2058 & ~n2117 ) ;
  assign n2214 = x80 & n2058 ;
  assign n2215 = ( n2063 & n2213 ) | ( n2063 & n2214 ) | ( n2213 & n2214 ) ;
  assign n2216 = ( ~n2063 & n2213 ) | ( ~n2063 & n2214 ) | ( n2213 & n2214 ) ;
  assign n2217 = ( n2063 & ~n2215 ) | ( n2063 & n2216 ) | ( ~n2215 & n2216 ) ;
  assign n2218 = ( x81 & n2212 ) | ( x81 & ~n2217 ) | ( n2212 & ~n2217 ) ;
  assign n2219 = ( x81 & n2064 ) | ( x81 & ~n2117 ) | ( n2064 & ~n2117 ) ;
  assign n2220 = x81 & n2064 ;
  assign n2221 = ( ~n2069 & n2219 ) | ( ~n2069 & n2220 ) | ( n2219 & n2220 ) ;
  assign n2222 = ( n2069 & n2219 ) | ( n2069 & n2220 ) | ( n2219 & n2220 ) ;
  assign n2223 = ( n2069 & n2221 ) | ( n2069 & ~n2222 ) | ( n2221 & ~n2222 ) ;
  assign n2224 = ( x82 & n2218 ) | ( x82 & ~n2223 ) | ( n2218 & ~n2223 ) ;
  assign n2225 = ( x82 & n2070 ) | ( x82 & ~n2117 ) | ( n2070 & ~n2117 ) ;
  assign n2226 = x82 & n2070 ;
  assign n2227 = ( n2075 & n2225 ) | ( n2075 & n2226 ) | ( n2225 & n2226 ) ;
  assign n2228 = ( ~n2075 & n2225 ) | ( ~n2075 & n2226 ) | ( n2225 & n2226 ) ;
  assign n2229 = ( n2075 & ~n2227 ) | ( n2075 & n2228 ) | ( ~n2227 & n2228 ) ;
  assign n2230 = ( x83 & n2224 ) | ( x83 & ~n2229 ) | ( n2224 & ~n2229 ) ;
  assign n2231 = ( x83 & n2076 ) | ( x83 & ~n2117 ) | ( n2076 & ~n2117 ) ;
  assign n2232 = x83 & n2076 ;
  assign n2233 = ( ~n2081 & n2231 ) | ( ~n2081 & n2232 ) | ( n2231 & n2232 ) ;
  assign n2234 = ( n2081 & n2231 ) | ( n2081 & n2232 ) | ( n2231 & n2232 ) ;
  assign n2235 = ( n2081 & n2233 ) | ( n2081 & ~n2234 ) | ( n2233 & ~n2234 ) ;
  assign n2236 = ( x84 & n2230 ) | ( x84 & ~n2235 ) | ( n2230 & ~n2235 ) ;
  assign n2237 = ( x84 & n2082 ) | ( x84 & ~n2117 ) | ( n2082 & ~n2117 ) ;
  assign n2238 = x84 & n2082 ;
  assign n2239 = ( n2087 & n2237 ) | ( n2087 & n2238 ) | ( n2237 & n2238 ) ;
  assign n2240 = ( ~n2087 & n2237 ) | ( ~n2087 & n2238 ) | ( n2237 & n2238 ) ;
  assign n2241 = ( n2087 & ~n2239 ) | ( n2087 & n2240 ) | ( ~n2239 & n2240 ) ;
  assign n2242 = ( x85 & n2236 ) | ( x85 & ~n2241 ) | ( n2236 & ~n2241 ) ;
  assign n2243 = ( x85 & n2088 ) | ( x85 & ~n2117 ) | ( n2088 & ~n2117 ) ;
  assign n2244 = x85 & n2088 ;
  assign n2245 = ( ~n2093 & n2243 ) | ( ~n2093 & n2244 ) | ( n2243 & n2244 ) ;
  assign n2246 = ( n2093 & n2243 ) | ( n2093 & n2244 ) | ( n2243 & n2244 ) ;
  assign n2247 = ( n2093 & n2245 ) | ( n2093 & ~n2246 ) | ( n2245 & ~n2246 ) ;
  assign n2248 = ( x86 & n2242 ) | ( x86 & ~n2247 ) | ( n2242 & ~n2247 ) ;
  assign n2249 = ( x86 & n2094 ) | ( x86 & ~n2117 ) | ( n2094 & ~n2117 ) ;
  assign n2250 = x86 & n2094 ;
  assign n2251 = ( n2099 & n2249 ) | ( n2099 & n2250 ) | ( n2249 & n2250 ) ;
  assign n2252 = ( ~n2099 & n2249 ) | ( ~n2099 & n2250 ) | ( n2249 & n2250 ) ;
  assign n2253 = ( n2099 & ~n2251 ) | ( n2099 & n2252 ) | ( ~n2251 & n2252 ) ;
  assign n2254 = ( x87 & n2248 ) | ( x87 & ~n2253 ) | ( n2248 & ~n2253 ) ;
  assign n2255 = ( x87 & n2100 ) | ( x87 & ~n2117 ) | ( n2100 & ~n2117 ) ;
  assign n2256 = x87 & n2100 ;
  assign n2257 = ( ~n2105 & n2255 ) | ( ~n2105 & n2256 ) | ( n2255 & n2256 ) ;
  assign n2258 = ( n2105 & n2255 ) | ( n2105 & n2256 ) | ( n2255 & n2256 ) ;
  assign n2259 = ( n2105 & n2257 ) | ( n2105 & ~n2258 ) | ( n2257 & ~n2258 ) ;
  assign n2260 = ( x88 & n2254 ) | ( x88 & ~n2259 ) | ( n2254 & ~n2259 ) ;
  assign n2261 = ( x88 & n2106 ) | ( x88 & ~n2117 ) | ( n2106 & ~n2117 ) ;
  assign n2262 = x88 & n2106 ;
  assign n2263 = ( ~n2111 & n2261 ) | ( ~n2111 & n2262 ) | ( n2261 & n2262 ) ;
  assign n2264 = ( n2111 & n2261 ) | ( n2111 & n2262 ) | ( n2261 & n2262 ) ;
  assign n2265 = ( n2111 & n2263 ) | ( n2111 & ~n2264 ) | ( n2263 & ~n2264 ) ;
  assign n2266 = ( x89 & n2260 ) | ( x89 & ~n2265 ) | ( n2260 & ~n2265 ) ;
  assign n2267 = x90 & n2266 ;
  assign n2268 = ( x90 & ~n167 ) | ( x90 & n2266 ) | ( ~n167 & n2266 ) ;
  assign n2269 = ( n2115 & n2267 ) | ( n2115 & ~n2268 ) | ( n2267 & ~n2268 ) ;
  assign n2270 = ( x90 & ~n2115 ) | ( x90 & n2266 ) | ( ~n2115 & n2266 ) ;
  assign n2271 = n167 | n2270 ;
  assign n2272 = ( x37 & ~x64 ) | ( x37 & n2271 ) | ( ~x64 & n2271 ) ;
  assign n2273 = ~x37 & n2271 ;
  assign n2274 = ( n2121 & n2272 ) | ( n2121 & ~n2273 ) | ( n2272 & ~n2273 ) ;
  assign n2275 = ~x36 & x64 ;
  assign n2276 = ( x65 & ~n2274 ) | ( x65 & n2275 ) | ( ~n2274 & n2275 ) ;
  assign n2277 = ( x65 & n2121 ) | ( x65 & ~n2271 ) | ( n2121 & ~n2271 ) ;
  assign n2278 = x65 & n2121 ;
  assign n2279 = ( n2120 & n2277 ) | ( n2120 & n2278 ) | ( n2277 & n2278 ) ;
  assign n2280 = ( ~n2120 & n2277 ) | ( ~n2120 & n2278 ) | ( n2277 & n2278 ) ;
  assign n2281 = ( n2120 & ~n2279 ) | ( n2120 & n2280 ) | ( ~n2279 & n2280 ) ;
  assign n2282 = ( x66 & n2276 ) | ( x66 & ~n2281 ) | ( n2276 & ~n2281 ) ;
  assign n2283 = ( x66 & n2122 ) | ( x66 & ~n2271 ) | ( n2122 & ~n2271 ) ;
  assign n2284 = x66 & n2122 ;
  assign n2285 = ( n2127 & n2283 ) | ( n2127 & n2284 ) | ( n2283 & n2284 ) ;
  assign n2286 = ( ~n2127 & n2283 ) | ( ~n2127 & n2284 ) | ( n2283 & n2284 ) ;
  assign n2287 = ( n2127 & ~n2285 ) | ( n2127 & n2286 ) | ( ~n2285 & n2286 ) ;
  assign n2288 = ( x67 & n2282 ) | ( x67 & ~n2287 ) | ( n2282 & ~n2287 ) ;
  assign n2289 = ( x67 & n2128 ) | ( x67 & ~n2271 ) | ( n2128 & ~n2271 ) ;
  assign n2290 = x67 & n2128 ;
  assign n2291 = ( ~n2133 & n2289 ) | ( ~n2133 & n2290 ) | ( n2289 & n2290 ) ;
  assign n2292 = ( n2133 & n2289 ) | ( n2133 & n2290 ) | ( n2289 & n2290 ) ;
  assign n2293 = ( n2133 & n2291 ) | ( n2133 & ~n2292 ) | ( n2291 & ~n2292 ) ;
  assign n2294 = ( x68 & n2288 ) | ( x68 & ~n2293 ) | ( n2288 & ~n2293 ) ;
  assign n2295 = ( x68 & n2134 ) | ( x68 & ~n2271 ) | ( n2134 & ~n2271 ) ;
  assign n2296 = x68 & n2134 ;
  assign n2297 = ( n2139 & n2295 ) | ( n2139 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2298 = ( ~n2139 & n2295 ) | ( ~n2139 & n2296 ) | ( n2295 & n2296 ) ;
  assign n2299 = ( n2139 & ~n2297 ) | ( n2139 & n2298 ) | ( ~n2297 & n2298 ) ;
  assign n2300 = ( x69 & n2294 ) | ( x69 & ~n2299 ) | ( n2294 & ~n2299 ) ;
  assign n2301 = ( x69 & n2140 ) | ( x69 & ~n2271 ) | ( n2140 & ~n2271 ) ;
  assign n2302 = x69 & n2140 ;
  assign n2303 = ( ~n2145 & n2301 ) | ( ~n2145 & n2302 ) | ( n2301 & n2302 ) ;
  assign n2304 = ( n2145 & n2301 ) | ( n2145 & n2302 ) | ( n2301 & n2302 ) ;
  assign n2305 = ( n2145 & n2303 ) | ( n2145 & ~n2304 ) | ( n2303 & ~n2304 ) ;
  assign n2306 = ( x70 & n2300 ) | ( x70 & ~n2305 ) | ( n2300 & ~n2305 ) ;
  assign n2307 = ( x70 & n2146 ) | ( x70 & ~n2271 ) | ( n2146 & ~n2271 ) ;
  assign n2308 = x70 & n2146 ;
  assign n2309 = ( n2151 & n2307 ) | ( n2151 & n2308 ) | ( n2307 & n2308 ) ;
  assign n2310 = ( ~n2151 & n2307 ) | ( ~n2151 & n2308 ) | ( n2307 & n2308 ) ;
  assign n2311 = ( n2151 & ~n2309 ) | ( n2151 & n2310 ) | ( ~n2309 & n2310 ) ;
  assign n2312 = ( x71 & n2306 ) | ( x71 & ~n2311 ) | ( n2306 & ~n2311 ) ;
  assign n2313 = ( x71 & n2152 ) | ( x71 & ~n2271 ) | ( n2152 & ~n2271 ) ;
  assign n2314 = x71 & n2152 ;
  assign n2315 = ( ~n2157 & n2313 ) | ( ~n2157 & n2314 ) | ( n2313 & n2314 ) ;
  assign n2316 = ( n2157 & n2313 ) | ( n2157 & n2314 ) | ( n2313 & n2314 ) ;
  assign n2317 = ( n2157 & n2315 ) | ( n2157 & ~n2316 ) | ( n2315 & ~n2316 ) ;
  assign n2318 = ( x72 & n2312 ) | ( x72 & ~n2317 ) | ( n2312 & ~n2317 ) ;
  assign n2319 = ( x72 & n2158 ) | ( x72 & ~n2271 ) | ( n2158 & ~n2271 ) ;
  assign n2320 = x72 & n2158 ;
  assign n2321 = ( n2163 & n2319 ) | ( n2163 & n2320 ) | ( n2319 & n2320 ) ;
  assign n2322 = ( ~n2163 & n2319 ) | ( ~n2163 & n2320 ) | ( n2319 & n2320 ) ;
  assign n2323 = ( n2163 & ~n2321 ) | ( n2163 & n2322 ) | ( ~n2321 & n2322 ) ;
  assign n2324 = ( x73 & n2318 ) | ( x73 & ~n2323 ) | ( n2318 & ~n2323 ) ;
  assign n2325 = ( x73 & n2164 ) | ( x73 & ~n2271 ) | ( n2164 & ~n2271 ) ;
  assign n2326 = x73 & n2164 ;
  assign n2327 = ( ~n2169 & n2325 ) | ( ~n2169 & n2326 ) | ( n2325 & n2326 ) ;
  assign n2328 = ( n2169 & n2325 ) | ( n2169 & n2326 ) | ( n2325 & n2326 ) ;
  assign n2329 = ( n2169 & n2327 ) | ( n2169 & ~n2328 ) | ( n2327 & ~n2328 ) ;
  assign n2330 = ( x74 & n2324 ) | ( x74 & ~n2329 ) | ( n2324 & ~n2329 ) ;
  assign n2331 = ( x74 & n2170 ) | ( x74 & ~n2271 ) | ( n2170 & ~n2271 ) ;
  assign n2332 = x74 & n2170 ;
  assign n2333 = ( n2175 & n2331 ) | ( n2175 & n2332 ) | ( n2331 & n2332 ) ;
  assign n2334 = ( ~n2175 & n2331 ) | ( ~n2175 & n2332 ) | ( n2331 & n2332 ) ;
  assign n2335 = ( n2175 & ~n2333 ) | ( n2175 & n2334 ) | ( ~n2333 & n2334 ) ;
  assign n2336 = ( x75 & n2330 ) | ( x75 & ~n2335 ) | ( n2330 & ~n2335 ) ;
  assign n2337 = ( x75 & n2176 ) | ( x75 & ~n2271 ) | ( n2176 & ~n2271 ) ;
  assign n2338 = x75 & n2176 ;
  assign n2339 = ( ~n2181 & n2337 ) | ( ~n2181 & n2338 ) | ( n2337 & n2338 ) ;
  assign n2340 = ( n2181 & n2337 ) | ( n2181 & n2338 ) | ( n2337 & n2338 ) ;
  assign n2341 = ( n2181 & n2339 ) | ( n2181 & ~n2340 ) | ( n2339 & ~n2340 ) ;
  assign n2342 = ( x76 & n2336 ) | ( x76 & ~n2341 ) | ( n2336 & ~n2341 ) ;
  assign n2343 = ( x76 & n2182 ) | ( x76 & ~n2271 ) | ( n2182 & ~n2271 ) ;
  assign n2344 = x76 & n2182 ;
  assign n2345 = ( n2187 & n2343 ) | ( n2187 & n2344 ) | ( n2343 & n2344 ) ;
  assign n2346 = ( ~n2187 & n2343 ) | ( ~n2187 & n2344 ) | ( n2343 & n2344 ) ;
  assign n2347 = ( n2187 & ~n2345 ) | ( n2187 & n2346 ) | ( ~n2345 & n2346 ) ;
  assign n2348 = ( x77 & n2342 ) | ( x77 & ~n2347 ) | ( n2342 & ~n2347 ) ;
  assign n2349 = ( x77 & n2188 ) | ( x77 & ~n2271 ) | ( n2188 & ~n2271 ) ;
  assign n2350 = x77 & n2188 ;
  assign n2351 = ( ~n2193 & n2349 ) | ( ~n2193 & n2350 ) | ( n2349 & n2350 ) ;
  assign n2352 = ( n2193 & n2349 ) | ( n2193 & n2350 ) | ( n2349 & n2350 ) ;
  assign n2353 = ( n2193 & n2351 ) | ( n2193 & ~n2352 ) | ( n2351 & ~n2352 ) ;
  assign n2354 = ( x78 & n2348 ) | ( x78 & ~n2353 ) | ( n2348 & ~n2353 ) ;
  assign n2355 = ( x78 & n2194 ) | ( x78 & ~n2271 ) | ( n2194 & ~n2271 ) ;
  assign n2356 = x78 & n2194 ;
  assign n2357 = ( n2199 & n2355 ) | ( n2199 & n2356 ) | ( n2355 & n2356 ) ;
  assign n2358 = ( ~n2199 & n2355 ) | ( ~n2199 & n2356 ) | ( n2355 & n2356 ) ;
  assign n2359 = ( n2199 & ~n2357 ) | ( n2199 & n2358 ) | ( ~n2357 & n2358 ) ;
  assign n2360 = ( x79 & n2354 ) | ( x79 & ~n2359 ) | ( n2354 & ~n2359 ) ;
  assign n2361 = ( x79 & n2200 ) | ( x79 & ~n2271 ) | ( n2200 & ~n2271 ) ;
  assign n2362 = x79 & n2200 ;
  assign n2363 = ( ~n2205 & n2361 ) | ( ~n2205 & n2362 ) | ( n2361 & n2362 ) ;
  assign n2364 = ( n2205 & n2361 ) | ( n2205 & n2362 ) | ( n2361 & n2362 ) ;
  assign n2365 = ( n2205 & n2363 ) | ( n2205 & ~n2364 ) | ( n2363 & ~n2364 ) ;
  assign n2366 = ( x80 & n2360 ) | ( x80 & ~n2365 ) | ( n2360 & ~n2365 ) ;
  assign n2367 = ( x80 & n2206 ) | ( x80 & ~n2271 ) | ( n2206 & ~n2271 ) ;
  assign n2368 = x80 & n2206 ;
  assign n2369 = ( n2211 & n2367 ) | ( n2211 & n2368 ) | ( n2367 & n2368 ) ;
  assign n2370 = ( ~n2211 & n2367 ) | ( ~n2211 & n2368 ) | ( n2367 & n2368 ) ;
  assign n2371 = ( n2211 & ~n2369 ) | ( n2211 & n2370 ) | ( ~n2369 & n2370 ) ;
  assign n2372 = ( x81 & n2366 ) | ( x81 & ~n2371 ) | ( n2366 & ~n2371 ) ;
  assign n2373 = ( x81 & n2212 ) | ( x81 & ~n2271 ) | ( n2212 & ~n2271 ) ;
  assign n2374 = x81 & n2212 ;
  assign n2375 = ( ~n2217 & n2373 ) | ( ~n2217 & n2374 ) | ( n2373 & n2374 ) ;
  assign n2376 = ( n2217 & n2373 ) | ( n2217 & n2374 ) | ( n2373 & n2374 ) ;
  assign n2377 = ( n2217 & n2375 ) | ( n2217 & ~n2376 ) | ( n2375 & ~n2376 ) ;
  assign n2378 = ( x82 & n2372 ) | ( x82 & ~n2377 ) | ( n2372 & ~n2377 ) ;
  assign n2379 = ( x82 & n2218 ) | ( x82 & ~n2271 ) | ( n2218 & ~n2271 ) ;
  assign n2380 = x82 & n2218 ;
  assign n2381 = ( n2223 & n2379 ) | ( n2223 & n2380 ) | ( n2379 & n2380 ) ;
  assign n2382 = ( ~n2223 & n2379 ) | ( ~n2223 & n2380 ) | ( n2379 & n2380 ) ;
  assign n2383 = ( n2223 & ~n2381 ) | ( n2223 & n2382 ) | ( ~n2381 & n2382 ) ;
  assign n2384 = ( x83 & n2378 ) | ( x83 & ~n2383 ) | ( n2378 & ~n2383 ) ;
  assign n2385 = ( x83 & n2224 ) | ( x83 & ~n2271 ) | ( n2224 & ~n2271 ) ;
  assign n2386 = x83 & n2224 ;
  assign n2387 = ( ~n2229 & n2385 ) | ( ~n2229 & n2386 ) | ( n2385 & n2386 ) ;
  assign n2388 = ( n2229 & n2385 ) | ( n2229 & n2386 ) | ( n2385 & n2386 ) ;
  assign n2389 = ( n2229 & n2387 ) | ( n2229 & ~n2388 ) | ( n2387 & ~n2388 ) ;
  assign n2390 = ( x84 & n2384 ) | ( x84 & ~n2389 ) | ( n2384 & ~n2389 ) ;
  assign n2391 = ( x84 & n2230 ) | ( x84 & ~n2271 ) | ( n2230 & ~n2271 ) ;
  assign n2392 = x84 & n2230 ;
  assign n2393 = ( n2235 & n2391 ) | ( n2235 & n2392 ) | ( n2391 & n2392 ) ;
  assign n2394 = ( ~n2235 & n2391 ) | ( ~n2235 & n2392 ) | ( n2391 & n2392 ) ;
  assign n2395 = ( n2235 & ~n2393 ) | ( n2235 & n2394 ) | ( ~n2393 & n2394 ) ;
  assign n2396 = ( x85 & n2390 ) | ( x85 & ~n2395 ) | ( n2390 & ~n2395 ) ;
  assign n2397 = ( x85 & n2236 ) | ( x85 & ~n2271 ) | ( n2236 & ~n2271 ) ;
  assign n2398 = x85 & n2236 ;
  assign n2399 = ( ~n2241 & n2397 ) | ( ~n2241 & n2398 ) | ( n2397 & n2398 ) ;
  assign n2400 = ( n2241 & n2397 ) | ( n2241 & n2398 ) | ( n2397 & n2398 ) ;
  assign n2401 = ( n2241 & n2399 ) | ( n2241 & ~n2400 ) | ( n2399 & ~n2400 ) ;
  assign n2402 = ( x86 & n2396 ) | ( x86 & ~n2401 ) | ( n2396 & ~n2401 ) ;
  assign n2403 = ( x86 & n2242 ) | ( x86 & ~n2271 ) | ( n2242 & ~n2271 ) ;
  assign n2404 = x86 & n2242 ;
  assign n2405 = ( n2247 & n2403 ) | ( n2247 & n2404 ) | ( n2403 & n2404 ) ;
  assign n2406 = ( ~n2247 & n2403 ) | ( ~n2247 & n2404 ) | ( n2403 & n2404 ) ;
  assign n2407 = ( n2247 & ~n2405 ) | ( n2247 & n2406 ) | ( ~n2405 & n2406 ) ;
  assign n2408 = ( x87 & n2402 ) | ( x87 & ~n2407 ) | ( n2402 & ~n2407 ) ;
  assign n2409 = ( x87 & n2248 ) | ( x87 & ~n2271 ) | ( n2248 & ~n2271 ) ;
  assign n2410 = x87 & n2248 ;
  assign n2411 = ( ~n2253 & n2409 ) | ( ~n2253 & n2410 ) | ( n2409 & n2410 ) ;
  assign n2412 = ( n2253 & n2409 ) | ( n2253 & n2410 ) | ( n2409 & n2410 ) ;
  assign n2413 = ( n2253 & n2411 ) | ( n2253 & ~n2412 ) | ( n2411 & ~n2412 ) ;
  assign n2414 = ( x88 & n2408 ) | ( x88 & ~n2413 ) | ( n2408 & ~n2413 ) ;
  assign n2415 = ( x88 & n2254 ) | ( x88 & ~n2271 ) | ( n2254 & ~n2271 ) ;
  assign n2416 = x88 & n2254 ;
  assign n2417 = ( n2259 & n2415 ) | ( n2259 & n2416 ) | ( n2415 & n2416 ) ;
  assign n2418 = ( ~n2259 & n2415 ) | ( ~n2259 & n2416 ) | ( n2415 & n2416 ) ;
  assign n2419 = ( n2259 & ~n2417 ) | ( n2259 & n2418 ) | ( ~n2417 & n2418 ) ;
  assign n2420 = ( x89 & n2414 ) | ( x89 & ~n2419 ) | ( n2414 & ~n2419 ) ;
  assign n2421 = ( x89 & n2260 ) | ( x89 & ~n2271 ) | ( n2260 & ~n2271 ) ;
  assign n2422 = x89 & n2260 ;
  assign n2423 = ( n2265 & n2421 ) | ( n2265 & n2422 ) | ( n2421 & n2422 ) ;
  assign n2424 = ( ~n2265 & n2421 ) | ( ~n2265 & n2422 ) | ( n2421 & n2422 ) ;
  assign n2425 = ( n2265 & ~n2423 ) | ( n2265 & n2424 ) | ( ~n2423 & n2424 ) ;
  assign n2426 = ( x90 & n2420 ) | ( x90 & ~n2425 ) | ( n2420 & ~n2425 ) ;
  assign n2427 = x91 | n2426 ;
  assign n2428 = ( x91 & n166 ) | ( x91 & n2426 ) | ( n166 & n2426 ) ;
  assign n2429 = ( n2269 & ~n2427 ) | ( n2269 & n2428 ) | ( ~n2427 & n2428 ) ;
  assign n2430 = ( x91 & ~n2269 ) | ( x91 & n2426 ) | ( ~n2269 & n2426 ) ;
  assign n2431 = n166 | n2430 ;
  assign n2432 = ( x36 & ~x64 ) | ( x36 & n2431 ) | ( ~x64 & n2431 ) ;
  assign n2433 = ~x36 & n2431 ;
  assign n2434 = ( n2275 & n2432 ) | ( n2275 & ~n2433 ) | ( n2432 & ~n2433 ) ;
  assign n2435 = ~x35 & x64 ;
  assign n2436 = ( x65 & ~n2434 ) | ( x65 & n2435 ) | ( ~n2434 & n2435 ) ;
  assign n2437 = ( x65 & n2275 ) | ( x65 & ~n2431 ) | ( n2275 & ~n2431 ) ;
  assign n2438 = x65 & n2275 ;
  assign n2439 = ( n2274 & n2437 ) | ( n2274 & n2438 ) | ( n2437 & n2438 ) ;
  assign n2440 = ( ~n2274 & n2437 ) | ( ~n2274 & n2438 ) | ( n2437 & n2438 ) ;
  assign n2441 = ( n2274 & ~n2439 ) | ( n2274 & n2440 ) | ( ~n2439 & n2440 ) ;
  assign n2442 = ( x66 & n2436 ) | ( x66 & ~n2441 ) | ( n2436 & ~n2441 ) ;
  assign n2443 = ( x66 & n2276 ) | ( x66 & ~n2431 ) | ( n2276 & ~n2431 ) ;
  assign n2444 = x66 & n2276 ;
  assign n2445 = ( n2281 & n2443 ) | ( n2281 & n2444 ) | ( n2443 & n2444 ) ;
  assign n2446 = ( ~n2281 & n2443 ) | ( ~n2281 & n2444 ) | ( n2443 & n2444 ) ;
  assign n2447 = ( n2281 & ~n2445 ) | ( n2281 & n2446 ) | ( ~n2445 & n2446 ) ;
  assign n2448 = ( x67 & n2442 ) | ( x67 & ~n2447 ) | ( n2442 & ~n2447 ) ;
  assign n2449 = ( x67 & n2282 ) | ( x67 & ~n2431 ) | ( n2282 & ~n2431 ) ;
  assign n2450 = x67 & n2282 ;
  assign n2451 = ( ~n2287 & n2449 ) | ( ~n2287 & n2450 ) | ( n2449 & n2450 ) ;
  assign n2452 = ( n2287 & n2449 ) | ( n2287 & n2450 ) | ( n2449 & n2450 ) ;
  assign n2453 = ( n2287 & n2451 ) | ( n2287 & ~n2452 ) | ( n2451 & ~n2452 ) ;
  assign n2454 = ( x68 & n2448 ) | ( x68 & ~n2453 ) | ( n2448 & ~n2453 ) ;
  assign n2455 = ( x68 & n2288 ) | ( x68 & ~n2431 ) | ( n2288 & ~n2431 ) ;
  assign n2456 = x68 & n2288 ;
  assign n2457 = ( n2293 & n2455 ) | ( n2293 & n2456 ) | ( n2455 & n2456 ) ;
  assign n2458 = ( ~n2293 & n2455 ) | ( ~n2293 & n2456 ) | ( n2455 & n2456 ) ;
  assign n2459 = ( n2293 & ~n2457 ) | ( n2293 & n2458 ) | ( ~n2457 & n2458 ) ;
  assign n2460 = ( x69 & n2454 ) | ( x69 & ~n2459 ) | ( n2454 & ~n2459 ) ;
  assign n2461 = ( x69 & n2294 ) | ( x69 & ~n2431 ) | ( n2294 & ~n2431 ) ;
  assign n2462 = x69 & n2294 ;
  assign n2463 = ( ~n2299 & n2461 ) | ( ~n2299 & n2462 ) | ( n2461 & n2462 ) ;
  assign n2464 = ( n2299 & n2461 ) | ( n2299 & n2462 ) | ( n2461 & n2462 ) ;
  assign n2465 = ( n2299 & n2463 ) | ( n2299 & ~n2464 ) | ( n2463 & ~n2464 ) ;
  assign n2466 = ( x70 & n2460 ) | ( x70 & ~n2465 ) | ( n2460 & ~n2465 ) ;
  assign n2467 = ( x70 & n2300 ) | ( x70 & ~n2431 ) | ( n2300 & ~n2431 ) ;
  assign n2468 = x70 & n2300 ;
  assign n2469 = ( n2305 & n2467 ) | ( n2305 & n2468 ) | ( n2467 & n2468 ) ;
  assign n2470 = ( ~n2305 & n2467 ) | ( ~n2305 & n2468 ) | ( n2467 & n2468 ) ;
  assign n2471 = ( n2305 & ~n2469 ) | ( n2305 & n2470 ) | ( ~n2469 & n2470 ) ;
  assign n2472 = ( x71 & n2466 ) | ( x71 & ~n2471 ) | ( n2466 & ~n2471 ) ;
  assign n2473 = ( x71 & n2306 ) | ( x71 & ~n2431 ) | ( n2306 & ~n2431 ) ;
  assign n2474 = x71 & n2306 ;
  assign n2475 = ( ~n2311 & n2473 ) | ( ~n2311 & n2474 ) | ( n2473 & n2474 ) ;
  assign n2476 = ( n2311 & n2473 ) | ( n2311 & n2474 ) | ( n2473 & n2474 ) ;
  assign n2477 = ( n2311 & n2475 ) | ( n2311 & ~n2476 ) | ( n2475 & ~n2476 ) ;
  assign n2478 = ( x72 & n2472 ) | ( x72 & ~n2477 ) | ( n2472 & ~n2477 ) ;
  assign n2479 = ( x72 & n2312 ) | ( x72 & ~n2431 ) | ( n2312 & ~n2431 ) ;
  assign n2480 = x72 & n2312 ;
  assign n2481 = ( n2317 & n2479 ) | ( n2317 & n2480 ) | ( n2479 & n2480 ) ;
  assign n2482 = ( ~n2317 & n2479 ) | ( ~n2317 & n2480 ) | ( n2479 & n2480 ) ;
  assign n2483 = ( n2317 & ~n2481 ) | ( n2317 & n2482 ) | ( ~n2481 & n2482 ) ;
  assign n2484 = ( x73 & n2478 ) | ( x73 & ~n2483 ) | ( n2478 & ~n2483 ) ;
  assign n2485 = ( x73 & n2318 ) | ( x73 & ~n2431 ) | ( n2318 & ~n2431 ) ;
  assign n2486 = x73 & n2318 ;
  assign n2487 = ( ~n2323 & n2485 ) | ( ~n2323 & n2486 ) | ( n2485 & n2486 ) ;
  assign n2488 = ( n2323 & n2485 ) | ( n2323 & n2486 ) | ( n2485 & n2486 ) ;
  assign n2489 = ( n2323 & n2487 ) | ( n2323 & ~n2488 ) | ( n2487 & ~n2488 ) ;
  assign n2490 = ( x74 & n2484 ) | ( x74 & ~n2489 ) | ( n2484 & ~n2489 ) ;
  assign n2491 = ( x74 & n2324 ) | ( x74 & ~n2431 ) | ( n2324 & ~n2431 ) ;
  assign n2492 = x74 & n2324 ;
  assign n2493 = ( n2329 & n2491 ) | ( n2329 & n2492 ) | ( n2491 & n2492 ) ;
  assign n2494 = ( ~n2329 & n2491 ) | ( ~n2329 & n2492 ) | ( n2491 & n2492 ) ;
  assign n2495 = ( n2329 & ~n2493 ) | ( n2329 & n2494 ) | ( ~n2493 & n2494 ) ;
  assign n2496 = ( x75 & n2490 ) | ( x75 & ~n2495 ) | ( n2490 & ~n2495 ) ;
  assign n2497 = ( x75 & n2330 ) | ( x75 & ~n2431 ) | ( n2330 & ~n2431 ) ;
  assign n2498 = x75 & n2330 ;
  assign n2499 = ( ~n2335 & n2497 ) | ( ~n2335 & n2498 ) | ( n2497 & n2498 ) ;
  assign n2500 = ( n2335 & n2497 ) | ( n2335 & n2498 ) | ( n2497 & n2498 ) ;
  assign n2501 = ( n2335 & n2499 ) | ( n2335 & ~n2500 ) | ( n2499 & ~n2500 ) ;
  assign n2502 = ( x76 & n2496 ) | ( x76 & ~n2501 ) | ( n2496 & ~n2501 ) ;
  assign n2503 = ( x76 & n2336 ) | ( x76 & ~n2431 ) | ( n2336 & ~n2431 ) ;
  assign n2504 = x76 & n2336 ;
  assign n2505 = ( n2341 & n2503 ) | ( n2341 & n2504 ) | ( n2503 & n2504 ) ;
  assign n2506 = ( ~n2341 & n2503 ) | ( ~n2341 & n2504 ) | ( n2503 & n2504 ) ;
  assign n2507 = ( n2341 & ~n2505 ) | ( n2341 & n2506 ) | ( ~n2505 & n2506 ) ;
  assign n2508 = ( x77 & n2502 ) | ( x77 & ~n2507 ) | ( n2502 & ~n2507 ) ;
  assign n2509 = ( x77 & n2342 ) | ( x77 & ~n2431 ) | ( n2342 & ~n2431 ) ;
  assign n2510 = x77 & n2342 ;
  assign n2511 = ( ~n2347 & n2509 ) | ( ~n2347 & n2510 ) | ( n2509 & n2510 ) ;
  assign n2512 = ( n2347 & n2509 ) | ( n2347 & n2510 ) | ( n2509 & n2510 ) ;
  assign n2513 = ( n2347 & n2511 ) | ( n2347 & ~n2512 ) | ( n2511 & ~n2512 ) ;
  assign n2514 = ( x78 & n2508 ) | ( x78 & ~n2513 ) | ( n2508 & ~n2513 ) ;
  assign n2515 = ( x78 & n2348 ) | ( x78 & ~n2431 ) | ( n2348 & ~n2431 ) ;
  assign n2516 = x78 & n2348 ;
  assign n2517 = ( n2353 & n2515 ) | ( n2353 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2518 = ( ~n2353 & n2515 ) | ( ~n2353 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2519 = ( n2353 & ~n2517 ) | ( n2353 & n2518 ) | ( ~n2517 & n2518 ) ;
  assign n2520 = ( x79 & n2514 ) | ( x79 & ~n2519 ) | ( n2514 & ~n2519 ) ;
  assign n2521 = ( x79 & n2354 ) | ( x79 & ~n2431 ) | ( n2354 & ~n2431 ) ;
  assign n2522 = x79 & n2354 ;
  assign n2523 = ( ~n2359 & n2521 ) | ( ~n2359 & n2522 ) | ( n2521 & n2522 ) ;
  assign n2524 = ( n2359 & n2521 ) | ( n2359 & n2522 ) | ( n2521 & n2522 ) ;
  assign n2525 = ( n2359 & n2523 ) | ( n2359 & ~n2524 ) | ( n2523 & ~n2524 ) ;
  assign n2526 = ( x80 & n2520 ) | ( x80 & ~n2525 ) | ( n2520 & ~n2525 ) ;
  assign n2527 = ( x80 & n2360 ) | ( x80 & ~n2431 ) | ( n2360 & ~n2431 ) ;
  assign n2528 = x80 & n2360 ;
  assign n2529 = ( n2365 & n2527 ) | ( n2365 & n2528 ) | ( n2527 & n2528 ) ;
  assign n2530 = ( ~n2365 & n2527 ) | ( ~n2365 & n2528 ) | ( n2527 & n2528 ) ;
  assign n2531 = ( n2365 & ~n2529 ) | ( n2365 & n2530 ) | ( ~n2529 & n2530 ) ;
  assign n2532 = ( x81 & n2526 ) | ( x81 & ~n2531 ) | ( n2526 & ~n2531 ) ;
  assign n2533 = ( x81 & n2366 ) | ( x81 & ~n2431 ) | ( n2366 & ~n2431 ) ;
  assign n2534 = x81 & n2366 ;
  assign n2535 = ( ~n2371 & n2533 ) | ( ~n2371 & n2534 ) | ( n2533 & n2534 ) ;
  assign n2536 = ( n2371 & n2533 ) | ( n2371 & n2534 ) | ( n2533 & n2534 ) ;
  assign n2537 = ( n2371 & n2535 ) | ( n2371 & ~n2536 ) | ( n2535 & ~n2536 ) ;
  assign n2538 = ( x82 & n2532 ) | ( x82 & ~n2537 ) | ( n2532 & ~n2537 ) ;
  assign n2539 = ( x82 & n2372 ) | ( x82 & ~n2431 ) | ( n2372 & ~n2431 ) ;
  assign n2540 = x82 & n2372 ;
  assign n2541 = ( n2377 & n2539 ) | ( n2377 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2542 = ( ~n2377 & n2539 ) | ( ~n2377 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2543 = ( n2377 & ~n2541 ) | ( n2377 & n2542 ) | ( ~n2541 & n2542 ) ;
  assign n2544 = ( x83 & n2538 ) | ( x83 & ~n2543 ) | ( n2538 & ~n2543 ) ;
  assign n2545 = ( x83 & n2378 ) | ( x83 & ~n2431 ) | ( n2378 & ~n2431 ) ;
  assign n2546 = x83 & n2378 ;
  assign n2547 = ( ~n2383 & n2545 ) | ( ~n2383 & n2546 ) | ( n2545 & n2546 ) ;
  assign n2548 = ( n2383 & n2545 ) | ( n2383 & n2546 ) | ( n2545 & n2546 ) ;
  assign n2549 = ( n2383 & n2547 ) | ( n2383 & ~n2548 ) | ( n2547 & ~n2548 ) ;
  assign n2550 = ( x84 & n2544 ) | ( x84 & ~n2549 ) | ( n2544 & ~n2549 ) ;
  assign n2551 = ( x84 & n2384 ) | ( x84 & ~n2431 ) | ( n2384 & ~n2431 ) ;
  assign n2552 = x84 & n2384 ;
  assign n2553 = ( n2389 & n2551 ) | ( n2389 & n2552 ) | ( n2551 & n2552 ) ;
  assign n2554 = ( ~n2389 & n2551 ) | ( ~n2389 & n2552 ) | ( n2551 & n2552 ) ;
  assign n2555 = ( n2389 & ~n2553 ) | ( n2389 & n2554 ) | ( ~n2553 & n2554 ) ;
  assign n2556 = ( x85 & n2550 ) | ( x85 & ~n2555 ) | ( n2550 & ~n2555 ) ;
  assign n2557 = ( x85 & n2390 ) | ( x85 & ~n2431 ) | ( n2390 & ~n2431 ) ;
  assign n2558 = x85 & n2390 ;
  assign n2559 = ( ~n2395 & n2557 ) | ( ~n2395 & n2558 ) | ( n2557 & n2558 ) ;
  assign n2560 = ( n2395 & n2557 ) | ( n2395 & n2558 ) | ( n2557 & n2558 ) ;
  assign n2561 = ( n2395 & n2559 ) | ( n2395 & ~n2560 ) | ( n2559 & ~n2560 ) ;
  assign n2562 = ( x86 & n2556 ) | ( x86 & ~n2561 ) | ( n2556 & ~n2561 ) ;
  assign n2563 = ( x86 & n2396 ) | ( x86 & ~n2431 ) | ( n2396 & ~n2431 ) ;
  assign n2564 = x86 & n2396 ;
  assign n2565 = ( n2401 & n2563 ) | ( n2401 & n2564 ) | ( n2563 & n2564 ) ;
  assign n2566 = ( ~n2401 & n2563 ) | ( ~n2401 & n2564 ) | ( n2563 & n2564 ) ;
  assign n2567 = ( n2401 & ~n2565 ) | ( n2401 & n2566 ) | ( ~n2565 & n2566 ) ;
  assign n2568 = ( x87 & n2562 ) | ( x87 & ~n2567 ) | ( n2562 & ~n2567 ) ;
  assign n2569 = ( x87 & n2402 ) | ( x87 & ~n2431 ) | ( n2402 & ~n2431 ) ;
  assign n2570 = x87 & n2402 ;
  assign n2571 = ( ~n2407 & n2569 ) | ( ~n2407 & n2570 ) | ( n2569 & n2570 ) ;
  assign n2572 = ( n2407 & n2569 ) | ( n2407 & n2570 ) | ( n2569 & n2570 ) ;
  assign n2573 = ( n2407 & n2571 ) | ( n2407 & ~n2572 ) | ( n2571 & ~n2572 ) ;
  assign n2574 = ( x88 & n2568 ) | ( x88 & ~n2573 ) | ( n2568 & ~n2573 ) ;
  assign n2575 = ( x88 & n2408 ) | ( x88 & ~n2431 ) | ( n2408 & ~n2431 ) ;
  assign n2576 = x88 & n2408 ;
  assign n2577 = ( n2413 & n2575 ) | ( n2413 & n2576 ) | ( n2575 & n2576 ) ;
  assign n2578 = ( ~n2413 & n2575 ) | ( ~n2413 & n2576 ) | ( n2575 & n2576 ) ;
  assign n2579 = ( n2413 & ~n2577 ) | ( n2413 & n2578 ) | ( ~n2577 & n2578 ) ;
  assign n2580 = ( x89 & n2574 ) | ( x89 & ~n2579 ) | ( n2574 & ~n2579 ) ;
  assign n2581 = ( x89 & n2414 ) | ( x89 & ~n2431 ) | ( n2414 & ~n2431 ) ;
  assign n2582 = x89 & n2414 ;
  assign n2583 = ( ~n2419 & n2581 ) | ( ~n2419 & n2582 ) | ( n2581 & n2582 ) ;
  assign n2584 = ( n2419 & n2581 ) | ( n2419 & n2582 ) | ( n2581 & n2582 ) ;
  assign n2585 = ( n2419 & n2583 ) | ( n2419 & ~n2584 ) | ( n2583 & ~n2584 ) ;
  assign n2586 = ( x90 & n2580 ) | ( x90 & ~n2585 ) | ( n2580 & ~n2585 ) ;
  assign n2587 = ( x90 & n2420 ) | ( x90 & ~n2431 ) | ( n2420 & ~n2431 ) ;
  assign n2588 = x90 & n2420 ;
  assign n2589 = ( ~n2425 & n2587 ) | ( ~n2425 & n2588 ) | ( n2587 & n2588 ) ;
  assign n2590 = ( n2425 & n2587 ) | ( n2425 & n2588 ) | ( n2587 & n2588 ) ;
  assign n2591 = ( n2425 & n2589 ) | ( n2425 & ~n2590 ) | ( n2589 & ~n2590 ) ;
  assign n2592 = ( x91 & n2586 ) | ( x91 & ~n2591 ) | ( n2586 & ~n2591 ) ;
  assign n2593 = x92 | n2592 ;
  assign n2594 = ( x92 & n165 ) | ( x92 & n2592 ) | ( n165 & n2592 ) ;
  assign n2595 = ( n2429 & ~n2593 ) | ( n2429 & n2594 ) | ( ~n2593 & n2594 ) ;
  assign n2596 = ( x92 & ~n2429 ) | ( x92 & n2592 ) | ( ~n2429 & n2592 ) ;
  assign n2597 = n165 | n2596 ;
  assign n2598 = ( x35 & ~x64 ) | ( x35 & n2597 ) | ( ~x64 & n2597 ) ;
  assign n2599 = ~x35 & n2597 ;
  assign n2600 = ( n2435 & n2598 ) | ( n2435 & ~n2599 ) | ( n2598 & ~n2599 ) ;
  assign n2601 = ~x34 & x64 ;
  assign n2602 = ( x65 & ~n2600 ) | ( x65 & n2601 ) | ( ~n2600 & n2601 ) ;
  assign n2603 = ( x65 & n2435 ) | ( x65 & ~n2597 ) | ( n2435 & ~n2597 ) ;
  assign n2604 = x65 & n2435 ;
  assign n2605 = ( n2434 & n2603 ) | ( n2434 & n2604 ) | ( n2603 & n2604 ) ;
  assign n2606 = ( ~n2434 & n2603 ) | ( ~n2434 & n2604 ) | ( n2603 & n2604 ) ;
  assign n2607 = ( n2434 & ~n2605 ) | ( n2434 & n2606 ) | ( ~n2605 & n2606 ) ;
  assign n2608 = ( x66 & n2602 ) | ( x66 & ~n2607 ) | ( n2602 & ~n2607 ) ;
  assign n2609 = ( x66 & n2436 ) | ( x66 & ~n2597 ) | ( n2436 & ~n2597 ) ;
  assign n2610 = x66 & n2436 ;
  assign n2611 = ( n2441 & n2609 ) | ( n2441 & n2610 ) | ( n2609 & n2610 ) ;
  assign n2612 = ( ~n2441 & n2609 ) | ( ~n2441 & n2610 ) | ( n2609 & n2610 ) ;
  assign n2613 = ( n2441 & ~n2611 ) | ( n2441 & n2612 ) | ( ~n2611 & n2612 ) ;
  assign n2614 = ( x67 & n2608 ) | ( x67 & ~n2613 ) | ( n2608 & ~n2613 ) ;
  assign n2615 = ( x67 & n2442 ) | ( x67 & ~n2597 ) | ( n2442 & ~n2597 ) ;
  assign n2616 = x67 & n2442 ;
  assign n2617 = ( ~n2447 & n2615 ) | ( ~n2447 & n2616 ) | ( n2615 & n2616 ) ;
  assign n2618 = ( n2447 & n2615 ) | ( n2447 & n2616 ) | ( n2615 & n2616 ) ;
  assign n2619 = ( n2447 & n2617 ) | ( n2447 & ~n2618 ) | ( n2617 & ~n2618 ) ;
  assign n2620 = ( x68 & n2614 ) | ( x68 & ~n2619 ) | ( n2614 & ~n2619 ) ;
  assign n2621 = ( x68 & n2448 ) | ( x68 & ~n2597 ) | ( n2448 & ~n2597 ) ;
  assign n2622 = x68 & n2448 ;
  assign n2623 = ( n2453 & n2621 ) | ( n2453 & n2622 ) | ( n2621 & n2622 ) ;
  assign n2624 = ( ~n2453 & n2621 ) | ( ~n2453 & n2622 ) | ( n2621 & n2622 ) ;
  assign n2625 = ( n2453 & ~n2623 ) | ( n2453 & n2624 ) | ( ~n2623 & n2624 ) ;
  assign n2626 = ( x69 & n2620 ) | ( x69 & ~n2625 ) | ( n2620 & ~n2625 ) ;
  assign n2627 = ( x69 & n2454 ) | ( x69 & ~n2597 ) | ( n2454 & ~n2597 ) ;
  assign n2628 = x69 & n2454 ;
  assign n2629 = ( ~n2459 & n2627 ) | ( ~n2459 & n2628 ) | ( n2627 & n2628 ) ;
  assign n2630 = ( n2459 & n2627 ) | ( n2459 & n2628 ) | ( n2627 & n2628 ) ;
  assign n2631 = ( n2459 & n2629 ) | ( n2459 & ~n2630 ) | ( n2629 & ~n2630 ) ;
  assign n2632 = ( x70 & n2626 ) | ( x70 & ~n2631 ) | ( n2626 & ~n2631 ) ;
  assign n2633 = ( x70 & n2460 ) | ( x70 & ~n2597 ) | ( n2460 & ~n2597 ) ;
  assign n2634 = x70 & n2460 ;
  assign n2635 = ( n2465 & n2633 ) | ( n2465 & n2634 ) | ( n2633 & n2634 ) ;
  assign n2636 = ( ~n2465 & n2633 ) | ( ~n2465 & n2634 ) | ( n2633 & n2634 ) ;
  assign n2637 = ( n2465 & ~n2635 ) | ( n2465 & n2636 ) | ( ~n2635 & n2636 ) ;
  assign n2638 = ( x71 & n2632 ) | ( x71 & ~n2637 ) | ( n2632 & ~n2637 ) ;
  assign n2639 = ( x71 & n2466 ) | ( x71 & ~n2597 ) | ( n2466 & ~n2597 ) ;
  assign n2640 = x71 & n2466 ;
  assign n2641 = ( ~n2471 & n2639 ) | ( ~n2471 & n2640 ) | ( n2639 & n2640 ) ;
  assign n2642 = ( n2471 & n2639 ) | ( n2471 & n2640 ) | ( n2639 & n2640 ) ;
  assign n2643 = ( n2471 & n2641 ) | ( n2471 & ~n2642 ) | ( n2641 & ~n2642 ) ;
  assign n2644 = ( x72 & n2638 ) | ( x72 & ~n2643 ) | ( n2638 & ~n2643 ) ;
  assign n2645 = ( x72 & n2472 ) | ( x72 & ~n2597 ) | ( n2472 & ~n2597 ) ;
  assign n2646 = x72 & n2472 ;
  assign n2647 = ( n2477 & n2645 ) | ( n2477 & n2646 ) | ( n2645 & n2646 ) ;
  assign n2648 = ( ~n2477 & n2645 ) | ( ~n2477 & n2646 ) | ( n2645 & n2646 ) ;
  assign n2649 = ( n2477 & ~n2647 ) | ( n2477 & n2648 ) | ( ~n2647 & n2648 ) ;
  assign n2650 = ( x73 & n2644 ) | ( x73 & ~n2649 ) | ( n2644 & ~n2649 ) ;
  assign n2651 = ( x73 & n2478 ) | ( x73 & ~n2597 ) | ( n2478 & ~n2597 ) ;
  assign n2652 = x73 & n2478 ;
  assign n2653 = ( ~n2483 & n2651 ) | ( ~n2483 & n2652 ) | ( n2651 & n2652 ) ;
  assign n2654 = ( n2483 & n2651 ) | ( n2483 & n2652 ) | ( n2651 & n2652 ) ;
  assign n2655 = ( n2483 & n2653 ) | ( n2483 & ~n2654 ) | ( n2653 & ~n2654 ) ;
  assign n2656 = ( x74 & n2650 ) | ( x74 & ~n2655 ) | ( n2650 & ~n2655 ) ;
  assign n2657 = ( x74 & n2484 ) | ( x74 & ~n2597 ) | ( n2484 & ~n2597 ) ;
  assign n2658 = x74 & n2484 ;
  assign n2659 = ( n2489 & n2657 ) | ( n2489 & n2658 ) | ( n2657 & n2658 ) ;
  assign n2660 = ( ~n2489 & n2657 ) | ( ~n2489 & n2658 ) | ( n2657 & n2658 ) ;
  assign n2661 = ( n2489 & ~n2659 ) | ( n2489 & n2660 ) | ( ~n2659 & n2660 ) ;
  assign n2662 = ( x75 & n2656 ) | ( x75 & ~n2661 ) | ( n2656 & ~n2661 ) ;
  assign n2663 = ( x75 & n2490 ) | ( x75 & ~n2597 ) | ( n2490 & ~n2597 ) ;
  assign n2664 = x75 & n2490 ;
  assign n2665 = ( ~n2495 & n2663 ) | ( ~n2495 & n2664 ) | ( n2663 & n2664 ) ;
  assign n2666 = ( n2495 & n2663 ) | ( n2495 & n2664 ) | ( n2663 & n2664 ) ;
  assign n2667 = ( n2495 & n2665 ) | ( n2495 & ~n2666 ) | ( n2665 & ~n2666 ) ;
  assign n2668 = ( x76 & n2662 ) | ( x76 & ~n2667 ) | ( n2662 & ~n2667 ) ;
  assign n2669 = ( x76 & n2496 ) | ( x76 & ~n2597 ) | ( n2496 & ~n2597 ) ;
  assign n2670 = x76 & n2496 ;
  assign n2671 = ( n2501 & n2669 ) | ( n2501 & n2670 ) | ( n2669 & n2670 ) ;
  assign n2672 = ( ~n2501 & n2669 ) | ( ~n2501 & n2670 ) | ( n2669 & n2670 ) ;
  assign n2673 = ( n2501 & ~n2671 ) | ( n2501 & n2672 ) | ( ~n2671 & n2672 ) ;
  assign n2674 = ( x77 & n2668 ) | ( x77 & ~n2673 ) | ( n2668 & ~n2673 ) ;
  assign n2675 = ( x77 & n2502 ) | ( x77 & ~n2597 ) | ( n2502 & ~n2597 ) ;
  assign n2676 = x77 & n2502 ;
  assign n2677 = ( ~n2507 & n2675 ) | ( ~n2507 & n2676 ) | ( n2675 & n2676 ) ;
  assign n2678 = ( n2507 & n2675 ) | ( n2507 & n2676 ) | ( n2675 & n2676 ) ;
  assign n2679 = ( n2507 & n2677 ) | ( n2507 & ~n2678 ) | ( n2677 & ~n2678 ) ;
  assign n2680 = ( x78 & n2674 ) | ( x78 & ~n2679 ) | ( n2674 & ~n2679 ) ;
  assign n2681 = ( x78 & n2508 ) | ( x78 & ~n2597 ) | ( n2508 & ~n2597 ) ;
  assign n2682 = x78 & n2508 ;
  assign n2683 = ( n2513 & n2681 ) | ( n2513 & n2682 ) | ( n2681 & n2682 ) ;
  assign n2684 = ( ~n2513 & n2681 ) | ( ~n2513 & n2682 ) | ( n2681 & n2682 ) ;
  assign n2685 = ( n2513 & ~n2683 ) | ( n2513 & n2684 ) | ( ~n2683 & n2684 ) ;
  assign n2686 = ( x79 & n2680 ) | ( x79 & ~n2685 ) | ( n2680 & ~n2685 ) ;
  assign n2687 = ( x79 & n2514 ) | ( x79 & ~n2597 ) | ( n2514 & ~n2597 ) ;
  assign n2688 = x79 & n2514 ;
  assign n2689 = ( ~n2519 & n2687 ) | ( ~n2519 & n2688 ) | ( n2687 & n2688 ) ;
  assign n2690 = ( n2519 & n2687 ) | ( n2519 & n2688 ) | ( n2687 & n2688 ) ;
  assign n2691 = ( n2519 & n2689 ) | ( n2519 & ~n2690 ) | ( n2689 & ~n2690 ) ;
  assign n2692 = ( x80 & n2686 ) | ( x80 & ~n2691 ) | ( n2686 & ~n2691 ) ;
  assign n2693 = ( x80 & n2520 ) | ( x80 & ~n2597 ) | ( n2520 & ~n2597 ) ;
  assign n2694 = x80 & n2520 ;
  assign n2695 = ( n2525 & n2693 ) | ( n2525 & n2694 ) | ( n2693 & n2694 ) ;
  assign n2696 = ( ~n2525 & n2693 ) | ( ~n2525 & n2694 ) | ( n2693 & n2694 ) ;
  assign n2697 = ( n2525 & ~n2695 ) | ( n2525 & n2696 ) | ( ~n2695 & n2696 ) ;
  assign n2698 = ( x81 & n2692 ) | ( x81 & ~n2697 ) | ( n2692 & ~n2697 ) ;
  assign n2699 = ( x81 & n2526 ) | ( x81 & ~n2597 ) | ( n2526 & ~n2597 ) ;
  assign n2700 = x81 & n2526 ;
  assign n2701 = ( ~n2531 & n2699 ) | ( ~n2531 & n2700 ) | ( n2699 & n2700 ) ;
  assign n2702 = ( n2531 & n2699 ) | ( n2531 & n2700 ) | ( n2699 & n2700 ) ;
  assign n2703 = ( n2531 & n2701 ) | ( n2531 & ~n2702 ) | ( n2701 & ~n2702 ) ;
  assign n2704 = ( x82 & n2698 ) | ( x82 & ~n2703 ) | ( n2698 & ~n2703 ) ;
  assign n2705 = ( x82 & n2532 ) | ( x82 & ~n2597 ) | ( n2532 & ~n2597 ) ;
  assign n2706 = x82 & n2532 ;
  assign n2707 = ( n2537 & n2705 ) | ( n2537 & n2706 ) | ( n2705 & n2706 ) ;
  assign n2708 = ( ~n2537 & n2705 ) | ( ~n2537 & n2706 ) | ( n2705 & n2706 ) ;
  assign n2709 = ( n2537 & ~n2707 ) | ( n2537 & n2708 ) | ( ~n2707 & n2708 ) ;
  assign n2710 = ( x83 & n2704 ) | ( x83 & ~n2709 ) | ( n2704 & ~n2709 ) ;
  assign n2711 = ( x83 & n2538 ) | ( x83 & ~n2597 ) | ( n2538 & ~n2597 ) ;
  assign n2712 = x83 & n2538 ;
  assign n2713 = ( ~n2543 & n2711 ) | ( ~n2543 & n2712 ) | ( n2711 & n2712 ) ;
  assign n2714 = ( n2543 & n2711 ) | ( n2543 & n2712 ) | ( n2711 & n2712 ) ;
  assign n2715 = ( n2543 & n2713 ) | ( n2543 & ~n2714 ) | ( n2713 & ~n2714 ) ;
  assign n2716 = ( x84 & n2710 ) | ( x84 & ~n2715 ) | ( n2710 & ~n2715 ) ;
  assign n2717 = ( x84 & n2544 ) | ( x84 & ~n2597 ) | ( n2544 & ~n2597 ) ;
  assign n2718 = x84 & n2544 ;
  assign n2719 = ( n2549 & n2717 ) | ( n2549 & n2718 ) | ( n2717 & n2718 ) ;
  assign n2720 = ( ~n2549 & n2717 ) | ( ~n2549 & n2718 ) | ( n2717 & n2718 ) ;
  assign n2721 = ( n2549 & ~n2719 ) | ( n2549 & n2720 ) | ( ~n2719 & n2720 ) ;
  assign n2722 = ( x85 & n2716 ) | ( x85 & ~n2721 ) | ( n2716 & ~n2721 ) ;
  assign n2723 = ( x85 & n2550 ) | ( x85 & ~n2597 ) | ( n2550 & ~n2597 ) ;
  assign n2724 = x85 & n2550 ;
  assign n2725 = ( ~n2555 & n2723 ) | ( ~n2555 & n2724 ) | ( n2723 & n2724 ) ;
  assign n2726 = ( n2555 & n2723 ) | ( n2555 & n2724 ) | ( n2723 & n2724 ) ;
  assign n2727 = ( n2555 & n2725 ) | ( n2555 & ~n2726 ) | ( n2725 & ~n2726 ) ;
  assign n2728 = ( x86 & n2722 ) | ( x86 & ~n2727 ) | ( n2722 & ~n2727 ) ;
  assign n2729 = ( x86 & n2556 ) | ( x86 & ~n2597 ) | ( n2556 & ~n2597 ) ;
  assign n2730 = x86 & n2556 ;
  assign n2731 = ( n2561 & n2729 ) | ( n2561 & n2730 ) | ( n2729 & n2730 ) ;
  assign n2732 = ( ~n2561 & n2729 ) | ( ~n2561 & n2730 ) | ( n2729 & n2730 ) ;
  assign n2733 = ( n2561 & ~n2731 ) | ( n2561 & n2732 ) | ( ~n2731 & n2732 ) ;
  assign n2734 = ( x87 & n2728 ) | ( x87 & ~n2733 ) | ( n2728 & ~n2733 ) ;
  assign n2735 = ( x87 & n2562 ) | ( x87 & ~n2597 ) | ( n2562 & ~n2597 ) ;
  assign n2736 = x87 & n2562 ;
  assign n2737 = ( ~n2567 & n2735 ) | ( ~n2567 & n2736 ) | ( n2735 & n2736 ) ;
  assign n2738 = ( n2567 & n2735 ) | ( n2567 & n2736 ) | ( n2735 & n2736 ) ;
  assign n2739 = ( n2567 & n2737 ) | ( n2567 & ~n2738 ) | ( n2737 & ~n2738 ) ;
  assign n2740 = ( x88 & n2734 ) | ( x88 & ~n2739 ) | ( n2734 & ~n2739 ) ;
  assign n2741 = ( x88 & n2568 ) | ( x88 & ~n2597 ) | ( n2568 & ~n2597 ) ;
  assign n2742 = x88 & n2568 ;
  assign n2743 = ( n2573 & n2741 ) | ( n2573 & n2742 ) | ( n2741 & n2742 ) ;
  assign n2744 = ( ~n2573 & n2741 ) | ( ~n2573 & n2742 ) | ( n2741 & n2742 ) ;
  assign n2745 = ( n2573 & ~n2743 ) | ( n2573 & n2744 ) | ( ~n2743 & n2744 ) ;
  assign n2746 = ( x89 & n2740 ) | ( x89 & ~n2745 ) | ( n2740 & ~n2745 ) ;
  assign n2747 = ( x89 & n2574 ) | ( x89 & ~n2597 ) | ( n2574 & ~n2597 ) ;
  assign n2748 = x89 & n2574 ;
  assign n2749 = ( ~n2579 & n2747 ) | ( ~n2579 & n2748 ) | ( n2747 & n2748 ) ;
  assign n2750 = ( n2579 & n2747 ) | ( n2579 & n2748 ) | ( n2747 & n2748 ) ;
  assign n2751 = ( n2579 & n2749 ) | ( n2579 & ~n2750 ) | ( n2749 & ~n2750 ) ;
  assign n2752 = ( x90 & n2746 ) | ( x90 & ~n2751 ) | ( n2746 & ~n2751 ) ;
  assign n2753 = ( x90 & n2580 ) | ( x90 & ~n2597 ) | ( n2580 & ~n2597 ) ;
  assign n2754 = x90 & n2580 ;
  assign n2755 = ( n2585 & n2753 ) | ( n2585 & n2754 ) | ( n2753 & n2754 ) ;
  assign n2756 = ( ~n2585 & n2753 ) | ( ~n2585 & n2754 ) | ( n2753 & n2754 ) ;
  assign n2757 = ( n2585 & ~n2755 ) | ( n2585 & n2756 ) | ( ~n2755 & n2756 ) ;
  assign n2758 = ( x91 & n2752 ) | ( x91 & ~n2757 ) | ( n2752 & ~n2757 ) ;
  assign n2759 = ( x91 & n2586 ) | ( x91 & ~n2597 ) | ( n2586 & ~n2597 ) ;
  assign n2760 = x91 & n2586 ;
  assign n2761 = ( n2591 & n2759 ) | ( n2591 & n2760 ) | ( n2759 & n2760 ) ;
  assign n2762 = ( ~n2591 & n2759 ) | ( ~n2591 & n2760 ) | ( n2759 & n2760 ) ;
  assign n2763 = ( n2591 & ~n2761 ) | ( n2591 & n2762 ) | ( ~n2761 & n2762 ) ;
  assign n2764 = ( x92 & n2758 ) | ( x92 & ~n2763 ) | ( n2758 & ~n2763 ) ;
  assign n2765 = ( x93 & ~n2595 ) | ( x93 & n2764 ) | ( ~n2595 & n2764 ) ;
  assign n2766 = n164 | n2765 ;
  assign n2767 = n2595 & n2766 ;
  assign n2768 = n280 | n2767 ;
  assign n2769 = ( x34 & ~x64 ) | ( x34 & n2766 ) | ( ~x64 & n2766 ) ;
  assign n2770 = ~x34 & n2766 ;
  assign n2771 = ( n2601 & n2769 ) | ( n2601 & ~n2770 ) | ( n2769 & ~n2770 ) ;
  assign n2772 = ~x33 & x64 ;
  assign n2773 = ( x65 & ~n2771 ) | ( x65 & n2772 ) | ( ~n2771 & n2772 ) ;
  assign n2774 = ( x65 & n2601 ) | ( x65 & ~n2766 ) | ( n2601 & ~n2766 ) ;
  assign n2775 = x65 & n2601 ;
  assign n2776 = ( n2600 & n2774 ) | ( n2600 & n2775 ) | ( n2774 & n2775 ) ;
  assign n2777 = ( ~n2600 & n2774 ) | ( ~n2600 & n2775 ) | ( n2774 & n2775 ) ;
  assign n2778 = ( n2600 & ~n2776 ) | ( n2600 & n2777 ) | ( ~n2776 & n2777 ) ;
  assign n2779 = ( x66 & n2773 ) | ( x66 & ~n2778 ) | ( n2773 & ~n2778 ) ;
  assign n2780 = ( x66 & n2602 ) | ( x66 & ~n2766 ) | ( n2602 & ~n2766 ) ;
  assign n2781 = x66 & n2602 ;
  assign n2782 = ( n2607 & n2780 ) | ( n2607 & n2781 ) | ( n2780 & n2781 ) ;
  assign n2783 = ( ~n2607 & n2780 ) | ( ~n2607 & n2781 ) | ( n2780 & n2781 ) ;
  assign n2784 = ( n2607 & ~n2782 ) | ( n2607 & n2783 ) | ( ~n2782 & n2783 ) ;
  assign n2785 = ( x67 & n2779 ) | ( x67 & ~n2784 ) | ( n2779 & ~n2784 ) ;
  assign n2786 = ( x67 & n2608 ) | ( x67 & ~n2766 ) | ( n2608 & ~n2766 ) ;
  assign n2787 = x67 & n2608 ;
  assign n2788 = ( ~n2613 & n2786 ) | ( ~n2613 & n2787 ) | ( n2786 & n2787 ) ;
  assign n2789 = ( n2613 & n2786 ) | ( n2613 & n2787 ) | ( n2786 & n2787 ) ;
  assign n2790 = ( n2613 & n2788 ) | ( n2613 & ~n2789 ) | ( n2788 & ~n2789 ) ;
  assign n2791 = ( x68 & n2785 ) | ( x68 & ~n2790 ) | ( n2785 & ~n2790 ) ;
  assign n2792 = ( x68 & n2614 ) | ( x68 & ~n2766 ) | ( n2614 & ~n2766 ) ;
  assign n2793 = x68 & n2614 ;
  assign n2794 = ( n2619 & n2792 ) | ( n2619 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2795 = ( ~n2619 & n2792 ) | ( ~n2619 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2796 = ( n2619 & ~n2794 ) | ( n2619 & n2795 ) | ( ~n2794 & n2795 ) ;
  assign n2797 = ( x69 & n2791 ) | ( x69 & ~n2796 ) | ( n2791 & ~n2796 ) ;
  assign n2798 = ( x69 & n2620 ) | ( x69 & ~n2766 ) | ( n2620 & ~n2766 ) ;
  assign n2799 = x69 & n2620 ;
  assign n2800 = ( ~n2625 & n2798 ) | ( ~n2625 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2801 = ( n2625 & n2798 ) | ( n2625 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2802 = ( n2625 & n2800 ) | ( n2625 & ~n2801 ) | ( n2800 & ~n2801 ) ;
  assign n2803 = ( x70 & n2797 ) | ( x70 & ~n2802 ) | ( n2797 & ~n2802 ) ;
  assign n2804 = ( x70 & n2626 ) | ( x70 & ~n2766 ) | ( n2626 & ~n2766 ) ;
  assign n2805 = x70 & n2626 ;
  assign n2806 = ( n2631 & n2804 ) | ( n2631 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2807 = ( ~n2631 & n2804 ) | ( ~n2631 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2808 = ( n2631 & ~n2806 ) | ( n2631 & n2807 ) | ( ~n2806 & n2807 ) ;
  assign n2809 = ( x71 & n2803 ) | ( x71 & ~n2808 ) | ( n2803 & ~n2808 ) ;
  assign n2810 = ( x71 & n2632 ) | ( x71 & ~n2766 ) | ( n2632 & ~n2766 ) ;
  assign n2811 = x71 & n2632 ;
  assign n2812 = ( ~n2637 & n2810 ) | ( ~n2637 & n2811 ) | ( n2810 & n2811 ) ;
  assign n2813 = ( n2637 & n2810 ) | ( n2637 & n2811 ) | ( n2810 & n2811 ) ;
  assign n2814 = ( n2637 & n2812 ) | ( n2637 & ~n2813 ) | ( n2812 & ~n2813 ) ;
  assign n2815 = ( x72 & n2809 ) | ( x72 & ~n2814 ) | ( n2809 & ~n2814 ) ;
  assign n2816 = ( x72 & n2638 ) | ( x72 & ~n2766 ) | ( n2638 & ~n2766 ) ;
  assign n2817 = x72 & n2638 ;
  assign n2818 = ( n2643 & n2816 ) | ( n2643 & n2817 ) | ( n2816 & n2817 ) ;
  assign n2819 = ( ~n2643 & n2816 ) | ( ~n2643 & n2817 ) | ( n2816 & n2817 ) ;
  assign n2820 = ( n2643 & ~n2818 ) | ( n2643 & n2819 ) | ( ~n2818 & n2819 ) ;
  assign n2821 = ( x73 & n2815 ) | ( x73 & ~n2820 ) | ( n2815 & ~n2820 ) ;
  assign n2822 = ( x73 & n2644 ) | ( x73 & ~n2766 ) | ( n2644 & ~n2766 ) ;
  assign n2823 = x73 & n2644 ;
  assign n2824 = ( ~n2649 & n2822 ) | ( ~n2649 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = ( n2649 & n2822 ) | ( n2649 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2826 = ( n2649 & n2824 ) | ( n2649 & ~n2825 ) | ( n2824 & ~n2825 ) ;
  assign n2827 = ( x74 & n2821 ) | ( x74 & ~n2826 ) | ( n2821 & ~n2826 ) ;
  assign n2828 = ( x74 & n2650 ) | ( x74 & ~n2766 ) | ( n2650 & ~n2766 ) ;
  assign n2829 = x74 & n2650 ;
  assign n2830 = ( n2655 & n2828 ) | ( n2655 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = ( ~n2655 & n2828 ) | ( ~n2655 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2832 = ( n2655 & ~n2830 ) | ( n2655 & n2831 ) | ( ~n2830 & n2831 ) ;
  assign n2833 = ( x75 & n2827 ) | ( x75 & ~n2832 ) | ( n2827 & ~n2832 ) ;
  assign n2834 = ( x75 & n2656 ) | ( x75 & ~n2766 ) | ( n2656 & ~n2766 ) ;
  assign n2835 = x75 & n2656 ;
  assign n2836 = ( ~n2661 & n2834 ) | ( ~n2661 & n2835 ) | ( n2834 & n2835 ) ;
  assign n2837 = ( n2661 & n2834 ) | ( n2661 & n2835 ) | ( n2834 & n2835 ) ;
  assign n2838 = ( n2661 & n2836 ) | ( n2661 & ~n2837 ) | ( n2836 & ~n2837 ) ;
  assign n2839 = ( x76 & n2833 ) | ( x76 & ~n2838 ) | ( n2833 & ~n2838 ) ;
  assign n2840 = ( x76 & n2662 ) | ( x76 & ~n2766 ) | ( n2662 & ~n2766 ) ;
  assign n2841 = x76 & n2662 ;
  assign n2842 = ( n2667 & n2840 ) | ( n2667 & n2841 ) | ( n2840 & n2841 ) ;
  assign n2843 = ( ~n2667 & n2840 ) | ( ~n2667 & n2841 ) | ( n2840 & n2841 ) ;
  assign n2844 = ( n2667 & ~n2842 ) | ( n2667 & n2843 ) | ( ~n2842 & n2843 ) ;
  assign n2845 = ( x77 & n2839 ) | ( x77 & ~n2844 ) | ( n2839 & ~n2844 ) ;
  assign n2846 = ( x77 & n2668 ) | ( x77 & ~n2766 ) | ( n2668 & ~n2766 ) ;
  assign n2847 = x77 & n2668 ;
  assign n2848 = ( ~n2673 & n2846 ) | ( ~n2673 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2849 = ( n2673 & n2846 ) | ( n2673 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2850 = ( n2673 & n2848 ) | ( n2673 & ~n2849 ) | ( n2848 & ~n2849 ) ;
  assign n2851 = ( x78 & n2845 ) | ( x78 & ~n2850 ) | ( n2845 & ~n2850 ) ;
  assign n2852 = ( x78 & n2674 ) | ( x78 & ~n2766 ) | ( n2674 & ~n2766 ) ;
  assign n2853 = x78 & n2674 ;
  assign n2854 = ( n2679 & n2852 ) | ( n2679 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2855 = ( ~n2679 & n2852 ) | ( ~n2679 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2856 = ( n2679 & ~n2854 ) | ( n2679 & n2855 ) | ( ~n2854 & n2855 ) ;
  assign n2857 = ( x79 & n2851 ) | ( x79 & ~n2856 ) | ( n2851 & ~n2856 ) ;
  assign n2858 = ( x79 & n2680 ) | ( x79 & ~n2766 ) | ( n2680 & ~n2766 ) ;
  assign n2859 = x79 & n2680 ;
  assign n2860 = ( ~n2685 & n2858 ) | ( ~n2685 & n2859 ) | ( n2858 & n2859 ) ;
  assign n2861 = ( n2685 & n2858 ) | ( n2685 & n2859 ) | ( n2858 & n2859 ) ;
  assign n2862 = ( n2685 & n2860 ) | ( n2685 & ~n2861 ) | ( n2860 & ~n2861 ) ;
  assign n2863 = ( x80 & n2857 ) | ( x80 & ~n2862 ) | ( n2857 & ~n2862 ) ;
  assign n2864 = ( x80 & n2686 ) | ( x80 & ~n2766 ) | ( n2686 & ~n2766 ) ;
  assign n2865 = x80 & n2686 ;
  assign n2866 = ( n2691 & n2864 ) | ( n2691 & n2865 ) | ( n2864 & n2865 ) ;
  assign n2867 = ( ~n2691 & n2864 ) | ( ~n2691 & n2865 ) | ( n2864 & n2865 ) ;
  assign n2868 = ( n2691 & ~n2866 ) | ( n2691 & n2867 ) | ( ~n2866 & n2867 ) ;
  assign n2869 = ( x81 & n2863 ) | ( x81 & ~n2868 ) | ( n2863 & ~n2868 ) ;
  assign n2870 = ( x81 & n2692 ) | ( x81 & ~n2766 ) | ( n2692 & ~n2766 ) ;
  assign n2871 = x81 & n2692 ;
  assign n2872 = ( ~n2697 & n2870 ) | ( ~n2697 & n2871 ) | ( n2870 & n2871 ) ;
  assign n2873 = ( n2697 & n2870 ) | ( n2697 & n2871 ) | ( n2870 & n2871 ) ;
  assign n2874 = ( n2697 & n2872 ) | ( n2697 & ~n2873 ) | ( n2872 & ~n2873 ) ;
  assign n2875 = ( x82 & n2869 ) | ( x82 & ~n2874 ) | ( n2869 & ~n2874 ) ;
  assign n2876 = ( x82 & n2698 ) | ( x82 & ~n2766 ) | ( n2698 & ~n2766 ) ;
  assign n2877 = x82 & n2698 ;
  assign n2878 = ( n2703 & n2876 ) | ( n2703 & n2877 ) | ( n2876 & n2877 ) ;
  assign n2879 = ( ~n2703 & n2876 ) | ( ~n2703 & n2877 ) | ( n2876 & n2877 ) ;
  assign n2880 = ( n2703 & ~n2878 ) | ( n2703 & n2879 ) | ( ~n2878 & n2879 ) ;
  assign n2881 = ( x83 & n2875 ) | ( x83 & ~n2880 ) | ( n2875 & ~n2880 ) ;
  assign n2882 = ( x83 & n2704 ) | ( x83 & ~n2766 ) | ( n2704 & ~n2766 ) ;
  assign n2883 = x83 & n2704 ;
  assign n2884 = ( ~n2709 & n2882 ) | ( ~n2709 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2885 = ( n2709 & n2882 ) | ( n2709 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2886 = ( n2709 & n2884 ) | ( n2709 & ~n2885 ) | ( n2884 & ~n2885 ) ;
  assign n2887 = ( x84 & n2881 ) | ( x84 & ~n2886 ) | ( n2881 & ~n2886 ) ;
  assign n2888 = ( x84 & n2710 ) | ( x84 & ~n2766 ) | ( n2710 & ~n2766 ) ;
  assign n2889 = x84 & n2710 ;
  assign n2890 = ( n2715 & n2888 ) | ( n2715 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2891 = ( ~n2715 & n2888 ) | ( ~n2715 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2892 = ( n2715 & ~n2890 ) | ( n2715 & n2891 ) | ( ~n2890 & n2891 ) ;
  assign n2893 = ( x85 & n2887 ) | ( x85 & ~n2892 ) | ( n2887 & ~n2892 ) ;
  assign n2894 = ( x85 & n2716 ) | ( x85 & ~n2766 ) | ( n2716 & ~n2766 ) ;
  assign n2895 = x85 & n2716 ;
  assign n2896 = ( ~n2721 & n2894 ) | ( ~n2721 & n2895 ) | ( n2894 & n2895 ) ;
  assign n2897 = ( n2721 & n2894 ) | ( n2721 & n2895 ) | ( n2894 & n2895 ) ;
  assign n2898 = ( n2721 & n2896 ) | ( n2721 & ~n2897 ) | ( n2896 & ~n2897 ) ;
  assign n2899 = ( x86 & n2893 ) | ( x86 & ~n2898 ) | ( n2893 & ~n2898 ) ;
  assign n2900 = ( x86 & n2722 ) | ( x86 & ~n2766 ) | ( n2722 & ~n2766 ) ;
  assign n2901 = x86 & n2722 ;
  assign n2902 = ( n2727 & n2900 ) | ( n2727 & n2901 ) | ( n2900 & n2901 ) ;
  assign n2903 = ( ~n2727 & n2900 ) | ( ~n2727 & n2901 ) | ( n2900 & n2901 ) ;
  assign n2904 = ( n2727 & ~n2902 ) | ( n2727 & n2903 ) | ( ~n2902 & n2903 ) ;
  assign n2905 = ( x87 & n2899 ) | ( x87 & ~n2904 ) | ( n2899 & ~n2904 ) ;
  assign n2906 = ( x87 & n2728 ) | ( x87 & ~n2766 ) | ( n2728 & ~n2766 ) ;
  assign n2907 = x87 & n2728 ;
  assign n2908 = ( ~n2733 & n2906 ) | ( ~n2733 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2909 = ( n2733 & n2906 ) | ( n2733 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2910 = ( n2733 & n2908 ) | ( n2733 & ~n2909 ) | ( n2908 & ~n2909 ) ;
  assign n2911 = ( x88 & n2905 ) | ( x88 & ~n2910 ) | ( n2905 & ~n2910 ) ;
  assign n2912 = ( x88 & n2734 ) | ( x88 & ~n2766 ) | ( n2734 & ~n2766 ) ;
  assign n2913 = x88 & n2734 ;
  assign n2914 = ( n2739 & n2912 ) | ( n2739 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2915 = ( ~n2739 & n2912 ) | ( ~n2739 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2916 = ( n2739 & ~n2914 ) | ( n2739 & n2915 ) | ( ~n2914 & n2915 ) ;
  assign n2917 = ( x89 & n2911 ) | ( x89 & ~n2916 ) | ( n2911 & ~n2916 ) ;
  assign n2918 = ( x89 & n2740 ) | ( x89 & ~n2766 ) | ( n2740 & ~n2766 ) ;
  assign n2919 = x89 & n2740 ;
  assign n2920 = ( ~n2745 & n2918 ) | ( ~n2745 & n2919 ) | ( n2918 & n2919 ) ;
  assign n2921 = ( n2745 & n2918 ) | ( n2745 & n2919 ) | ( n2918 & n2919 ) ;
  assign n2922 = ( n2745 & n2920 ) | ( n2745 & ~n2921 ) | ( n2920 & ~n2921 ) ;
  assign n2923 = ( x90 & n2917 ) | ( x90 & ~n2922 ) | ( n2917 & ~n2922 ) ;
  assign n2924 = ( x90 & n2746 ) | ( x90 & ~n2766 ) | ( n2746 & ~n2766 ) ;
  assign n2925 = x90 & n2746 ;
  assign n2926 = ( n2751 & n2924 ) | ( n2751 & n2925 ) | ( n2924 & n2925 ) ;
  assign n2927 = ( ~n2751 & n2924 ) | ( ~n2751 & n2925 ) | ( n2924 & n2925 ) ;
  assign n2928 = ( n2751 & ~n2926 ) | ( n2751 & n2927 ) | ( ~n2926 & n2927 ) ;
  assign n2929 = ( x91 & n2923 ) | ( x91 & ~n2928 ) | ( n2923 & ~n2928 ) ;
  assign n2930 = ( x91 & n2752 ) | ( x91 & ~n2766 ) | ( n2752 & ~n2766 ) ;
  assign n2931 = x91 & n2752 ;
  assign n2932 = ( ~n2757 & n2930 ) | ( ~n2757 & n2931 ) | ( n2930 & n2931 ) ;
  assign n2933 = ( n2757 & n2930 ) | ( n2757 & n2931 ) | ( n2930 & n2931 ) ;
  assign n2934 = ( n2757 & n2932 ) | ( n2757 & ~n2933 ) | ( n2932 & ~n2933 ) ;
  assign n2935 = ( x92 & n2929 ) | ( x92 & ~n2934 ) | ( n2929 & ~n2934 ) ;
  assign n2936 = ( x92 & n2758 ) | ( x92 & ~n2766 ) | ( n2758 & ~n2766 ) ;
  assign n2937 = x92 & n2758 ;
  assign n2938 = ( ~n2763 & n2936 ) | ( ~n2763 & n2937 ) | ( n2936 & n2937 ) ;
  assign n2939 = ( n2763 & n2936 ) | ( n2763 & n2937 ) | ( n2936 & n2937 ) ;
  assign n2940 = ( n2763 & n2938 ) | ( n2763 & ~n2939 ) | ( n2938 & ~n2939 ) ;
  assign n2941 = ( x93 & n2935 ) | ( x93 & ~n2940 ) | ( n2935 & ~n2940 ) ;
  assign n2942 = x94 | n2941 ;
  assign n2943 = ( x94 & n163 ) | ( x94 & n2941 ) | ( n163 & n2941 ) ;
  assign n2944 = ( n2768 & ~n2942 ) | ( n2768 & n2943 ) | ( ~n2942 & n2943 ) ;
  assign n2945 = ( x94 & ~n2768 ) | ( x94 & n2941 ) | ( ~n2768 & n2941 ) ;
  assign n2946 = n163 | n2945 ;
  assign n2947 = ( x33 & ~x64 ) | ( x33 & n2946 ) | ( ~x64 & n2946 ) ;
  assign n2948 = ~x33 & n2946 ;
  assign n2949 = ( n2772 & n2947 ) | ( n2772 & ~n2948 ) | ( n2947 & ~n2948 ) ;
  assign n2950 = ~x32 & x64 ;
  assign n2951 = ( x65 & ~n2949 ) | ( x65 & n2950 ) | ( ~n2949 & n2950 ) ;
  assign n2952 = ( x65 & n2772 ) | ( x65 & ~n2946 ) | ( n2772 & ~n2946 ) ;
  assign n2953 = x65 & n2772 ;
  assign n2954 = ( n2771 & n2952 ) | ( n2771 & n2953 ) | ( n2952 & n2953 ) ;
  assign n2955 = ( ~n2771 & n2952 ) | ( ~n2771 & n2953 ) | ( n2952 & n2953 ) ;
  assign n2956 = ( n2771 & ~n2954 ) | ( n2771 & n2955 ) | ( ~n2954 & n2955 ) ;
  assign n2957 = ( x66 & n2951 ) | ( x66 & ~n2956 ) | ( n2951 & ~n2956 ) ;
  assign n2958 = ( x66 & n2773 ) | ( x66 & ~n2946 ) | ( n2773 & ~n2946 ) ;
  assign n2959 = x66 & n2773 ;
  assign n2960 = ( n2778 & n2958 ) | ( n2778 & n2959 ) | ( n2958 & n2959 ) ;
  assign n2961 = ( ~n2778 & n2958 ) | ( ~n2778 & n2959 ) | ( n2958 & n2959 ) ;
  assign n2962 = ( n2778 & ~n2960 ) | ( n2778 & n2961 ) | ( ~n2960 & n2961 ) ;
  assign n2963 = ( x67 & n2957 ) | ( x67 & ~n2962 ) | ( n2957 & ~n2962 ) ;
  assign n2964 = ( x67 & n2779 ) | ( x67 & ~n2946 ) | ( n2779 & ~n2946 ) ;
  assign n2965 = x67 & n2779 ;
  assign n2966 = ( ~n2784 & n2964 ) | ( ~n2784 & n2965 ) | ( n2964 & n2965 ) ;
  assign n2967 = ( n2784 & n2964 ) | ( n2784 & n2965 ) | ( n2964 & n2965 ) ;
  assign n2968 = ( n2784 & n2966 ) | ( n2784 & ~n2967 ) | ( n2966 & ~n2967 ) ;
  assign n2969 = ( x68 & n2963 ) | ( x68 & ~n2968 ) | ( n2963 & ~n2968 ) ;
  assign n2970 = ( x68 & n2785 ) | ( x68 & ~n2946 ) | ( n2785 & ~n2946 ) ;
  assign n2971 = x68 & n2785 ;
  assign n2972 = ( n2790 & n2970 ) | ( n2790 & n2971 ) | ( n2970 & n2971 ) ;
  assign n2973 = ( ~n2790 & n2970 ) | ( ~n2790 & n2971 ) | ( n2970 & n2971 ) ;
  assign n2974 = ( n2790 & ~n2972 ) | ( n2790 & n2973 ) | ( ~n2972 & n2973 ) ;
  assign n2975 = ( x69 & n2969 ) | ( x69 & ~n2974 ) | ( n2969 & ~n2974 ) ;
  assign n2976 = ( x69 & n2791 ) | ( x69 & ~n2946 ) | ( n2791 & ~n2946 ) ;
  assign n2977 = x69 & n2791 ;
  assign n2978 = ( ~n2796 & n2976 ) | ( ~n2796 & n2977 ) | ( n2976 & n2977 ) ;
  assign n2979 = ( n2796 & n2976 ) | ( n2796 & n2977 ) | ( n2976 & n2977 ) ;
  assign n2980 = ( n2796 & n2978 ) | ( n2796 & ~n2979 ) | ( n2978 & ~n2979 ) ;
  assign n2981 = ( x70 & n2975 ) | ( x70 & ~n2980 ) | ( n2975 & ~n2980 ) ;
  assign n2982 = ( x70 & n2797 ) | ( x70 & ~n2946 ) | ( n2797 & ~n2946 ) ;
  assign n2983 = x70 & n2797 ;
  assign n2984 = ( n2802 & n2982 ) | ( n2802 & n2983 ) | ( n2982 & n2983 ) ;
  assign n2985 = ( ~n2802 & n2982 ) | ( ~n2802 & n2983 ) | ( n2982 & n2983 ) ;
  assign n2986 = ( n2802 & ~n2984 ) | ( n2802 & n2985 ) | ( ~n2984 & n2985 ) ;
  assign n2987 = ( x71 & n2981 ) | ( x71 & ~n2986 ) | ( n2981 & ~n2986 ) ;
  assign n2988 = ( x71 & n2803 ) | ( x71 & ~n2946 ) | ( n2803 & ~n2946 ) ;
  assign n2989 = x71 & n2803 ;
  assign n2990 = ( ~n2808 & n2988 ) | ( ~n2808 & n2989 ) | ( n2988 & n2989 ) ;
  assign n2991 = ( n2808 & n2988 ) | ( n2808 & n2989 ) | ( n2988 & n2989 ) ;
  assign n2992 = ( n2808 & n2990 ) | ( n2808 & ~n2991 ) | ( n2990 & ~n2991 ) ;
  assign n2993 = ( x72 & n2987 ) | ( x72 & ~n2992 ) | ( n2987 & ~n2992 ) ;
  assign n2994 = ( x72 & n2809 ) | ( x72 & ~n2946 ) | ( n2809 & ~n2946 ) ;
  assign n2995 = x72 & n2809 ;
  assign n2996 = ( n2814 & n2994 ) | ( n2814 & n2995 ) | ( n2994 & n2995 ) ;
  assign n2997 = ( ~n2814 & n2994 ) | ( ~n2814 & n2995 ) | ( n2994 & n2995 ) ;
  assign n2998 = ( n2814 & ~n2996 ) | ( n2814 & n2997 ) | ( ~n2996 & n2997 ) ;
  assign n2999 = ( x73 & n2993 ) | ( x73 & ~n2998 ) | ( n2993 & ~n2998 ) ;
  assign n3000 = ( x73 & n2815 ) | ( x73 & ~n2946 ) | ( n2815 & ~n2946 ) ;
  assign n3001 = x73 & n2815 ;
  assign n3002 = ( ~n2820 & n3000 ) | ( ~n2820 & n3001 ) | ( n3000 & n3001 ) ;
  assign n3003 = ( n2820 & n3000 ) | ( n2820 & n3001 ) | ( n3000 & n3001 ) ;
  assign n3004 = ( n2820 & n3002 ) | ( n2820 & ~n3003 ) | ( n3002 & ~n3003 ) ;
  assign n3005 = ( x74 & n2999 ) | ( x74 & ~n3004 ) | ( n2999 & ~n3004 ) ;
  assign n3006 = ( x74 & n2821 ) | ( x74 & ~n2946 ) | ( n2821 & ~n2946 ) ;
  assign n3007 = x74 & n2821 ;
  assign n3008 = ( n2826 & n3006 ) | ( n2826 & n3007 ) | ( n3006 & n3007 ) ;
  assign n3009 = ( ~n2826 & n3006 ) | ( ~n2826 & n3007 ) | ( n3006 & n3007 ) ;
  assign n3010 = ( n2826 & ~n3008 ) | ( n2826 & n3009 ) | ( ~n3008 & n3009 ) ;
  assign n3011 = ( x75 & n3005 ) | ( x75 & ~n3010 ) | ( n3005 & ~n3010 ) ;
  assign n3012 = ( x75 & n2827 ) | ( x75 & ~n2946 ) | ( n2827 & ~n2946 ) ;
  assign n3013 = x75 & n2827 ;
  assign n3014 = ( ~n2832 & n3012 ) | ( ~n2832 & n3013 ) | ( n3012 & n3013 ) ;
  assign n3015 = ( n2832 & n3012 ) | ( n2832 & n3013 ) | ( n3012 & n3013 ) ;
  assign n3016 = ( n2832 & n3014 ) | ( n2832 & ~n3015 ) | ( n3014 & ~n3015 ) ;
  assign n3017 = ( x76 & n3011 ) | ( x76 & ~n3016 ) | ( n3011 & ~n3016 ) ;
  assign n3018 = ( x76 & n2833 ) | ( x76 & ~n2946 ) | ( n2833 & ~n2946 ) ;
  assign n3019 = x76 & n2833 ;
  assign n3020 = ( n2838 & n3018 ) | ( n2838 & n3019 ) | ( n3018 & n3019 ) ;
  assign n3021 = ( ~n2838 & n3018 ) | ( ~n2838 & n3019 ) | ( n3018 & n3019 ) ;
  assign n3022 = ( n2838 & ~n3020 ) | ( n2838 & n3021 ) | ( ~n3020 & n3021 ) ;
  assign n3023 = ( x77 & n3017 ) | ( x77 & ~n3022 ) | ( n3017 & ~n3022 ) ;
  assign n3024 = ( x77 & n2839 ) | ( x77 & ~n2946 ) | ( n2839 & ~n2946 ) ;
  assign n3025 = x77 & n2839 ;
  assign n3026 = ( ~n2844 & n3024 ) | ( ~n2844 & n3025 ) | ( n3024 & n3025 ) ;
  assign n3027 = ( n2844 & n3024 ) | ( n2844 & n3025 ) | ( n3024 & n3025 ) ;
  assign n3028 = ( n2844 & n3026 ) | ( n2844 & ~n3027 ) | ( n3026 & ~n3027 ) ;
  assign n3029 = ( x78 & n3023 ) | ( x78 & ~n3028 ) | ( n3023 & ~n3028 ) ;
  assign n3030 = ( x78 & n2845 ) | ( x78 & ~n2946 ) | ( n2845 & ~n2946 ) ;
  assign n3031 = x78 & n2845 ;
  assign n3032 = ( n2850 & n3030 ) | ( n2850 & n3031 ) | ( n3030 & n3031 ) ;
  assign n3033 = ( ~n2850 & n3030 ) | ( ~n2850 & n3031 ) | ( n3030 & n3031 ) ;
  assign n3034 = ( n2850 & ~n3032 ) | ( n2850 & n3033 ) | ( ~n3032 & n3033 ) ;
  assign n3035 = ( x79 & n3029 ) | ( x79 & ~n3034 ) | ( n3029 & ~n3034 ) ;
  assign n3036 = ( x79 & n2851 ) | ( x79 & ~n2946 ) | ( n2851 & ~n2946 ) ;
  assign n3037 = x79 & n2851 ;
  assign n3038 = ( ~n2856 & n3036 ) | ( ~n2856 & n3037 ) | ( n3036 & n3037 ) ;
  assign n3039 = ( n2856 & n3036 ) | ( n2856 & n3037 ) | ( n3036 & n3037 ) ;
  assign n3040 = ( n2856 & n3038 ) | ( n2856 & ~n3039 ) | ( n3038 & ~n3039 ) ;
  assign n3041 = ( x80 & n3035 ) | ( x80 & ~n3040 ) | ( n3035 & ~n3040 ) ;
  assign n3042 = ( x80 & n2857 ) | ( x80 & ~n2946 ) | ( n2857 & ~n2946 ) ;
  assign n3043 = x80 & n2857 ;
  assign n3044 = ( n2862 & n3042 ) | ( n2862 & n3043 ) | ( n3042 & n3043 ) ;
  assign n3045 = ( ~n2862 & n3042 ) | ( ~n2862 & n3043 ) | ( n3042 & n3043 ) ;
  assign n3046 = ( n2862 & ~n3044 ) | ( n2862 & n3045 ) | ( ~n3044 & n3045 ) ;
  assign n3047 = ( x81 & n3041 ) | ( x81 & ~n3046 ) | ( n3041 & ~n3046 ) ;
  assign n3048 = ( x81 & n2863 ) | ( x81 & ~n2946 ) | ( n2863 & ~n2946 ) ;
  assign n3049 = x81 & n2863 ;
  assign n3050 = ( ~n2868 & n3048 ) | ( ~n2868 & n3049 ) | ( n3048 & n3049 ) ;
  assign n3051 = ( n2868 & n3048 ) | ( n2868 & n3049 ) | ( n3048 & n3049 ) ;
  assign n3052 = ( n2868 & n3050 ) | ( n2868 & ~n3051 ) | ( n3050 & ~n3051 ) ;
  assign n3053 = ( x82 & n3047 ) | ( x82 & ~n3052 ) | ( n3047 & ~n3052 ) ;
  assign n3054 = ( x82 & n2869 ) | ( x82 & ~n2946 ) | ( n2869 & ~n2946 ) ;
  assign n3055 = x82 & n2869 ;
  assign n3056 = ( n2874 & n3054 ) | ( n2874 & n3055 ) | ( n3054 & n3055 ) ;
  assign n3057 = ( ~n2874 & n3054 ) | ( ~n2874 & n3055 ) | ( n3054 & n3055 ) ;
  assign n3058 = ( n2874 & ~n3056 ) | ( n2874 & n3057 ) | ( ~n3056 & n3057 ) ;
  assign n3059 = ( x83 & n3053 ) | ( x83 & ~n3058 ) | ( n3053 & ~n3058 ) ;
  assign n3060 = ( x83 & n2875 ) | ( x83 & ~n2946 ) | ( n2875 & ~n2946 ) ;
  assign n3061 = x83 & n2875 ;
  assign n3062 = ( ~n2880 & n3060 ) | ( ~n2880 & n3061 ) | ( n3060 & n3061 ) ;
  assign n3063 = ( n2880 & n3060 ) | ( n2880 & n3061 ) | ( n3060 & n3061 ) ;
  assign n3064 = ( n2880 & n3062 ) | ( n2880 & ~n3063 ) | ( n3062 & ~n3063 ) ;
  assign n3065 = ( x84 & n3059 ) | ( x84 & ~n3064 ) | ( n3059 & ~n3064 ) ;
  assign n3066 = ( x84 & n2881 ) | ( x84 & ~n2946 ) | ( n2881 & ~n2946 ) ;
  assign n3067 = x84 & n2881 ;
  assign n3068 = ( n2886 & n3066 ) | ( n2886 & n3067 ) | ( n3066 & n3067 ) ;
  assign n3069 = ( ~n2886 & n3066 ) | ( ~n2886 & n3067 ) | ( n3066 & n3067 ) ;
  assign n3070 = ( n2886 & ~n3068 ) | ( n2886 & n3069 ) | ( ~n3068 & n3069 ) ;
  assign n3071 = ( x85 & n3065 ) | ( x85 & ~n3070 ) | ( n3065 & ~n3070 ) ;
  assign n3072 = ( x85 & n2887 ) | ( x85 & ~n2946 ) | ( n2887 & ~n2946 ) ;
  assign n3073 = x85 & n2887 ;
  assign n3074 = ( ~n2892 & n3072 ) | ( ~n2892 & n3073 ) | ( n3072 & n3073 ) ;
  assign n3075 = ( n2892 & n3072 ) | ( n2892 & n3073 ) | ( n3072 & n3073 ) ;
  assign n3076 = ( n2892 & n3074 ) | ( n2892 & ~n3075 ) | ( n3074 & ~n3075 ) ;
  assign n3077 = ( x86 & n3071 ) | ( x86 & ~n3076 ) | ( n3071 & ~n3076 ) ;
  assign n3078 = ( x86 & n2893 ) | ( x86 & ~n2946 ) | ( n2893 & ~n2946 ) ;
  assign n3079 = x86 & n2893 ;
  assign n3080 = ( n2898 & n3078 ) | ( n2898 & n3079 ) | ( n3078 & n3079 ) ;
  assign n3081 = ( ~n2898 & n3078 ) | ( ~n2898 & n3079 ) | ( n3078 & n3079 ) ;
  assign n3082 = ( n2898 & ~n3080 ) | ( n2898 & n3081 ) | ( ~n3080 & n3081 ) ;
  assign n3083 = ( x87 & n3077 ) | ( x87 & ~n3082 ) | ( n3077 & ~n3082 ) ;
  assign n3084 = ( x87 & n2899 ) | ( x87 & ~n2946 ) | ( n2899 & ~n2946 ) ;
  assign n3085 = x87 & n2899 ;
  assign n3086 = ( ~n2904 & n3084 ) | ( ~n2904 & n3085 ) | ( n3084 & n3085 ) ;
  assign n3087 = ( n2904 & n3084 ) | ( n2904 & n3085 ) | ( n3084 & n3085 ) ;
  assign n3088 = ( n2904 & n3086 ) | ( n2904 & ~n3087 ) | ( n3086 & ~n3087 ) ;
  assign n3089 = ( x88 & n3083 ) | ( x88 & ~n3088 ) | ( n3083 & ~n3088 ) ;
  assign n3090 = ( x88 & n2905 ) | ( x88 & ~n2946 ) | ( n2905 & ~n2946 ) ;
  assign n3091 = x88 & n2905 ;
  assign n3092 = ( n2910 & n3090 ) | ( n2910 & n3091 ) | ( n3090 & n3091 ) ;
  assign n3093 = ( ~n2910 & n3090 ) | ( ~n2910 & n3091 ) | ( n3090 & n3091 ) ;
  assign n3094 = ( n2910 & ~n3092 ) | ( n2910 & n3093 ) | ( ~n3092 & n3093 ) ;
  assign n3095 = ( x89 & n3089 ) | ( x89 & ~n3094 ) | ( n3089 & ~n3094 ) ;
  assign n3096 = ( x89 & n2911 ) | ( x89 & ~n2946 ) | ( n2911 & ~n2946 ) ;
  assign n3097 = x89 & n2911 ;
  assign n3098 = ( ~n2916 & n3096 ) | ( ~n2916 & n3097 ) | ( n3096 & n3097 ) ;
  assign n3099 = ( n2916 & n3096 ) | ( n2916 & n3097 ) | ( n3096 & n3097 ) ;
  assign n3100 = ( n2916 & n3098 ) | ( n2916 & ~n3099 ) | ( n3098 & ~n3099 ) ;
  assign n3101 = ( x90 & n3095 ) | ( x90 & ~n3100 ) | ( n3095 & ~n3100 ) ;
  assign n3102 = ( x90 & n2917 ) | ( x90 & ~n2946 ) | ( n2917 & ~n2946 ) ;
  assign n3103 = x90 & n2917 ;
  assign n3104 = ( n2922 & n3102 ) | ( n2922 & n3103 ) | ( n3102 & n3103 ) ;
  assign n3105 = ( ~n2922 & n3102 ) | ( ~n2922 & n3103 ) | ( n3102 & n3103 ) ;
  assign n3106 = ( n2922 & ~n3104 ) | ( n2922 & n3105 ) | ( ~n3104 & n3105 ) ;
  assign n3107 = ( x91 & n3101 ) | ( x91 & ~n3106 ) | ( n3101 & ~n3106 ) ;
  assign n3108 = ( x91 & n2923 ) | ( x91 & ~n2946 ) | ( n2923 & ~n2946 ) ;
  assign n3109 = x91 & n2923 ;
  assign n3110 = ( ~n2928 & n3108 ) | ( ~n2928 & n3109 ) | ( n3108 & n3109 ) ;
  assign n3111 = ( n2928 & n3108 ) | ( n2928 & n3109 ) | ( n3108 & n3109 ) ;
  assign n3112 = ( n2928 & n3110 ) | ( n2928 & ~n3111 ) | ( n3110 & ~n3111 ) ;
  assign n3113 = ( x92 & n3107 ) | ( x92 & ~n3112 ) | ( n3107 & ~n3112 ) ;
  assign n3114 = ( x92 & n2929 ) | ( x92 & ~n2946 ) | ( n2929 & ~n2946 ) ;
  assign n3115 = x92 & n2929 ;
  assign n3116 = ( n2934 & n3114 ) | ( n2934 & n3115 ) | ( n3114 & n3115 ) ;
  assign n3117 = ( ~n2934 & n3114 ) | ( ~n2934 & n3115 ) | ( n3114 & n3115 ) ;
  assign n3118 = ( n2934 & ~n3116 ) | ( n2934 & n3117 ) | ( ~n3116 & n3117 ) ;
  assign n3119 = ( x93 & n3113 ) | ( x93 & ~n3118 ) | ( n3113 & ~n3118 ) ;
  assign n3120 = ( x93 & n2935 ) | ( x93 & ~n2946 ) | ( n2935 & ~n2946 ) ;
  assign n3121 = x93 & n2935 ;
  assign n3122 = ( n2940 & n3120 ) | ( n2940 & n3121 ) | ( n3120 & n3121 ) ;
  assign n3123 = ( ~n2940 & n3120 ) | ( ~n2940 & n3121 ) | ( n3120 & n3121 ) ;
  assign n3124 = ( n2940 & ~n3122 ) | ( n2940 & n3123 ) | ( ~n3122 & n3123 ) ;
  assign n3125 = ( x94 & n3119 ) | ( x94 & ~n3124 ) | ( n3119 & ~n3124 ) ;
  assign n3126 = x95 | n3125 ;
  assign n3127 = ( x95 & n162 ) | ( x95 & n3125 ) | ( n162 & n3125 ) ;
  assign n3128 = ( n2944 & ~n3126 ) | ( n2944 & n3127 ) | ( ~n3126 & n3127 ) ;
  assign n3129 = ( x95 & ~n2944 ) | ( x95 & n3125 ) | ( ~n2944 & n3125 ) ;
  assign n3130 = n162 | n3129 ;
  assign n3131 = ( x32 & ~x64 ) | ( x32 & n3130 ) | ( ~x64 & n3130 ) ;
  assign n3132 = ~x32 & n3130 ;
  assign n3133 = ( n2950 & n3131 ) | ( n2950 & ~n3132 ) | ( n3131 & ~n3132 ) ;
  assign n3134 = ~x31 & x64 ;
  assign n3135 = ( x65 & ~n3133 ) | ( x65 & n3134 ) | ( ~n3133 & n3134 ) ;
  assign n3136 = ( x65 & n2950 ) | ( x65 & ~n3130 ) | ( n2950 & ~n3130 ) ;
  assign n3137 = x65 & n2950 ;
  assign n3138 = ( n2949 & n3136 ) | ( n2949 & n3137 ) | ( n3136 & n3137 ) ;
  assign n3139 = ( ~n2949 & n3136 ) | ( ~n2949 & n3137 ) | ( n3136 & n3137 ) ;
  assign n3140 = ( n2949 & ~n3138 ) | ( n2949 & n3139 ) | ( ~n3138 & n3139 ) ;
  assign n3141 = ( x66 & n3135 ) | ( x66 & ~n3140 ) | ( n3135 & ~n3140 ) ;
  assign n3142 = ( x66 & n2951 ) | ( x66 & ~n3130 ) | ( n2951 & ~n3130 ) ;
  assign n3143 = x66 & n2951 ;
  assign n3144 = ( n2956 & n3142 ) | ( n2956 & n3143 ) | ( n3142 & n3143 ) ;
  assign n3145 = ( ~n2956 & n3142 ) | ( ~n2956 & n3143 ) | ( n3142 & n3143 ) ;
  assign n3146 = ( n2956 & ~n3144 ) | ( n2956 & n3145 ) | ( ~n3144 & n3145 ) ;
  assign n3147 = ( x67 & n3141 ) | ( x67 & ~n3146 ) | ( n3141 & ~n3146 ) ;
  assign n3148 = ( x67 & n2957 ) | ( x67 & ~n3130 ) | ( n2957 & ~n3130 ) ;
  assign n3149 = x67 & n2957 ;
  assign n3150 = ( ~n2962 & n3148 ) | ( ~n2962 & n3149 ) | ( n3148 & n3149 ) ;
  assign n3151 = ( n2962 & n3148 ) | ( n2962 & n3149 ) | ( n3148 & n3149 ) ;
  assign n3152 = ( n2962 & n3150 ) | ( n2962 & ~n3151 ) | ( n3150 & ~n3151 ) ;
  assign n3153 = ( x68 & n3147 ) | ( x68 & ~n3152 ) | ( n3147 & ~n3152 ) ;
  assign n3154 = ( x68 & n2963 ) | ( x68 & ~n3130 ) | ( n2963 & ~n3130 ) ;
  assign n3155 = x68 & n2963 ;
  assign n3156 = ( n2968 & n3154 ) | ( n2968 & n3155 ) | ( n3154 & n3155 ) ;
  assign n3157 = ( ~n2968 & n3154 ) | ( ~n2968 & n3155 ) | ( n3154 & n3155 ) ;
  assign n3158 = ( n2968 & ~n3156 ) | ( n2968 & n3157 ) | ( ~n3156 & n3157 ) ;
  assign n3159 = ( x69 & n3153 ) | ( x69 & ~n3158 ) | ( n3153 & ~n3158 ) ;
  assign n3160 = ( x69 & n2969 ) | ( x69 & ~n3130 ) | ( n2969 & ~n3130 ) ;
  assign n3161 = x69 & n2969 ;
  assign n3162 = ( ~n2974 & n3160 ) | ( ~n2974 & n3161 ) | ( n3160 & n3161 ) ;
  assign n3163 = ( n2974 & n3160 ) | ( n2974 & n3161 ) | ( n3160 & n3161 ) ;
  assign n3164 = ( n2974 & n3162 ) | ( n2974 & ~n3163 ) | ( n3162 & ~n3163 ) ;
  assign n3165 = ( x70 & n3159 ) | ( x70 & ~n3164 ) | ( n3159 & ~n3164 ) ;
  assign n3166 = ( x70 & n2975 ) | ( x70 & ~n3130 ) | ( n2975 & ~n3130 ) ;
  assign n3167 = x70 & n2975 ;
  assign n3168 = ( n2980 & n3166 ) | ( n2980 & n3167 ) | ( n3166 & n3167 ) ;
  assign n3169 = ( ~n2980 & n3166 ) | ( ~n2980 & n3167 ) | ( n3166 & n3167 ) ;
  assign n3170 = ( n2980 & ~n3168 ) | ( n2980 & n3169 ) | ( ~n3168 & n3169 ) ;
  assign n3171 = ( x71 & n3165 ) | ( x71 & ~n3170 ) | ( n3165 & ~n3170 ) ;
  assign n3172 = ( x71 & n2981 ) | ( x71 & ~n3130 ) | ( n2981 & ~n3130 ) ;
  assign n3173 = x71 & n2981 ;
  assign n3174 = ( ~n2986 & n3172 ) | ( ~n2986 & n3173 ) | ( n3172 & n3173 ) ;
  assign n3175 = ( n2986 & n3172 ) | ( n2986 & n3173 ) | ( n3172 & n3173 ) ;
  assign n3176 = ( n2986 & n3174 ) | ( n2986 & ~n3175 ) | ( n3174 & ~n3175 ) ;
  assign n3177 = ( x72 & n3171 ) | ( x72 & ~n3176 ) | ( n3171 & ~n3176 ) ;
  assign n3178 = ( x72 & n2987 ) | ( x72 & ~n3130 ) | ( n2987 & ~n3130 ) ;
  assign n3179 = x72 & n2987 ;
  assign n3180 = ( n2992 & n3178 ) | ( n2992 & n3179 ) | ( n3178 & n3179 ) ;
  assign n3181 = ( ~n2992 & n3178 ) | ( ~n2992 & n3179 ) | ( n3178 & n3179 ) ;
  assign n3182 = ( n2992 & ~n3180 ) | ( n2992 & n3181 ) | ( ~n3180 & n3181 ) ;
  assign n3183 = ( x73 & n3177 ) | ( x73 & ~n3182 ) | ( n3177 & ~n3182 ) ;
  assign n3184 = ( x73 & n2993 ) | ( x73 & ~n3130 ) | ( n2993 & ~n3130 ) ;
  assign n3185 = x73 & n2993 ;
  assign n3186 = ( ~n2998 & n3184 ) | ( ~n2998 & n3185 ) | ( n3184 & n3185 ) ;
  assign n3187 = ( n2998 & n3184 ) | ( n2998 & n3185 ) | ( n3184 & n3185 ) ;
  assign n3188 = ( n2998 & n3186 ) | ( n2998 & ~n3187 ) | ( n3186 & ~n3187 ) ;
  assign n3189 = ( x74 & n3183 ) | ( x74 & ~n3188 ) | ( n3183 & ~n3188 ) ;
  assign n3190 = ( x74 & n2999 ) | ( x74 & ~n3130 ) | ( n2999 & ~n3130 ) ;
  assign n3191 = x74 & n2999 ;
  assign n3192 = ( n3004 & n3190 ) | ( n3004 & n3191 ) | ( n3190 & n3191 ) ;
  assign n3193 = ( ~n3004 & n3190 ) | ( ~n3004 & n3191 ) | ( n3190 & n3191 ) ;
  assign n3194 = ( n3004 & ~n3192 ) | ( n3004 & n3193 ) | ( ~n3192 & n3193 ) ;
  assign n3195 = ( x75 & n3189 ) | ( x75 & ~n3194 ) | ( n3189 & ~n3194 ) ;
  assign n3196 = ( x75 & n3005 ) | ( x75 & ~n3130 ) | ( n3005 & ~n3130 ) ;
  assign n3197 = x75 & n3005 ;
  assign n3198 = ( ~n3010 & n3196 ) | ( ~n3010 & n3197 ) | ( n3196 & n3197 ) ;
  assign n3199 = ( n3010 & n3196 ) | ( n3010 & n3197 ) | ( n3196 & n3197 ) ;
  assign n3200 = ( n3010 & n3198 ) | ( n3010 & ~n3199 ) | ( n3198 & ~n3199 ) ;
  assign n3201 = ( x76 & n3195 ) | ( x76 & ~n3200 ) | ( n3195 & ~n3200 ) ;
  assign n3202 = ( x76 & n3011 ) | ( x76 & ~n3130 ) | ( n3011 & ~n3130 ) ;
  assign n3203 = x76 & n3011 ;
  assign n3204 = ( n3016 & n3202 ) | ( n3016 & n3203 ) | ( n3202 & n3203 ) ;
  assign n3205 = ( ~n3016 & n3202 ) | ( ~n3016 & n3203 ) | ( n3202 & n3203 ) ;
  assign n3206 = ( n3016 & ~n3204 ) | ( n3016 & n3205 ) | ( ~n3204 & n3205 ) ;
  assign n3207 = ( x77 & n3201 ) | ( x77 & ~n3206 ) | ( n3201 & ~n3206 ) ;
  assign n3208 = ( x77 & n3017 ) | ( x77 & ~n3130 ) | ( n3017 & ~n3130 ) ;
  assign n3209 = x77 & n3017 ;
  assign n3210 = ( ~n3022 & n3208 ) | ( ~n3022 & n3209 ) | ( n3208 & n3209 ) ;
  assign n3211 = ( n3022 & n3208 ) | ( n3022 & n3209 ) | ( n3208 & n3209 ) ;
  assign n3212 = ( n3022 & n3210 ) | ( n3022 & ~n3211 ) | ( n3210 & ~n3211 ) ;
  assign n3213 = ( x78 & n3207 ) | ( x78 & ~n3212 ) | ( n3207 & ~n3212 ) ;
  assign n3214 = ( x78 & n3023 ) | ( x78 & ~n3130 ) | ( n3023 & ~n3130 ) ;
  assign n3215 = x78 & n3023 ;
  assign n3216 = ( n3028 & n3214 ) | ( n3028 & n3215 ) | ( n3214 & n3215 ) ;
  assign n3217 = ( ~n3028 & n3214 ) | ( ~n3028 & n3215 ) | ( n3214 & n3215 ) ;
  assign n3218 = ( n3028 & ~n3216 ) | ( n3028 & n3217 ) | ( ~n3216 & n3217 ) ;
  assign n3219 = ( x79 & n3213 ) | ( x79 & ~n3218 ) | ( n3213 & ~n3218 ) ;
  assign n3220 = ( x79 & n3029 ) | ( x79 & ~n3130 ) | ( n3029 & ~n3130 ) ;
  assign n3221 = x79 & n3029 ;
  assign n3222 = ( ~n3034 & n3220 ) | ( ~n3034 & n3221 ) | ( n3220 & n3221 ) ;
  assign n3223 = ( n3034 & n3220 ) | ( n3034 & n3221 ) | ( n3220 & n3221 ) ;
  assign n3224 = ( n3034 & n3222 ) | ( n3034 & ~n3223 ) | ( n3222 & ~n3223 ) ;
  assign n3225 = ( x80 & n3219 ) | ( x80 & ~n3224 ) | ( n3219 & ~n3224 ) ;
  assign n3226 = ( x80 & n3035 ) | ( x80 & ~n3130 ) | ( n3035 & ~n3130 ) ;
  assign n3227 = x80 & n3035 ;
  assign n3228 = ( n3040 & n3226 ) | ( n3040 & n3227 ) | ( n3226 & n3227 ) ;
  assign n3229 = ( ~n3040 & n3226 ) | ( ~n3040 & n3227 ) | ( n3226 & n3227 ) ;
  assign n3230 = ( n3040 & ~n3228 ) | ( n3040 & n3229 ) | ( ~n3228 & n3229 ) ;
  assign n3231 = ( x81 & n3225 ) | ( x81 & ~n3230 ) | ( n3225 & ~n3230 ) ;
  assign n3232 = ( x81 & n3041 ) | ( x81 & ~n3130 ) | ( n3041 & ~n3130 ) ;
  assign n3233 = x81 & n3041 ;
  assign n3234 = ( ~n3046 & n3232 ) | ( ~n3046 & n3233 ) | ( n3232 & n3233 ) ;
  assign n3235 = ( n3046 & n3232 ) | ( n3046 & n3233 ) | ( n3232 & n3233 ) ;
  assign n3236 = ( n3046 & n3234 ) | ( n3046 & ~n3235 ) | ( n3234 & ~n3235 ) ;
  assign n3237 = ( x82 & n3231 ) | ( x82 & ~n3236 ) | ( n3231 & ~n3236 ) ;
  assign n3238 = ( x82 & n3047 ) | ( x82 & ~n3130 ) | ( n3047 & ~n3130 ) ;
  assign n3239 = x82 & n3047 ;
  assign n3240 = ( n3052 & n3238 ) | ( n3052 & n3239 ) | ( n3238 & n3239 ) ;
  assign n3241 = ( ~n3052 & n3238 ) | ( ~n3052 & n3239 ) | ( n3238 & n3239 ) ;
  assign n3242 = ( n3052 & ~n3240 ) | ( n3052 & n3241 ) | ( ~n3240 & n3241 ) ;
  assign n3243 = ( x83 & n3237 ) | ( x83 & ~n3242 ) | ( n3237 & ~n3242 ) ;
  assign n3244 = ( x83 & n3053 ) | ( x83 & ~n3130 ) | ( n3053 & ~n3130 ) ;
  assign n3245 = x83 & n3053 ;
  assign n3246 = ( ~n3058 & n3244 ) | ( ~n3058 & n3245 ) | ( n3244 & n3245 ) ;
  assign n3247 = ( n3058 & n3244 ) | ( n3058 & n3245 ) | ( n3244 & n3245 ) ;
  assign n3248 = ( n3058 & n3246 ) | ( n3058 & ~n3247 ) | ( n3246 & ~n3247 ) ;
  assign n3249 = ( x84 & n3243 ) | ( x84 & ~n3248 ) | ( n3243 & ~n3248 ) ;
  assign n3250 = ( x84 & n3059 ) | ( x84 & ~n3130 ) | ( n3059 & ~n3130 ) ;
  assign n3251 = x84 & n3059 ;
  assign n3252 = ( n3064 & n3250 ) | ( n3064 & n3251 ) | ( n3250 & n3251 ) ;
  assign n3253 = ( ~n3064 & n3250 ) | ( ~n3064 & n3251 ) | ( n3250 & n3251 ) ;
  assign n3254 = ( n3064 & ~n3252 ) | ( n3064 & n3253 ) | ( ~n3252 & n3253 ) ;
  assign n3255 = ( x85 & n3249 ) | ( x85 & ~n3254 ) | ( n3249 & ~n3254 ) ;
  assign n3256 = ( x85 & n3065 ) | ( x85 & ~n3130 ) | ( n3065 & ~n3130 ) ;
  assign n3257 = x85 & n3065 ;
  assign n3258 = ( ~n3070 & n3256 ) | ( ~n3070 & n3257 ) | ( n3256 & n3257 ) ;
  assign n3259 = ( n3070 & n3256 ) | ( n3070 & n3257 ) | ( n3256 & n3257 ) ;
  assign n3260 = ( n3070 & n3258 ) | ( n3070 & ~n3259 ) | ( n3258 & ~n3259 ) ;
  assign n3261 = ( x86 & n3255 ) | ( x86 & ~n3260 ) | ( n3255 & ~n3260 ) ;
  assign n3262 = ( x86 & n3071 ) | ( x86 & ~n3130 ) | ( n3071 & ~n3130 ) ;
  assign n3263 = x86 & n3071 ;
  assign n3264 = ( n3076 & n3262 ) | ( n3076 & n3263 ) | ( n3262 & n3263 ) ;
  assign n3265 = ( ~n3076 & n3262 ) | ( ~n3076 & n3263 ) | ( n3262 & n3263 ) ;
  assign n3266 = ( n3076 & ~n3264 ) | ( n3076 & n3265 ) | ( ~n3264 & n3265 ) ;
  assign n3267 = ( x87 & n3261 ) | ( x87 & ~n3266 ) | ( n3261 & ~n3266 ) ;
  assign n3268 = ( x87 & n3077 ) | ( x87 & ~n3130 ) | ( n3077 & ~n3130 ) ;
  assign n3269 = x87 & n3077 ;
  assign n3270 = ( ~n3082 & n3268 ) | ( ~n3082 & n3269 ) | ( n3268 & n3269 ) ;
  assign n3271 = ( n3082 & n3268 ) | ( n3082 & n3269 ) | ( n3268 & n3269 ) ;
  assign n3272 = ( n3082 & n3270 ) | ( n3082 & ~n3271 ) | ( n3270 & ~n3271 ) ;
  assign n3273 = ( x88 & n3267 ) | ( x88 & ~n3272 ) | ( n3267 & ~n3272 ) ;
  assign n3274 = ( x88 & n3083 ) | ( x88 & ~n3130 ) | ( n3083 & ~n3130 ) ;
  assign n3275 = x88 & n3083 ;
  assign n3276 = ( n3088 & n3274 ) | ( n3088 & n3275 ) | ( n3274 & n3275 ) ;
  assign n3277 = ( ~n3088 & n3274 ) | ( ~n3088 & n3275 ) | ( n3274 & n3275 ) ;
  assign n3278 = ( n3088 & ~n3276 ) | ( n3088 & n3277 ) | ( ~n3276 & n3277 ) ;
  assign n3279 = ( x89 & n3273 ) | ( x89 & ~n3278 ) | ( n3273 & ~n3278 ) ;
  assign n3280 = ( x89 & n3089 ) | ( x89 & ~n3130 ) | ( n3089 & ~n3130 ) ;
  assign n3281 = x89 & n3089 ;
  assign n3282 = ( ~n3094 & n3280 ) | ( ~n3094 & n3281 ) | ( n3280 & n3281 ) ;
  assign n3283 = ( n3094 & n3280 ) | ( n3094 & n3281 ) | ( n3280 & n3281 ) ;
  assign n3284 = ( n3094 & n3282 ) | ( n3094 & ~n3283 ) | ( n3282 & ~n3283 ) ;
  assign n3285 = ( x90 & n3279 ) | ( x90 & ~n3284 ) | ( n3279 & ~n3284 ) ;
  assign n3286 = ( x90 & n3095 ) | ( x90 & ~n3130 ) | ( n3095 & ~n3130 ) ;
  assign n3287 = x90 & n3095 ;
  assign n3288 = ( n3100 & n3286 ) | ( n3100 & n3287 ) | ( n3286 & n3287 ) ;
  assign n3289 = ( ~n3100 & n3286 ) | ( ~n3100 & n3287 ) | ( n3286 & n3287 ) ;
  assign n3290 = ( n3100 & ~n3288 ) | ( n3100 & n3289 ) | ( ~n3288 & n3289 ) ;
  assign n3291 = ( x91 & n3285 ) | ( x91 & ~n3290 ) | ( n3285 & ~n3290 ) ;
  assign n3292 = ( x91 & n3101 ) | ( x91 & ~n3130 ) | ( n3101 & ~n3130 ) ;
  assign n3293 = x91 & n3101 ;
  assign n3294 = ( ~n3106 & n3292 ) | ( ~n3106 & n3293 ) | ( n3292 & n3293 ) ;
  assign n3295 = ( n3106 & n3292 ) | ( n3106 & n3293 ) | ( n3292 & n3293 ) ;
  assign n3296 = ( n3106 & n3294 ) | ( n3106 & ~n3295 ) | ( n3294 & ~n3295 ) ;
  assign n3297 = ( x92 & n3291 ) | ( x92 & ~n3296 ) | ( n3291 & ~n3296 ) ;
  assign n3298 = ( x92 & n3107 ) | ( x92 & ~n3130 ) | ( n3107 & ~n3130 ) ;
  assign n3299 = x92 & n3107 ;
  assign n3300 = ( n3112 & n3298 ) | ( n3112 & n3299 ) | ( n3298 & n3299 ) ;
  assign n3301 = ( ~n3112 & n3298 ) | ( ~n3112 & n3299 ) | ( n3298 & n3299 ) ;
  assign n3302 = ( n3112 & ~n3300 ) | ( n3112 & n3301 ) | ( ~n3300 & n3301 ) ;
  assign n3303 = ( x93 & n3297 ) | ( x93 & ~n3302 ) | ( n3297 & ~n3302 ) ;
  assign n3304 = ( x93 & n3113 ) | ( x93 & ~n3130 ) | ( n3113 & ~n3130 ) ;
  assign n3305 = x93 & n3113 ;
  assign n3306 = ( ~n3118 & n3304 ) | ( ~n3118 & n3305 ) | ( n3304 & n3305 ) ;
  assign n3307 = ( n3118 & n3304 ) | ( n3118 & n3305 ) | ( n3304 & n3305 ) ;
  assign n3308 = ( n3118 & n3306 ) | ( n3118 & ~n3307 ) | ( n3306 & ~n3307 ) ;
  assign n3309 = ( x94 & n3303 ) | ( x94 & ~n3308 ) | ( n3303 & ~n3308 ) ;
  assign n3310 = ( x94 & n3119 ) | ( x94 & ~n3130 ) | ( n3119 & ~n3130 ) ;
  assign n3311 = x94 & n3119 ;
  assign n3312 = ( ~n3124 & n3310 ) | ( ~n3124 & n3311 ) | ( n3310 & n3311 ) ;
  assign n3313 = ( n3124 & n3310 ) | ( n3124 & n3311 ) | ( n3310 & n3311 ) ;
  assign n3314 = ( n3124 & n3312 ) | ( n3124 & ~n3313 ) | ( n3312 & ~n3313 ) ;
  assign n3315 = ( x95 & n3309 ) | ( x95 & ~n3314 ) | ( n3309 & ~n3314 ) ;
  assign n3316 = ( x96 & ~n3128 ) | ( x96 & n3315 ) | ( ~n3128 & n3315 ) ;
  assign n3317 = n161 | n3316 ;
  assign n3318 = n3128 & n3317 ;
  assign n3319 = n280 | n3318 ;
  assign n3320 = ( x31 & ~x64 ) | ( x31 & n3317 ) | ( ~x64 & n3317 ) ;
  assign n3321 = ~x31 & n3317 ;
  assign n3322 = ( n3134 & n3320 ) | ( n3134 & ~n3321 ) | ( n3320 & ~n3321 ) ;
  assign n3323 = ~x30 & x64 ;
  assign n3324 = ( x65 & ~n3322 ) | ( x65 & n3323 ) | ( ~n3322 & n3323 ) ;
  assign n3325 = ( x65 & n3134 ) | ( x65 & ~n3317 ) | ( n3134 & ~n3317 ) ;
  assign n3326 = x65 & n3134 ;
  assign n3327 = ( n3133 & n3325 ) | ( n3133 & n3326 ) | ( n3325 & n3326 ) ;
  assign n3328 = ( ~n3133 & n3325 ) | ( ~n3133 & n3326 ) | ( n3325 & n3326 ) ;
  assign n3329 = ( n3133 & ~n3327 ) | ( n3133 & n3328 ) | ( ~n3327 & n3328 ) ;
  assign n3330 = ( x66 & n3324 ) | ( x66 & ~n3329 ) | ( n3324 & ~n3329 ) ;
  assign n3331 = ( x66 & n3135 ) | ( x66 & ~n3317 ) | ( n3135 & ~n3317 ) ;
  assign n3332 = x66 & n3135 ;
  assign n3333 = ( n3140 & n3331 ) | ( n3140 & n3332 ) | ( n3331 & n3332 ) ;
  assign n3334 = ( ~n3140 & n3331 ) | ( ~n3140 & n3332 ) | ( n3331 & n3332 ) ;
  assign n3335 = ( n3140 & ~n3333 ) | ( n3140 & n3334 ) | ( ~n3333 & n3334 ) ;
  assign n3336 = ( x67 & n3330 ) | ( x67 & ~n3335 ) | ( n3330 & ~n3335 ) ;
  assign n3337 = ( x67 & n3141 ) | ( x67 & ~n3317 ) | ( n3141 & ~n3317 ) ;
  assign n3338 = x67 & n3141 ;
  assign n3339 = ( ~n3146 & n3337 ) | ( ~n3146 & n3338 ) | ( n3337 & n3338 ) ;
  assign n3340 = ( n3146 & n3337 ) | ( n3146 & n3338 ) | ( n3337 & n3338 ) ;
  assign n3341 = ( n3146 & n3339 ) | ( n3146 & ~n3340 ) | ( n3339 & ~n3340 ) ;
  assign n3342 = ( x68 & n3336 ) | ( x68 & ~n3341 ) | ( n3336 & ~n3341 ) ;
  assign n3343 = ( x68 & n3147 ) | ( x68 & ~n3317 ) | ( n3147 & ~n3317 ) ;
  assign n3344 = x68 & n3147 ;
  assign n3345 = ( n3152 & n3343 ) | ( n3152 & n3344 ) | ( n3343 & n3344 ) ;
  assign n3346 = ( ~n3152 & n3343 ) | ( ~n3152 & n3344 ) | ( n3343 & n3344 ) ;
  assign n3347 = ( n3152 & ~n3345 ) | ( n3152 & n3346 ) | ( ~n3345 & n3346 ) ;
  assign n3348 = ( x69 & n3342 ) | ( x69 & ~n3347 ) | ( n3342 & ~n3347 ) ;
  assign n3349 = ( x69 & n3153 ) | ( x69 & ~n3317 ) | ( n3153 & ~n3317 ) ;
  assign n3350 = x69 & n3153 ;
  assign n3351 = ( ~n3158 & n3349 ) | ( ~n3158 & n3350 ) | ( n3349 & n3350 ) ;
  assign n3352 = ( n3158 & n3349 ) | ( n3158 & n3350 ) | ( n3349 & n3350 ) ;
  assign n3353 = ( n3158 & n3351 ) | ( n3158 & ~n3352 ) | ( n3351 & ~n3352 ) ;
  assign n3354 = ( x70 & n3348 ) | ( x70 & ~n3353 ) | ( n3348 & ~n3353 ) ;
  assign n3355 = ( x70 & n3159 ) | ( x70 & ~n3317 ) | ( n3159 & ~n3317 ) ;
  assign n3356 = x70 & n3159 ;
  assign n3357 = ( n3164 & n3355 ) | ( n3164 & n3356 ) | ( n3355 & n3356 ) ;
  assign n3358 = ( ~n3164 & n3355 ) | ( ~n3164 & n3356 ) | ( n3355 & n3356 ) ;
  assign n3359 = ( n3164 & ~n3357 ) | ( n3164 & n3358 ) | ( ~n3357 & n3358 ) ;
  assign n3360 = ( x71 & n3354 ) | ( x71 & ~n3359 ) | ( n3354 & ~n3359 ) ;
  assign n3361 = ( x71 & n3165 ) | ( x71 & ~n3317 ) | ( n3165 & ~n3317 ) ;
  assign n3362 = x71 & n3165 ;
  assign n3363 = ( ~n3170 & n3361 ) | ( ~n3170 & n3362 ) | ( n3361 & n3362 ) ;
  assign n3364 = ( n3170 & n3361 ) | ( n3170 & n3362 ) | ( n3361 & n3362 ) ;
  assign n3365 = ( n3170 & n3363 ) | ( n3170 & ~n3364 ) | ( n3363 & ~n3364 ) ;
  assign n3366 = ( x72 & n3360 ) | ( x72 & ~n3365 ) | ( n3360 & ~n3365 ) ;
  assign n3367 = ( x72 & n3171 ) | ( x72 & ~n3317 ) | ( n3171 & ~n3317 ) ;
  assign n3368 = x72 & n3171 ;
  assign n3369 = ( n3176 & n3367 ) | ( n3176 & n3368 ) | ( n3367 & n3368 ) ;
  assign n3370 = ( ~n3176 & n3367 ) | ( ~n3176 & n3368 ) | ( n3367 & n3368 ) ;
  assign n3371 = ( n3176 & ~n3369 ) | ( n3176 & n3370 ) | ( ~n3369 & n3370 ) ;
  assign n3372 = ( x73 & n3366 ) | ( x73 & ~n3371 ) | ( n3366 & ~n3371 ) ;
  assign n3373 = ( x73 & n3177 ) | ( x73 & ~n3317 ) | ( n3177 & ~n3317 ) ;
  assign n3374 = x73 & n3177 ;
  assign n3375 = ( ~n3182 & n3373 ) | ( ~n3182 & n3374 ) | ( n3373 & n3374 ) ;
  assign n3376 = ( n3182 & n3373 ) | ( n3182 & n3374 ) | ( n3373 & n3374 ) ;
  assign n3377 = ( n3182 & n3375 ) | ( n3182 & ~n3376 ) | ( n3375 & ~n3376 ) ;
  assign n3378 = ( x74 & n3372 ) | ( x74 & ~n3377 ) | ( n3372 & ~n3377 ) ;
  assign n3379 = ( x74 & n3183 ) | ( x74 & ~n3317 ) | ( n3183 & ~n3317 ) ;
  assign n3380 = x74 & n3183 ;
  assign n3381 = ( n3188 & n3379 ) | ( n3188 & n3380 ) | ( n3379 & n3380 ) ;
  assign n3382 = ( ~n3188 & n3379 ) | ( ~n3188 & n3380 ) | ( n3379 & n3380 ) ;
  assign n3383 = ( n3188 & ~n3381 ) | ( n3188 & n3382 ) | ( ~n3381 & n3382 ) ;
  assign n3384 = ( x75 & n3378 ) | ( x75 & ~n3383 ) | ( n3378 & ~n3383 ) ;
  assign n3385 = ( x75 & n3189 ) | ( x75 & ~n3317 ) | ( n3189 & ~n3317 ) ;
  assign n3386 = x75 & n3189 ;
  assign n3387 = ( ~n3194 & n3385 ) | ( ~n3194 & n3386 ) | ( n3385 & n3386 ) ;
  assign n3388 = ( n3194 & n3385 ) | ( n3194 & n3386 ) | ( n3385 & n3386 ) ;
  assign n3389 = ( n3194 & n3387 ) | ( n3194 & ~n3388 ) | ( n3387 & ~n3388 ) ;
  assign n3390 = ( x76 & n3384 ) | ( x76 & ~n3389 ) | ( n3384 & ~n3389 ) ;
  assign n3391 = ( x76 & n3195 ) | ( x76 & ~n3317 ) | ( n3195 & ~n3317 ) ;
  assign n3392 = x76 & n3195 ;
  assign n3393 = ( n3200 & n3391 ) | ( n3200 & n3392 ) | ( n3391 & n3392 ) ;
  assign n3394 = ( ~n3200 & n3391 ) | ( ~n3200 & n3392 ) | ( n3391 & n3392 ) ;
  assign n3395 = ( n3200 & ~n3393 ) | ( n3200 & n3394 ) | ( ~n3393 & n3394 ) ;
  assign n3396 = ( x77 & n3390 ) | ( x77 & ~n3395 ) | ( n3390 & ~n3395 ) ;
  assign n3397 = ( x77 & n3201 ) | ( x77 & ~n3317 ) | ( n3201 & ~n3317 ) ;
  assign n3398 = x77 & n3201 ;
  assign n3399 = ( ~n3206 & n3397 ) | ( ~n3206 & n3398 ) | ( n3397 & n3398 ) ;
  assign n3400 = ( n3206 & n3397 ) | ( n3206 & n3398 ) | ( n3397 & n3398 ) ;
  assign n3401 = ( n3206 & n3399 ) | ( n3206 & ~n3400 ) | ( n3399 & ~n3400 ) ;
  assign n3402 = ( x78 & n3396 ) | ( x78 & ~n3401 ) | ( n3396 & ~n3401 ) ;
  assign n3403 = ( x78 & n3207 ) | ( x78 & ~n3317 ) | ( n3207 & ~n3317 ) ;
  assign n3404 = x78 & n3207 ;
  assign n3405 = ( n3212 & n3403 ) | ( n3212 & n3404 ) | ( n3403 & n3404 ) ;
  assign n3406 = ( ~n3212 & n3403 ) | ( ~n3212 & n3404 ) | ( n3403 & n3404 ) ;
  assign n3407 = ( n3212 & ~n3405 ) | ( n3212 & n3406 ) | ( ~n3405 & n3406 ) ;
  assign n3408 = ( x79 & n3402 ) | ( x79 & ~n3407 ) | ( n3402 & ~n3407 ) ;
  assign n3409 = ( x79 & n3213 ) | ( x79 & ~n3317 ) | ( n3213 & ~n3317 ) ;
  assign n3410 = x79 & n3213 ;
  assign n3411 = ( ~n3218 & n3409 ) | ( ~n3218 & n3410 ) | ( n3409 & n3410 ) ;
  assign n3412 = ( n3218 & n3409 ) | ( n3218 & n3410 ) | ( n3409 & n3410 ) ;
  assign n3413 = ( n3218 & n3411 ) | ( n3218 & ~n3412 ) | ( n3411 & ~n3412 ) ;
  assign n3414 = ( x80 & n3408 ) | ( x80 & ~n3413 ) | ( n3408 & ~n3413 ) ;
  assign n3415 = ( x80 & n3219 ) | ( x80 & ~n3317 ) | ( n3219 & ~n3317 ) ;
  assign n3416 = x80 & n3219 ;
  assign n3417 = ( n3224 & n3415 ) | ( n3224 & n3416 ) | ( n3415 & n3416 ) ;
  assign n3418 = ( ~n3224 & n3415 ) | ( ~n3224 & n3416 ) | ( n3415 & n3416 ) ;
  assign n3419 = ( n3224 & ~n3417 ) | ( n3224 & n3418 ) | ( ~n3417 & n3418 ) ;
  assign n3420 = ( x81 & n3414 ) | ( x81 & ~n3419 ) | ( n3414 & ~n3419 ) ;
  assign n3421 = ( x81 & n3225 ) | ( x81 & ~n3317 ) | ( n3225 & ~n3317 ) ;
  assign n3422 = x81 & n3225 ;
  assign n3423 = ( ~n3230 & n3421 ) | ( ~n3230 & n3422 ) | ( n3421 & n3422 ) ;
  assign n3424 = ( n3230 & n3421 ) | ( n3230 & n3422 ) | ( n3421 & n3422 ) ;
  assign n3425 = ( n3230 & n3423 ) | ( n3230 & ~n3424 ) | ( n3423 & ~n3424 ) ;
  assign n3426 = ( x82 & n3420 ) | ( x82 & ~n3425 ) | ( n3420 & ~n3425 ) ;
  assign n3427 = ( x82 & n3231 ) | ( x82 & ~n3317 ) | ( n3231 & ~n3317 ) ;
  assign n3428 = x82 & n3231 ;
  assign n3429 = ( n3236 & n3427 ) | ( n3236 & n3428 ) | ( n3427 & n3428 ) ;
  assign n3430 = ( ~n3236 & n3427 ) | ( ~n3236 & n3428 ) | ( n3427 & n3428 ) ;
  assign n3431 = ( n3236 & ~n3429 ) | ( n3236 & n3430 ) | ( ~n3429 & n3430 ) ;
  assign n3432 = ( x83 & n3426 ) | ( x83 & ~n3431 ) | ( n3426 & ~n3431 ) ;
  assign n3433 = ( x83 & n3237 ) | ( x83 & ~n3317 ) | ( n3237 & ~n3317 ) ;
  assign n3434 = x83 & n3237 ;
  assign n3435 = ( ~n3242 & n3433 ) | ( ~n3242 & n3434 ) | ( n3433 & n3434 ) ;
  assign n3436 = ( n3242 & n3433 ) | ( n3242 & n3434 ) | ( n3433 & n3434 ) ;
  assign n3437 = ( n3242 & n3435 ) | ( n3242 & ~n3436 ) | ( n3435 & ~n3436 ) ;
  assign n3438 = ( x84 & n3432 ) | ( x84 & ~n3437 ) | ( n3432 & ~n3437 ) ;
  assign n3439 = ( x84 & n3243 ) | ( x84 & ~n3317 ) | ( n3243 & ~n3317 ) ;
  assign n3440 = x84 & n3243 ;
  assign n3441 = ( n3248 & n3439 ) | ( n3248 & n3440 ) | ( n3439 & n3440 ) ;
  assign n3442 = ( ~n3248 & n3439 ) | ( ~n3248 & n3440 ) | ( n3439 & n3440 ) ;
  assign n3443 = ( n3248 & ~n3441 ) | ( n3248 & n3442 ) | ( ~n3441 & n3442 ) ;
  assign n3444 = ( x85 & n3438 ) | ( x85 & ~n3443 ) | ( n3438 & ~n3443 ) ;
  assign n3445 = ( x85 & n3249 ) | ( x85 & ~n3317 ) | ( n3249 & ~n3317 ) ;
  assign n3446 = x85 & n3249 ;
  assign n3447 = ( ~n3254 & n3445 ) | ( ~n3254 & n3446 ) | ( n3445 & n3446 ) ;
  assign n3448 = ( n3254 & n3445 ) | ( n3254 & n3446 ) | ( n3445 & n3446 ) ;
  assign n3449 = ( n3254 & n3447 ) | ( n3254 & ~n3448 ) | ( n3447 & ~n3448 ) ;
  assign n3450 = ( x86 & n3444 ) | ( x86 & ~n3449 ) | ( n3444 & ~n3449 ) ;
  assign n3451 = ( x86 & n3255 ) | ( x86 & ~n3317 ) | ( n3255 & ~n3317 ) ;
  assign n3452 = x86 & n3255 ;
  assign n3453 = ( n3260 & n3451 ) | ( n3260 & n3452 ) | ( n3451 & n3452 ) ;
  assign n3454 = ( ~n3260 & n3451 ) | ( ~n3260 & n3452 ) | ( n3451 & n3452 ) ;
  assign n3455 = ( n3260 & ~n3453 ) | ( n3260 & n3454 ) | ( ~n3453 & n3454 ) ;
  assign n3456 = ( x87 & n3450 ) | ( x87 & ~n3455 ) | ( n3450 & ~n3455 ) ;
  assign n3457 = ( x87 & n3261 ) | ( x87 & ~n3317 ) | ( n3261 & ~n3317 ) ;
  assign n3458 = x87 & n3261 ;
  assign n3459 = ( ~n3266 & n3457 ) | ( ~n3266 & n3458 ) | ( n3457 & n3458 ) ;
  assign n3460 = ( n3266 & n3457 ) | ( n3266 & n3458 ) | ( n3457 & n3458 ) ;
  assign n3461 = ( n3266 & n3459 ) | ( n3266 & ~n3460 ) | ( n3459 & ~n3460 ) ;
  assign n3462 = ( x88 & n3456 ) | ( x88 & ~n3461 ) | ( n3456 & ~n3461 ) ;
  assign n3463 = ( x88 & n3267 ) | ( x88 & ~n3317 ) | ( n3267 & ~n3317 ) ;
  assign n3464 = x88 & n3267 ;
  assign n3465 = ( n3272 & n3463 ) | ( n3272 & n3464 ) | ( n3463 & n3464 ) ;
  assign n3466 = ( ~n3272 & n3463 ) | ( ~n3272 & n3464 ) | ( n3463 & n3464 ) ;
  assign n3467 = ( n3272 & ~n3465 ) | ( n3272 & n3466 ) | ( ~n3465 & n3466 ) ;
  assign n3468 = ( x89 & n3462 ) | ( x89 & ~n3467 ) | ( n3462 & ~n3467 ) ;
  assign n3469 = ( x89 & n3273 ) | ( x89 & ~n3317 ) | ( n3273 & ~n3317 ) ;
  assign n3470 = x89 & n3273 ;
  assign n3471 = ( ~n3278 & n3469 ) | ( ~n3278 & n3470 ) | ( n3469 & n3470 ) ;
  assign n3472 = ( n3278 & n3469 ) | ( n3278 & n3470 ) | ( n3469 & n3470 ) ;
  assign n3473 = ( n3278 & n3471 ) | ( n3278 & ~n3472 ) | ( n3471 & ~n3472 ) ;
  assign n3474 = ( x90 & n3468 ) | ( x90 & ~n3473 ) | ( n3468 & ~n3473 ) ;
  assign n3475 = ( x90 & n3279 ) | ( x90 & ~n3317 ) | ( n3279 & ~n3317 ) ;
  assign n3476 = x90 & n3279 ;
  assign n3477 = ( n3284 & n3475 ) | ( n3284 & n3476 ) | ( n3475 & n3476 ) ;
  assign n3478 = ( ~n3284 & n3475 ) | ( ~n3284 & n3476 ) | ( n3475 & n3476 ) ;
  assign n3479 = ( n3284 & ~n3477 ) | ( n3284 & n3478 ) | ( ~n3477 & n3478 ) ;
  assign n3480 = ( x91 & n3474 ) | ( x91 & ~n3479 ) | ( n3474 & ~n3479 ) ;
  assign n3481 = ( x91 & n3285 ) | ( x91 & ~n3317 ) | ( n3285 & ~n3317 ) ;
  assign n3482 = x91 & n3285 ;
  assign n3483 = ( ~n3290 & n3481 ) | ( ~n3290 & n3482 ) | ( n3481 & n3482 ) ;
  assign n3484 = ( n3290 & n3481 ) | ( n3290 & n3482 ) | ( n3481 & n3482 ) ;
  assign n3485 = ( n3290 & n3483 ) | ( n3290 & ~n3484 ) | ( n3483 & ~n3484 ) ;
  assign n3486 = ( x92 & n3480 ) | ( x92 & ~n3485 ) | ( n3480 & ~n3485 ) ;
  assign n3487 = ( x92 & n3291 ) | ( x92 & ~n3317 ) | ( n3291 & ~n3317 ) ;
  assign n3488 = x92 & n3291 ;
  assign n3489 = ( n3296 & n3487 ) | ( n3296 & n3488 ) | ( n3487 & n3488 ) ;
  assign n3490 = ( ~n3296 & n3487 ) | ( ~n3296 & n3488 ) | ( n3487 & n3488 ) ;
  assign n3491 = ( n3296 & ~n3489 ) | ( n3296 & n3490 ) | ( ~n3489 & n3490 ) ;
  assign n3492 = ( x93 & n3486 ) | ( x93 & ~n3491 ) | ( n3486 & ~n3491 ) ;
  assign n3493 = ( x93 & n3297 ) | ( x93 & ~n3317 ) | ( n3297 & ~n3317 ) ;
  assign n3494 = x93 & n3297 ;
  assign n3495 = ( ~n3302 & n3493 ) | ( ~n3302 & n3494 ) | ( n3493 & n3494 ) ;
  assign n3496 = ( n3302 & n3493 ) | ( n3302 & n3494 ) | ( n3493 & n3494 ) ;
  assign n3497 = ( n3302 & n3495 ) | ( n3302 & ~n3496 ) | ( n3495 & ~n3496 ) ;
  assign n3498 = ( x94 & n3492 ) | ( x94 & ~n3497 ) | ( n3492 & ~n3497 ) ;
  assign n3499 = ( x94 & n3303 ) | ( x94 & ~n3317 ) | ( n3303 & ~n3317 ) ;
  assign n3500 = x94 & n3303 ;
  assign n3501 = ( n3308 & n3499 ) | ( n3308 & n3500 ) | ( n3499 & n3500 ) ;
  assign n3502 = ( ~n3308 & n3499 ) | ( ~n3308 & n3500 ) | ( n3499 & n3500 ) ;
  assign n3503 = ( n3308 & ~n3501 ) | ( n3308 & n3502 ) | ( ~n3501 & n3502 ) ;
  assign n3504 = ( x95 & n3498 ) | ( x95 & ~n3503 ) | ( n3498 & ~n3503 ) ;
  assign n3505 = ( x95 & n3309 ) | ( x95 & ~n3317 ) | ( n3309 & ~n3317 ) ;
  assign n3506 = x95 & n3309 ;
  assign n3507 = ( n3314 & n3505 ) | ( n3314 & n3506 ) | ( n3505 & n3506 ) ;
  assign n3508 = ( ~n3314 & n3505 ) | ( ~n3314 & n3506 ) | ( n3505 & n3506 ) ;
  assign n3509 = ( n3314 & ~n3507 ) | ( n3314 & n3508 ) | ( ~n3507 & n3508 ) ;
  assign n3510 = ( x96 & n3504 ) | ( x96 & ~n3509 ) | ( n3504 & ~n3509 ) ;
  assign n3511 = x97 | n3510 ;
  assign n3512 = x98 | n159 ;
  assign n3513 = ( x97 & n3510 ) | ( x97 & n3512 ) | ( n3510 & n3512 ) ;
  assign n3514 = ( n3319 & ~n3511 ) | ( n3319 & n3513 ) | ( ~n3511 & n3513 ) ;
  assign n3515 = ( x97 & ~n3319 ) | ( x97 & n3510 ) | ( ~n3319 & n3510 ) ;
  assign n3516 = n3512 | n3515 ;
  assign n3517 = ( x30 & ~x64 ) | ( x30 & n3516 ) | ( ~x64 & n3516 ) ;
  assign n3518 = ~x30 & n3516 ;
  assign n3519 = ( n3323 & n3517 ) | ( n3323 & ~n3518 ) | ( n3517 & ~n3518 ) ;
  assign n3520 = ~x29 & x64 ;
  assign n3521 = ( x65 & ~n3519 ) | ( x65 & n3520 ) | ( ~n3519 & n3520 ) ;
  assign n3522 = ( x65 & n3323 ) | ( x65 & ~n3516 ) | ( n3323 & ~n3516 ) ;
  assign n3523 = x65 & n3323 ;
  assign n3524 = ( n3322 & n3522 ) | ( n3322 & n3523 ) | ( n3522 & n3523 ) ;
  assign n3525 = ( ~n3322 & n3522 ) | ( ~n3322 & n3523 ) | ( n3522 & n3523 ) ;
  assign n3526 = ( n3322 & ~n3524 ) | ( n3322 & n3525 ) | ( ~n3524 & n3525 ) ;
  assign n3527 = ( x66 & n3521 ) | ( x66 & ~n3526 ) | ( n3521 & ~n3526 ) ;
  assign n3528 = ( x66 & n3324 ) | ( x66 & ~n3516 ) | ( n3324 & ~n3516 ) ;
  assign n3529 = x66 & n3324 ;
  assign n3530 = ( n3329 & n3528 ) | ( n3329 & n3529 ) | ( n3528 & n3529 ) ;
  assign n3531 = ( ~n3329 & n3528 ) | ( ~n3329 & n3529 ) | ( n3528 & n3529 ) ;
  assign n3532 = ( n3329 & ~n3530 ) | ( n3329 & n3531 ) | ( ~n3530 & n3531 ) ;
  assign n3533 = ( x67 & n3527 ) | ( x67 & ~n3532 ) | ( n3527 & ~n3532 ) ;
  assign n3534 = ( x67 & n3330 ) | ( x67 & ~n3516 ) | ( n3330 & ~n3516 ) ;
  assign n3535 = x67 & n3330 ;
  assign n3536 = ( ~n3335 & n3534 ) | ( ~n3335 & n3535 ) | ( n3534 & n3535 ) ;
  assign n3537 = ( n3335 & n3534 ) | ( n3335 & n3535 ) | ( n3534 & n3535 ) ;
  assign n3538 = ( n3335 & n3536 ) | ( n3335 & ~n3537 ) | ( n3536 & ~n3537 ) ;
  assign n3539 = ( x68 & n3533 ) | ( x68 & ~n3538 ) | ( n3533 & ~n3538 ) ;
  assign n3540 = ( x68 & n3336 ) | ( x68 & ~n3516 ) | ( n3336 & ~n3516 ) ;
  assign n3541 = x68 & n3336 ;
  assign n3542 = ( n3341 & n3540 ) | ( n3341 & n3541 ) | ( n3540 & n3541 ) ;
  assign n3543 = ( ~n3341 & n3540 ) | ( ~n3341 & n3541 ) | ( n3540 & n3541 ) ;
  assign n3544 = ( n3341 & ~n3542 ) | ( n3341 & n3543 ) | ( ~n3542 & n3543 ) ;
  assign n3545 = ( x69 & n3539 ) | ( x69 & ~n3544 ) | ( n3539 & ~n3544 ) ;
  assign n3546 = ( x69 & n3342 ) | ( x69 & ~n3516 ) | ( n3342 & ~n3516 ) ;
  assign n3547 = x69 & n3342 ;
  assign n3548 = ( ~n3347 & n3546 ) | ( ~n3347 & n3547 ) | ( n3546 & n3547 ) ;
  assign n3549 = ( n3347 & n3546 ) | ( n3347 & n3547 ) | ( n3546 & n3547 ) ;
  assign n3550 = ( n3347 & n3548 ) | ( n3347 & ~n3549 ) | ( n3548 & ~n3549 ) ;
  assign n3551 = ( x70 & n3545 ) | ( x70 & ~n3550 ) | ( n3545 & ~n3550 ) ;
  assign n3552 = ( x70 & n3348 ) | ( x70 & ~n3516 ) | ( n3348 & ~n3516 ) ;
  assign n3553 = x70 & n3348 ;
  assign n3554 = ( n3353 & n3552 ) | ( n3353 & n3553 ) | ( n3552 & n3553 ) ;
  assign n3555 = ( ~n3353 & n3552 ) | ( ~n3353 & n3553 ) | ( n3552 & n3553 ) ;
  assign n3556 = ( n3353 & ~n3554 ) | ( n3353 & n3555 ) | ( ~n3554 & n3555 ) ;
  assign n3557 = ( x71 & n3551 ) | ( x71 & ~n3556 ) | ( n3551 & ~n3556 ) ;
  assign n3558 = ( x71 & n3354 ) | ( x71 & ~n3516 ) | ( n3354 & ~n3516 ) ;
  assign n3559 = x71 & n3354 ;
  assign n3560 = ( ~n3359 & n3558 ) | ( ~n3359 & n3559 ) | ( n3558 & n3559 ) ;
  assign n3561 = ( n3359 & n3558 ) | ( n3359 & n3559 ) | ( n3558 & n3559 ) ;
  assign n3562 = ( n3359 & n3560 ) | ( n3359 & ~n3561 ) | ( n3560 & ~n3561 ) ;
  assign n3563 = ( x72 & n3557 ) | ( x72 & ~n3562 ) | ( n3557 & ~n3562 ) ;
  assign n3564 = ( x72 & n3360 ) | ( x72 & ~n3516 ) | ( n3360 & ~n3516 ) ;
  assign n3565 = x72 & n3360 ;
  assign n3566 = ( n3365 & n3564 ) | ( n3365 & n3565 ) | ( n3564 & n3565 ) ;
  assign n3567 = ( ~n3365 & n3564 ) | ( ~n3365 & n3565 ) | ( n3564 & n3565 ) ;
  assign n3568 = ( n3365 & ~n3566 ) | ( n3365 & n3567 ) | ( ~n3566 & n3567 ) ;
  assign n3569 = ( x73 & n3563 ) | ( x73 & ~n3568 ) | ( n3563 & ~n3568 ) ;
  assign n3570 = ( x73 & n3366 ) | ( x73 & ~n3516 ) | ( n3366 & ~n3516 ) ;
  assign n3571 = x73 & n3366 ;
  assign n3572 = ( ~n3371 & n3570 ) | ( ~n3371 & n3571 ) | ( n3570 & n3571 ) ;
  assign n3573 = ( n3371 & n3570 ) | ( n3371 & n3571 ) | ( n3570 & n3571 ) ;
  assign n3574 = ( n3371 & n3572 ) | ( n3371 & ~n3573 ) | ( n3572 & ~n3573 ) ;
  assign n3575 = ( x74 & n3569 ) | ( x74 & ~n3574 ) | ( n3569 & ~n3574 ) ;
  assign n3576 = ( x74 & n3372 ) | ( x74 & ~n3516 ) | ( n3372 & ~n3516 ) ;
  assign n3577 = x74 & n3372 ;
  assign n3578 = ( n3377 & n3576 ) | ( n3377 & n3577 ) | ( n3576 & n3577 ) ;
  assign n3579 = ( ~n3377 & n3576 ) | ( ~n3377 & n3577 ) | ( n3576 & n3577 ) ;
  assign n3580 = ( n3377 & ~n3578 ) | ( n3377 & n3579 ) | ( ~n3578 & n3579 ) ;
  assign n3581 = ( x75 & n3575 ) | ( x75 & ~n3580 ) | ( n3575 & ~n3580 ) ;
  assign n3582 = ( x75 & n3378 ) | ( x75 & ~n3516 ) | ( n3378 & ~n3516 ) ;
  assign n3583 = x75 & n3378 ;
  assign n3584 = ( ~n3383 & n3582 ) | ( ~n3383 & n3583 ) | ( n3582 & n3583 ) ;
  assign n3585 = ( n3383 & n3582 ) | ( n3383 & n3583 ) | ( n3582 & n3583 ) ;
  assign n3586 = ( n3383 & n3584 ) | ( n3383 & ~n3585 ) | ( n3584 & ~n3585 ) ;
  assign n3587 = ( x76 & n3581 ) | ( x76 & ~n3586 ) | ( n3581 & ~n3586 ) ;
  assign n3588 = ( x76 & n3384 ) | ( x76 & ~n3516 ) | ( n3384 & ~n3516 ) ;
  assign n3589 = x76 & n3384 ;
  assign n3590 = ( n3389 & n3588 ) | ( n3389 & n3589 ) | ( n3588 & n3589 ) ;
  assign n3591 = ( ~n3389 & n3588 ) | ( ~n3389 & n3589 ) | ( n3588 & n3589 ) ;
  assign n3592 = ( n3389 & ~n3590 ) | ( n3389 & n3591 ) | ( ~n3590 & n3591 ) ;
  assign n3593 = ( x77 & n3587 ) | ( x77 & ~n3592 ) | ( n3587 & ~n3592 ) ;
  assign n3594 = ( x77 & n3390 ) | ( x77 & ~n3516 ) | ( n3390 & ~n3516 ) ;
  assign n3595 = x77 & n3390 ;
  assign n3596 = ( ~n3395 & n3594 ) | ( ~n3395 & n3595 ) | ( n3594 & n3595 ) ;
  assign n3597 = ( n3395 & n3594 ) | ( n3395 & n3595 ) | ( n3594 & n3595 ) ;
  assign n3598 = ( n3395 & n3596 ) | ( n3395 & ~n3597 ) | ( n3596 & ~n3597 ) ;
  assign n3599 = ( x78 & n3593 ) | ( x78 & ~n3598 ) | ( n3593 & ~n3598 ) ;
  assign n3600 = ( x78 & n3396 ) | ( x78 & ~n3516 ) | ( n3396 & ~n3516 ) ;
  assign n3601 = x78 & n3396 ;
  assign n3602 = ( n3401 & n3600 ) | ( n3401 & n3601 ) | ( n3600 & n3601 ) ;
  assign n3603 = ( ~n3401 & n3600 ) | ( ~n3401 & n3601 ) | ( n3600 & n3601 ) ;
  assign n3604 = ( n3401 & ~n3602 ) | ( n3401 & n3603 ) | ( ~n3602 & n3603 ) ;
  assign n3605 = ( x79 & n3599 ) | ( x79 & ~n3604 ) | ( n3599 & ~n3604 ) ;
  assign n3606 = ( x79 & n3402 ) | ( x79 & ~n3516 ) | ( n3402 & ~n3516 ) ;
  assign n3607 = x79 & n3402 ;
  assign n3608 = ( ~n3407 & n3606 ) | ( ~n3407 & n3607 ) | ( n3606 & n3607 ) ;
  assign n3609 = ( n3407 & n3606 ) | ( n3407 & n3607 ) | ( n3606 & n3607 ) ;
  assign n3610 = ( n3407 & n3608 ) | ( n3407 & ~n3609 ) | ( n3608 & ~n3609 ) ;
  assign n3611 = ( x80 & n3605 ) | ( x80 & ~n3610 ) | ( n3605 & ~n3610 ) ;
  assign n3612 = ( x80 & n3408 ) | ( x80 & ~n3516 ) | ( n3408 & ~n3516 ) ;
  assign n3613 = x80 & n3408 ;
  assign n3614 = ( n3413 & n3612 ) | ( n3413 & n3613 ) | ( n3612 & n3613 ) ;
  assign n3615 = ( ~n3413 & n3612 ) | ( ~n3413 & n3613 ) | ( n3612 & n3613 ) ;
  assign n3616 = ( n3413 & ~n3614 ) | ( n3413 & n3615 ) | ( ~n3614 & n3615 ) ;
  assign n3617 = ( x81 & n3611 ) | ( x81 & ~n3616 ) | ( n3611 & ~n3616 ) ;
  assign n3618 = ( x81 & n3414 ) | ( x81 & ~n3516 ) | ( n3414 & ~n3516 ) ;
  assign n3619 = x81 & n3414 ;
  assign n3620 = ( ~n3419 & n3618 ) | ( ~n3419 & n3619 ) | ( n3618 & n3619 ) ;
  assign n3621 = ( n3419 & n3618 ) | ( n3419 & n3619 ) | ( n3618 & n3619 ) ;
  assign n3622 = ( n3419 & n3620 ) | ( n3419 & ~n3621 ) | ( n3620 & ~n3621 ) ;
  assign n3623 = ( x82 & n3617 ) | ( x82 & ~n3622 ) | ( n3617 & ~n3622 ) ;
  assign n3624 = ( x82 & n3420 ) | ( x82 & ~n3516 ) | ( n3420 & ~n3516 ) ;
  assign n3625 = x82 & n3420 ;
  assign n3626 = ( n3425 & n3624 ) | ( n3425 & n3625 ) | ( n3624 & n3625 ) ;
  assign n3627 = ( ~n3425 & n3624 ) | ( ~n3425 & n3625 ) | ( n3624 & n3625 ) ;
  assign n3628 = ( n3425 & ~n3626 ) | ( n3425 & n3627 ) | ( ~n3626 & n3627 ) ;
  assign n3629 = ( x83 & n3623 ) | ( x83 & ~n3628 ) | ( n3623 & ~n3628 ) ;
  assign n3630 = ( x83 & n3426 ) | ( x83 & ~n3516 ) | ( n3426 & ~n3516 ) ;
  assign n3631 = x83 & n3426 ;
  assign n3632 = ( ~n3431 & n3630 ) | ( ~n3431 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3633 = ( n3431 & n3630 ) | ( n3431 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3634 = ( n3431 & n3632 ) | ( n3431 & ~n3633 ) | ( n3632 & ~n3633 ) ;
  assign n3635 = ( x84 & n3629 ) | ( x84 & ~n3634 ) | ( n3629 & ~n3634 ) ;
  assign n3636 = ( x84 & n3432 ) | ( x84 & ~n3516 ) | ( n3432 & ~n3516 ) ;
  assign n3637 = x84 & n3432 ;
  assign n3638 = ( n3437 & n3636 ) | ( n3437 & n3637 ) | ( n3636 & n3637 ) ;
  assign n3639 = ( ~n3437 & n3636 ) | ( ~n3437 & n3637 ) | ( n3636 & n3637 ) ;
  assign n3640 = ( n3437 & ~n3638 ) | ( n3437 & n3639 ) | ( ~n3638 & n3639 ) ;
  assign n3641 = ( x85 & n3635 ) | ( x85 & ~n3640 ) | ( n3635 & ~n3640 ) ;
  assign n3642 = ( x85 & n3438 ) | ( x85 & ~n3516 ) | ( n3438 & ~n3516 ) ;
  assign n3643 = x85 & n3438 ;
  assign n3644 = ( ~n3443 & n3642 ) | ( ~n3443 & n3643 ) | ( n3642 & n3643 ) ;
  assign n3645 = ( n3443 & n3642 ) | ( n3443 & n3643 ) | ( n3642 & n3643 ) ;
  assign n3646 = ( n3443 & n3644 ) | ( n3443 & ~n3645 ) | ( n3644 & ~n3645 ) ;
  assign n3647 = ( x86 & n3641 ) | ( x86 & ~n3646 ) | ( n3641 & ~n3646 ) ;
  assign n3648 = ( x86 & n3444 ) | ( x86 & ~n3516 ) | ( n3444 & ~n3516 ) ;
  assign n3649 = x86 & n3444 ;
  assign n3650 = ( n3449 & n3648 ) | ( n3449 & n3649 ) | ( n3648 & n3649 ) ;
  assign n3651 = ( ~n3449 & n3648 ) | ( ~n3449 & n3649 ) | ( n3648 & n3649 ) ;
  assign n3652 = ( n3449 & ~n3650 ) | ( n3449 & n3651 ) | ( ~n3650 & n3651 ) ;
  assign n3653 = ( x87 & n3647 ) | ( x87 & ~n3652 ) | ( n3647 & ~n3652 ) ;
  assign n3654 = ( x87 & n3450 ) | ( x87 & ~n3516 ) | ( n3450 & ~n3516 ) ;
  assign n3655 = x87 & n3450 ;
  assign n3656 = ( ~n3455 & n3654 ) | ( ~n3455 & n3655 ) | ( n3654 & n3655 ) ;
  assign n3657 = ( n3455 & n3654 ) | ( n3455 & n3655 ) | ( n3654 & n3655 ) ;
  assign n3658 = ( n3455 & n3656 ) | ( n3455 & ~n3657 ) | ( n3656 & ~n3657 ) ;
  assign n3659 = ( x88 & n3653 ) | ( x88 & ~n3658 ) | ( n3653 & ~n3658 ) ;
  assign n3660 = ( x88 & n3456 ) | ( x88 & ~n3516 ) | ( n3456 & ~n3516 ) ;
  assign n3661 = x88 & n3456 ;
  assign n3662 = ( n3461 & n3660 ) | ( n3461 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3663 = ( ~n3461 & n3660 ) | ( ~n3461 & n3661 ) | ( n3660 & n3661 ) ;
  assign n3664 = ( n3461 & ~n3662 ) | ( n3461 & n3663 ) | ( ~n3662 & n3663 ) ;
  assign n3665 = ( x89 & n3659 ) | ( x89 & ~n3664 ) | ( n3659 & ~n3664 ) ;
  assign n3666 = ( x89 & n3462 ) | ( x89 & ~n3516 ) | ( n3462 & ~n3516 ) ;
  assign n3667 = x89 & n3462 ;
  assign n3668 = ( ~n3467 & n3666 ) | ( ~n3467 & n3667 ) | ( n3666 & n3667 ) ;
  assign n3669 = ( n3467 & n3666 ) | ( n3467 & n3667 ) | ( n3666 & n3667 ) ;
  assign n3670 = ( n3467 & n3668 ) | ( n3467 & ~n3669 ) | ( n3668 & ~n3669 ) ;
  assign n3671 = ( x90 & n3665 ) | ( x90 & ~n3670 ) | ( n3665 & ~n3670 ) ;
  assign n3672 = ( x90 & n3468 ) | ( x90 & ~n3516 ) | ( n3468 & ~n3516 ) ;
  assign n3673 = x90 & n3468 ;
  assign n3674 = ( n3473 & n3672 ) | ( n3473 & n3673 ) | ( n3672 & n3673 ) ;
  assign n3675 = ( ~n3473 & n3672 ) | ( ~n3473 & n3673 ) | ( n3672 & n3673 ) ;
  assign n3676 = ( n3473 & ~n3674 ) | ( n3473 & n3675 ) | ( ~n3674 & n3675 ) ;
  assign n3677 = ( x91 & n3671 ) | ( x91 & ~n3676 ) | ( n3671 & ~n3676 ) ;
  assign n3678 = ( x91 & n3474 ) | ( x91 & ~n3516 ) | ( n3474 & ~n3516 ) ;
  assign n3679 = x91 & n3474 ;
  assign n3680 = ( ~n3479 & n3678 ) | ( ~n3479 & n3679 ) | ( n3678 & n3679 ) ;
  assign n3681 = ( n3479 & n3678 ) | ( n3479 & n3679 ) | ( n3678 & n3679 ) ;
  assign n3682 = ( n3479 & n3680 ) | ( n3479 & ~n3681 ) | ( n3680 & ~n3681 ) ;
  assign n3683 = ( x92 & n3677 ) | ( x92 & ~n3682 ) | ( n3677 & ~n3682 ) ;
  assign n3684 = ( x92 & n3480 ) | ( x92 & ~n3516 ) | ( n3480 & ~n3516 ) ;
  assign n3685 = x92 & n3480 ;
  assign n3686 = ( n3485 & n3684 ) | ( n3485 & n3685 ) | ( n3684 & n3685 ) ;
  assign n3687 = ( ~n3485 & n3684 ) | ( ~n3485 & n3685 ) | ( n3684 & n3685 ) ;
  assign n3688 = ( n3485 & ~n3686 ) | ( n3485 & n3687 ) | ( ~n3686 & n3687 ) ;
  assign n3689 = ( x93 & n3683 ) | ( x93 & ~n3688 ) | ( n3683 & ~n3688 ) ;
  assign n3690 = ( x93 & n3486 ) | ( x93 & ~n3516 ) | ( n3486 & ~n3516 ) ;
  assign n3691 = x93 & n3486 ;
  assign n3692 = ( ~n3491 & n3690 ) | ( ~n3491 & n3691 ) | ( n3690 & n3691 ) ;
  assign n3693 = ( n3491 & n3690 ) | ( n3491 & n3691 ) | ( n3690 & n3691 ) ;
  assign n3694 = ( n3491 & n3692 ) | ( n3491 & ~n3693 ) | ( n3692 & ~n3693 ) ;
  assign n3695 = ( x94 & n3689 ) | ( x94 & ~n3694 ) | ( n3689 & ~n3694 ) ;
  assign n3696 = ( x94 & n3492 ) | ( x94 & ~n3516 ) | ( n3492 & ~n3516 ) ;
  assign n3697 = x94 & n3492 ;
  assign n3698 = ( n3497 & n3696 ) | ( n3497 & n3697 ) | ( n3696 & n3697 ) ;
  assign n3699 = ( ~n3497 & n3696 ) | ( ~n3497 & n3697 ) | ( n3696 & n3697 ) ;
  assign n3700 = ( n3497 & ~n3698 ) | ( n3497 & n3699 ) | ( ~n3698 & n3699 ) ;
  assign n3701 = ( x95 & n3695 ) | ( x95 & ~n3700 ) | ( n3695 & ~n3700 ) ;
  assign n3702 = ( x95 & n3498 ) | ( x95 & ~n3516 ) | ( n3498 & ~n3516 ) ;
  assign n3703 = x95 & n3498 ;
  assign n3704 = ( ~n3503 & n3702 ) | ( ~n3503 & n3703 ) | ( n3702 & n3703 ) ;
  assign n3705 = ( n3503 & n3702 ) | ( n3503 & n3703 ) | ( n3702 & n3703 ) ;
  assign n3706 = ( n3503 & n3704 ) | ( n3503 & ~n3705 ) | ( n3704 & ~n3705 ) ;
  assign n3707 = ( x96 & n3701 ) | ( x96 & ~n3706 ) | ( n3701 & ~n3706 ) ;
  assign n3708 = ( x96 & n3504 ) | ( x96 & ~n3516 ) | ( n3504 & ~n3516 ) ;
  assign n3709 = x96 & n3504 ;
  assign n3710 = ( ~n3509 & n3708 ) | ( ~n3509 & n3709 ) | ( n3708 & n3709 ) ;
  assign n3711 = ( n3509 & n3708 ) | ( n3509 & n3709 ) | ( n3708 & n3709 ) ;
  assign n3712 = ( n3509 & n3710 ) | ( n3509 & ~n3711 ) | ( n3710 & ~n3711 ) ;
  assign n3713 = ( x97 & n3707 ) | ( x97 & ~n3712 ) | ( n3707 & ~n3712 ) ;
  assign n3714 = x98 | n3713 ;
  assign n3715 = ( x98 & n159 ) | ( x98 & n3713 ) | ( n159 & n3713 ) ;
  assign n3716 = ( n3514 & ~n3714 ) | ( n3514 & n3715 ) | ( ~n3714 & n3715 ) ;
  assign n3717 = ( x98 & ~n3514 ) | ( x98 & n3713 ) | ( ~n3514 & n3713 ) ;
  assign n3718 = n159 | n3717 ;
  assign n3719 = ( x29 & ~x64 ) | ( x29 & n3718 ) | ( ~x64 & n3718 ) ;
  assign n3720 = ~x29 & n3718 ;
  assign n3721 = ( n3520 & n3719 ) | ( n3520 & ~n3720 ) | ( n3719 & ~n3720 ) ;
  assign n3722 = ~x28 & x64 ;
  assign n3723 = ( x65 & ~n3721 ) | ( x65 & n3722 ) | ( ~n3721 & n3722 ) ;
  assign n3724 = ( x65 & n3520 ) | ( x65 & ~n3718 ) | ( n3520 & ~n3718 ) ;
  assign n3725 = x65 & n3520 ;
  assign n3726 = ( n3519 & n3724 ) | ( n3519 & n3725 ) | ( n3724 & n3725 ) ;
  assign n3727 = ( ~n3519 & n3724 ) | ( ~n3519 & n3725 ) | ( n3724 & n3725 ) ;
  assign n3728 = ( n3519 & ~n3726 ) | ( n3519 & n3727 ) | ( ~n3726 & n3727 ) ;
  assign n3729 = ( x66 & n3723 ) | ( x66 & ~n3728 ) | ( n3723 & ~n3728 ) ;
  assign n3730 = ( x66 & n3521 ) | ( x66 & ~n3718 ) | ( n3521 & ~n3718 ) ;
  assign n3731 = x66 & n3521 ;
  assign n3732 = ( n3526 & n3730 ) | ( n3526 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3733 = ( ~n3526 & n3730 ) | ( ~n3526 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3734 = ( n3526 & ~n3732 ) | ( n3526 & n3733 ) | ( ~n3732 & n3733 ) ;
  assign n3735 = ( x67 & n3729 ) | ( x67 & ~n3734 ) | ( n3729 & ~n3734 ) ;
  assign n3736 = ( x67 & n3527 ) | ( x67 & ~n3718 ) | ( n3527 & ~n3718 ) ;
  assign n3737 = x67 & n3527 ;
  assign n3738 = ( ~n3532 & n3736 ) | ( ~n3532 & n3737 ) | ( n3736 & n3737 ) ;
  assign n3739 = ( n3532 & n3736 ) | ( n3532 & n3737 ) | ( n3736 & n3737 ) ;
  assign n3740 = ( n3532 & n3738 ) | ( n3532 & ~n3739 ) | ( n3738 & ~n3739 ) ;
  assign n3741 = ( x68 & n3735 ) | ( x68 & ~n3740 ) | ( n3735 & ~n3740 ) ;
  assign n3742 = ( x68 & n3533 ) | ( x68 & ~n3718 ) | ( n3533 & ~n3718 ) ;
  assign n3743 = x68 & n3533 ;
  assign n3744 = ( n3538 & n3742 ) | ( n3538 & n3743 ) | ( n3742 & n3743 ) ;
  assign n3745 = ( ~n3538 & n3742 ) | ( ~n3538 & n3743 ) | ( n3742 & n3743 ) ;
  assign n3746 = ( n3538 & ~n3744 ) | ( n3538 & n3745 ) | ( ~n3744 & n3745 ) ;
  assign n3747 = ( x69 & n3741 ) | ( x69 & ~n3746 ) | ( n3741 & ~n3746 ) ;
  assign n3748 = ( x69 & n3539 ) | ( x69 & ~n3718 ) | ( n3539 & ~n3718 ) ;
  assign n3749 = x69 & n3539 ;
  assign n3750 = ( ~n3544 & n3748 ) | ( ~n3544 & n3749 ) | ( n3748 & n3749 ) ;
  assign n3751 = ( n3544 & n3748 ) | ( n3544 & n3749 ) | ( n3748 & n3749 ) ;
  assign n3752 = ( n3544 & n3750 ) | ( n3544 & ~n3751 ) | ( n3750 & ~n3751 ) ;
  assign n3753 = ( x70 & n3747 ) | ( x70 & ~n3752 ) | ( n3747 & ~n3752 ) ;
  assign n3754 = ( x70 & n3545 ) | ( x70 & ~n3718 ) | ( n3545 & ~n3718 ) ;
  assign n3755 = x70 & n3545 ;
  assign n3756 = ( n3550 & n3754 ) | ( n3550 & n3755 ) | ( n3754 & n3755 ) ;
  assign n3757 = ( ~n3550 & n3754 ) | ( ~n3550 & n3755 ) | ( n3754 & n3755 ) ;
  assign n3758 = ( n3550 & ~n3756 ) | ( n3550 & n3757 ) | ( ~n3756 & n3757 ) ;
  assign n3759 = ( x71 & n3753 ) | ( x71 & ~n3758 ) | ( n3753 & ~n3758 ) ;
  assign n3760 = ( x71 & n3551 ) | ( x71 & ~n3718 ) | ( n3551 & ~n3718 ) ;
  assign n3761 = x71 & n3551 ;
  assign n3762 = ( ~n3556 & n3760 ) | ( ~n3556 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3763 = ( n3556 & n3760 ) | ( n3556 & n3761 ) | ( n3760 & n3761 ) ;
  assign n3764 = ( n3556 & n3762 ) | ( n3556 & ~n3763 ) | ( n3762 & ~n3763 ) ;
  assign n3765 = ( x72 & n3759 ) | ( x72 & ~n3764 ) | ( n3759 & ~n3764 ) ;
  assign n3766 = ( x72 & n3557 ) | ( x72 & ~n3718 ) | ( n3557 & ~n3718 ) ;
  assign n3767 = x72 & n3557 ;
  assign n3768 = ( n3562 & n3766 ) | ( n3562 & n3767 ) | ( n3766 & n3767 ) ;
  assign n3769 = ( ~n3562 & n3766 ) | ( ~n3562 & n3767 ) | ( n3766 & n3767 ) ;
  assign n3770 = ( n3562 & ~n3768 ) | ( n3562 & n3769 ) | ( ~n3768 & n3769 ) ;
  assign n3771 = ( x73 & n3765 ) | ( x73 & ~n3770 ) | ( n3765 & ~n3770 ) ;
  assign n3772 = ( x73 & n3563 ) | ( x73 & ~n3718 ) | ( n3563 & ~n3718 ) ;
  assign n3773 = x73 & n3563 ;
  assign n3774 = ( ~n3568 & n3772 ) | ( ~n3568 & n3773 ) | ( n3772 & n3773 ) ;
  assign n3775 = ( n3568 & n3772 ) | ( n3568 & n3773 ) | ( n3772 & n3773 ) ;
  assign n3776 = ( n3568 & n3774 ) | ( n3568 & ~n3775 ) | ( n3774 & ~n3775 ) ;
  assign n3777 = ( x74 & n3771 ) | ( x74 & ~n3776 ) | ( n3771 & ~n3776 ) ;
  assign n3778 = ( x74 & n3569 ) | ( x74 & ~n3718 ) | ( n3569 & ~n3718 ) ;
  assign n3779 = x74 & n3569 ;
  assign n3780 = ( n3574 & n3778 ) | ( n3574 & n3779 ) | ( n3778 & n3779 ) ;
  assign n3781 = ( ~n3574 & n3778 ) | ( ~n3574 & n3779 ) | ( n3778 & n3779 ) ;
  assign n3782 = ( n3574 & ~n3780 ) | ( n3574 & n3781 ) | ( ~n3780 & n3781 ) ;
  assign n3783 = ( x75 & n3777 ) | ( x75 & ~n3782 ) | ( n3777 & ~n3782 ) ;
  assign n3784 = ( x75 & n3575 ) | ( x75 & ~n3718 ) | ( n3575 & ~n3718 ) ;
  assign n3785 = x75 & n3575 ;
  assign n3786 = ( ~n3580 & n3784 ) | ( ~n3580 & n3785 ) | ( n3784 & n3785 ) ;
  assign n3787 = ( n3580 & n3784 ) | ( n3580 & n3785 ) | ( n3784 & n3785 ) ;
  assign n3788 = ( n3580 & n3786 ) | ( n3580 & ~n3787 ) | ( n3786 & ~n3787 ) ;
  assign n3789 = ( x76 & n3783 ) | ( x76 & ~n3788 ) | ( n3783 & ~n3788 ) ;
  assign n3790 = ( x76 & n3581 ) | ( x76 & ~n3718 ) | ( n3581 & ~n3718 ) ;
  assign n3791 = x76 & n3581 ;
  assign n3792 = ( n3586 & n3790 ) | ( n3586 & n3791 ) | ( n3790 & n3791 ) ;
  assign n3793 = ( ~n3586 & n3790 ) | ( ~n3586 & n3791 ) | ( n3790 & n3791 ) ;
  assign n3794 = ( n3586 & ~n3792 ) | ( n3586 & n3793 ) | ( ~n3792 & n3793 ) ;
  assign n3795 = ( x77 & n3789 ) | ( x77 & ~n3794 ) | ( n3789 & ~n3794 ) ;
  assign n3796 = ( x77 & n3587 ) | ( x77 & ~n3718 ) | ( n3587 & ~n3718 ) ;
  assign n3797 = x77 & n3587 ;
  assign n3798 = ( ~n3592 & n3796 ) | ( ~n3592 & n3797 ) | ( n3796 & n3797 ) ;
  assign n3799 = ( n3592 & n3796 ) | ( n3592 & n3797 ) | ( n3796 & n3797 ) ;
  assign n3800 = ( n3592 & n3798 ) | ( n3592 & ~n3799 ) | ( n3798 & ~n3799 ) ;
  assign n3801 = ( x78 & n3795 ) | ( x78 & ~n3800 ) | ( n3795 & ~n3800 ) ;
  assign n3802 = ( x78 & n3593 ) | ( x78 & ~n3718 ) | ( n3593 & ~n3718 ) ;
  assign n3803 = x78 & n3593 ;
  assign n3804 = ( n3598 & n3802 ) | ( n3598 & n3803 ) | ( n3802 & n3803 ) ;
  assign n3805 = ( ~n3598 & n3802 ) | ( ~n3598 & n3803 ) | ( n3802 & n3803 ) ;
  assign n3806 = ( n3598 & ~n3804 ) | ( n3598 & n3805 ) | ( ~n3804 & n3805 ) ;
  assign n3807 = ( x79 & n3801 ) | ( x79 & ~n3806 ) | ( n3801 & ~n3806 ) ;
  assign n3808 = ( x79 & n3599 ) | ( x79 & ~n3718 ) | ( n3599 & ~n3718 ) ;
  assign n3809 = x79 & n3599 ;
  assign n3810 = ( ~n3604 & n3808 ) | ( ~n3604 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3811 = ( n3604 & n3808 ) | ( n3604 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3812 = ( n3604 & n3810 ) | ( n3604 & ~n3811 ) | ( n3810 & ~n3811 ) ;
  assign n3813 = ( x80 & n3807 ) | ( x80 & ~n3812 ) | ( n3807 & ~n3812 ) ;
  assign n3814 = ( x80 & n3605 ) | ( x80 & ~n3718 ) | ( n3605 & ~n3718 ) ;
  assign n3815 = x80 & n3605 ;
  assign n3816 = ( n3610 & n3814 ) | ( n3610 & n3815 ) | ( n3814 & n3815 ) ;
  assign n3817 = ( ~n3610 & n3814 ) | ( ~n3610 & n3815 ) | ( n3814 & n3815 ) ;
  assign n3818 = ( n3610 & ~n3816 ) | ( n3610 & n3817 ) | ( ~n3816 & n3817 ) ;
  assign n3819 = ( x81 & n3813 ) | ( x81 & ~n3818 ) | ( n3813 & ~n3818 ) ;
  assign n3820 = ( x81 & n3611 ) | ( x81 & ~n3718 ) | ( n3611 & ~n3718 ) ;
  assign n3821 = x81 & n3611 ;
  assign n3822 = ( ~n3616 & n3820 ) | ( ~n3616 & n3821 ) | ( n3820 & n3821 ) ;
  assign n3823 = ( n3616 & n3820 ) | ( n3616 & n3821 ) | ( n3820 & n3821 ) ;
  assign n3824 = ( n3616 & n3822 ) | ( n3616 & ~n3823 ) | ( n3822 & ~n3823 ) ;
  assign n3825 = ( x82 & n3819 ) | ( x82 & ~n3824 ) | ( n3819 & ~n3824 ) ;
  assign n3826 = ( x82 & n3617 ) | ( x82 & ~n3718 ) | ( n3617 & ~n3718 ) ;
  assign n3827 = x82 & n3617 ;
  assign n3828 = ( n3622 & n3826 ) | ( n3622 & n3827 ) | ( n3826 & n3827 ) ;
  assign n3829 = ( ~n3622 & n3826 ) | ( ~n3622 & n3827 ) | ( n3826 & n3827 ) ;
  assign n3830 = ( n3622 & ~n3828 ) | ( n3622 & n3829 ) | ( ~n3828 & n3829 ) ;
  assign n3831 = ( x83 & n3825 ) | ( x83 & ~n3830 ) | ( n3825 & ~n3830 ) ;
  assign n3832 = ( x83 & n3623 ) | ( x83 & ~n3718 ) | ( n3623 & ~n3718 ) ;
  assign n3833 = x83 & n3623 ;
  assign n3834 = ( ~n3628 & n3832 ) | ( ~n3628 & n3833 ) | ( n3832 & n3833 ) ;
  assign n3835 = ( n3628 & n3832 ) | ( n3628 & n3833 ) | ( n3832 & n3833 ) ;
  assign n3836 = ( n3628 & n3834 ) | ( n3628 & ~n3835 ) | ( n3834 & ~n3835 ) ;
  assign n3837 = ( x84 & n3831 ) | ( x84 & ~n3836 ) | ( n3831 & ~n3836 ) ;
  assign n3838 = ( x84 & n3629 ) | ( x84 & ~n3718 ) | ( n3629 & ~n3718 ) ;
  assign n3839 = x84 & n3629 ;
  assign n3840 = ( n3634 & n3838 ) | ( n3634 & n3839 ) | ( n3838 & n3839 ) ;
  assign n3841 = ( ~n3634 & n3838 ) | ( ~n3634 & n3839 ) | ( n3838 & n3839 ) ;
  assign n3842 = ( n3634 & ~n3840 ) | ( n3634 & n3841 ) | ( ~n3840 & n3841 ) ;
  assign n3843 = ( x85 & n3837 ) | ( x85 & ~n3842 ) | ( n3837 & ~n3842 ) ;
  assign n3844 = ( x85 & n3635 ) | ( x85 & ~n3718 ) | ( n3635 & ~n3718 ) ;
  assign n3845 = x85 & n3635 ;
  assign n3846 = ( ~n3640 & n3844 ) | ( ~n3640 & n3845 ) | ( n3844 & n3845 ) ;
  assign n3847 = ( n3640 & n3844 ) | ( n3640 & n3845 ) | ( n3844 & n3845 ) ;
  assign n3848 = ( n3640 & n3846 ) | ( n3640 & ~n3847 ) | ( n3846 & ~n3847 ) ;
  assign n3849 = ( x86 & n3843 ) | ( x86 & ~n3848 ) | ( n3843 & ~n3848 ) ;
  assign n3850 = ( x86 & n3641 ) | ( x86 & ~n3718 ) | ( n3641 & ~n3718 ) ;
  assign n3851 = x86 & n3641 ;
  assign n3852 = ( n3646 & n3850 ) | ( n3646 & n3851 ) | ( n3850 & n3851 ) ;
  assign n3853 = ( ~n3646 & n3850 ) | ( ~n3646 & n3851 ) | ( n3850 & n3851 ) ;
  assign n3854 = ( n3646 & ~n3852 ) | ( n3646 & n3853 ) | ( ~n3852 & n3853 ) ;
  assign n3855 = ( x87 & n3849 ) | ( x87 & ~n3854 ) | ( n3849 & ~n3854 ) ;
  assign n3856 = ( x87 & n3647 ) | ( x87 & ~n3718 ) | ( n3647 & ~n3718 ) ;
  assign n3857 = x87 & n3647 ;
  assign n3858 = ( ~n3652 & n3856 ) | ( ~n3652 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3859 = ( n3652 & n3856 ) | ( n3652 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3860 = ( n3652 & n3858 ) | ( n3652 & ~n3859 ) | ( n3858 & ~n3859 ) ;
  assign n3861 = ( x88 & n3855 ) | ( x88 & ~n3860 ) | ( n3855 & ~n3860 ) ;
  assign n3862 = ( x88 & n3653 ) | ( x88 & ~n3718 ) | ( n3653 & ~n3718 ) ;
  assign n3863 = x88 & n3653 ;
  assign n3864 = ( n3658 & n3862 ) | ( n3658 & n3863 ) | ( n3862 & n3863 ) ;
  assign n3865 = ( ~n3658 & n3862 ) | ( ~n3658 & n3863 ) | ( n3862 & n3863 ) ;
  assign n3866 = ( n3658 & ~n3864 ) | ( n3658 & n3865 ) | ( ~n3864 & n3865 ) ;
  assign n3867 = ( x89 & n3861 ) | ( x89 & ~n3866 ) | ( n3861 & ~n3866 ) ;
  assign n3868 = ( x89 & n3659 ) | ( x89 & ~n3718 ) | ( n3659 & ~n3718 ) ;
  assign n3869 = x89 & n3659 ;
  assign n3870 = ( ~n3664 & n3868 ) | ( ~n3664 & n3869 ) | ( n3868 & n3869 ) ;
  assign n3871 = ( n3664 & n3868 ) | ( n3664 & n3869 ) | ( n3868 & n3869 ) ;
  assign n3872 = ( n3664 & n3870 ) | ( n3664 & ~n3871 ) | ( n3870 & ~n3871 ) ;
  assign n3873 = ( x90 & n3867 ) | ( x90 & ~n3872 ) | ( n3867 & ~n3872 ) ;
  assign n3874 = ( x90 & n3665 ) | ( x90 & ~n3718 ) | ( n3665 & ~n3718 ) ;
  assign n3875 = x90 & n3665 ;
  assign n3876 = ( n3670 & n3874 ) | ( n3670 & n3875 ) | ( n3874 & n3875 ) ;
  assign n3877 = ( ~n3670 & n3874 ) | ( ~n3670 & n3875 ) | ( n3874 & n3875 ) ;
  assign n3878 = ( n3670 & ~n3876 ) | ( n3670 & n3877 ) | ( ~n3876 & n3877 ) ;
  assign n3879 = ( x91 & n3873 ) | ( x91 & ~n3878 ) | ( n3873 & ~n3878 ) ;
  assign n3880 = ( x91 & n3671 ) | ( x91 & ~n3718 ) | ( n3671 & ~n3718 ) ;
  assign n3881 = x91 & n3671 ;
  assign n3882 = ( ~n3676 & n3880 ) | ( ~n3676 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3883 = ( n3676 & n3880 ) | ( n3676 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3884 = ( n3676 & n3882 ) | ( n3676 & ~n3883 ) | ( n3882 & ~n3883 ) ;
  assign n3885 = ( x92 & n3879 ) | ( x92 & ~n3884 ) | ( n3879 & ~n3884 ) ;
  assign n3886 = ( x92 & n3677 ) | ( x92 & ~n3718 ) | ( n3677 & ~n3718 ) ;
  assign n3887 = x92 & n3677 ;
  assign n3888 = ( n3682 & n3886 ) | ( n3682 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3889 = ( ~n3682 & n3886 ) | ( ~n3682 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3890 = ( n3682 & ~n3888 ) | ( n3682 & n3889 ) | ( ~n3888 & n3889 ) ;
  assign n3891 = ( x93 & n3885 ) | ( x93 & ~n3890 ) | ( n3885 & ~n3890 ) ;
  assign n3892 = ( x93 & n3683 ) | ( x93 & ~n3718 ) | ( n3683 & ~n3718 ) ;
  assign n3893 = x93 & n3683 ;
  assign n3894 = ( ~n3688 & n3892 ) | ( ~n3688 & n3893 ) | ( n3892 & n3893 ) ;
  assign n3895 = ( n3688 & n3892 ) | ( n3688 & n3893 ) | ( n3892 & n3893 ) ;
  assign n3896 = ( n3688 & n3894 ) | ( n3688 & ~n3895 ) | ( n3894 & ~n3895 ) ;
  assign n3897 = ( x94 & n3891 ) | ( x94 & ~n3896 ) | ( n3891 & ~n3896 ) ;
  assign n3898 = ( x94 & n3689 ) | ( x94 & ~n3718 ) | ( n3689 & ~n3718 ) ;
  assign n3899 = x94 & n3689 ;
  assign n3900 = ( n3694 & n3898 ) | ( n3694 & n3899 ) | ( n3898 & n3899 ) ;
  assign n3901 = ( ~n3694 & n3898 ) | ( ~n3694 & n3899 ) | ( n3898 & n3899 ) ;
  assign n3902 = ( n3694 & ~n3900 ) | ( n3694 & n3901 ) | ( ~n3900 & n3901 ) ;
  assign n3903 = ( x95 & n3897 ) | ( x95 & ~n3902 ) | ( n3897 & ~n3902 ) ;
  assign n3904 = ( x95 & n3695 ) | ( x95 & ~n3718 ) | ( n3695 & ~n3718 ) ;
  assign n3905 = x95 & n3695 ;
  assign n3906 = ( ~n3700 & n3904 ) | ( ~n3700 & n3905 ) | ( n3904 & n3905 ) ;
  assign n3907 = ( n3700 & n3904 ) | ( n3700 & n3905 ) | ( n3904 & n3905 ) ;
  assign n3908 = ( n3700 & n3906 ) | ( n3700 & ~n3907 ) | ( n3906 & ~n3907 ) ;
  assign n3909 = ( x96 & n3903 ) | ( x96 & ~n3908 ) | ( n3903 & ~n3908 ) ;
  assign n3910 = ( x96 & n3701 ) | ( x96 & ~n3718 ) | ( n3701 & ~n3718 ) ;
  assign n3911 = x96 & n3701 ;
  assign n3912 = ( n3706 & n3910 ) | ( n3706 & n3911 ) | ( n3910 & n3911 ) ;
  assign n3913 = ( ~n3706 & n3910 ) | ( ~n3706 & n3911 ) | ( n3910 & n3911 ) ;
  assign n3914 = ( n3706 & ~n3912 ) | ( n3706 & n3913 ) | ( ~n3912 & n3913 ) ;
  assign n3915 = ( x97 & n3909 ) | ( x97 & ~n3914 ) | ( n3909 & ~n3914 ) ;
  assign n3916 = ( x97 & n3707 ) | ( x97 & ~n3718 ) | ( n3707 & ~n3718 ) ;
  assign n3917 = x97 & n3707 ;
  assign n3918 = ( n3712 & n3916 ) | ( n3712 & n3917 ) | ( n3916 & n3917 ) ;
  assign n3919 = ( ~n3712 & n3916 ) | ( ~n3712 & n3917 ) | ( n3916 & n3917 ) ;
  assign n3920 = ( n3712 & ~n3918 ) | ( n3712 & n3919 ) | ( ~n3918 & n3919 ) ;
  assign n3921 = ( x98 & n3915 ) | ( x98 & ~n3920 ) | ( n3915 & ~n3920 ) ;
  assign n3922 = x99 | n3921 ;
  assign n3923 = ( x99 & n158 ) | ( x99 & n3921 ) | ( n158 & n3921 ) ;
  assign n3924 = ( n3716 & ~n3922 ) | ( n3716 & n3923 ) | ( ~n3922 & n3923 ) ;
  assign n3925 = ( x99 & ~n3716 ) | ( x99 & n3921 ) | ( ~n3716 & n3921 ) ;
  assign n3926 = n158 | n3925 ;
  assign n3927 = ( x28 & ~x64 ) | ( x28 & n3926 ) | ( ~x64 & n3926 ) ;
  assign n3928 = ~x28 & n3926 ;
  assign n3929 = ( n3722 & n3927 ) | ( n3722 & ~n3928 ) | ( n3927 & ~n3928 ) ;
  assign n3930 = ~x27 & x64 ;
  assign n3931 = ( x65 & ~n3929 ) | ( x65 & n3930 ) | ( ~n3929 & n3930 ) ;
  assign n3932 = ( x65 & n3722 ) | ( x65 & ~n3926 ) | ( n3722 & ~n3926 ) ;
  assign n3933 = x65 & n3722 ;
  assign n3934 = ( n3721 & n3932 ) | ( n3721 & n3933 ) | ( n3932 & n3933 ) ;
  assign n3935 = ( ~n3721 & n3932 ) | ( ~n3721 & n3933 ) | ( n3932 & n3933 ) ;
  assign n3936 = ( n3721 & ~n3934 ) | ( n3721 & n3935 ) | ( ~n3934 & n3935 ) ;
  assign n3937 = ( x66 & n3931 ) | ( x66 & ~n3936 ) | ( n3931 & ~n3936 ) ;
  assign n3938 = ( x66 & n3723 ) | ( x66 & ~n3926 ) | ( n3723 & ~n3926 ) ;
  assign n3939 = x66 & n3723 ;
  assign n3940 = ( n3728 & n3938 ) | ( n3728 & n3939 ) | ( n3938 & n3939 ) ;
  assign n3941 = ( ~n3728 & n3938 ) | ( ~n3728 & n3939 ) | ( n3938 & n3939 ) ;
  assign n3942 = ( n3728 & ~n3940 ) | ( n3728 & n3941 ) | ( ~n3940 & n3941 ) ;
  assign n3943 = ( x67 & n3937 ) | ( x67 & ~n3942 ) | ( n3937 & ~n3942 ) ;
  assign n3944 = ( x67 & n3729 ) | ( x67 & ~n3926 ) | ( n3729 & ~n3926 ) ;
  assign n3945 = x67 & n3729 ;
  assign n3946 = ( ~n3734 & n3944 ) | ( ~n3734 & n3945 ) | ( n3944 & n3945 ) ;
  assign n3947 = ( n3734 & n3944 ) | ( n3734 & n3945 ) | ( n3944 & n3945 ) ;
  assign n3948 = ( n3734 & n3946 ) | ( n3734 & ~n3947 ) | ( n3946 & ~n3947 ) ;
  assign n3949 = ( x68 & n3943 ) | ( x68 & ~n3948 ) | ( n3943 & ~n3948 ) ;
  assign n3950 = ( x68 & n3735 ) | ( x68 & ~n3926 ) | ( n3735 & ~n3926 ) ;
  assign n3951 = x68 & n3735 ;
  assign n3952 = ( n3740 & n3950 ) | ( n3740 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3953 = ( ~n3740 & n3950 ) | ( ~n3740 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3954 = ( n3740 & ~n3952 ) | ( n3740 & n3953 ) | ( ~n3952 & n3953 ) ;
  assign n3955 = ( x69 & n3949 ) | ( x69 & ~n3954 ) | ( n3949 & ~n3954 ) ;
  assign n3956 = ( x69 & n3741 ) | ( x69 & ~n3926 ) | ( n3741 & ~n3926 ) ;
  assign n3957 = x69 & n3741 ;
  assign n3958 = ( ~n3746 & n3956 ) | ( ~n3746 & n3957 ) | ( n3956 & n3957 ) ;
  assign n3959 = ( n3746 & n3956 ) | ( n3746 & n3957 ) | ( n3956 & n3957 ) ;
  assign n3960 = ( n3746 & n3958 ) | ( n3746 & ~n3959 ) | ( n3958 & ~n3959 ) ;
  assign n3961 = ( x70 & n3955 ) | ( x70 & ~n3960 ) | ( n3955 & ~n3960 ) ;
  assign n3962 = ( x70 & n3747 ) | ( x70 & ~n3926 ) | ( n3747 & ~n3926 ) ;
  assign n3963 = x70 & n3747 ;
  assign n3964 = ( n3752 & n3962 ) | ( n3752 & n3963 ) | ( n3962 & n3963 ) ;
  assign n3965 = ( ~n3752 & n3962 ) | ( ~n3752 & n3963 ) | ( n3962 & n3963 ) ;
  assign n3966 = ( n3752 & ~n3964 ) | ( n3752 & n3965 ) | ( ~n3964 & n3965 ) ;
  assign n3967 = ( x71 & n3961 ) | ( x71 & ~n3966 ) | ( n3961 & ~n3966 ) ;
  assign n3968 = ( x71 & n3753 ) | ( x71 & ~n3926 ) | ( n3753 & ~n3926 ) ;
  assign n3969 = x71 & n3753 ;
  assign n3970 = ( ~n3758 & n3968 ) | ( ~n3758 & n3969 ) | ( n3968 & n3969 ) ;
  assign n3971 = ( n3758 & n3968 ) | ( n3758 & n3969 ) | ( n3968 & n3969 ) ;
  assign n3972 = ( n3758 & n3970 ) | ( n3758 & ~n3971 ) | ( n3970 & ~n3971 ) ;
  assign n3973 = ( x72 & n3967 ) | ( x72 & ~n3972 ) | ( n3967 & ~n3972 ) ;
  assign n3974 = ( x72 & n3759 ) | ( x72 & ~n3926 ) | ( n3759 & ~n3926 ) ;
  assign n3975 = x72 & n3759 ;
  assign n3976 = ( n3764 & n3974 ) | ( n3764 & n3975 ) | ( n3974 & n3975 ) ;
  assign n3977 = ( ~n3764 & n3974 ) | ( ~n3764 & n3975 ) | ( n3974 & n3975 ) ;
  assign n3978 = ( n3764 & ~n3976 ) | ( n3764 & n3977 ) | ( ~n3976 & n3977 ) ;
  assign n3979 = ( x73 & n3973 ) | ( x73 & ~n3978 ) | ( n3973 & ~n3978 ) ;
  assign n3980 = ( x73 & n3765 ) | ( x73 & ~n3926 ) | ( n3765 & ~n3926 ) ;
  assign n3981 = x73 & n3765 ;
  assign n3982 = ( ~n3770 & n3980 ) | ( ~n3770 & n3981 ) | ( n3980 & n3981 ) ;
  assign n3983 = ( n3770 & n3980 ) | ( n3770 & n3981 ) | ( n3980 & n3981 ) ;
  assign n3984 = ( n3770 & n3982 ) | ( n3770 & ~n3983 ) | ( n3982 & ~n3983 ) ;
  assign n3985 = ( x74 & n3979 ) | ( x74 & ~n3984 ) | ( n3979 & ~n3984 ) ;
  assign n3986 = ( x74 & n3771 ) | ( x74 & ~n3926 ) | ( n3771 & ~n3926 ) ;
  assign n3987 = x74 & n3771 ;
  assign n3988 = ( n3776 & n3986 ) | ( n3776 & n3987 ) | ( n3986 & n3987 ) ;
  assign n3989 = ( ~n3776 & n3986 ) | ( ~n3776 & n3987 ) | ( n3986 & n3987 ) ;
  assign n3990 = ( n3776 & ~n3988 ) | ( n3776 & n3989 ) | ( ~n3988 & n3989 ) ;
  assign n3991 = ( x75 & n3985 ) | ( x75 & ~n3990 ) | ( n3985 & ~n3990 ) ;
  assign n3992 = ( x75 & n3777 ) | ( x75 & ~n3926 ) | ( n3777 & ~n3926 ) ;
  assign n3993 = x75 & n3777 ;
  assign n3994 = ( ~n3782 & n3992 ) | ( ~n3782 & n3993 ) | ( n3992 & n3993 ) ;
  assign n3995 = ( n3782 & n3992 ) | ( n3782 & n3993 ) | ( n3992 & n3993 ) ;
  assign n3996 = ( n3782 & n3994 ) | ( n3782 & ~n3995 ) | ( n3994 & ~n3995 ) ;
  assign n3997 = ( x76 & n3991 ) | ( x76 & ~n3996 ) | ( n3991 & ~n3996 ) ;
  assign n3998 = ( x76 & n3783 ) | ( x76 & ~n3926 ) | ( n3783 & ~n3926 ) ;
  assign n3999 = x76 & n3783 ;
  assign n4000 = ( n3788 & n3998 ) | ( n3788 & n3999 ) | ( n3998 & n3999 ) ;
  assign n4001 = ( ~n3788 & n3998 ) | ( ~n3788 & n3999 ) | ( n3998 & n3999 ) ;
  assign n4002 = ( n3788 & ~n4000 ) | ( n3788 & n4001 ) | ( ~n4000 & n4001 ) ;
  assign n4003 = ( x77 & n3997 ) | ( x77 & ~n4002 ) | ( n3997 & ~n4002 ) ;
  assign n4004 = ( x77 & n3789 ) | ( x77 & ~n3926 ) | ( n3789 & ~n3926 ) ;
  assign n4005 = x77 & n3789 ;
  assign n4006 = ( ~n3794 & n4004 ) | ( ~n3794 & n4005 ) | ( n4004 & n4005 ) ;
  assign n4007 = ( n3794 & n4004 ) | ( n3794 & n4005 ) | ( n4004 & n4005 ) ;
  assign n4008 = ( n3794 & n4006 ) | ( n3794 & ~n4007 ) | ( n4006 & ~n4007 ) ;
  assign n4009 = ( x78 & n4003 ) | ( x78 & ~n4008 ) | ( n4003 & ~n4008 ) ;
  assign n4010 = ( x78 & n3795 ) | ( x78 & ~n3926 ) | ( n3795 & ~n3926 ) ;
  assign n4011 = x78 & n3795 ;
  assign n4012 = ( n3800 & n4010 ) | ( n3800 & n4011 ) | ( n4010 & n4011 ) ;
  assign n4013 = ( ~n3800 & n4010 ) | ( ~n3800 & n4011 ) | ( n4010 & n4011 ) ;
  assign n4014 = ( n3800 & ~n4012 ) | ( n3800 & n4013 ) | ( ~n4012 & n4013 ) ;
  assign n4015 = ( x79 & n4009 ) | ( x79 & ~n4014 ) | ( n4009 & ~n4014 ) ;
  assign n4016 = ( x79 & n3801 ) | ( x79 & ~n3926 ) | ( n3801 & ~n3926 ) ;
  assign n4017 = x79 & n3801 ;
  assign n4018 = ( ~n3806 & n4016 ) | ( ~n3806 & n4017 ) | ( n4016 & n4017 ) ;
  assign n4019 = ( n3806 & n4016 ) | ( n3806 & n4017 ) | ( n4016 & n4017 ) ;
  assign n4020 = ( n3806 & n4018 ) | ( n3806 & ~n4019 ) | ( n4018 & ~n4019 ) ;
  assign n4021 = ( x80 & n4015 ) | ( x80 & ~n4020 ) | ( n4015 & ~n4020 ) ;
  assign n4022 = ( x80 & n3807 ) | ( x80 & ~n3926 ) | ( n3807 & ~n3926 ) ;
  assign n4023 = x80 & n3807 ;
  assign n4024 = ( n3812 & n4022 ) | ( n3812 & n4023 ) | ( n4022 & n4023 ) ;
  assign n4025 = ( ~n3812 & n4022 ) | ( ~n3812 & n4023 ) | ( n4022 & n4023 ) ;
  assign n4026 = ( n3812 & ~n4024 ) | ( n3812 & n4025 ) | ( ~n4024 & n4025 ) ;
  assign n4027 = ( x81 & n4021 ) | ( x81 & ~n4026 ) | ( n4021 & ~n4026 ) ;
  assign n4028 = ( x81 & n3813 ) | ( x81 & ~n3926 ) | ( n3813 & ~n3926 ) ;
  assign n4029 = x81 & n3813 ;
  assign n4030 = ( ~n3818 & n4028 ) | ( ~n3818 & n4029 ) | ( n4028 & n4029 ) ;
  assign n4031 = ( n3818 & n4028 ) | ( n3818 & n4029 ) | ( n4028 & n4029 ) ;
  assign n4032 = ( n3818 & n4030 ) | ( n3818 & ~n4031 ) | ( n4030 & ~n4031 ) ;
  assign n4033 = ( x82 & n4027 ) | ( x82 & ~n4032 ) | ( n4027 & ~n4032 ) ;
  assign n4034 = ( x82 & n3819 ) | ( x82 & ~n3926 ) | ( n3819 & ~n3926 ) ;
  assign n4035 = x82 & n3819 ;
  assign n4036 = ( n3824 & n4034 ) | ( n3824 & n4035 ) | ( n4034 & n4035 ) ;
  assign n4037 = ( ~n3824 & n4034 ) | ( ~n3824 & n4035 ) | ( n4034 & n4035 ) ;
  assign n4038 = ( n3824 & ~n4036 ) | ( n3824 & n4037 ) | ( ~n4036 & n4037 ) ;
  assign n4039 = ( x83 & n4033 ) | ( x83 & ~n4038 ) | ( n4033 & ~n4038 ) ;
  assign n4040 = ( x83 & n3825 ) | ( x83 & ~n3926 ) | ( n3825 & ~n3926 ) ;
  assign n4041 = x83 & n3825 ;
  assign n4042 = ( ~n3830 & n4040 ) | ( ~n3830 & n4041 ) | ( n4040 & n4041 ) ;
  assign n4043 = ( n3830 & n4040 ) | ( n3830 & n4041 ) | ( n4040 & n4041 ) ;
  assign n4044 = ( n3830 & n4042 ) | ( n3830 & ~n4043 ) | ( n4042 & ~n4043 ) ;
  assign n4045 = ( x84 & n4039 ) | ( x84 & ~n4044 ) | ( n4039 & ~n4044 ) ;
  assign n4046 = ( x84 & n3831 ) | ( x84 & ~n3926 ) | ( n3831 & ~n3926 ) ;
  assign n4047 = x84 & n3831 ;
  assign n4048 = ( n3836 & n4046 ) | ( n3836 & n4047 ) | ( n4046 & n4047 ) ;
  assign n4049 = ( ~n3836 & n4046 ) | ( ~n3836 & n4047 ) | ( n4046 & n4047 ) ;
  assign n4050 = ( n3836 & ~n4048 ) | ( n3836 & n4049 ) | ( ~n4048 & n4049 ) ;
  assign n4051 = ( x85 & n4045 ) | ( x85 & ~n4050 ) | ( n4045 & ~n4050 ) ;
  assign n4052 = ( x85 & n3837 ) | ( x85 & ~n3926 ) | ( n3837 & ~n3926 ) ;
  assign n4053 = x85 & n3837 ;
  assign n4054 = ( ~n3842 & n4052 ) | ( ~n3842 & n4053 ) | ( n4052 & n4053 ) ;
  assign n4055 = ( n3842 & n4052 ) | ( n3842 & n4053 ) | ( n4052 & n4053 ) ;
  assign n4056 = ( n3842 & n4054 ) | ( n3842 & ~n4055 ) | ( n4054 & ~n4055 ) ;
  assign n4057 = ( x86 & n4051 ) | ( x86 & ~n4056 ) | ( n4051 & ~n4056 ) ;
  assign n4058 = ( x86 & n3843 ) | ( x86 & ~n3926 ) | ( n3843 & ~n3926 ) ;
  assign n4059 = x86 & n3843 ;
  assign n4060 = ( n3848 & n4058 ) | ( n3848 & n4059 ) | ( n4058 & n4059 ) ;
  assign n4061 = ( ~n3848 & n4058 ) | ( ~n3848 & n4059 ) | ( n4058 & n4059 ) ;
  assign n4062 = ( n3848 & ~n4060 ) | ( n3848 & n4061 ) | ( ~n4060 & n4061 ) ;
  assign n4063 = ( x87 & n4057 ) | ( x87 & ~n4062 ) | ( n4057 & ~n4062 ) ;
  assign n4064 = ( x87 & n3849 ) | ( x87 & ~n3926 ) | ( n3849 & ~n3926 ) ;
  assign n4065 = x87 & n3849 ;
  assign n4066 = ( ~n3854 & n4064 ) | ( ~n3854 & n4065 ) | ( n4064 & n4065 ) ;
  assign n4067 = ( n3854 & n4064 ) | ( n3854 & n4065 ) | ( n4064 & n4065 ) ;
  assign n4068 = ( n3854 & n4066 ) | ( n3854 & ~n4067 ) | ( n4066 & ~n4067 ) ;
  assign n4069 = ( x88 & n4063 ) | ( x88 & ~n4068 ) | ( n4063 & ~n4068 ) ;
  assign n4070 = ( x88 & n3855 ) | ( x88 & ~n3926 ) | ( n3855 & ~n3926 ) ;
  assign n4071 = x88 & n3855 ;
  assign n4072 = ( n3860 & n4070 ) | ( n3860 & n4071 ) | ( n4070 & n4071 ) ;
  assign n4073 = ( ~n3860 & n4070 ) | ( ~n3860 & n4071 ) | ( n4070 & n4071 ) ;
  assign n4074 = ( n3860 & ~n4072 ) | ( n3860 & n4073 ) | ( ~n4072 & n4073 ) ;
  assign n4075 = ( x89 & n4069 ) | ( x89 & ~n4074 ) | ( n4069 & ~n4074 ) ;
  assign n4076 = ( x89 & n3861 ) | ( x89 & ~n3926 ) | ( n3861 & ~n3926 ) ;
  assign n4077 = x89 & n3861 ;
  assign n4078 = ( ~n3866 & n4076 ) | ( ~n3866 & n4077 ) | ( n4076 & n4077 ) ;
  assign n4079 = ( n3866 & n4076 ) | ( n3866 & n4077 ) | ( n4076 & n4077 ) ;
  assign n4080 = ( n3866 & n4078 ) | ( n3866 & ~n4079 ) | ( n4078 & ~n4079 ) ;
  assign n4081 = ( x90 & n4075 ) | ( x90 & ~n4080 ) | ( n4075 & ~n4080 ) ;
  assign n4082 = ( x90 & n3867 ) | ( x90 & ~n3926 ) | ( n3867 & ~n3926 ) ;
  assign n4083 = x90 & n3867 ;
  assign n4084 = ( n3872 & n4082 ) | ( n3872 & n4083 ) | ( n4082 & n4083 ) ;
  assign n4085 = ( ~n3872 & n4082 ) | ( ~n3872 & n4083 ) | ( n4082 & n4083 ) ;
  assign n4086 = ( n3872 & ~n4084 ) | ( n3872 & n4085 ) | ( ~n4084 & n4085 ) ;
  assign n4087 = ( x91 & n4081 ) | ( x91 & ~n4086 ) | ( n4081 & ~n4086 ) ;
  assign n4088 = ( x91 & n3873 ) | ( x91 & ~n3926 ) | ( n3873 & ~n3926 ) ;
  assign n4089 = x91 & n3873 ;
  assign n4090 = ( ~n3878 & n4088 ) | ( ~n3878 & n4089 ) | ( n4088 & n4089 ) ;
  assign n4091 = ( n3878 & n4088 ) | ( n3878 & n4089 ) | ( n4088 & n4089 ) ;
  assign n4092 = ( n3878 & n4090 ) | ( n3878 & ~n4091 ) | ( n4090 & ~n4091 ) ;
  assign n4093 = ( x92 & n4087 ) | ( x92 & ~n4092 ) | ( n4087 & ~n4092 ) ;
  assign n4094 = ( x92 & n3879 ) | ( x92 & ~n3926 ) | ( n3879 & ~n3926 ) ;
  assign n4095 = x92 & n3879 ;
  assign n4096 = ( n3884 & n4094 ) | ( n3884 & n4095 ) | ( n4094 & n4095 ) ;
  assign n4097 = ( ~n3884 & n4094 ) | ( ~n3884 & n4095 ) | ( n4094 & n4095 ) ;
  assign n4098 = ( n3884 & ~n4096 ) | ( n3884 & n4097 ) | ( ~n4096 & n4097 ) ;
  assign n4099 = ( x93 & n4093 ) | ( x93 & ~n4098 ) | ( n4093 & ~n4098 ) ;
  assign n4100 = ( x93 & n3885 ) | ( x93 & ~n3926 ) | ( n3885 & ~n3926 ) ;
  assign n4101 = x93 & n3885 ;
  assign n4102 = ( ~n3890 & n4100 ) | ( ~n3890 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4103 = ( n3890 & n4100 ) | ( n3890 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4104 = ( n3890 & n4102 ) | ( n3890 & ~n4103 ) | ( n4102 & ~n4103 ) ;
  assign n4105 = ( x94 & n4099 ) | ( x94 & ~n4104 ) | ( n4099 & ~n4104 ) ;
  assign n4106 = ( x94 & n3891 ) | ( x94 & ~n3926 ) | ( n3891 & ~n3926 ) ;
  assign n4107 = x94 & n3891 ;
  assign n4108 = ( n3896 & n4106 ) | ( n3896 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4109 = ( ~n3896 & n4106 ) | ( ~n3896 & n4107 ) | ( n4106 & n4107 ) ;
  assign n4110 = ( n3896 & ~n4108 ) | ( n3896 & n4109 ) | ( ~n4108 & n4109 ) ;
  assign n4111 = ( x95 & n4105 ) | ( x95 & ~n4110 ) | ( n4105 & ~n4110 ) ;
  assign n4112 = ( x95 & n3897 ) | ( x95 & ~n3926 ) | ( n3897 & ~n3926 ) ;
  assign n4113 = x95 & n3897 ;
  assign n4114 = ( ~n3902 & n4112 ) | ( ~n3902 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4115 = ( n3902 & n4112 ) | ( n3902 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4116 = ( n3902 & n4114 ) | ( n3902 & ~n4115 ) | ( n4114 & ~n4115 ) ;
  assign n4117 = ( x96 & n4111 ) | ( x96 & ~n4116 ) | ( n4111 & ~n4116 ) ;
  assign n4118 = ( x96 & n3903 ) | ( x96 & ~n3926 ) | ( n3903 & ~n3926 ) ;
  assign n4119 = x96 & n3903 ;
  assign n4120 = ( n3908 & n4118 ) | ( n3908 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4121 = ( ~n3908 & n4118 ) | ( ~n3908 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4122 = ( n3908 & ~n4120 ) | ( n3908 & n4121 ) | ( ~n4120 & n4121 ) ;
  assign n4123 = ( x97 & n4117 ) | ( x97 & ~n4122 ) | ( n4117 & ~n4122 ) ;
  assign n4124 = ( x97 & n3909 ) | ( x97 & ~n3926 ) | ( n3909 & ~n3926 ) ;
  assign n4125 = x97 & n3909 ;
  assign n4126 = ( ~n3914 & n4124 ) | ( ~n3914 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4127 = ( n3914 & n4124 ) | ( n3914 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4128 = ( n3914 & n4126 ) | ( n3914 & ~n4127 ) | ( n4126 & ~n4127 ) ;
  assign n4129 = ( x98 & n4123 ) | ( x98 & ~n4128 ) | ( n4123 & ~n4128 ) ;
  assign n4130 = ( x98 & n3915 ) | ( x98 & ~n3926 ) | ( n3915 & ~n3926 ) ;
  assign n4131 = x98 & n3915 ;
  assign n4132 = ( ~n3920 & n4130 ) | ( ~n3920 & n4131 ) | ( n4130 & n4131 ) ;
  assign n4133 = ( n3920 & n4130 ) | ( n3920 & n4131 ) | ( n4130 & n4131 ) ;
  assign n4134 = ( n3920 & n4132 ) | ( n3920 & ~n4133 ) | ( n4132 & ~n4133 ) ;
  assign n4135 = ( x99 & n4129 ) | ( x99 & ~n4134 ) | ( n4129 & ~n4134 ) ;
  assign n4136 = x100 | n4135 ;
  assign n4137 = ( x100 & n157 ) | ( x100 & n4135 ) | ( n157 & n4135 ) ;
  assign n4138 = ( n3924 & ~n4136 ) | ( n3924 & n4137 ) | ( ~n4136 & n4137 ) ;
  assign n4139 = ( x100 & ~n3924 ) | ( x100 & n4135 ) | ( ~n3924 & n4135 ) ;
  assign n4140 = n157 | n4139 ;
  assign n4141 = ( x27 & ~x64 ) | ( x27 & n4140 ) | ( ~x64 & n4140 ) ;
  assign n4142 = ~x27 & n4140 ;
  assign n4143 = ( n3930 & n4141 ) | ( n3930 & ~n4142 ) | ( n4141 & ~n4142 ) ;
  assign n4144 = ~x26 & x64 ;
  assign n4145 = ( x65 & ~n4143 ) | ( x65 & n4144 ) | ( ~n4143 & n4144 ) ;
  assign n4146 = ( x65 & n3930 ) | ( x65 & ~n4140 ) | ( n3930 & ~n4140 ) ;
  assign n4147 = x65 & n3930 ;
  assign n4148 = ( n3929 & n4146 ) | ( n3929 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4149 = ( ~n3929 & n4146 ) | ( ~n3929 & n4147 ) | ( n4146 & n4147 ) ;
  assign n4150 = ( n3929 & ~n4148 ) | ( n3929 & n4149 ) | ( ~n4148 & n4149 ) ;
  assign n4151 = ( x66 & n4145 ) | ( x66 & ~n4150 ) | ( n4145 & ~n4150 ) ;
  assign n4152 = ( x66 & n3931 ) | ( x66 & ~n4140 ) | ( n3931 & ~n4140 ) ;
  assign n4153 = x66 & n3931 ;
  assign n4154 = ( n3936 & n4152 ) | ( n3936 & n4153 ) | ( n4152 & n4153 ) ;
  assign n4155 = ( ~n3936 & n4152 ) | ( ~n3936 & n4153 ) | ( n4152 & n4153 ) ;
  assign n4156 = ( n3936 & ~n4154 ) | ( n3936 & n4155 ) | ( ~n4154 & n4155 ) ;
  assign n4157 = ( x67 & n4151 ) | ( x67 & ~n4156 ) | ( n4151 & ~n4156 ) ;
  assign n4158 = ( x67 & n3937 ) | ( x67 & ~n4140 ) | ( n3937 & ~n4140 ) ;
  assign n4159 = x67 & n3937 ;
  assign n4160 = ( ~n3942 & n4158 ) | ( ~n3942 & n4159 ) | ( n4158 & n4159 ) ;
  assign n4161 = ( n3942 & n4158 ) | ( n3942 & n4159 ) | ( n4158 & n4159 ) ;
  assign n4162 = ( n3942 & n4160 ) | ( n3942 & ~n4161 ) | ( n4160 & ~n4161 ) ;
  assign n4163 = ( x68 & n4157 ) | ( x68 & ~n4162 ) | ( n4157 & ~n4162 ) ;
  assign n4164 = ( x68 & n3943 ) | ( x68 & ~n4140 ) | ( n3943 & ~n4140 ) ;
  assign n4165 = x68 & n3943 ;
  assign n4166 = ( n3948 & n4164 ) | ( n3948 & n4165 ) | ( n4164 & n4165 ) ;
  assign n4167 = ( ~n3948 & n4164 ) | ( ~n3948 & n4165 ) | ( n4164 & n4165 ) ;
  assign n4168 = ( n3948 & ~n4166 ) | ( n3948 & n4167 ) | ( ~n4166 & n4167 ) ;
  assign n4169 = ( x69 & n4163 ) | ( x69 & ~n4168 ) | ( n4163 & ~n4168 ) ;
  assign n4170 = ( x69 & n3949 ) | ( x69 & ~n4140 ) | ( n3949 & ~n4140 ) ;
  assign n4171 = x69 & n3949 ;
  assign n4172 = ( ~n3954 & n4170 ) | ( ~n3954 & n4171 ) | ( n4170 & n4171 ) ;
  assign n4173 = ( n3954 & n4170 ) | ( n3954 & n4171 ) | ( n4170 & n4171 ) ;
  assign n4174 = ( n3954 & n4172 ) | ( n3954 & ~n4173 ) | ( n4172 & ~n4173 ) ;
  assign n4175 = ( x70 & n4169 ) | ( x70 & ~n4174 ) | ( n4169 & ~n4174 ) ;
  assign n4176 = ( x70 & n3955 ) | ( x70 & ~n4140 ) | ( n3955 & ~n4140 ) ;
  assign n4177 = x70 & n3955 ;
  assign n4178 = ( n3960 & n4176 ) | ( n3960 & n4177 ) | ( n4176 & n4177 ) ;
  assign n4179 = ( ~n3960 & n4176 ) | ( ~n3960 & n4177 ) | ( n4176 & n4177 ) ;
  assign n4180 = ( n3960 & ~n4178 ) | ( n3960 & n4179 ) | ( ~n4178 & n4179 ) ;
  assign n4181 = ( x71 & n4175 ) | ( x71 & ~n4180 ) | ( n4175 & ~n4180 ) ;
  assign n4182 = ( x71 & n3961 ) | ( x71 & ~n4140 ) | ( n3961 & ~n4140 ) ;
  assign n4183 = x71 & n3961 ;
  assign n4184 = ( ~n3966 & n4182 ) | ( ~n3966 & n4183 ) | ( n4182 & n4183 ) ;
  assign n4185 = ( n3966 & n4182 ) | ( n3966 & n4183 ) | ( n4182 & n4183 ) ;
  assign n4186 = ( n3966 & n4184 ) | ( n3966 & ~n4185 ) | ( n4184 & ~n4185 ) ;
  assign n4187 = ( x72 & n4181 ) | ( x72 & ~n4186 ) | ( n4181 & ~n4186 ) ;
  assign n4188 = ( x72 & n3967 ) | ( x72 & ~n4140 ) | ( n3967 & ~n4140 ) ;
  assign n4189 = x72 & n3967 ;
  assign n4190 = ( n3972 & n4188 ) | ( n3972 & n4189 ) | ( n4188 & n4189 ) ;
  assign n4191 = ( ~n3972 & n4188 ) | ( ~n3972 & n4189 ) | ( n4188 & n4189 ) ;
  assign n4192 = ( n3972 & ~n4190 ) | ( n3972 & n4191 ) | ( ~n4190 & n4191 ) ;
  assign n4193 = ( x73 & n4187 ) | ( x73 & ~n4192 ) | ( n4187 & ~n4192 ) ;
  assign n4194 = ( x73 & n3973 ) | ( x73 & ~n4140 ) | ( n3973 & ~n4140 ) ;
  assign n4195 = x73 & n3973 ;
  assign n4196 = ( ~n3978 & n4194 ) | ( ~n3978 & n4195 ) | ( n4194 & n4195 ) ;
  assign n4197 = ( n3978 & n4194 ) | ( n3978 & n4195 ) | ( n4194 & n4195 ) ;
  assign n4198 = ( n3978 & n4196 ) | ( n3978 & ~n4197 ) | ( n4196 & ~n4197 ) ;
  assign n4199 = ( x74 & n4193 ) | ( x74 & ~n4198 ) | ( n4193 & ~n4198 ) ;
  assign n4200 = ( x74 & n3979 ) | ( x74 & ~n4140 ) | ( n3979 & ~n4140 ) ;
  assign n4201 = x74 & n3979 ;
  assign n4202 = ( n3984 & n4200 ) | ( n3984 & n4201 ) | ( n4200 & n4201 ) ;
  assign n4203 = ( ~n3984 & n4200 ) | ( ~n3984 & n4201 ) | ( n4200 & n4201 ) ;
  assign n4204 = ( n3984 & ~n4202 ) | ( n3984 & n4203 ) | ( ~n4202 & n4203 ) ;
  assign n4205 = ( x75 & n4199 ) | ( x75 & ~n4204 ) | ( n4199 & ~n4204 ) ;
  assign n4206 = ( x75 & n3985 ) | ( x75 & ~n4140 ) | ( n3985 & ~n4140 ) ;
  assign n4207 = x75 & n3985 ;
  assign n4208 = ( ~n3990 & n4206 ) | ( ~n3990 & n4207 ) | ( n4206 & n4207 ) ;
  assign n4209 = ( n3990 & n4206 ) | ( n3990 & n4207 ) | ( n4206 & n4207 ) ;
  assign n4210 = ( n3990 & n4208 ) | ( n3990 & ~n4209 ) | ( n4208 & ~n4209 ) ;
  assign n4211 = ( x76 & n4205 ) | ( x76 & ~n4210 ) | ( n4205 & ~n4210 ) ;
  assign n4212 = ( x76 & n3991 ) | ( x76 & ~n4140 ) | ( n3991 & ~n4140 ) ;
  assign n4213 = x76 & n3991 ;
  assign n4214 = ( n3996 & n4212 ) | ( n3996 & n4213 ) | ( n4212 & n4213 ) ;
  assign n4215 = ( ~n3996 & n4212 ) | ( ~n3996 & n4213 ) | ( n4212 & n4213 ) ;
  assign n4216 = ( n3996 & ~n4214 ) | ( n3996 & n4215 ) | ( ~n4214 & n4215 ) ;
  assign n4217 = ( x77 & n4211 ) | ( x77 & ~n4216 ) | ( n4211 & ~n4216 ) ;
  assign n4218 = ( x77 & n3997 ) | ( x77 & ~n4140 ) | ( n3997 & ~n4140 ) ;
  assign n4219 = x77 & n3997 ;
  assign n4220 = ( ~n4002 & n4218 ) | ( ~n4002 & n4219 ) | ( n4218 & n4219 ) ;
  assign n4221 = ( n4002 & n4218 ) | ( n4002 & n4219 ) | ( n4218 & n4219 ) ;
  assign n4222 = ( n4002 & n4220 ) | ( n4002 & ~n4221 ) | ( n4220 & ~n4221 ) ;
  assign n4223 = ( x78 & n4217 ) | ( x78 & ~n4222 ) | ( n4217 & ~n4222 ) ;
  assign n4224 = ( x78 & n4003 ) | ( x78 & ~n4140 ) | ( n4003 & ~n4140 ) ;
  assign n4225 = x78 & n4003 ;
  assign n4226 = ( n4008 & n4224 ) | ( n4008 & n4225 ) | ( n4224 & n4225 ) ;
  assign n4227 = ( ~n4008 & n4224 ) | ( ~n4008 & n4225 ) | ( n4224 & n4225 ) ;
  assign n4228 = ( n4008 & ~n4226 ) | ( n4008 & n4227 ) | ( ~n4226 & n4227 ) ;
  assign n4229 = ( x79 & n4223 ) | ( x79 & ~n4228 ) | ( n4223 & ~n4228 ) ;
  assign n4230 = ( x79 & n4009 ) | ( x79 & ~n4140 ) | ( n4009 & ~n4140 ) ;
  assign n4231 = x79 & n4009 ;
  assign n4232 = ( ~n4014 & n4230 ) | ( ~n4014 & n4231 ) | ( n4230 & n4231 ) ;
  assign n4233 = ( n4014 & n4230 ) | ( n4014 & n4231 ) | ( n4230 & n4231 ) ;
  assign n4234 = ( n4014 & n4232 ) | ( n4014 & ~n4233 ) | ( n4232 & ~n4233 ) ;
  assign n4235 = ( x80 & n4229 ) | ( x80 & ~n4234 ) | ( n4229 & ~n4234 ) ;
  assign n4236 = ( x80 & n4015 ) | ( x80 & ~n4140 ) | ( n4015 & ~n4140 ) ;
  assign n4237 = x80 & n4015 ;
  assign n4238 = ( n4020 & n4236 ) | ( n4020 & n4237 ) | ( n4236 & n4237 ) ;
  assign n4239 = ( ~n4020 & n4236 ) | ( ~n4020 & n4237 ) | ( n4236 & n4237 ) ;
  assign n4240 = ( n4020 & ~n4238 ) | ( n4020 & n4239 ) | ( ~n4238 & n4239 ) ;
  assign n4241 = ( x81 & n4235 ) | ( x81 & ~n4240 ) | ( n4235 & ~n4240 ) ;
  assign n4242 = ( x81 & n4021 ) | ( x81 & ~n4140 ) | ( n4021 & ~n4140 ) ;
  assign n4243 = x81 & n4021 ;
  assign n4244 = ( ~n4026 & n4242 ) | ( ~n4026 & n4243 ) | ( n4242 & n4243 ) ;
  assign n4245 = ( n4026 & n4242 ) | ( n4026 & n4243 ) | ( n4242 & n4243 ) ;
  assign n4246 = ( n4026 & n4244 ) | ( n4026 & ~n4245 ) | ( n4244 & ~n4245 ) ;
  assign n4247 = ( x82 & n4241 ) | ( x82 & ~n4246 ) | ( n4241 & ~n4246 ) ;
  assign n4248 = ( x82 & n4027 ) | ( x82 & ~n4140 ) | ( n4027 & ~n4140 ) ;
  assign n4249 = x82 & n4027 ;
  assign n4250 = ( n4032 & n4248 ) | ( n4032 & n4249 ) | ( n4248 & n4249 ) ;
  assign n4251 = ( ~n4032 & n4248 ) | ( ~n4032 & n4249 ) | ( n4248 & n4249 ) ;
  assign n4252 = ( n4032 & ~n4250 ) | ( n4032 & n4251 ) | ( ~n4250 & n4251 ) ;
  assign n4253 = ( x83 & n4247 ) | ( x83 & ~n4252 ) | ( n4247 & ~n4252 ) ;
  assign n4254 = ( x83 & n4033 ) | ( x83 & ~n4140 ) | ( n4033 & ~n4140 ) ;
  assign n4255 = x83 & n4033 ;
  assign n4256 = ( ~n4038 & n4254 ) | ( ~n4038 & n4255 ) | ( n4254 & n4255 ) ;
  assign n4257 = ( n4038 & n4254 ) | ( n4038 & n4255 ) | ( n4254 & n4255 ) ;
  assign n4258 = ( n4038 & n4256 ) | ( n4038 & ~n4257 ) | ( n4256 & ~n4257 ) ;
  assign n4259 = ( x84 & n4253 ) | ( x84 & ~n4258 ) | ( n4253 & ~n4258 ) ;
  assign n4260 = ( x84 & n4039 ) | ( x84 & ~n4140 ) | ( n4039 & ~n4140 ) ;
  assign n4261 = x84 & n4039 ;
  assign n4262 = ( n4044 & n4260 ) | ( n4044 & n4261 ) | ( n4260 & n4261 ) ;
  assign n4263 = ( ~n4044 & n4260 ) | ( ~n4044 & n4261 ) | ( n4260 & n4261 ) ;
  assign n4264 = ( n4044 & ~n4262 ) | ( n4044 & n4263 ) | ( ~n4262 & n4263 ) ;
  assign n4265 = ( x85 & n4259 ) | ( x85 & ~n4264 ) | ( n4259 & ~n4264 ) ;
  assign n4266 = ( x85 & n4045 ) | ( x85 & ~n4140 ) | ( n4045 & ~n4140 ) ;
  assign n4267 = x85 & n4045 ;
  assign n4268 = ( ~n4050 & n4266 ) | ( ~n4050 & n4267 ) | ( n4266 & n4267 ) ;
  assign n4269 = ( n4050 & n4266 ) | ( n4050 & n4267 ) | ( n4266 & n4267 ) ;
  assign n4270 = ( n4050 & n4268 ) | ( n4050 & ~n4269 ) | ( n4268 & ~n4269 ) ;
  assign n4271 = ( x86 & n4265 ) | ( x86 & ~n4270 ) | ( n4265 & ~n4270 ) ;
  assign n4272 = ( x86 & n4051 ) | ( x86 & ~n4140 ) | ( n4051 & ~n4140 ) ;
  assign n4273 = x86 & n4051 ;
  assign n4274 = ( n4056 & n4272 ) | ( n4056 & n4273 ) | ( n4272 & n4273 ) ;
  assign n4275 = ( ~n4056 & n4272 ) | ( ~n4056 & n4273 ) | ( n4272 & n4273 ) ;
  assign n4276 = ( n4056 & ~n4274 ) | ( n4056 & n4275 ) | ( ~n4274 & n4275 ) ;
  assign n4277 = ( x87 & n4271 ) | ( x87 & ~n4276 ) | ( n4271 & ~n4276 ) ;
  assign n4278 = ( x87 & n4057 ) | ( x87 & ~n4140 ) | ( n4057 & ~n4140 ) ;
  assign n4279 = x87 & n4057 ;
  assign n4280 = ( ~n4062 & n4278 ) | ( ~n4062 & n4279 ) | ( n4278 & n4279 ) ;
  assign n4281 = ( n4062 & n4278 ) | ( n4062 & n4279 ) | ( n4278 & n4279 ) ;
  assign n4282 = ( n4062 & n4280 ) | ( n4062 & ~n4281 ) | ( n4280 & ~n4281 ) ;
  assign n4283 = ( x88 & n4277 ) | ( x88 & ~n4282 ) | ( n4277 & ~n4282 ) ;
  assign n4284 = ( x88 & n4063 ) | ( x88 & ~n4140 ) | ( n4063 & ~n4140 ) ;
  assign n4285 = x88 & n4063 ;
  assign n4286 = ( n4068 & n4284 ) | ( n4068 & n4285 ) | ( n4284 & n4285 ) ;
  assign n4287 = ( ~n4068 & n4284 ) | ( ~n4068 & n4285 ) | ( n4284 & n4285 ) ;
  assign n4288 = ( n4068 & ~n4286 ) | ( n4068 & n4287 ) | ( ~n4286 & n4287 ) ;
  assign n4289 = ( x89 & n4283 ) | ( x89 & ~n4288 ) | ( n4283 & ~n4288 ) ;
  assign n4290 = ( x89 & n4069 ) | ( x89 & ~n4140 ) | ( n4069 & ~n4140 ) ;
  assign n4291 = x89 & n4069 ;
  assign n4292 = ( ~n4074 & n4290 ) | ( ~n4074 & n4291 ) | ( n4290 & n4291 ) ;
  assign n4293 = ( n4074 & n4290 ) | ( n4074 & n4291 ) | ( n4290 & n4291 ) ;
  assign n4294 = ( n4074 & n4292 ) | ( n4074 & ~n4293 ) | ( n4292 & ~n4293 ) ;
  assign n4295 = ( x90 & n4289 ) | ( x90 & ~n4294 ) | ( n4289 & ~n4294 ) ;
  assign n4296 = ( x90 & n4075 ) | ( x90 & ~n4140 ) | ( n4075 & ~n4140 ) ;
  assign n4297 = x90 & n4075 ;
  assign n4298 = ( n4080 & n4296 ) | ( n4080 & n4297 ) | ( n4296 & n4297 ) ;
  assign n4299 = ( ~n4080 & n4296 ) | ( ~n4080 & n4297 ) | ( n4296 & n4297 ) ;
  assign n4300 = ( n4080 & ~n4298 ) | ( n4080 & n4299 ) | ( ~n4298 & n4299 ) ;
  assign n4301 = ( x91 & n4295 ) | ( x91 & ~n4300 ) | ( n4295 & ~n4300 ) ;
  assign n4302 = ( x91 & n4081 ) | ( x91 & ~n4140 ) | ( n4081 & ~n4140 ) ;
  assign n4303 = x91 & n4081 ;
  assign n4304 = ( ~n4086 & n4302 ) | ( ~n4086 & n4303 ) | ( n4302 & n4303 ) ;
  assign n4305 = ( n4086 & n4302 ) | ( n4086 & n4303 ) | ( n4302 & n4303 ) ;
  assign n4306 = ( n4086 & n4304 ) | ( n4086 & ~n4305 ) | ( n4304 & ~n4305 ) ;
  assign n4307 = ( x92 & n4301 ) | ( x92 & ~n4306 ) | ( n4301 & ~n4306 ) ;
  assign n4308 = ( x92 & n4087 ) | ( x92 & ~n4140 ) | ( n4087 & ~n4140 ) ;
  assign n4309 = x92 & n4087 ;
  assign n4310 = ( n4092 & n4308 ) | ( n4092 & n4309 ) | ( n4308 & n4309 ) ;
  assign n4311 = ( ~n4092 & n4308 ) | ( ~n4092 & n4309 ) | ( n4308 & n4309 ) ;
  assign n4312 = ( n4092 & ~n4310 ) | ( n4092 & n4311 ) | ( ~n4310 & n4311 ) ;
  assign n4313 = ( x93 & n4307 ) | ( x93 & ~n4312 ) | ( n4307 & ~n4312 ) ;
  assign n4314 = ( x93 & n4093 ) | ( x93 & ~n4140 ) | ( n4093 & ~n4140 ) ;
  assign n4315 = x93 & n4093 ;
  assign n4316 = ( ~n4098 & n4314 ) | ( ~n4098 & n4315 ) | ( n4314 & n4315 ) ;
  assign n4317 = ( n4098 & n4314 ) | ( n4098 & n4315 ) | ( n4314 & n4315 ) ;
  assign n4318 = ( n4098 & n4316 ) | ( n4098 & ~n4317 ) | ( n4316 & ~n4317 ) ;
  assign n4319 = ( x94 & n4313 ) | ( x94 & ~n4318 ) | ( n4313 & ~n4318 ) ;
  assign n4320 = ( x94 & n4099 ) | ( x94 & ~n4140 ) | ( n4099 & ~n4140 ) ;
  assign n4321 = x94 & n4099 ;
  assign n4322 = ( n4104 & n4320 ) | ( n4104 & n4321 ) | ( n4320 & n4321 ) ;
  assign n4323 = ( ~n4104 & n4320 ) | ( ~n4104 & n4321 ) | ( n4320 & n4321 ) ;
  assign n4324 = ( n4104 & ~n4322 ) | ( n4104 & n4323 ) | ( ~n4322 & n4323 ) ;
  assign n4325 = ( x95 & n4319 ) | ( x95 & ~n4324 ) | ( n4319 & ~n4324 ) ;
  assign n4326 = ( x95 & n4105 ) | ( x95 & ~n4140 ) | ( n4105 & ~n4140 ) ;
  assign n4327 = x95 & n4105 ;
  assign n4328 = ( ~n4110 & n4326 ) | ( ~n4110 & n4327 ) | ( n4326 & n4327 ) ;
  assign n4329 = ( n4110 & n4326 ) | ( n4110 & n4327 ) | ( n4326 & n4327 ) ;
  assign n4330 = ( n4110 & n4328 ) | ( n4110 & ~n4329 ) | ( n4328 & ~n4329 ) ;
  assign n4331 = ( x96 & n4325 ) | ( x96 & ~n4330 ) | ( n4325 & ~n4330 ) ;
  assign n4332 = ( x96 & n4111 ) | ( x96 & ~n4140 ) | ( n4111 & ~n4140 ) ;
  assign n4333 = x96 & n4111 ;
  assign n4334 = ( n4116 & n4332 ) | ( n4116 & n4333 ) | ( n4332 & n4333 ) ;
  assign n4335 = ( ~n4116 & n4332 ) | ( ~n4116 & n4333 ) | ( n4332 & n4333 ) ;
  assign n4336 = ( n4116 & ~n4334 ) | ( n4116 & n4335 ) | ( ~n4334 & n4335 ) ;
  assign n4337 = ( x97 & n4331 ) | ( x97 & ~n4336 ) | ( n4331 & ~n4336 ) ;
  assign n4338 = ( x97 & n4117 ) | ( x97 & ~n4140 ) | ( n4117 & ~n4140 ) ;
  assign n4339 = x97 & n4117 ;
  assign n4340 = ( ~n4122 & n4338 ) | ( ~n4122 & n4339 ) | ( n4338 & n4339 ) ;
  assign n4341 = ( n4122 & n4338 ) | ( n4122 & n4339 ) | ( n4338 & n4339 ) ;
  assign n4342 = ( n4122 & n4340 ) | ( n4122 & ~n4341 ) | ( n4340 & ~n4341 ) ;
  assign n4343 = ( x98 & n4337 ) | ( x98 & ~n4342 ) | ( n4337 & ~n4342 ) ;
  assign n4344 = ( x98 & n4123 ) | ( x98 & ~n4140 ) | ( n4123 & ~n4140 ) ;
  assign n4345 = x98 & n4123 ;
  assign n4346 = ( n4128 & n4344 ) | ( n4128 & n4345 ) | ( n4344 & n4345 ) ;
  assign n4347 = ( ~n4128 & n4344 ) | ( ~n4128 & n4345 ) | ( n4344 & n4345 ) ;
  assign n4348 = ( n4128 & ~n4346 ) | ( n4128 & n4347 ) | ( ~n4346 & n4347 ) ;
  assign n4349 = ( x99 & n4343 ) | ( x99 & ~n4348 ) | ( n4343 & ~n4348 ) ;
  assign n4350 = ( x99 & n4129 ) | ( x99 & ~n4140 ) | ( n4129 & ~n4140 ) ;
  assign n4351 = x99 & n4129 ;
  assign n4352 = ( n4134 & n4350 ) | ( n4134 & n4351 ) | ( n4350 & n4351 ) ;
  assign n4353 = ( ~n4134 & n4350 ) | ( ~n4134 & n4351 ) | ( n4350 & n4351 ) ;
  assign n4354 = ( n4134 & ~n4352 ) | ( n4134 & n4353 ) | ( ~n4352 & n4353 ) ;
  assign n4355 = ( x100 & n4349 ) | ( x100 & ~n4354 ) | ( n4349 & ~n4354 ) ;
  assign n4356 = x101 | n4355 ;
  assign n4357 = x102 | n155 ;
  assign n4358 = ( x101 & n4355 ) | ( x101 & n4357 ) | ( n4355 & n4357 ) ;
  assign n4359 = ( n4138 & ~n4356 ) | ( n4138 & n4358 ) | ( ~n4356 & n4358 ) ;
  assign n4360 = ( x101 & ~n4138 ) | ( x101 & n4355 ) | ( ~n4138 & n4355 ) ;
  assign n4361 = n4357 | n4360 ;
  assign n4362 = ( x26 & ~x64 ) | ( x26 & n4361 ) | ( ~x64 & n4361 ) ;
  assign n4363 = ~x26 & n4361 ;
  assign n4364 = ( n4144 & n4362 ) | ( n4144 & ~n4363 ) | ( n4362 & ~n4363 ) ;
  assign n4365 = ~x25 & x64 ;
  assign n4366 = ( x65 & ~n4364 ) | ( x65 & n4365 ) | ( ~n4364 & n4365 ) ;
  assign n4367 = ( x65 & n4144 ) | ( x65 & ~n4361 ) | ( n4144 & ~n4361 ) ;
  assign n4368 = x65 & n4144 ;
  assign n4369 = ( n4143 & n4367 ) | ( n4143 & n4368 ) | ( n4367 & n4368 ) ;
  assign n4370 = ( ~n4143 & n4367 ) | ( ~n4143 & n4368 ) | ( n4367 & n4368 ) ;
  assign n4371 = ( n4143 & ~n4369 ) | ( n4143 & n4370 ) | ( ~n4369 & n4370 ) ;
  assign n4372 = ( x66 & n4366 ) | ( x66 & ~n4371 ) | ( n4366 & ~n4371 ) ;
  assign n4373 = ( x66 & n4145 ) | ( x66 & ~n4361 ) | ( n4145 & ~n4361 ) ;
  assign n4374 = x66 & n4145 ;
  assign n4375 = ( n4150 & n4373 ) | ( n4150 & n4374 ) | ( n4373 & n4374 ) ;
  assign n4376 = ( ~n4150 & n4373 ) | ( ~n4150 & n4374 ) | ( n4373 & n4374 ) ;
  assign n4377 = ( n4150 & ~n4375 ) | ( n4150 & n4376 ) | ( ~n4375 & n4376 ) ;
  assign n4378 = ( x67 & n4372 ) | ( x67 & ~n4377 ) | ( n4372 & ~n4377 ) ;
  assign n4379 = ( x67 & n4151 ) | ( x67 & ~n4361 ) | ( n4151 & ~n4361 ) ;
  assign n4380 = x67 & n4151 ;
  assign n4381 = ( ~n4156 & n4379 ) | ( ~n4156 & n4380 ) | ( n4379 & n4380 ) ;
  assign n4382 = ( n4156 & n4379 ) | ( n4156 & n4380 ) | ( n4379 & n4380 ) ;
  assign n4383 = ( n4156 & n4381 ) | ( n4156 & ~n4382 ) | ( n4381 & ~n4382 ) ;
  assign n4384 = ( x68 & n4378 ) | ( x68 & ~n4383 ) | ( n4378 & ~n4383 ) ;
  assign n4385 = ( x68 & n4157 ) | ( x68 & ~n4361 ) | ( n4157 & ~n4361 ) ;
  assign n4386 = x68 & n4157 ;
  assign n4387 = ( n4162 & n4385 ) | ( n4162 & n4386 ) | ( n4385 & n4386 ) ;
  assign n4388 = ( ~n4162 & n4385 ) | ( ~n4162 & n4386 ) | ( n4385 & n4386 ) ;
  assign n4389 = ( n4162 & ~n4387 ) | ( n4162 & n4388 ) | ( ~n4387 & n4388 ) ;
  assign n4390 = ( x69 & n4384 ) | ( x69 & ~n4389 ) | ( n4384 & ~n4389 ) ;
  assign n4391 = ( x69 & n4163 ) | ( x69 & ~n4361 ) | ( n4163 & ~n4361 ) ;
  assign n4392 = x69 & n4163 ;
  assign n4393 = ( ~n4168 & n4391 ) | ( ~n4168 & n4392 ) | ( n4391 & n4392 ) ;
  assign n4394 = ( n4168 & n4391 ) | ( n4168 & n4392 ) | ( n4391 & n4392 ) ;
  assign n4395 = ( n4168 & n4393 ) | ( n4168 & ~n4394 ) | ( n4393 & ~n4394 ) ;
  assign n4396 = ( x70 & n4390 ) | ( x70 & ~n4395 ) | ( n4390 & ~n4395 ) ;
  assign n4397 = ( x70 & n4169 ) | ( x70 & ~n4361 ) | ( n4169 & ~n4361 ) ;
  assign n4398 = x70 & n4169 ;
  assign n4399 = ( n4174 & n4397 ) | ( n4174 & n4398 ) | ( n4397 & n4398 ) ;
  assign n4400 = ( ~n4174 & n4397 ) | ( ~n4174 & n4398 ) | ( n4397 & n4398 ) ;
  assign n4401 = ( n4174 & ~n4399 ) | ( n4174 & n4400 ) | ( ~n4399 & n4400 ) ;
  assign n4402 = ( x71 & n4396 ) | ( x71 & ~n4401 ) | ( n4396 & ~n4401 ) ;
  assign n4403 = ( x71 & n4175 ) | ( x71 & ~n4361 ) | ( n4175 & ~n4361 ) ;
  assign n4404 = x71 & n4175 ;
  assign n4405 = ( ~n4180 & n4403 ) | ( ~n4180 & n4404 ) | ( n4403 & n4404 ) ;
  assign n4406 = ( n4180 & n4403 ) | ( n4180 & n4404 ) | ( n4403 & n4404 ) ;
  assign n4407 = ( n4180 & n4405 ) | ( n4180 & ~n4406 ) | ( n4405 & ~n4406 ) ;
  assign n4408 = ( x72 & n4402 ) | ( x72 & ~n4407 ) | ( n4402 & ~n4407 ) ;
  assign n4409 = ( x72 & n4181 ) | ( x72 & ~n4361 ) | ( n4181 & ~n4361 ) ;
  assign n4410 = x72 & n4181 ;
  assign n4411 = ( n4186 & n4409 ) | ( n4186 & n4410 ) | ( n4409 & n4410 ) ;
  assign n4412 = ( ~n4186 & n4409 ) | ( ~n4186 & n4410 ) | ( n4409 & n4410 ) ;
  assign n4413 = ( n4186 & ~n4411 ) | ( n4186 & n4412 ) | ( ~n4411 & n4412 ) ;
  assign n4414 = ( x73 & n4408 ) | ( x73 & ~n4413 ) | ( n4408 & ~n4413 ) ;
  assign n4415 = ( x73 & n4187 ) | ( x73 & ~n4361 ) | ( n4187 & ~n4361 ) ;
  assign n4416 = x73 & n4187 ;
  assign n4417 = ( ~n4192 & n4415 ) | ( ~n4192 & n4416 ) | ( n4415 & n4416 ) ;
  assign n4418 = ( n4192 & n4415 ) | ( n4192 & n4416 ) | ( n4415 & n4416 ) ;
  assign n4419 = ( n4192 & n4417 ) | ( n4192 & ~n4418 ) | ( n4417 & ~n4418 ) ;
  assign n4420 = ( x74 & n4414 ) | ( x74 & ~n4419 ) | ( n4414 & ~n4419 ) ;
  assign n4421 = ( x74 & n4193 ) | ( x74 & ~n4361 ) | ( n4193 & ~n4361 ) ;
  assign n4422 = x74 & n4193 ;
  assign n4423 = ( n4198 & n4421 ) | ( n4198 & n4422 ) | ( n4421 & n4422 ) ;
  assign n4424 = ( ~n4198 & n4421 ) | ( ~n4198 & n4422 ) | ( n4421 & n4422 ) ;
  assign n4425 = ( n4198 & ~n4423 ) | ( n4198 & n4424 ) | ( ~n4423 & n4424 ) ;
  assign n4426 = ( x75 & n4420 ) | ( x75 & ~n4425 ) | ( n4420 & ~n4425 ) ;
  assign n4427 = ( x75 & n4199 ) | ( x75 & ~n4361 ) | ( n4199 & ~n4361 ) ;
  assign n4428 = x75 & n4199 ;
  assign n4429 = ( ~n4204 & n4427 ) | ( ~n4204 & n4428 ) | ( n4427 & n4428 ) ;
  assign n4430 = ( n4204 & n4427 ) | ( n4204 & n4428 ) | ( n4427 & n4428 ) ;
  assign n4431 = ( n4204 & n4429 ) | ( n4204 & ~n4430 ) | ( n4429 & ~n4430 ) ;
  assign n4432 = ( x76 & n4426 ) | ( x76 & ~n4431 ) | ( n4426 & ~n4431 ) ;
  assign n4433 = ( x76 & n4205 ) | ( x76 & ~n4361 ) | ( n4205 & ~n4361 ) ;
  assign n4434 = x76 & n4205 ;
  assign n4435 = ( n4210 & n4433 ) | ( n4210 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4436 = ( ~n4210 & n4433 ) | ( ~n4210 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4437 = ( n4210 & ~n4435 ) | ( n4210 & n4436 ) | ( ~n4435 & n4436 ) ;
  assign n4438 = ( x77 & n4432 ) | ( x77 & ~n4437 ) | ( n4432 & ~n4437 ) ;
  assign n4439 = ( x77 & n4211 ) | ( x77 & ~n4361 ) | ( n4211 & ~n4361 ) ;
  assign n4440 = x77 & n4211 ;
  assign n4441 = ( ~n4216 & n4439 ) | ( ~n4216 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4442 = ( n4216 & n4439 ) | ( n4216 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4443 = ( n4216 & n4441 ) | ( n4216 & ~n4442 ) | ( n4441 & ~n4442 ) ;
  assign n4444 = ( x78 & n4438 ) | ( x78 & ~n4443 ) | ( n4438 & ~n4443 ) ;
  assign n4445 = ( x78 & n4217 ) | ( x78 & ~n4361 ) | ( n4217 & ~n4361 ) ;
  assign n4446 = x78 & n4217 ;
  assign n4447 = ( n4222 & n4445 ) | ( n4222 & n4446 ) | ( n4445 & n4446 ) ;
  assign n4448 = ( ~n4222 & n4445 ) | ( ~n4222 & n4446 ) | ( n4445 & n4446 ) ;
  assign n4449 = ( n4222 & ~n4447 ) | ( n4222 & n4448 ) | ( ~n4447 & n4448 ) ;
  assign n4450 = ( x79 & n4444 ) | ( x79 & ~n4449 ) | ( n4444 & ~n4449 ) ;
  assign n4451 = ( x79 & n4223 ) | ( x79 & ~n4361 ) | ( n4223 & ~n4361 ) ;
  assign n4452 = x79 & n4223 ;
  assign n4453 = ( ~n4228 & n4451 ) | ( ~n4228 & n4452 ) | ( n4451 & n4452 ) ;
  assign n4454 = ( n4228 & n4451 ) | ( n4228 & n4452 ) | ( n4451 & n4452 ) ;
  assign n4455 = ( n4228 & n4453 ) | ( n4228 & ~n4454 ) | ( n4453 & ~n4454 ) ;
  assign n4456 = ( x80 & n4450 ) | ( x80 & ~n4455 ) | ( n4450 & ~n4455 ) ;
  assign n4457 = ( x80 & n4229 ) | ( x80 & ~n4361 ) | ( n4229 & ~n4361 ) ;
  assign n4458 = x80 & n4229 ;
  assign n4459 = ( n4234 & n4457 ) | ( n4234 & n4458 ) | ( n4457 & n4458 ) ;
  assign n4460 = ( ~n4234 & n4457 ) | ( ~n4234 & n4458 ) | ( n4457 & n4458 ) ;
  assign n4461 = ( n4234 & ~n4459 ) | ( n4234 & n4460 ) | ( ~n4459 & n4460 ) ;
  assign n4462 = ( x81 & n4456 ) | ( x81 & ~n4461 ) | ( n4456 & ~n4461 ) ;
  assign n4463 = ( x81 & n4235 ) | ( x81 & ~n4361 ) | ( n4235 & ~n4361 ) ;
  assign n4464 = x81 & n4235 ;
  assign n4465 = ( ~n4240 & n4463 ) | ( ~n4240 & n4464 ) | ( n4463 & n4464 ) ;
  assign n4466 = ( n4240 & n4463 ) | ( n4240 & n4464 ) | ( n4463 & n4464 ) ;
  assign n4467 = ( n4240 & n4465 ) | ( n4240 & ~n4466 ) | ( n4465 & ~n4466 ) ;
  assign n4468 = ( x82 & n4462 ) | ( x82 & ~n4467 ) | ( n4462 & ~n4467 ) ;
  assign n4469 = ( x82 & n4241 ) | ( x82 & ~n4361 ) | ( n4241 & ~n4361 ) ;
  assign n4470 = x82 & n4241 ;
  assign n4471 = ( n4246 & n4469 ) | ( n4246 & n4470 ) | ( n4469 & n4470 ) ;
  assign n4472 = ( ~n4246 & n4469 ) | ( ~n4246 & n4470 ) | ( n4469 & n4470 ) ;
  assign n4473 = ( n4246 & ~n4471 ) | ( n4246 & n4472 ) | ( ~n4471 & n4472 ) ;
  assign n4474 = ( x83 & n4468 ) | ( x83 & ~n4473 ) | ( n4468 & ~n4473 ) ;
  assign n4475 = ( x83 & n4247 ) | ( x83 & ~n4361 ) | ( n4247 & ~n4361 ) ;
  assign n4476 = x83 & n4247 ;
  assign n4477 = ( ~n4252 & n4475 ) | ( ~n4252 & n4476 ) | ( n4475 & n4476 ) ;
  assign n4478 = ( n4252 & n4475 ) | ( n4252 & n4476 ) | ( n4475 & n4476 ) ;
  assign n4479 = ( n4252 & n4477 ) | ( n4252 & ~n4478 ) | ( n4477 & ~n4478 ) ;
  assign n4480 = ( x84 & n4474 ) | ( x84 & ~n4479 ) | ( n4474 & ~n4479 ) ;
  assign n4481 = ( x84 & n4253 ) | ( x84 & ~n4361 ) | ( n4253 & ~n4361 ) ;
  assign n4482 = x84 & n4253 ;
  assign n4483 = ( n4258 & n4481 ) | ( n4258 & n4482 ) | ( n4481 & n4482 ) ;
  assign n4484 = ( ~n4258 & n4481 ) | ( ~n4258 & n4482 ) | ( n4481 & n4482 ) ;
  assign n4485 = ( n4258 & ~n4483 ) | ( n4258 & n4484 ) | ( ~n4483 & n4484 ) ;
  assign n4486 = ( x85 & n4480 ) | ( x85 & ~n4485 ) | ( n4480 & ~n4485 ) ;
  assign n4487 = ( x85 & n4259 ) | ( x85 & ~n4361 ) | ( n4259 & ~n4361 ) ;
  assign n4488 = x85 & n4259 ;
  assign n4489 = ( ~n4264 & n4487 ) | ( ~n4264 & n4488 ) | ( n4487 & n4488 ) ;
  assign n4490 = ( n4264 & n4487 ) | ( n4264 & n4488 ) | ( n4487 & n4488 ) ;
  assign n4491 = ( n4264 & n4489 ) | ( n4264 & ~n4490 ) | ( n4489 & ~n4490 ) ;
  assign n4492 = ( x86 & n4486 ) | ( x86 & ~n4491 ) | ( n4486 & ~n4491 ) ;
  assign n4493 = ( x86 & n4265 ) | ( x86 & ~n4361 ) | ( n4265 & ~n4361 ) ;
  assign n4494 = x86 & n4265 ;
  assign n4495 = ( n4270 & n4493 ) | ( n4270 & n4494 ) | ( n4493 & n4494 ) ;
  assign n4496 = ( ~n4270 & n4493 ) | ( ~n4270 & n4494 ) | ( n4493 & n4494 ) ;
  assign n4497 = ( n4270 & ~n4495 ) | ( n4270 & n4496 ) | ( ~n4495 & n4496 ) ;
  assign n4498 = ( x87 & n4492 ) | ( x87 & ~n4497 ) | ( n4492 & ~n4497 ) ;
  assign n4499 = ( x87 & n4271 ) | ( x87 & ~n4361 ) | ( n4271 & ~n4361 ) ;
  assign n4500 = x87 & n4271 ;
  assign n4501 = ( ~n4276 & n4499 ) | ( ~n4276 & n4500 ) | ( n4499 & n4500 ) ;
  assign n4502 = ( n4276 & n4499 ) | ( n4276 & n4500 ) | ( n4499 & n4500 ) ;
  assign n4503 = ( n4276 & n4501 ) | ( n4276 & ~n4502 ) | ( n4501 & ~n4502 ) ;
  assign n4504 = ( x88 & n4498 ) | ( x88 & ~n4503 ) | ( n4498 & ~n4503 ) ;
  assign n4505 = ( x88 & n4277 ) | ( x88 & ~n4361 ) | ( n4277 & ~n4361 ) ;
  assign n4506 = x88 & n4277 ;
  assign n4507 = ( n4282 & n4505 ) | ( n4282 & n4506 ) | ( n4505 & n4506 ) ;
  assign n4508 = ( ~n4282 & n4505 ) | ( ~n4282 & n4506 ) | ( n4505 & n4506 ) ;
  assign n4509 = ( n4282 & ~n4507 ) | ( n4282 & n4508 ) | ( ~n4507 & n4508 ) ;
  assign n4510 = ( x89 & n4504 ) | ( x89 & ~n4509 ) | ( n4504 & ~n4509 ) ;
  assign n4511 = ( x89 & n4283 ) | ( x89 & ~n4361 ) | ( n4283 & ~n4361 ) ;
  assign n4512 = x89 & n4283 ;
  assign n4513 = ( ~n4288 & n4511 ) | ( ~n4288 & n4512 ) | ( n4511 & n4512 ) ;
  assign n4514 = ( n4288 & n4511 ) | ( n4288 & n4512 ) | ( n4511 & n4512 ) ;
  assign n4515 = ( n4288 & n4513 ) | ( n4288 & ~n4514 ) | ( n4513 & ~n4514 ) ;
  assign n4516 = ( x90 & n4510 ) | ( x90 & ~n4515 ) | ( n4510 & ~n4515 ) ;
  assign n4517 = ( x90 & n4289 ) | ( x90 & ~n4361 ) | ( n4289 & ~n4361 ) ;
  assign n4518 = x90 & n4289 ;
  assign n4519 = ( n4294 & n4517 ) | ( n4294 & n4518 ) | ( n4517 & n4518 ) ;
  assign n4520 = ( ~n4294 & n4517 ) | ( ~n4294 & n4518 ) | ( n4517 & n4518 ) ;
  assign n4521 = ( n4294 & ~n4519 ) | ( n4294 & n4520 ) | ( ~n4519 & n4520 ) ;
  assign n4522 = ( x91 & n4516 ) | ( x91 & ~n4521 ) | ( n4516 & ~n4521 ) ;
  assign n4523 = ( x91 & n4295 ) | ( x91 & ~n4361 ) | ( n4295 & ~n4361 ) ;
  assign n4524 = x91 & n4295 ;
  assign n4525 = ( ~n4300 & n4523 ) | ( ~n4300 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4526 = ( n4300 & n4523 ) | ( n4300 & n4524 ) | ( n4523 & n4524 ) ;
  assign n4527 = ( n4300 & n4525 ) | ( n4300 & ~n4526 ) | ( n4525 & ~n4526 ) ;
  assign n4528 = ( x92 & n4522 ) | ( x92 & ~n4527 ) | ( n4522 & ~n4527 ) ;
  assign n4529 = ( x92 & n4301 ) | ( x92 & ~n4361 ) | ( n4301 & ~n4361 ) ;
  assign n4530 = x92 & n4301 ;
  assign n4531 = ( n4306 & n4529 ) | ( n4306 & n4530 ) | ( n4529 & n4530 ) ;
  assign n4532 = ( ~n4306 & n4529 ) | ( ~n4306 & n4530 ) | ( n4529 & n4530 ) ;
  assign n4533 = ( n4306 & ~n4531 ) | ( n4306 & n4532 ) | ( ~n4531 & n4532 ) ;
  assign n4534 = ( x93 & n4528 ) | ( x93 & ~n4533 ) | ( n4528 & ~n4533 ) ;
  assign n4535 = ( x93 & n4307 ) | ( x93 & ~n4361 ) | ( n4307 & ~n4361 ) ;
  assign n4536 = x93 & n4307 ;
  assign n4537 = ( ~n4312 & n4535 ) | ( ~n4312 & n4536 ) | ( n4535 & n4536 ) ;
  assign n4538 = ( n4312 & n4535 ) | ( n4312 & n4536 ) | ( n4535 & n4536 ) ;
  assign n4539 = ( n4312 & n4537 ) | ( n4312 & ~n4538 ) | ( n4537 & ~n4538 ) ;
  assign n4540 = ( x94 & n4534 ) | ( x94 & ~n4539 ) | ( n4534 & ~n4539 ) ;
  assign n4541 = ( x94 & n4313 ) | ( x94 & ~n4361 ) | ( n4313 & ~n4361 ) ;
  assign n4542 = x94 & n4313 ;
  assign n4543 = ( n4318 & n4541 ) | ( n4318 & n4542 ) | ( n4541 & n4542 ) ;
  assign n4544 = ( ~n4318 & n4541 ) | ( ~n4318 & n4542 ) | ( n4541 & n4542 ) ;
  assign n4545 = ( n4318 & ~n4543 ) | ( n4318 & n4544 ) | ( ~n4543 & n4544 ) ;
  assign n4546 = ( x95 & n4540 ) | ( x95 & ~n4545 ) | ( n4540 & ~n4545 ) ;
  assign n4547 = ( x95 & n4319 ) | ( x95 & ~n4361 ) | ( n4319 & ~n4361 ) ;
  assign n4548 = x95 & n4319 ;
  assign n4549 = ( ~n4324 & n4547 ) | ( ~n4324 & n4548 ) | ( n4547 & n4548 ) ;
  assign n4550 = ( n4324 & n4547 ) | ( n4324 & n4548 ) | ( n4547 & n4548 ) ;
  assign n4551 = ( n4324 & n4549 ) | ( n4324 & ~n4550 ) | ( n4549 & ~n4550 ) ;
  assign n4552 = ( x96 & n4546 ) | ( x96 & ~n4551 ) | ( n4546 & ~n4551 ) ;
  assign n4553 = ( x96 & n4325 ) | ( x96 & ~n4361 ) | ( n4325 & ~n4361 ) ;
  assign n4554 = x96 & n4325 ;
  assign n4555 = ( n4330 & n4553 ) | ( n4330 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4556 = ( ~n4330 & n4553 ) | ( ~n4330 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4557 = ( n4330 & ~n4555 ) | ( n4330 & n4556 ) | ( ~n4555 & n4556 ) ;
  assign n4558 = ( x97 & n4552 ) | ( x97 & ~n4557 ) | ( n4552 & ~n4557 ) ;
  assign n4559 = ( x97 & n4331 ) | ( x97 & ~n4361 ) | ( n4331 & ~n4361 ) ;
  assign n4560 = x97 & n4331 ;
  assign n4561 = ( ~n4336 & n4559 ) | ( ~n4336 & n4560 ) | ( n4559 & n4560 ) ;
  assign n4562 = ( n4336 & n4559 ) | ( n4336 & n4560 ) | ( n4559 & n4560 ) ;
  assign n4563 = ( n4336 & n4561 ) | ( n4336 & ~n4562 ) | ( n4561 & ~n4562 ) ;
  assign n4564 = ( x98 & n4558 ) | ( x98 & ~n4563 ) | ( n4558 & ~n4563 ) ;
  assign n4565 = ( x98 & n4337 ) | ( x98 & ~n4361 ) | ( n4337 & ~n4361 ) ;
  assign n4566 = x98 & n4337 ;
  assign n4567 = ( n4342 & n4565 ) | ( n4342 & n4566 ) | ( n4565 & n4566 ) ;
  assign n4568 = ( ~n4342 & n4565 ) | ( ~n4342 & n4566 ) | ( n4565 & n4566 ) ;
  assign n4569 = ( n4342 & ~n4567 ) | ( n4342 & n4568 ) | ( ~n4567 & n4568 ) ;
  assign n4570 = ( x99 & n4564 ) | ( x99 & ~n4569 ) | ( n4564 & ~n4569 ) ;
  assign n4571 = ( x99 & n4343 ) | ( x99 & ~n4361 ) | ( n4343 & ~n4361 ) ;
  assign n4572 = x99 & n4343 ;
  assign n4573 = ( ~n4348 & n4571 ) | ( ~n4348 & n4572 ) | ( n4571 & n4572 ) ;
  assign n4574 = ( n4348 & n4571 ) | ( n4348 & n4572 ) | ( n4571 & n4572 ) ;
  assign n4575 = ( n4348 & n4573 ) | ( n4348 & ~n4574 ) | ( n4573 & ~n4574 ) ;
  assign n4576 = ( x100 & n4570 ) | ( x100 & ~n4575 ) | ( n4570 & ~n4575 ) ;
  assign n4577 = ( x100 & n4349 ) | ( x100 & ~n4361 ) | ( n4349 & ~n4361 ) ;
  assign n4578 = x100 & n4349 ;
  assign n4579 = ( ~n4354 & n4577 ) | ( ~n4354 & n4578 ) | ( n4577 & n4578 ) ;
  assign n4580 = ( n4354 & n4577 ) | ( n4354 & n4578 ) | ( n4577 & n4578 ) ;
  assign n4581 = ( n4354 & n4579 ) | ( n4354 & ~n4580 ) | ( n4579 & ~n4580 ) ;
  assign n4582 = ( x101 & n4576 ) | ( x101 & ~n4581 ) | ( n4576 & ~n4581 ) ;
  assign n4583 = x102 | n4582 ;
  assign n4584 = ( x102 & n155 ) | ( x102 & n4582 ) | ( n155 & n4582 ) ;
  assign n4585 = ( n4359 & ~n4583 ) | ( n4359 & n4584 ) | ( ~n4583 & n4584 ) ;
  assign n4586 = ( x102 & ~n4359 ) | ( x102 & n4582 ) | ( ~n4359 & n4582 ) ;
  assign n4587 = n155 | n4586 ;
  assign n4588 = ( x25 & ~x64 ) | ( x25 & n4587 ) | ( ~x64 & n4587 ) ;
  assign n4589 = ~x25 & n4587 ;
  assign n4590 = ( n4365 & n4588 ) | ( n4365 & ~n4589 ) | ( n4588 & ~n4589 ) ;
  assign n4591 = ~x24 & x64 ;
  assign n4592 = ( x65 & ~n4590 ) | ( x65 & n4591 ) | ( ~n4590 & n4591 ) ;
  assign n4593 = ( x65 & n4365 ) | ( x65 & ~n4587 ) | ( n4365 & ~n4587 ) ;
  assign n4594 = x65 & n4365 ;
  assign n4595 = ( n4364 & n4593 ) | ( n4364 & n4594 ) | ( n4593 & n4594 ) ;
  assign n4596 = ( ~n4364 & n4593 ) | ( ~n4364 & n4594 ) | ( n4593 & n4594 ) ;
  assign n4597 = ( n4364 & ~n4595 ) | ( n4364 & n4596 ) | ( ~n4595 & n4596 ) ;
  assign n4598 = ( x66 & n4592 ) | ( x66 & ~n4597 ) | ( n4592 & ~n4597 ) ;
  assign n4599 = ( x66 & n4366 ) | ( x66 & ~n4587 ) | ( n4366 & ~n4587 ) ;
  assign n4600 = x66 & n4366 ;
  assign n4601 = ( n4371 & n4599 ) | ( n4371 & n4600 ) | ( n4599 & n4600 ) ;
  assign n4602 = ( ~n4371 & n4599 ) | ( ~n4371 & n4600 ) | ( n4599 & n4600 ) ;
  assign n4603 = ( n4371 & ~n4601 ) | ( n4371 & n4602 ) | ( ~n4601 & n4602 ) ;
  assign n4604 = ( x67 & n4598 ) | ( x67 & ~n4603 ) | ( n4598 & ~n4603 ) ;
  assign n4605 = ( x67 & n4372 ) | ( x67 & ~n4587 ) | ( n4372 & ~n4587 ) ;
  assign n4606 = x67 & n4372 ;
  assign n4607 = ( ~n4377 & n4605 ) | ( ~n4377 & n4606 ) | ( n4605 & n4606 ) ;
  assign n4608 = ( n4377 & n4605 ) | ( n4377 & n4606 ) | ( n4605 & n4606 ) ;
  assign n4609 = ( n4377 & n4607 ) | ( n4377 & ~n4608 ) | ( n4607 & ~n4608 ) ;
  assign n4610 = ( x68 & n4604 ) | ( x68 & ~n4609 ) | ( n4604 & ~n4609 ) ;
  assign n4611 = ( x68 & n4378 ) | ( x68 & ~n4587 ) | ( n4378 & ~n4587 ) ;
  assign n4612 = x68 & n4378 ;
  assign n4613 = ( n4383 & n4611 ) | ( n4383 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4614 = ( ~n4383 & n4611 ) | ( ~n4383 & n4612 ) | ( n4611 & n4612 ) ;
  assign n4615 = ( n4383 & ~n4613 ) | ( n4383 & n4614 ) | ( ~n4613 & n4614 ) ;
  assign n4616 = ( x69 & n4610 ) | ( x69 & ~n4615 ) | ( n4610 & ~n4615 ) ;
  assign n4617 = ( x69 & n4384 ) | ( x69 & ~n4587 ) | ( n4384 & ~n4587 ) ;
  assign n4618 = x69 & n4384 ;
  assign n4619 = ( ~n4389 & n4617 ) | ( ~n4389 & n4618 ) | ( n4617 & n4618 ) ;
  assign n4620 = ( n4389 & n4617 ) | ( n4389 & n4618 ) | ( n4617 & n4618 ) ;
  assign n4621 = ( n4389 & n4619 ) | ( n4389 & ~n4620 ) | ( n4619 & ~n4620 ) ;
  assign n4622 = ( x70 & n4616 ) | ( x70 & ~n4621 ) | ( n4616 & ~n4621 ) ;
  assign n4623 = ( x70 & n4390 ) | ( x70 & ~n4587 ) | ( n4390 & ~n4587 ) ;
  assign n4624 = x70 & n4390 ;
  assign n4625 = ( n4395 & n4623 ) | ( n4395 & n4624 ) | ( n4623 & n4624 ) ;
  assign n4626 = ( ~n4395 & n4623 ) | ( ~n4395 & n4624 ) | ( n4623 & n4624 ) ;
  assign n4627 = ( n4395 & ~n4625 ) | ( n4395 & n4626 ) | ( ~n4625 & n4626 ) ;
  assign n4628 = ( x71 & n4622 ) | ( x71 & ~n4627 ) | ( n4622 & ~n4627 ) ;
  assign n4629 = ( x71 & n4396 ) | ( x71 & ~n4587 ) | ( n4396 & ~n4587 ) ;
  assign n4630 = x71 & n4396 ;
  assign n4631 = ( ~n4401 & n4629 ) | ( ~n4401 & n4630 ) | ( n4629 & n4630 ) ;
  assign n4632 = ( n4401 & n4629 ) | ( n4401 & n4630 ) | ( n4629 & n4630 ) ;
  assign n4633 = ( n4401 & n4631 ) | ( n4401 & ~n4632 ) | ( n4631 & ~n4632 ) ;
  assign n4634 = ( x72 & n4628 ) | ( x72 & ~n4633 ) | ( n4628 & ~n4633 ) ;
  assign n4635 = ( x72 & n4402 ) | ( x72 & ~n4587 ) | ( n4402 & ~n4587 ) ;
  assign n4636 = x72 & n4402 ;
  assign n4637 = ( n4407 & n4635 ) | ( n4407 & n4636 ) | ( n4635 & n4636 ) ;
  assign n4638 = ( ~n4407 & n4635 ) | ( ~n4407 & n4636 ) | ( n4635 & n4636 ) ;
  assign n4639 = ( n4407 & ~n4637 ) | ( n4407 & n4638 ) | ( ~n4637 & n4638 ) ;
  assign n4640 = ( x73 & n4634 ) | ( x73 & ~n4639 ) | ( n4634 & ~n4639 ) ;
  assign n4641 = ( x73 & n4408 ) | ( x73 & ~n4587 ) | ( n4408 & ~n4587 ) ;
  assign n4642 = x73 & n4408 ;
  assign n4643 = ( ~n4413 & n4641 ) | ( ~n4413 & n4642 ) | ( n4641 & n4642 ) ;
  assign n4644 = ( n4413 & n4641 ) | ( n4413 & n4642 ) | ( n4641 & n4642 ) ;
  assign n4645 = ( n4413 & n4643 ) | ( n4413 & ~n4644 ) | ( n4643 & ~n4644 ) ;
  assign n4646 = ( x74 & n4640 ) | ( x74 & ~n4645 ) | ( n4640 & ~n4645 ) ;
  assign n4647 = ( x74 & n4414 ) | ( x74 & ~n4587 ) | ( n4414 & ~n4587 ) ;
  assign n4648 = x74 & n4414 ;
  assign n4649 = ( n4419 & n4647 ) | ( n4419 & n4648 ) | ( n4647 & n4648 ) ;
  assign n4650 = ( ~n4419 & n4647 ) | ( ~n4419 & n4648 ) | ( n4647 & n4648 ) ;
  assign n4651 = ( n4419 & ~n4649 ) | ( n4419 & n4650 ) | ( ~n4649 & n4650 ) ;
  assign n4652 = ( x75 & n4646 ) | ( x75 & ~n4651 ) | ( n4646 & ~n4651 ) ;
  assign n4653 = ( x75 & n4420 ) | ( x75 & ~n4587 ) | ( n4420 & ~n4587 ) ;
  assign n4654 = x75 & n4420 ;
  assign n4655 = ( ~n4425 & n4653 ) | ( ~n4425 & n4654 ) | ( n4653 & n4654 ) ;
  assign n4656 = ( n4425 & n4653 ) | ( n4425 & n4654 ) | ( n4653 & n4654 ) ;
  assign n4657 = ( n4425 & n4655 ) | ( n4425 & ~n4656 ) | ( n4655 & ~n4656 ) ;
  assign n4658 = ( x76 & n4652 ) | ( x76 & ~n4657 ) | ( n4652 & ~n4657 ) ;
  assign n4659 = ( x76 & n4426 ) | ( x76 & ~n4587 ) | ( n4426 & ~n4587 ) ;
  assign n4660 = x76 & n4426 ;
  assign n4661 = ( n4431 & n4659 ) | ( n4431 & n4660 ) | ( n4659 & n4660 ) ;
  assign n4662 = ( ~n4431 & n4659 ) | ( ~n4431 & n4660 ) | ( n4659 & n4660 ) ;
  assign n4663 = ( n4431 & ~n4661 ) | ( n4431 & n4662 ) | ( ~n4661 & n4662 ) ;
  assign n4664 = ( x77 & n4658 ) | ( x77 & ~n4663 ) | ( n4658 & ~n4663 ) ;
  assign n4665 = ( x77 & n4432 ) | ( x77 & ~n4587 ) | ( n4432 & ~n4587 ) ;
  assign n4666 = x77 & n4432 ;
  assign n4667 = ( ~n4437 & n4665 ) | ( ~n4437 & n4666 ) | ( n4665 & n4666 ) ;
  assign n4668 = ( n4437 & n4665 ) | ( n4437 & n4666 ) | ( n4665 & n4666 ) ;
  assign n4669 = ( n4437 & n4667 ) | ( n4437 & ~n4668 ) | ( n4667 & ~n4668 ) ;
  assign n4670 = ( x78 & n4664 ) | ( x78 & ~n4669 ) | ( n4664 & ~n4669 ) ;
  assign n4671 = ( x78 & n4438 ) | ( x78 & ~n4587 ) | ( n4438 & ~n4587 ) ;
  assign n4672 = x78 & n4438 ;
  assign n4673 = ( n4443 & n4671 ) | ( n4443 & n4672 ) | ( n4671 & n4672 ) ;
  assign n4674 = ( ~n4443 & n4671 ) | ( ~n4443 & n4672 ) | ( n4671 & n4672 ) ;
  assign n4675 = ( n4443 & ~n4673 ) | ( n4443 & n4674 ) | ( ~n4673 & n4674 ) ;
  assign n4676 = ( x79 & n4670 ) | ( x79 & ~n4675 ) | ( n4670 & ~n4675 ) ;
  assign n4677 = ( x79 & n4444 ) | ( x79 & ~n4587 ) | ( n4444 & ~n4587 ) ;
  assign n4678 = x79 & n4444 ;
  assign n4679 = ( ~n4449 & n4677 ) | ( ~n4449 & n4678 ) | ( n4677 & n4678 ) ;
  assign n4680 = ( n4449 & n4677 ) | ( n4449 & n4678 ) | ( n4677 & n4678 ) ;
  assign n4681 = ( n4449 & n4679 ) | ( n4449 & ~n4680 ) | ( n4679 & ~n4680 ) ;
  assign n4682 = ( x80 & n4676 ) | ( x80 & ~n4681 ) | ( n4676 & ~n4681 ) ;
  assign n4683 = ( x80 & n4450 ) | ( x80 & ~n4587 ) | ( n4450 & ~n4587 ) ;
  assign n4684 = x80 & n4450 ;
  assign n4685 = ( n4455 & n4683 ) | ( n4455 & n4684 ) | ( n4683 & n4684 ) ;
  assign n4686 = ( ~n4455 & n4683 ) | ( ~n4455 & n4684 ) | ( n4683 & n4684 ) ;
  assign n4687 = ( n4455 & ~n4685 ) | ( n4455 & n4686 ) | ( ~n4685 & n4686 ) ;
  assign n4688 = ( x81 & n4682 ) | ( x81 & ~n4687 ) | ( n4682 & ~n4687 ) ;
  assign n4689 = ( x81 & n4456 ) | ( x81 & ~n4587 ) | ( n4456 & ~n4587 ) ;
  assign n4690 = x81 & n4456 ;
  assign n4691 = ( ~n4461 & n4689 ) | ( ~n4461 & n4690 ) | ( n4689 & n4690 ) ;
  assign n4692 = ( n4461 & n4689 ) | ( n4461 & n4690 ) | ( n4689 & n4690 ) ;
  assign n4693 = ( n4461 & n4691 ) | ( n4461 & ~n4692 ) | ( n4691 & ~n4692 ) ;
  assign n4694 = ( x82 & n4688 ) | ( x82 & ~n4693 ) | ( n4688 & ~n4693 ) ;
  assign n4695 = ( x82 & n4462 ) | ( x82 & ~n4587 ) | ( n4462 & ~n4587 ) ;
  assign n4696 = x82 & n4462 ;
  assign n4697 = ( n4467 & n4695 ) | ( n4467 & n4696 ) | ( n4695 & n4696 ) ;
  assign n4698 = ( ~n4467 & n4695 ) | ( ~n4467 & n4696 ) | ( n4695 & n4696 ) ;
  assign n4699 = ( n4467 & ~n4697 ) | ( n4467 & n4698 ) | ( ~n4697 & n4698 ) ;
  assign n4700 = ( x83 & n4694 ) | ( x83 & ~n4699 ) | ( n4694 & ~n4699 ) ;
  assign n4701 = ( x83 & n4468 ) | ( x83 & ~n4587 ) | ( n4468 & ~n4587 ) ;
  assign n4702 = x83 & n4468 ;
  assign n4703 = ( ~n4473 & n4701 ) | ( ~n4473 & n4702 ) | ( n4701 & n4702 ) ;
  assign n4704 = ( n4473 & n4701 ) | ( n4473 & n4702 ) | ( n4701 & n4702 ) ;
  assign n4705 = ( n4473 & n4703 ) | ( n4473 & ~n4704 ) | ( n4703 & ~n4704 ) ;
  assign n4706 = ( x84 & n4700 ) | ( x84 & ~n4705 ) | ( n4700 & ~n4705 ) ;
  assign n4707 = ( x84 & n4474 ) | ( x84 & ~n4587 ) | ( n4474 & ~n4587 ) ;
  assign n4708 = x84 & n4474 ;
  assign n4709 = ( n4479 & n4707 ) | ( n4479 & n4708 ) | ( n4707 & n4708 ) ;
  assign n4710 = ( ~n4479 & n4707 ) | ( ~n4479 & n4708 ) | ( n4707 & n4708 ) ;
  assign n4711 = ( n4479 & ~n4709 ) | ( n4479 & n4710 ) | ( ~n4709 & n4710 ) ;
  assign n4712 = ( x85 & n4706 ) | ( x85 & ~n4711 ) | ( n4706 & ~n4711 ) ;
  assign n4713 = ( x85 & n4480 ) | ( x85 & ~n4587 ) | ( n4480 & ~n4587 ) ;
  assign n4714 = x85 & n4480 ;
  assign n4715 = ( ~n4485 & n4713 ) | ( ~n4485 & n4714 ) | ( n4713 & n4714 ) ;
  assign n4716 = ( n4485 & n4713 ) | ( n4485 & n4714 ) | ( n4713 & n4714 ) ;
  assign n4717 = ( n4485 & n4715 ) | ( n4485 & ~n4716 ) | ( n4715 & ~n4716 ) ;
  assign n4718 = ( x86 & n4712 ) | ( x86 & ~n4717 ) | ( n4712 & ~n4717 ) ;
  assign n4719 = ( x86 & n4486 ) | ( x86 & ~n4587 ) | ( n4486 & ~n4587 ) ;
  assign n4720 = x86 & n4486 ;
  assign n4721 = ( n4491 & n4719 ) | ( n4491 & n4720 ) | ( n4719 & n4720 ) ;
  assign n4722 = ( ~n4491 & n4719 ) | ( ~n4491 & n4720 ) | ( n4719 & n4720 ) ;
  assign n4723 = ( n4491 & ~n4721 ) | ( n4491 & n4722 ) | ( ~n4721 & n4722 ) ;
  assign n4724 = ( x87 & n4718 ) | ( x87 & ~n4723 ) | ( n4718 & ~n4723 ) ;
  assign n4725 = ( x87 & n4492 ) | ( x87 & ~n4587 ) | ( n4492 & ~n4587 ) ;
  assign n4726 = x87 & n4492 ;
  assign n4727 = ( ~n4497 & n4725 ) | ( ~n4497 & n4726 ) | ( n4725 & n4726 ) ;
  assign n4728 = ( n4497 & n4725 ) | ( n4497 & n4726 ) | ( n4725 & n4726 ) ;
  assign n4729 = ( n4497 & n4727 ) | ( n4497 & ~n4728 ) | ( n4727 & ~n4728 ) ;
  assign n4730 = ( x88 & n4724 ) | ( x88 & ~n4729 ) | ( n4724 & ~n4729 ) ;
  assign n4731 = ( x88 & n4498 ) | ( x88 & ~n4587 ) | ( n4498 & ~n4587 ) ;
  assign n4732 = x88 & n4498 ;
  assign n4733 = ( n4503 & n4731 ) | ( n4503 & n4732 ) | ( n4731 & n4732 ) ;
  assign n4734 = ( ~n4503 & n4731 ) | ( ~n4503 & n4732 ) | ( n4731 & n4732 ) ;
  assign n4735 = ( n4503 & ~n4733 ) | ( n4503 & n4734 ) | ( ~n4733 & n4734 ) ;
  assign n4736 = ( x89 & n4730 ) | ( x89 & ~n4735 ) | ( n4730 & ~n4735 ) ;
  assign n4737 = ( x89 & n4504 ) | ( x89 & ~n4587 ) | ( n4504 & ~n4587 ) ;
  assign n4738 = x89 & n4504 ;
  assign n4739 = ( ~n4509 & n4737 ) | ( ~n4509 & n4738 ) | ( n4737 & n4738 ) ;
  assign n4740 = ( n4509 & n4737 ) | ( n4509 & n4738 ) | ( n4737 & n4738 ) ;
  assign n4741 = ( n4509 & n4739 ) | ( n4509 & ~n4740 ) | ( n4739 & ~n4740 ) ;
  assign n4742 = ( x90 & n4736 ) | ( x90 & ~n4741 ) | ( n4736 & ~n4741 ) ;
  assign n4743 = ( x90 & n4510 ) | ( x90 & ~n4587 ) | ( n4510 & ~n4587 ) ;
  assign n4744 = x90 & n4510 ;
  assign n4745 = ( n4515 & n4743 ) | ( n4515 & n4744 ) | ( n4743 & n4744 ) ;
  assign n4746 = ( ~n4515 & n4743 ) | ( ~n4515 & n4744 ) | ( n4743 & n4744 ) ;
  assign n4747 = ( n4515 & ~n4745 ) | ( n4515 & n4746 ) | ( ~n4745 & n4746 ) ;
  assign n4748 = ( x91 & n4742 ) | ( x91 & ~n4747 ) | ( n4742 & ~n4747 ) ;
  assign n4749 = ( x91 & n4516 ) | ( x91 & ~n4587 ) | ( n4516 & ~n4587 ) ;
  assign n4750 = x91 & n4516 ;
  assign n4751 = ( ~n4521 & n4749 ) | ( ~n4521 & n4750 ) | ( n4749 & n4750 ) ;
  assign n4752 = ( n4521 & n4749 ) | ( n4521 & n4750 ) | ( n4749 & n4750 ) ;
  assign n4753 = ( n4521 & n4751 ) | ( n4521 & ~n4752 ) | ( n4751 & ~n4752 ) ;
  assign n4754 = ( x92 & n4748 ) | ( x92 & ~n4753 ) | ( n4748 & ~n4753 ) ;
  assign n4755 = ( x92 & n4522 ) | ( x92 & ~n4587 ) | ( n4522 & ~n4587 ) ;
  assign n4756 = x92 & n4522 ;
  assign n4757 = ( n4527 & n4755 ) | ( n4527 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4758 = ( ~n4527 & n4755 ) | ( ~n4527 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4759 = ( n4527 & ~n4757 ) | ( n4527 & n4758 ) | ( ~n4757 & n4758 ) ;
  assign n4760 = ( x93 & n4754 ) | ( x93 & ~n4759 ) | ( n4754 & ~n4759 ) ;
  assign n4761 = ( x93 & n4528 ) | ( x93 & ~n4587 ) | ( n4528 & ~n4587 ) ;
  assign n4762 = x93 & n4528 ;
  assign n4763 = ( ~n4533 & n4761 ) | ( ~n4533 & n4762 ) | ( n4761 & n4762 ) ;
  assign n4764 = ( n4533 & n4761 ) | ( n4533 & n4762 ) | ( n4761 & n4762 ) ;
  assign n4765 = ( n4533 & n4763 ) | ( n4533 & ~n4764 ) | ( n4763 & ~n4764 ) ;
  assign n4766 = ( x94 & n4760 ) | ( x94 & ~n4765 ) | ( n4760 & ~n4765 ) ;
  assign n4767 = ( x94 & n4534 ) | ( x94 & ~n4587 ) | ( n4534 & ~n4587 ) ;
  assign n4768 = x94 & n4534 ;
  assign n4769 = ( n4539 & n4767 ) | ( n4539 & n4768 ) | ( n4767 & n4768 ) ;
  assign n4770 = ( ~n4539 & n4767 ) | ( ~n4539 & n4768 ) | ( n4767 & n4768 ) ;
  assign n4771 = ( n4539 & ~n4769 ) | ( n4539 & n4770 ) | ( ~n4769 & n4770 ) ;
  assign n4772 = ( x95 & n4766 ) | ( x95 & ~n4771 ) | ( n4766 & ~n4771 ) ;
  assign n4773 = ( x95 & n4540 ) | ( x95 & ~n4587 ) | ( n4540 & ~n4587 ) ;
  assign n4774 = x95 & n4540 ;
  assign n4775 = ( ~n4545 & n4773 ) | ( ~n4545 & n4774 ) | ( n4773 & n4774 ) ;
  assign n4776 = ( n4545 & n4773 ) | ( n4545 & n4774 ) | ( n4773 & n4774 ) ;
  assign n4777 = ( n4545 & n4775 ) | ( n4545 & ~n4776 ) | ( n4775 & ~n4776 ) ;
  assign n4778 = ( x96 & n4772 ) | ( x96 & ~n4777 ) | ( n4772 & ~n4777 ) ;
  assign n4779 = ( x96 & n4546 ) | ( x96 & ~n4587 ) | ( n4546 & ~n4587 ) ;
  assign n4780 = x96 & n4546 ;
  assign n4781 = ( n4551 & n4779 ) | ( n4551 & n4780 ) | ( n4779 & n4780 ) ;
  assign n4782 = ( ~n4551 & n4779 ) | ( ~n4551 & n4780 ) | ( n4779 & n4780 ) ;
  assign n4783 = ( n4551 & ~n4781 ) | ( n4551 & n4782 ) | ( ~n4781 & n4782 ) ;
  assign n4784 = ( x97 & n4778 ) | ( x97 & ~n4783 ) | ( n4778 & ~n4783 ) ;
  assign n4785 = ( x97 & n4552 ) | ( x97 & ~n4587 ) | ( n4552 & ~n4587 ) ;
  assign n4786 = x97 & n4552 ;
  assign n4787 = ( ~n4557 & n4785 ) | ( ~n4557 & n4786 ) | ( n4785 & n4786 ) ;
  assign n4788 = ( n4557 & n4785 ) | ( n4557 & n4786 ) | ( n4785 & n4786 ) ;
  assign n4789 = ( n4557 & n4787 ) | ( n4557 & ~n4788 ) | ( n4787 & ~n4788 ) ;
  assign n4790 = ( x98 & n4784 ) | ( x98 & ~n4789 ) | ( n4784 & ~n4789 ) ;
  assign n4791 = ( x98 & n4558 ) | ( x98 & ~n4587 ) | ( n4558 & ~n4587 ) ;
  assign n4792 = x98 & n4558 ;
  assign n4793 = ( n4563 & n4791 ) | ( n4563 & n4792 ) | ( n4791 & n4792 ) ;
  assign n4794 = ( ~n4563 & n4791 ) | ( ~n4563 & n4792 ) | ( n4791 & n4792 ) ;
  assign n4795 = ( n4563 & ~n4793 ) | ( n4563 & n4794 ) | ( ~n4793 & n4794 ) ;
  assign n4796 = ( x99 & n4790 ) | ( x99 & ~n4795 ) | ( n4790 & ~n4795 ) ;
  assign n4797 = ( x99 & n4564 ) | ( x99 & ~n4587 ) | ( n4564 & ~n4587 ) ;
  assign n4798 = x99 & n4564 ;
  assign n4799 = ( ~n4569 & n4797 ) | ( ~n4569 & n4798 ) | ( n4797 & n4798 ) ;
  assign n4800 = ( n4569 & n4797 ) | ( n4569 & n4798 ) | ( n4797 & n4798 ) ;
  assign n4801 = ( n4569 & n4799 ) | ( n4569 & ~n4800 ) | ( n4799 & ~n4800 ) ;
  assign n4802 = ( x100 & n4796 ) | ( x100 & ~n4801 ) | ( n4796 & ~n4801 ) ;
  assign n4803 = ( x100 & n4570 ) | ( x100 & ~n4587 ) | ( n4570 & ~n4587 ) ;
  assign n4804 = x100 & n4570 ;
  assign n4805 = ( n4575 & n4803 ) | ( n4575 & n4804 ) | ( n4803 & n4804 ) ;
  assign n4806 = ( ~n4575 & n4803 ) | ( ~n4575 & n4804 ) | ( n4803 & n4804 ) ;
  assign n4807 = ( n4575 & ~n4805 ) | ( n4575 & n4806 ) | ( ~n4805 & n4806 ) ;
  assign n4808 = ( x101 & n4802 ) | ( x101 & ~n4807 ) | ( n4802 & ~n4807 ) ;
  assign n4809 = ( x101 & n4576 ) | ( x101 & ~n4587 ) | ( n4576 & ~n4587 ) ;
  assign n4810 = x101 & n4576 ;
  assign n4811 = ( n4581 & n4809 ) | ( n4581 & n4810 ) | ( n4809 & n4810 ) ;
  assign n4812 = ( ~n4581 & n4809 ) | ( ~n4581 & n4810 ) | ( n4809 & n4810 ) ;
  assign n4813 = ( n4581 & ~n4811 ) | ( n4581 & n4812 ) | ( ~n4811 & n4812 ) ;
  assign n4814 = ( x102 & n4808 ) | ( x102 & ~n4813 ) | ( n4808 & ~n4813 ) ;
  assign n4815 = x103 | n4814 ;
  assign n4816 = ( x103 & n154 ) | ( x103 & n4814 ) | ( n154 & n4814 ) ;
  assign n4817 = ( n4585 & ~n4815 ) | ( n4585 & n4816 ) | ( ~n4815 & n4816 ) ;
  assign n4818 = ( x103 & ~n4585 ) | ( x103 & n4814 ) | ( ~n4585 & n4814 ) ;
  assign n4819 = n154 | n4818 ;
  assign n4820 = ( x24 & ~x64 ) | ( x24 & n4819 ) | ( ~x64 & n4819 ) ;
  assign n4821 = ~x24 & n4819 ;
  assign n4822 = ( n4591 & n4820 ) | ( n4591 & ~n4821 ) | ( n4820 & ~n4821 ) ;
  assign n4823 = ~x23 & x64 ;
  assign n4824 = ( x65 & ~n4822 ) | ( x65 & n4823 ) | ( ~n4822 & n4823 ) ;
  assign n4825 = ( x65 & n4591 ) | ( x65 & ~n4819 ) | ( n4591 & ~n4819 ) ;
  assign n4826 = x65 & n4591 ;
  assign n4827 = ( n4590 & n4825 ) | ( n4590 & n4826 ) | ( n4825 & n4826 ) ;
  assign n4828 = ( ~n4590 & n4825 ) | ( ~n4590 & n4826 ) | ( n4825 & n4826 ) ;
  assign n4829 = ( n4590 & ~n4827 ) | ( n4590 & n4828 ) | ( ~n4827 & n4828 ) ;
  assign n4830 = ( x66 & n4824 ) | ( x66 & ~n4829 ) | ( n4824 & ~n4829 ) ;
  assign n4831 = ( x66 & n4592 ) | ( x66 & ~n4819 ) | ( n4592 & ~n4819 ) ;
  assign n4832 = x66 & n4592 ;
  assign n4833 = ( n4597 & n4831 ) | ( n4597 & n4832 ) | ( n4831 & n4832 ) ;
  assign n4834 = ( ~n4597 & n4831 ) | ( ~n4597 & n4832 ) | ( n4831 & n4832 ) ;
  assign n4835 = ( n4597 & ~n4833 ) | ( n4597 & n4834 ) | ( ~n4833 & n4834 ) ;
  assign n4836 = ( x67 & n4830 ) | ( x67 & ~n4835 ) | ( n4830 & ~n4835 ) ;
  assign n4837 = ( x67 & n4598 ) | ( x67 & ~n4819 ) | ( n4598 & ~n4819 ) ;
  assign n4838 = x67 & n4598 ;
  assign n4839 = ( ~n4603 & n4837 ) | ( ~n4603 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4840 = ( n4603 & n4837 ) | ( n4603 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4841 = ( n4603 & n4839 ) | ( n4603 & ~n4840 ) | ( n4839 & ~n4840 ) ;
  assign n4842 = ( x68 & n4836 ) | ( x68 & ~n4841 ) | ( n4836 & ~n4841 ) ;
  assign n4843 = ( x68 & n4604 ) | ( x68 & ~n4819 ) | ( n4604 & ~n4819 ) ;
  assign n4844 = x68 & n4604 ;
  assign n4845 = ( n4609 & n4843 ) | ( n4609 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4846 = ( ~n4609 & n4843 ) | ( ~n4609 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4847 = ( n4609 & ~n4845 ) | ( n4609 & n4846 ) | ( ~n4845 & n4846 ) ;
  assign n4848 = ( x69 & n4842 ) | ( x69 & ~n4847 ) | ( n4842 & ~n4847 ) ;
  assign n4849 = ( x69 & n4610 ) | ( x69 & ~n4819 ) | ( n4610 & ~n4819 ) ;
  assign n4850 = x69 & n4610 ;
  assign n4851 = ( ~n4615 & n4849 ) | ( ~n4615 & n4850 ) | ( n4849 & n4850 ) ;
  assign n4852 = ( n4615 & n4849 ) | ( n4615 & n4850 ) | ( n4849 & n4850 ) ;
  assign n4853 = ( n4615 & n4851 ) | ( n4615 & ~n4852 ) | ( n4851 & ~n4852 ) ;
  assign n4854 = ( x70 & n4848 ) | ( x70 & ~n4853 ) | ( n4848 & ~n4853 ) ;
  assign n4855 = ( x70 & n4616 ) | ( x70 & ~n4819 ) | ( n4616 & ~n4819 ) ;
  assign n4856 = x70 & n4616 ;
  assign n4857 = ( n4621 & n4855 ) | ( n4621 & n4856 ) | ( n4855 & n4856 ) ;
  assign n4858 = ( ~n4621 & n4855 ) | ( ~n4621 & n4856 ) | ( n4855 & n4856 ) ;
  assign n4859 = ( n4621 & ~n4857 ) | ( n4621 & n4858 ) | ( ~n4857 & n4858 ) ;
  assign n4860 = ( x71 & n4854 ) | ( x71 & ~n4859 ) | ( n4854 & ~n4859 ) ;
  assign n4861 = ( x71 & n4622 ) | ( x71 & ~n4819 ) | ( n4622 & ~n4819 ) ;
  assign n4862 = x71 & n4622 ;
  assign n4863 = ( ~n4627 & n4861 ) | ( ~n4627 & n4862 ) | ( n4861 & n4862 ) ;
  assign n4864 = ( n4627 & n4861 ) | ( n4627 & n4862 ) | ( n4861 & n4862 ) ;
  assign n4865 = ( n4627 & n4863 ) | ( n4627 & ~n4864 ) | ( n4863 & ~n4864 ) ;
  assign n4866 = ( x72 & n4860 ) | ( x72 & ~n4865 ) | ( n4860 & ~n4865 ) ;
  assign n4867 = ( x72 & n4628 ) | ( x72 & ~n4819 ) | ( n4628 & ~n4819 ) ;
  assign n4868 = x72 & n4628 ;
  assign n4869 = ( n4633 & n4867 ) | ( n4633 & n4868 ) | ( n4867 & n4868 ) ;
  assign n4870 = ( ~n4633 & n4867 ) | ( ~n4633 & n4868 ) | ( n4867 & n4868 ) ;
  assign n4871 = ( n4633 & ~n4869 ) | ( n4633 & n4870 ) | ( ~n4869 & n4870 ) ;
  assign n4872 = ( x73 & n4866 ) | ( x73 & ~n4871 ) | ( n4866 & ~n4871 ) ;
  assign n4873 = ( x73 & n4634 ) | ( x73 & ~n4819 ) | ( n4634 & ~n4819 ) ;
  assign n4874 = x73 & n4634 ;
  assign n4875 = ( ~n4639 & n4873 ) | ( ~n4639 & n4874 ) | ( n4873 & n4874 ) ;
  assign n4876 = ( n4639 & n4873 ) | ( n4639 & n4874 ) | ( n4873 & n4874 ) ;
  assign n4877 = ( n4639 & n4875 ) | ( n4639 & ~n4876 ) | ( n4875 & ~n4876 ) ;
  assign n4878 = ( x74 & n4872 ) | ( x74 & ~n4877 ) | ( n4872 & ~n4877 ) ;
  assign n4879 = ( x74 & n4640 ) | ( x74 & ~n4819 ) | ( n4640 & ~n4819 ) ;
  assign n4880 = x74 & n4640 ;
  assign n4881 = ( n4645 & n4879 ) | ( n4645 & n4880 ) | ( n4879 & n4880 ) ;
  assign n4882 = ( ~n4645 & n4879 ) | ( ~n4645 & n4880 ) | ( n4879 & n4880 ) ;
  assign n4883 = ( n4645 & ~n4881 ) | ( n4645 & n4882 ) | ( ~n4881 & n4882 ) ;
  assign n4884 = ( x75 & n4878 ) | ( x75 & ~n4883 ) | ( n4878 & ~n4883 ) ;
  assign n4885 = ( x75 & n4646 ) | ( x75 & ~n4819 ) | ( n4646 & ~n4819 ) ;
  assign n4886 = x75 & n4646 ;
  assign n4887 = ( ~n4651 & n4885 ) | ( ~n4651 & n4886 ) | ( n4885 & n4886 ) ;
  assign n4888 = ( n4651 & n4885 ) | ( n4651 & n4886 ) | ( n4885 & n4886 ) ;
  assign n4889 = ( n4651 & n4887 ) | ( n4651 & ~n4888 ) | ( n4887 & ~n4888 ) ;
  assign n4890 = ( x76 & n4884 ) | ( x76 & ~n4889 ) | ( n4884 & ~n4889 ) ;
  assign n4891 = ( x76 & n4652 ) | ( x76 & ~n4819 ) | ( n4652 & ~n4819 ) ;
  assign n4892 = x76 & n4652 ;
  assign n4893 = ( n4657 & n4891 ) | ( n4657 & n4892 ) | ( n4891 & n4892 ) ;
  assign n4894 = ( ~n4657 & n4891 ) | ( ~n4657 & n4892 ) | ( n4891 & n4892 ) ;
  assign n4895 = ( n4657 & ~n4893 ) | ( n4657 & n4894 ) | ( ~n4893 & n4894 ) ;
  assign n4896 = ( x77 & n4890 ) | ( x77 & ~n4895 ) | ( n4890 & ~n4895 ) ;
  assign n4897 = ( x77 & n4658 ) | ( x77 & ~n4819 ) | ( n4658 & ~n4819 ) ;
  assign n4898 = x77 & n4658 ;
  assign n4899 = ( ~n4663 & n4897 ) | ( ~n4663 & n4898 ) | ( n4897 & n4898 ) ;
  assign n4900 = ( n4663 & n4897 ) | ( n4663 & n4898 ) | ( n4897 & n4898 ) ;
  assign n4901 = ( n4663 & n4899 ) | ( n4663 & ~n4900 ) | ( n4899 & ~n4900 ) ;
  assign n4902 = ( x78 & n4896 ) | ( x78 & ~n4901 ) | ( n4896 & ~n4901 ) ;
  assign n4903 = ( x78 & n4664 ) | ( x78 & ~n4819 ) | ( n4664 & ~n4819 ) ;
  assign n4904 = x78 & n4664 ;
  assign n4905 = ( n4669 & n4903 ) | ( n4669 & n4904 ) | ( n4903 & n4904 ) ;
  assign n4906 = ( ~n4669 & n4903 ) | ( ~n4669 & n4904 ) | ( n4903 & n4904 ) ;
  assign n4907 = ( n4669 & ~n4905 ) | ( n4669 & n4906 ) | ( ~n4905 & n4906 ) ;
  assign n4908 = ( x79 & n4902 ) | ( x79 & ~n4907 ) | ( n4902 & ~n4907 ) ;
  assign n4909 = ( x79 & n4670 ) | ( x79 & ~n4819 ) | ( n4670 & ~n4819 ) ;
  assign n4910 = x79 & n4670 ;
  assign n4911 = ( ~n4675 & n4909 ) | ( ~n4675 & n4910 ) | ( n4909 & n4910 ) ;
  assign n4912 = ( n4675 & n4909 ) | ( n4675 & n4910 ) | ( n4909 & n4910 ) ;
  assign n4913 = ( n4675 & n4911 ) | ( n4675 & ~n4912 ) | ( n4911 & ~n4912 ) ;
  assign n4914 = ( x80 & n4908 ) | ( x80 & ~n4913 ) | ( n4908 & ~n4913 ) ;
  assign n4915 = ( x80 & n4676 ) | ( x80 & ~n4819 ) | ( n4676 & ~n4819 ) ;
  assign n4916 = x80 & n4676 ;
  assign n4917 = ( n4681 & n4915 ) | ( n4681 & n4916 ) | ( n4915 & n4916 ) ;
  assign n4918 = ( ~n4681 & n4915 ) | ( ~n4681 & n4916 ) | ( n4915 & n4916 ) ;
  assign n4919 = ( n4681 & ~n4917 ) | ( n4681 & n4918 ) | ( ~n4917 & n4918 ) ;
  assign n4920 = ( x81 & n4914 ) | ( x81 & ~n4919 ) | ( n4914 & ~n4919 ) ;
  assign n4921 = ( x81 & n4682 ) | ( x81 & ~n4819 ) | ( n4682 & ~n4819 ) ;
  assign n4922 = x81 & n4682 ;
  assign n4923 = ( ~n4687 & n4921 ) | ( ~n4687 & n4922 ) | ( n4921 & n4922 ) ;
  assign n4924 = ( n4687 & n4921 ) | ( n4687 & n4922 ) | ( n4921 & n4922 ) ;
  assign n4925 = ( n4687 & n4923 ) | ( n4687 & ~n4924 ) | ( n4923 & ~n4924 ) ;
  assign n4926 = ( x82 & n4920 ) | ( x82 & ~n4925 ) | ( n4920 & ~n4925 ) ;
  assign n4927 = ( x82 & n4688 ) | ( x82 & ~n4819 ) | ( n4688 & ~n4819 ) ;
  assign n4928 = x82 & n4688 ;
  assign n4929 = ( n4693 & n4927 ) | ( n4693 & n4928 ) | ( n4927 & n4928 ) ;
  assign n4930 = ( ~n4693 & n4927 ) | ( ~n4693 & n4928 ) | ( n4927 & n4928 ) ;
  assign n4931 = ( n4693 & ~n4929 ) | ( n4693 & n4930 ) | ( ~n4929 & n4930 ) ;
  assign n4932 = ( x83 & n4926 ) | ( x83 & ~n4931 ) | ( n4926 & ~n4931 ) ;
  assign n4933 = ( x83 & n4694 ) | ( x83 & ~n4819 ) | ( n4694 & ~n4819 ) ;
  assign n4934 = x83 & n4694 ;
  assign n4935 = ( ~n4699 & n4933 ) | ( ~n4699 & n4934 ) | ( n4933 & n4934 ) ;
  assign n4936 = ( n4699 & n4933 ) | ( n4699 & n4934 ) | ( n4933 & n4934 ) ;
  assign n4937 = ( n4699 & n4935 ) | ( n4699 & ~n4936 ) | ( n4935 & ~n4936 ) ;
  assign n4938 = ( x84 & n4932 ) | ( x84 & ~n4937 ) | ( n4932 & ~n4937 ) ;
  assign n4939 = ( x84 & n4700 ) | ( x84 & ~n4819 ) | ( n4700 & ~n4819 ) ;
  assign n4940 = x84 & n4700 ;
  assign n4941 = ( n4705 & n4939 ) | ( n4705 & n4940 ) | ( n4939 & n4940 ) ;
  assign n4942 = ( ~n4705 & n4939 ) | ( ~n4705 & n4940 ) | ( n4939 & n4940 ) ;
  assign n4943 = ( n4705 & ~n4941 ) | ( n4705 & n4942 ) | ( ~n4941 & n4942 ) ;
  assign n4944 = ( x85 & n4938 ) | ( x85 & ~n4943 ) | ( n4938 & ~n4943 ) ;
  assign n4945 = ( x85 & n4706 ) | ( x85 & ~n4819 ) | ( n4706 & ~n4819 ) ;
  assign n4946 = x85 & n4706 ;
  assign n4947 = ( ~n4711 & n4945 ) | ( ~n4711 & n4946 ) | ( n4945 & n4946 ) ;
  assign n4948 = ( n4711 & n4945 ) | ( n4711 & n4946 ) | ( n4945 & n4946 ) ;
  assign n4949 = ( n4711 & n4947 ) | ( n4711 & ~n4948 ) | ( n4947 & ~n4948 ) ;
  assign n4950 = ( x86 & n4944 ) | ( x86 & ~n4949 ) | ( n4944 & ~n4949 ) ;
  assign n4951 = ( x86 & n4712 ) | ( x86 & ~n4819 ) | ( n4712 & ~n4819 ) ;
  assign n4952 = x86 & n4712 ;
  assign n4953 = ( n4717 & n4951 ) | ( n4717 & n4952 ) | ( n4951 & n4952 ) ;
  assign n4954 = ( ~n4717 & n4951 ) | ( ~n4717 & n4952 ) | ( n4951 & n4952 ) ;
  assign n4955 = ( n4717 & ~n4953 ) | ( n4717 & n4954 ) | ( ~n4953 & n4954 ) ;
  assign n4956 = ( x87 & n4950 ) | ( x87 & ~n4955 ) | ( n4950 & ~n4955 ) ;
  assign n4957 = ( x87 & n4718 ) | ( x87 & ~n4819 ) | ( n4718 & ~n4819 ) ;
  assign n4958 = x87 & n4718 ;
  assign n4959 = ( ~n4723 & n4957 ) | ( ~n4723 & n4958 ) | ( n4957 & n4958 ) ;
  assign n4960 = ( n4723 & n4957 ) | ( n4723 & n4958 ) | ( n4957 & n4958 ) ;
  assign n4961 = ( n4723 & n4959 ) | ( n4723 & ~n4960 ) | ( n4959 & ~n4960 ) ;
  assign n4962 = ( x88 & n4956 ) | ( x88 & ~n4961 ) | ( n4956 & ~n4961 ) ;
  assign n4963 = ( x88 & n4724 ) | ( x88 & ~n4819 ) | ( n4724 & ~n4819 ) ;
  assign n4964 = x88 & n4724 ;
  assign n4965 = ( n4729 & n4963 ) | ( n4729 & n4964 ) | ( n4963 & n4964 ) ;
  assign n4966 = ( ~n4729 & n4963 ) | ( ~n4729 & n4964 ) | ( n4963 & n4964 ) ;
  assign n4967 = ( n4729 & ~n4965 ) | ( n4729 & n4966 ) | ( ~n4965 & n4966 ) ;
  assign n4968 = ( x89 & n4962 ) | ( x89 & ~n4967 ) | ( n4962 & ~n4967 ) ;
  assign n4969 = ( x89 & n4730 ) | ( x89 & ~n4819 ) | ( n4730 & ~n4819 ) ;
  assign n4970 = x89 & n4730 ;
  assign n4971 = ( ~n4735 & n4969 ) | ( ~n4735 & n4970 ) | ( n4969 & n4970 ) ;
  assign n4972 = ( n4735 & n4969 ) | ( n4735 & n4970 ) | ( n4969 & n4970 ) ;
  assign n4973 = ( n4735 & n4971 ) | ( n4735 & ~n4972 ) | ( n4971 & ~n4972 ) ;
  assign n4974 = ( x90 & n4968 ) | ( x90 & ~n4973 ) | ( n4968 & ~n4973 ) ;
  assign n4975 = ( x90 & n4736 ) | ( x90 & ~n4819 ) | ( n4736 & ~n4819 ) ;
  assign n4976 = x90 & n4736 ;
  assign n4977 = ( n4741 & n4975 ) | ( n4741 & n4976 ) | ( n4975 & n4976 ) ;
  assign n4978 = ( ~n4741 & n4975 ) | ( ~n4741 & n4976 ) | ( n4975 & n4976 ) ;
  assign n4979 = ( n4741 & ~n4977 ) | ( n4741 & n4978 ) | ( ~n4977 & n4978 ) ;
  assign n4980 = ( x91 & n4974 ) | ( x91 & ~n4979 ) | ( n4974 & ~n4979 ) ;
  assign n4981 = ( x91 & n4742 ) | ( x91 & ~n4819 ) | ( n4742 & ~n4819 ) ;
  assign n4982 = x91 & n4742 ;
  assign n4983 = ( ~n4747 & n4981 ) | ( ~n4747 & n4982 ) | ( n4981 & n4982 ) ;
  assign n4984 = ( n4747 & n4981 ) | ( n4747 & n4982 ) | ( n4981 & n4982 ) ;
  assign n4985 = ( n4747 & n4983 ) | ( n4747 & ~n4984 ) | ( n4983 & ~n4984 ) ;
  assign n4986 = ( x92 & n4980 ) | ( x92 & ~n4985 ) | ( n4980 & ~n4985 ) ;
  assign n4987 = ( x92 & n4748 ) | ( x92 & ~n4819 ) | ( n4748 & ~n4819 ) ;
  assign n4988 = x92 & n4748 ;
  assign n4989 = ( n4753 & n4987 ) | ( n4753 & n4988 ) | ( n4987 & n4988 ) ;
  assign n4990 = ( ~n4753 & n4987 ) | ( ~n4753 & n4988 ) | ( n4987 & n4988 ) ;
  assign n4991 = ( n4753 & ~n4989 ) | ( n4753 & n4990 ) | ( ~n4989 & n4990 ) ;
  assign n4992 = ( x93 & n4986 ) | ( x93 & ~n4991 ) | ( n4986 & ~n4991 ) ;
  assign n4993 = ( x93 & n4754 ) | ( x93 & ~n4819 ) | ( n4754 & ~n4819 ) ;
  assign n4994 = x93 & n4754 ;
  assign n4995 = ( ~n4759 & n4993 ) | ( ~n4759 & n4994 ) | ( n4993 & n4994 ) ;
  assign n4996 = ( n4759 & n4993 ) | ( n4759 & n4994 ) | ( n4993 & n4994 ) ;
  assign n4997 = ( n4759 & n4995 ) | ( n4759 & ~n4996 ) | ( n4995 & ~n4996 ) ;
  assign n4998 = ( x94 & n4992 ) | ( x94 & ~n4997 ) | ( n4992 & ~n4997 ) ;
  assign n4999 = ( x94 & n4760 ) | ( x94 & ~n4819 ) | ( n4760 & ~n4819 ) ;
  assign n5000 = x94 & n4760 ;
  assign n5001 = ( n4765 & n4999 ) | ( n4765 & n5000 ) | ( n4999 & n5000 ) ;
  assign n5002 = ( ~n4765 & n4999 ) | ( ~n4765 & n5000 ) | ( n4999 & n5000 ) ;
  assign n5003 = ( n4765 & ~n5001 ) | ( n4765 & n5002 ) | ( ~n5001 & n5002 ) ;
  assign n5004 = ( x95 & n4998 ) | ( x95 & ~n5003 ) | ( n4998 & ~n5003 ) ;
  assign n5005 = ( x95 & n4766 ) | ( x95 & ~n4819 ) | ( n4766 & ~n4819 ) ;
  assign n5006 = x95 & n4766 ;
  assign n5007 = ( ~n4771 & n5005 ) | ( ~n4771 & n5006 ) | ( n5005 & n5006 ) ;
  assign n5008 = ( n4771 & n5005 ) | ( n4771 & n5006 ) | ( n5005 & n5006 ) ;
  assign n5009 = ( n4771 & n5007 ) | ( n4771 & ~n5008 ) | ( n5007 & ~n5008 ) ;
  assign n5010 = ( x96 & n5004 ) | ( x96 & ~n5009 ) | ( n5004 & ~n5009 ) ;
  assign n5011 = ( x96 & n4772 ) | ( x96 & ~n4819 ) | ( n4772 & ~n4819 ) ;
  assign n5012 = x96 & n4772 ;
  assign n5013 = ( n4777 & n5011 ) | ( n4777 & n5012 ) | ( n5011 & n5012 ) ;
  assign n5014 = ( ~n4777 & n5011 ) | ( ~n4777 & n5012 ) | ( n5011 & n5012 ) ;
  assign n5015 = ( n4777 & ~n5013 ) | ( n4777 & n5014 ) | ( ~n5013 & n5014 ) ;
  assign n5016 = ( x97 & n5010 ) | ( x97 & ~n5015 ) | ( n5010 & ~n5015 ) ;
  assign n5017 = ( x97 & n4778 ) | ( x97 & ~n4819 ) | ( n4778 & ~n4819 ) ;
  assign n5018 = x97 & n4778 ;
  assign n5019 = ( ~n4783 & n5017 ) | ( ~n4783 & n5018 ) | ( n5017 & n5018 ) ;
  assign n5020 = ( n4783 & n5017 ) | ( n4783 & n5018 ) | ( n5017 & n5018 ) ;
  assign n5021 = ( n4783 & n5019 ) | ( n4783 & ~n5020 ) | ( n5019 & ~n5020 ) ;
  assign n5022 = ( x98 & n5016 ) | ( x98 & ~n5021 ) | ( n5016 & ~n5021 ) ;
  assign n5023 = ( x98 & n4784 ) | ( x98 & ~n4819 ) | ( n4784 & ~n4819 ) ;
  assign n5024 = x98 & n4784 ;
  assign n5025 = ( n4789 & n5023 ) | ( n4789 & n5024 ) | ( n5023 & n5024 ) ;
  assign n5026 = ( ~n4789 & n5023 ) | ( ~n4789 & n5024 ) | ( n5023 & n5024 ) ;
  assign n5027 = ( n4789 & ~n5025 ) | ( n4789 & n5026 ) | ( ~n5025 & n5026 ) ;
  assign n5028 = ( x99 & n5022 ) | ( x99 & ~n5027 ) | ( n5022 & ~n5027 ) ;
  assign n5029 = ( x99 & n4790 ) | ( x99 & ~n4819 ) | ( n4790 & ~n4819 ) ;
  assign n5030 = x99 & n4790 ;
  assign n5031 = ( ~n4795 & n5029 ) | ( ~n4795 & n5030 ) | ( n5029 & n5030 ) ;
  assign n5032 = ( n4795 & n5029 ) | ( n4795 & n5030 ) | ( n5029 & n5030 ) ;
  assign n5033 = ( n4795 & n5031 ) | ( n4795 & ~n5032 ) | ( n5031 & ~n5032 ) ;
  assign n5034 = ( x100 & n5028 ) | ( x100 & ~n5033 ) | ( n5028 & ~n5033 ) ;
  assign n5035 = ( x100 & n4796 ) | ( x100 & ~n4819 ) | ( n4796 & ~n4819 ) ;
  assign n5036 = x100 & n4796 ;
  assign n5037 = ( n4801 & n5035 ) | ( n4801 & n5036 ) | ( n5035 & n5036 ) ;
  assign n5038 = ( ~n4801 & n5035 ) | ( ~n4801 & n5036 ) | ( n5035 & n5036 ) ;
  assign n5039 = ( n4801 & ~n5037 ) | ( n4801 & n5038 ) | ( ~n5037 & n5038 ) ;
  assign n5040 = ( x101 & n5034 ) | ( x101 & ~n5039 ) | ( n5034 & ~n5039 ) ;
  assign n5041 = ( x101 & n4802 ) | ( x101 & ~n4819 ) | ( n4802 & ~n4819 ) ;
  assign n5042 = x101 & n4802 ;
  assign n5043 = ( ~n4807 & n5041 ) | ( ~n4807 & n5042 ) | ( n5041 & n5042 ) ;
  assign n5044 = ( n4807 & n5041 ) | ( n4807 & n5042 ) | ( n5041 & n5042 ) ;
  assign n5045 = ( n4807 & n5043 ) | ( n4807 & ~n5044 ) | ( n5043 & ~n5044 ) ;
  assign n5046 = ( x102 & n5040 ) | ( x102 & ~n5045 ) | ( n5040 & ~n5045 ) ;
  assign n5047 = ( x102 & n4808 ) | ( x102 & ~n4819 ) | ( n4808 & ~n4819 ) ;
  assign n5048 = x102 & n4808 ;
  assign n5049 = ( ~n4813 & n5047 ) | ( ~n4813 & n5048 ) | ( n5047 & n5048 ) ;
  assign n5050 = ( n4813 & n5047 ) | ( n4813 & n5048 ) | ( n5047 & n5048 ) ;
  assign n5051 = ( n4813 & n5049 ) | ( n4813 & ~n5050 ) | ( n5049 & ~n5050 ) ;
  assign n5052 = ( x103 & n5046 ) | ( x103 & ~n5051 ) | ( n5046 & ~n5051 ) ;
  assign n5053 = x104 | n5052 ;
  assign n5054 = ( x104 & n153 ) | ( x104 & n5052 ) | ( n153 & n5052 ) ;
  assign n5055 = ( n4817 & ~n5053 ) | ( n4817 & n5054 ) | ( ~n5053 & n5054 ) ;
  assign n5056 = ( x104 & ~n4817 ) | ( x104 & n5052 ) | ( ~n4817 & n5052 ) ;
  assign n5057 = n153 | n5056 ;
  assign n5058 = ( x23 & ~x64 ) | ( x23 & n5057 ) | ( ~x64 & n5057 ) ;
  assign n5059 = ~x23 & n5057 ;
  assign n5060 = ( n4823 & n5058 ) | ( n4823 & ~n5059 ) | ( n5058 & ~n5059 ) ;
  assign n5061 = ~x22 & x64 ;
  assign n5062 = ( x65 & ~n5060 ) | ( x65 & n5061 ) | ( ~n5060 & n5061 ) ;
  assign n5063 = ( x65 & n4823 ) | ( x65 & ~n5057 ) | ( n4823 & ~n5057 ) ;
  assign n5064 = x65 & n4823 ;
  assign n5065 = ( n4822 & n5063 ) | ( n4822 & n5064 ) | ( n5063 & n5064 ) ;
  assign n5066 = ( ~n4822 & n5063 ) | ( ~n4822 & n5064 ) | ( n5063 & n5064 ) ;
  assign n5067 = ( n4822 & ~n5065 ) | ( n4822 & n5066 ) | ( ~n5065 & n5066 ) ;
  assign n5068 = ( x66 & n5062 ) | ( x66 & ~n5067 ) | ( n5062 & ~n5067 ) ;
  assign n5069 = ( x66 & n4824 ) | ( x66 & ~n5057 ) | ( n4824 & ~n5057 ) ;
  assign n5070 = x66 & n4824 ;
  assign n5071 = ( n4829 & n5069 ) | ( n4829 & n5070 ) | ( n5069 & n5070 ) ;
  assign n5072 = ( ~n4829 & n5069 ) | ( ~n4829 & n5070 ) | ( n5069 & n5070 ) ;
  assign n5073 = ( n4829 & ~n5071 ) | ( n4829 & n5072 ) | ( ~n5071 & n5072 ) ;
  assign n5074 = ( x67 & n5068 ) | ( x67 & ~n5073 ) | ( n5068 & ~n5073 ) ;
  assign n5075 = ( x67 & n4830 ) | ( x67 & ~n5057 ) | ( n4830 & ~n5057 ) ;
  assign n5076 = x67 & n4830 ;
  assign n5077 = ( ~n4835 & n5075 ) | ( ~n4835 & n5076 ) | ( n5075 & n5076 ) ;
  assign n5078 = ( n4835 & n5075 ) | ( n4835 & n5076 ) | ( n5075 & n5076 ) ;
  assign n5079 = ( n4835 & n5077 ) | ( n4835 & ~n5078 ) | ( n5077 & ~n5078 ) ;
  assign n5080 = ( x68 & n5074 ) | ( x68 & ~n5079 ) | ( n5074 & ~n5079 ) ;
  assign n5081 = ( x68 & n4836 ) | ( x68 & ~n5057 ) | ( n4836 & ~n5057 ) ;
  assign n5082 = x68 & n4836 ;
  assign n5083 = ( n4841 & n5081 ) | ( n4841 & n5082 ) | ( n5081 & n5082 ) ;
  assign n5084 = ( ~n4841 & n5081 ) | ( ~n4841 & n5082 ) | ( n5081 & n5082 ) ;
  assign n5085 = ( n4841 & ~n5083 ) | ( n4841 & n5084 ) | ( ~n5083 & n5084 ) ;
  assign n5086 = ( x69 & n5080 ) | ( x69 & ~n5085 ) | ( n5080 & ~n5085 ) ;
  assign n5087 = ( x69 & n4842 ) | ( x69 & ~n5057 ) | ( n4842 & ~n5057 ) ;
  assign n5088 = x69 & n4842 ;
  assign n5089 = ( ~n4847 & n5087 ) | ( ~n4847 & n5088 ) | ( n5087 & n5088 ) ;
  assign n5090 = ( n4847 & n5087 ) | ( n4847 & n5088 ) | ( n5087 & n5088 ) ;
  assign n5091 = ( n4847 & n5089 ) | ( n4847 & ~n5090 ) | ( n5089 & ~n5090 ) ;
  assign n5092 = ( x70 & n5086 ) | ( x70 & ~n5091 ) | ( n5086 & ~n5091 ) ;
  assign n5093 = ( x70 & n4848 ) | ( x70 & ~n5057 ) | ( n4848 & ~n5057 ) ;
  assign n5094 = x70 & n4848 ;
  assign n5095 = ( n4853 & n5093 ) | ( n4853 & n5094 ) | ( n5093 & n5094 ) ;
  assign n5096 = ( ~n4853 & n5093 ) | ( ~n4853 & n5094 ) | ( n5093 & n5094 ) ;
  assign n5097 = ( n4853 & ~n5095 ) | ( n4853 & n5096 ) | ( ~n5095 & n5096 ) ;
  assign n5098 = ( x71 & n5092 ) | ( x71 & ~n5097 ) | ( n5092 & ~n5097 ) ;
  assign n5099 = ( x71 & n4854 ) | ( x71 & ~n5057 ) | ( n4854 & ~n5057 ) ;
  assign n5100 = x71 & n4854 ;
  assign n5101 = ( ~n4859 & n5099 ) | ( ~n4859 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5102 = ( n4859 & n5099 ) | ( n4859 & n5100 ) | ( n5099 & n5100 ) ;
  assign n5103 = ( n4859 & n5101 ) | ( n4859 & ~n5102 ) | ( n5101 & ~n5102 ) ;
  assign n5104 = ( x72 & n5098 ) | ( x72 & ~n5103 ) | ( n5098 & ~n5103 ) ;
  assign n5105 = ( x72 & n4860 ) | ( x72 & ~n5057 ) | ( n4860 & ~n5057 ) ;
  assign n5106 = x72 & n4860 ;
  assign n5107 = ( n4865 & n5105 ) | ( n4865 & n5106 ) | ( n5105 & n5106 ) ;
  assign n5108 = ( ~n4865 & n5105 ) | ( ~n4865 & n5106 ) | ( n5105 & n5106 ) ;
  assign n5109 = ( n4865 & ~n5107 ) | ( n4865 & n5108 ) | ( ~n5107 & n5108 ) ;
  assign n5110 = ( x73 & n5104 ) | ( x73 & ~n5109 ) | ( n5104 & ~n5109 ) ;
  assign n5111 = ( x73 & n4866 ) | ( x73 & ~n5057 ) | ( n4866 & ~n5057 ) ;
  assign n5112 = x73 & n4866 ;
  assign n5113 = ( ~n4871 & n5111 ) | ( ~n4871 & n5112 ) | ( n5111 & n5112 ) ;
  assign n5114 = ( n4871 & n5111 ) | ( n4871 & n5112 ) | ( n5111 & n5112 ) ;
  assign n5115 = ( n4871 & n5113 ) | ( n4871 & ~n5114 ) | ( n5113 & ~n5114 ) ;
  assign n5116 = ( x74 & n5110 ) | ( x74 & ~n5115 ) | ( n5110 & ~n5115 ) ;
  assign n5117 = ( x74 & n4872 ) | ( x74 & ~n5057 ) | ( n4872 & ~n5057 ) ;
  assign n5118 = x74 & n4872 ;
  assign n5119 = ( n4877 & n5117 ) | ( n4877 & n5118 ) | ( n5117 & n5118 ) ;
  assign n5120 = ( ~n4877 & n5117 ) | ( ~n4877 & n5118 ) | ( n5117 & n5118 ) ;
  assign n5121 = ( n4877 & ~n5119 ) | ( n4877 & n5120 ) | ( ~n5119 & n5120 ) ;
  assign n5122 = ( x75 & n5116 ) | ( x75 & ~n5121 ) | ( n5116 & ~n5121 ) ;
  assign n5123 = ( x75 & n4878 ) | ( x75 & ~n5057 ) | ( n4878 & ~n5057 ) ;
  assign n5124 = x75 & n4878 ;
  assign n5125 = ( ~n4883 & n5123 ) | ( ~n4883 & n5124 ) | ( n5123 & n5124 ) ;
  assign n5126 = ( n4883 & n5123 ) | ( n4883 & n5124 ) | ( n5123 & n5124 ) ;
  assign n5127 = ( n4883 & n5125 ) | ( n4883 & ~n5126 ) | ( n5125 & ~n5126 ) ;
  assign n5128 = ( x76 & n5122 ) | ( x76 & ~n5127 ) | ( n5122 & ~n5127 ) ;
  assign n5129 = ( x76 & n4884 ) | ( x76 & ~n5057 ) | ( n4884 & ~n5057 ) ;
  assign n5130 = x76 & n4884 ;
  assign n5131 = ( n4889 & n5129 ) | ( n4889 & n5130 ) | ( n5129 & n5130 ) ;
  assign n5132 = ( ~n4889 & n5129 ) | ( ~n4889 & n5130 ) | ( n5129 & n5130 ) ;
  assign n5133 = ( n4889 & ~n5131 ) | ( n4889 & n5132 ) | ( ~n5131 & n5132 ) ;
  assign n5134 = ( x77 & n5128 ) | ( x77 & ~n5133 ) | ( n5128 & ~n5133 ) ;
  assign n5135 = ( x77 & n4890 ) | ( x77 & ~n5057 ) | ( n4890 & ~n5057 ) ;
  assign n5136 = x77 & n4890 ;
  assign n5137 = ( ~n4895 & n5135 ) | ( ~n4895 & n5136 ) | ( n5135 & n5136 ) ;
  assign n5138 = ( n4895 & n5135 ) | ( n4895 & n5136 ) | ( n5135 & n5136 ) ;
  assign n5139 = ( n4895 & n5137 ) | ( n4895 & ~n5138 ) | ( n5137 & ~n5138 ) ;
  assign n5140 = ( x78 & n5134 ) | ( x78 & ~n5139 ) | ( n5134 & ~n5139 ) ;
  assign n5141 = ( x78 & n4896 ) | ( x78 & ~n5057 ) | ( n4896 & ~n5057 ) ;
  assign n5142 = x78 & n4896 ;
  assign n5143 = ( n4901 & n5141 ) | ( n4901 & n5142 ) | ( n5141 & n5142 ) ;
  assign n5144 = ( ~n4901 & n5141 ) | ( ~n4901 & n5142 ) | ( n5141 & n5142 ) ;
  assign n5145 = ( n4901 & ~n5143 ) | ( n4901 & n5144 ) | ( ~n5143 & n5144 ) ;
  assign n5146 = ( x79 & n5140 ) | ( x79 & ~n5145 ) | ( n5140 & ~n5145 ) ;
  assign n5147 = ( x79 & n4902 ) | ( x79 & ~n5057 ) | ( n4902 & ~n5057 ) ;
  assign n5148 = x79 & n4902 ;
  assign n5149 = ( ~n4907 & n5147 ) | ( ~n4907 & n5148 ) | ( n5147 & n5148 ) ;
  assign n5150 = ( n4907 & n5147 ) | ( n4907 & n5148 ) | ( n5147 & n5148 ) ;
  assign n5151 = ( n4907 & n5149 ) | ( n4907 & ~n5150 ) | ( n5149 & ~n5150 ) ;
  assign n5152 = ( x80 & n5146 ) | ( x80 & ~n5151 ) | ( n5146 & ~n5151 ) ;
  assign n5153 = ( x80 & n4908 ) | ( x80 & ~n5057 ) | ( n4908 & ~n5057 ) ;
  assign n5154 = x80 & n4908 ;
  assign n5155 = ( n4913 & n5153 ) | ( n4913 & n5154 ) | ( n5153 & n5154 ) ;
  assign n5156 = ( ~n4913 & n5153 ) | ( ~n4913 & n5154 ) | ( n5153 & n5154 ) ;
  assign n5157 = ( n4913 & ~n5155 ) | ( n4913 & n5156 ) | ( ~n5155 & n5156 ) ;
  assign n5158 = ( x81 & n5152 ) | ( x81 & ~n5157 ) | ( n5152 & ~n5157 ) ;
  assign n5159 = ( x81 & n4914 ) | ( x81 & ~n5057 ) | ( n4914 & ~n5057 ) ;
  assign n5160 = x81 & n4914 ;
  assign n5161 = ( ~n4919 & n5159 ) | ( ~n4919 & n5160 ) | ( n5159 & n5160 ) ;
  assign n5162 = ( n4919 & n5159 ) | ( n4919 & n5160 ) | ( n5159 & n5160 ) ;
  assign n5163 = ( n4919 & n5161 ) | ( n4919 & ~n5162 ) | ( n5161 & ~n5162 ) ;
  assign n5164 = ( x82 & n5158 ) | ( x82 & ~n5163 ) | ( n5158 & ~n5163 ) ;
  assign n5165 = ( x82 & n4920 ) | ( x82 & ~n5057 ) | ( n4920 & ~n5057 ) ;
  assign n5166 = x82 & n4920 ;
  assign n5167 = ( n4925 & n5165 ) | ( n4925 & n5166 ) | ( n5165 & n5166 ) ;
  assign n5168 = ( ~n4925 & n5165 ) | ( ~n4925 & n5166 ) | ( n5165 & n5166 ) ;
  assign n5169 = ( n4925 & ~n5167 ) | ( n4925 & n5168 ) | ( ~n5167 & n5168 ) ;
  assign n5170 = ( x83 & n5164 ) | ( x83 & ~n5169 ) | ( n5164 & ~n5169 ) ;
  assign n5171 = ( x83 & n4926 ) | ( x83 & ~n5057 ) | ( n4926 & ~n5057 ) ;
  assign n5172 = x83 & n4926 ;
  assign n5173 = ( ~n4931 & n5171 ) | ( ~n4931 & n5172 ) | ( n5171 & n5172 ) ;
  assign n5174 = ( n4931 & n5171 ) | ( n4931 & n5172 ) | ( n5171 & n5172 ) ;
  assign n5175 = ( n4931 & n5173 ) | ( n4931 & ~n5174 ) | ( n5173 & ~n5174 ) ;
  assign n5176 = ( x84 & n5170 ) | ( x84 & ~n5175 ) | ( n5170 & ~n5175 ) ;
  assign n5177 = ( x84 & n4932 ) | ( x84 & ~n5057 ) | ( n4932 & ~n5057 ) ;
  assign n5178 = x84 & n4932 ;
  assign n5179 = ( n4937 & n5177 ) | ( n4937 & n5178 ) | ( n5177 & n5178 ) ;
  assign n5180 = ( ~n4937 & n5177 ) | ( ~n4937 & n5178 ) | ( n5177 & n5178 ) ;
  assign n5181 = ( n4937 & ~n5179 ) | ( n4937 & n5180 ) | ( ~n5179 & n5180 ) ;
  assign n5182 = ( x85 & n5176 ) | ( x85 & ~n5181 ) | ( n5176 & ~n5181 ) ;
  assign n5183 = ( x85 & n4938 ) | ( x85 & ~n5057 ) | ( n4938 & ~n5057 ) ;
  assign n5184 = x85 & n4938 ;
  assign n5185 = ( ~n4943 & n5183 ) | ( ~n4943 & n5184 ) | ( n5183 & n5184 ) ;
  assign n5186 = ( n4943 & n5183 ) | ( n4943 & n5184 ) | ( n5183 & n5184 ) ;
  assign n5187 = ( n4943 & n5185 ) | ( n4943 & ~n5186 ) | ( n5185 & ~n5186 ) ;
  assign n5188 = ( x86 & n5182 ) | ( x86 & ~n5187 ) | ( n5182 & ~n5187 ) ;
  assign n5189 = ( x86 & n4944 ) | ( x86 & ~n5057 ) | ( n4944 & ~n5057 ) ;
  assign n5190 = x86 & n4944 ;
  assign n5191 = ( n4949 & n5189 ) | ( n4949 & n5190 ) | ( n5189 & n5190 ) ;
  assign n5192 = ( ~n4949 & n5189 ) | ( ~n4949 & n5190 ) | ( n5189 & n5190 ) ;
  assign n5193 = ( n4949 & ~n5191 ) | ( n4949 & n5192 ) | ( ~n5191 & n5192 ) ;
  assign n5194 = ( x87 & n5188 ) | ( x87 & ~n5193 ) | ( n5188 & ~n5193 ) ;
  assign n5195 = ( x87 & n4950 ) | ( x87 & ~n5057 ) | ( n4950 & ~n5057 ) ;
  assign n5196 = x87 & n4950 ;
  assign n5197 = ( ~n4955 & n5195 ) | ( ~n4955 & n5196 ) | ( n5195 & n5196 ) ;
  assign n5198 = ( n4955 & n5195 ) | ( n4955 & n5196 ) | ( n5195 & n5196 ) ;
  assign n5199 = ( n4955 & n5197 ) | ( n4955 & ~n5198 ) | ( n5197 & ~n5198 ) ;
  assign n5200 = ( x88 & n5194 ) | ( x88 & ~n5199 ) | ( n5194 & ~n5199 ) ;
  assign n5201 = ( x88 & n4956 ) | ( x88 & ~n5057 ) | ( n4956 & ~n5057 ) ;
  assign n5202 = x88 & n4956 ;
  assign n5203 = ( n4961 & n5201 ) | ( n4961 & n5202 ) | ( n5201 & n5202 ) ;
  assign n5204 = ( ~n4961 & n5201 ) | ( ~n4961 & n5202 ) | ( n5201 & n5202 ) ;
  assign n5205 = ( n4961 & ~n5203 ) | ( n4961 & n5204 ) | ( ~n5203 & n5204 ) ;
  assign n5206 = ( x89 & n5200 ) | ( x89 & ~n5205 ) | ( n5200 & ~n5205 ) ;
  assign n5207 = ( x89 & n4962 ) | ( x89 & ~n5057 ) | ( n4962 & ~n5057 ) ;
  assign n5208 = x89 & n4962 ;
  assign n5209 = ( ~n4967 & n5207 ) | ( ~n4967 & n5208 ) | ( n5207 & n5208 ) ;
  assign n5210 = ( n4967 & n5207 ) | ( n4967 & n5208 ) | ( n5207 & n5208 ) ;
  assign n5211 = ( n4967 & n5209 ) | ( n4967 & ~n5210 ) | ( n5209 & ~n5210 ) ;
  assign n5212 = ( x90 & n5206 ) | ( x90 & ~n5211 ) | ( n5206 & ~n5211 ) ;
  assign n5213 = ( x90 & n4968 ) | ( x90 & ~n5057 ) | ( n4968 & ~n5057 ) ;
  assign n5214 = x90 & n4968 ;
  assign n5215 = ( n4973 & n5213 ) | ( n4973 & n5214 ) | ( n5213 & n5214 ) ;
  assign n5216 = ( ~n4973 & n5213 ) | ( ~n4973 & n5214 ) | ( n5213 & n5214 ) ;
  assign n5217 = ( n4973 & ~n5215 ) | ( n4973 & n5216 ) | ( ~n5215 & n5216 ) ;
  assign n5218 = ( x91 & n5212 ) | ( x91 & ~n5217 ) | ( n5212 & ~n5217 ) ;
  assign n5219 = ( x91 & n4974 ) | ( x91 & ~n5057 ) | ( n4974 & ~n5057 ) ;
  assign n5220 = x91 & n4974 ;
  assign n5221 = ( ~n4979 & n5219 ) | ( ~n4979 & n5220 ) | ( n5219 & n5220 ) ;
  assign n5222 = ( n4979 & n5219 ) | ( n4979 & n5220 ) | ( n5219 & n5220 ) ;
  assign n5223 = ( n4979 & n5221 ) | ( n4979 & ~n5222 ) | ( n5221 & ~n5222 ) ;
  assign n5224 = ( x92 & n5218 ) | ( x92 & ~n5223 ) | ( n5218 & ~n5223 ) ;
  assign n5225 = ( x92 & n4980 ) | ( x92 & ~n5057 ) | ( n4980 & ~n5057 ) ;
  assign n5226 = x92 & n4980 ;
  assign n5227 = ( n4985 & n5225 ) | ( n4985 & n5226 ) | ( n5225 & n5226 ) ;
  assign n5228 = ( ~n4985 & n5225 ) | ( ~n4985 & n5226 ) | ( n5225 & n5226 ) ;
  assign n5229 = ( n4985 & ~n5227 ) | ( n4985 & n5228 ) | ( ~n5227 & n5228 ) ;
  assign n5230 = ( x93 & n5224 ) | ( x93 & ~n5229 ) | ( n5224 & ~n5229 ) ;
  assign n5231 = ( x93 & n4986 ) | ( x93 & ~n5057 ) | ( n4986 & ~n5057 ) ;
  assign n5232 = x93 & n4986 ;
  assign n5233 = ( ~n4991 & n5231 ) | ( ~n4991 & n5232 ) | ( n5231 & n5232 ) ;
  assign n5234 = ( n4991 & n5231 ) | ( n4991 & n5232 ) | ( n5231 & n5232 ) ;
  assign n5235 = ( n4991 & n5233 ) | ( n4991 & ~n5234 ) | ( n5233 & ~n5234 ) ;
  assign n5236 = ( x94 & n5230 ) | ( x94 & ~n5235 ) | ( n5230 & ~n5235 ) ;
  assign n5237 = ( x94 & n4992 ) | ( x94 & ~n5057 ) | ( n4992 & ~n5057 ) ;
  assign n5238 = x94 & n4992 ;
  assign n5239 = ( n4997 & n5237 ) | ( n4997 & n5238 ) | ( n5237 & n5238 ) ;
  assign n5240 = ( ~n4997 & n5237 ) | ( ~n4997 & n5238 ) | ( n5237 & n5238 ) ;
  assign n5241 = ( n4997 & ~n5239 ) | ( n4997 & n5240 ) | ( ~n5239 & n5240 ) ;
  assign n5242 = ( x95 & n5236 ) | ( x95 & ~n5241 ) | ( n5236 & ~n5241 ) ;
  assign n5243 = ( x95 & n4998 ) | ( x95 & ~n5057 ) | ( n4998 & ~n5057 ) ;
  assign n5244 = x95 & n4998 ;
  assign n5245 = ( ~n5003 & n5243 ) | ( ~n5003 & n5244 ) | ( n5243 & n5244 ) ;
  assign n5246 = ( n5003 & n5243 ) | ( n5003 & n5244 ) | ( n5243 & n5244 ) ;
  assign n5247 = ( n5003 & n5245 ) | ( n5003 & ~n5246 ) | ( n5245 & ~n5246 ) ;
  assign n5248 = ( x96 & n5242 ) | ( x96 & ~n5247 ) | ( n5242 & ~n5247 ) ;
  assign n5249 = ( x96 & n5004 ) | ( x96 & ~n5057 ) | ( n5004 & ~n5057 ) ;
  assign n5250 = x96 & n5004 ;
  assign n5251 = ( n5009 & n5249 ) | ( n5009 & n5250 ) | ( n5249 & n5250 ) ;
  assign n5252 = ( ~n5009 & n5249 ) | ( ~n5009 & n5250 ) | ( n5249 & n5250 ) ;
  assign n5253 = ( n5009 & ~n5251 ) | ( n5009 & n5252 ) | ( ~n5251 & n5252 ) ;
  assign n5254 = ( x97 & n5248 ) | ( x97 & ~n5253 ) | ( n5248 & ~n5253 ) ;
  assign n5255 = ( x97 & n5010 ) | ( x97 & ~n5057 ) | ( n5010 & ~n5057 ) ;
  assign n5256 = x97 & n5010 ;
  assign n5257 = ( ~n5015 & n5255 ) | ( ~n5015 & n5256 ) | ( n5255 & n5256 ) ;
  assign n5258 = ( n5015 & n5255 ) | ( n5015 & n5256 ) | ( n5255 & n5256 ) ;
  assign n5259 = ( n5015 & n5257 ) | ( n5015 & ~n5258 ) | ( n5257 & ~n5258 ) ;
  assign n5260 = ( x98 & n5254 ) | ( x98 & ~n5259 ) | ( n5254 & ~n5259 ) ;
  assign n5261 = ( x98 & n5016 ) | ( x98 & ~n5057 ) | ( n5016 & ~n5057 ) ;
  assign n5262 = x98 & n5016 ;
  assign n5263 = ( n5021 & n5261 ) | ( n5021 & n5262 ) | ( n5261 & n5262 ) ;
  assign n5264 = ( ~n5021 & n5261 ) | ( ~n5021 & n5262 ) | ( n5261 & n5262 ) ;
  assign n5265 = ( n5021 & ~n5263 ) | ( n5021 & n5264 ) | ( ~n5263 & n5264 ) ;
  assign n5266 = ( x99 & n5260 ) | ( x99 & ~n5265 ) | ( n5260 & ~n5265 ) ;
  assign n5267 = ( x99 & n5022 ) | ( x99 & ~n5057 ) | ( n5022 & ~n5057 ) ;
  assign n5268 = x99 & n5022 ;
  assign n5269 = ( ~n5027 & n5267 ) | ( ~n5027 & n5268 ) | ( n5267 & n5268 ) ;
  assign n5270 = ( n5027 & n5267 ) | ( n5027 & n5268 ) | ( n5267 & n5268 ) ;
  assign n5271 = ( n5027 & n5269 ) | ( n5027 & ~n5270 ) | ( n5269 & ~n5270 ) ;
  assign n5272 = ( x100 & n5266 ) | ( x100 & ~n5271 ) | ( n5266 & ~n5271 ) ;
  assign n5273 = ( x100 & n5028 ) | ( x100 & ~n5057 ) | ( n5028 & ~n5057 ) ;
  assign n5274 = x100 & n5028 ;
  assign n5275 = ( n5033 & n5273 ) | ( n5033 & n5274 ) | ( n5273 & n5274 ) ;
  assign n5276 = ( ~n5033 & n5273 ) | ( ~n5033 & n5274 ) | ( n5273 & n5274 ) ;
  assign n5277 = ( n5033 & ~n5275 ) | ( n5033 & n5276 ) | ( ~n5275 & n5276 ) ;
  assign n5278 = ( x101 & n5272 ) | ( x101 & ~n5277 ) | ( n5272 & ~n5277 ) ;
  assign n5279 = ( x101 & n5034 ) | ( x101 & ~n5057 ) | ( n5034 & ~n5057 ) ;
  assign n5280 = x101 & n5034 ;
  assign n5281 = ( ~n5039 & n5279 ) | ( ~n5039 & n5280 ) | ( n5279 & n5280 ) ;
  assign n5282 = ( n5039 & n5279 ) | ( n5039 & n5280 ) | ( n5279 & n5280 ) ;
  assign n5283 = ( n5039 & n5281 ) | ( n5039 & ~n5282 ) | ( n5281 & ~n5282 ) ;
  assign n5284 = ( x102 & n5278 ) | ( x102 & ~n5283 ) | ( n5278 & ~n5283 ) ;
  assign n5285 = ( x102 & n5040 ) | ( x102 & ~n5057 ) | ( n5040 & ~n5057 ) ;
  assign n5286 = x102 & n5040 ;
  assign n5287 = ( n5045 & n5285 ) | ( n5045 & n5286 ) | ( n5285 & n5286 ) ;
  assign n5288 = ( ~n5045 & n5285 ) | ( ~n5045 & n5286 ) | ( n5285 & n5286 ) ;
  assign n5289 = ( n5045 & ~n5287 ) | ( n5045 & n5288 ) | ( ~n5287 & n5288 ) ;
  assign n5290 = ( x103 & n5284 ) | ( x103 & ~n5289 ) | ( n5284 & ~n5289 ) ;
  assign n5291 = ( x103 & n5046 ) | ( x103 & ~n5057 ) | ( n5046 & ~n5057 ) ;
  assign n5292 = x103 & n5046 ;
  assign n5293 = ( n5051 & n5291 ) | ( n5051 & n5292 ) | ( n5291 & n5292 ) ;
  assign n5294 = ( ~n5051 & n5291 ) | ( ~n5051 & n5292 ) | ( n5291 & n5292 ) ;
  assign n5295 = ( n5051 & ~n5293 ) | ( n5051 & n5294 ) | ( ~n5293 & n5294 ) ;
  assign n5296 = ( x104 & n5290 ) | ( x104 & ~n5295 ) | ( n5290 & ~n5295 ) ;
  assign n5297 = x105 | n5296 ;
  assign n5298 = ( x105 & n152 ) | ( x105 & n5296 ) | ( n152 & n5296 ) ;
  assign n5299 = ( n5055 & ~n5297 ) | ( n5055 & n5298 ) | ( ~n5297 & n5298 ) ;
  assign n5300 = ( x105 & ~n5055 ) | ( x105 & n5296 ) | ( ~n5055 & n5296 ) ;
  assign n5301 = n152 | n5300 ;
  assign n5302 = ( x22 & ~x64 ) | ( x22 & n5301 ) | ( ~x64 & n5301 ) ;
  assign n5303 = ~x22 & n5301 ;
  assign n5304 = ( n5061 & n5302 ) | ( n5061 & ~n5303 ) | ( n5302 & ~n5303 ) ;
  assign n5305 = ~x21 & x64 ;
  assign n5306 = ( x65 & ~n5304 ) | ( x65 & n5305 ) | ( ~n5304 & n5305 ) ;
  assign n5307 = ( x65 & n5061 ) | ( x65 & ~n5301 ) | ( n5061 & ~n5301 ) ;
  assign n5308 = x65 & n5061 ;
  assign n5309 = ( n5060 & n5307 ) | ( n5060 & n5308 ) | ( n5307 & n5308 ) ;
  assign n5310 = ( ~n5060 & n5307 ) | ( ~n5060 & n5308 ) | ( n5307 & n5308 ) ;
  assign n5311 = ( n5060 & ~n5309 ) | ( n5060 & n5310 ) | ( ~n5309 & n5310 ) ;
  assign n5312 = ( x66 & n5306 ) | ( x66 & ~n5311 ) | ( n5306 & ~n5311 ) ;
  assign n5313 = ( x66 & n5062 ) | ( x66 & ~n5301 ) | ( n5062 & ~n5301 ) ;
  assign n5314 = x66 & n5062 ;
  assign n5315 = ( n5067 & n5313 ) | ( n5067 & n5314 ) | ( n5313 & n5314 ) ;
  assign n5316 = ( ~n5067 & n5313 ) | ( ~n5067 & n5314 ) | ( n5313 & n5314 ) ;
  assign n5317 = ( n5067 & ~n5315 ) | ( n5067 & n5316 ) | ( ~n5315 & n5316 ) ;
  assign n5318 = ( x67 & n5312 ) | ( x67 & ~n5317 ) | ( n5312 & ~n5317 ) ;
  assign n5319 = ( x67 & n5068 ) | ( x67 & ~n5301 ) | ( n5068 & ~n5301 ) ;
  assign n5320 = x67 & n5068 ;
  assign n5321 = ( ~n5073 & n5319 ) | ( ~n5073 & n5320 ) | ( n5319 & n5320 ) ;
  assign n5322 = ( n5073 & n5319 ) | ( n5073 & n5320 ) | ( n5319 & n5320 ) ;
  assign n5323 = ( n5073 & n5321 ) | ( n5073 & ~n5322 ) | ( n5321 & ~n5322 ) ;
  assign n5324 = ( x68 & n5318 ) | ( x68 & ~n5323 ) | ( n5318 & ~n5323 ) ;
  assign n5325 = ( x68 & n5074 ) | ( x68 & ~n5301 ) | ( n5074 & ~n5301 ) ;
  assign n5326 = x68 & n5074 ;
  assign n5327 = ( n5079 & n5325 ) | ( n5079 & n5326 ) | ( n5325 & n5326 ) ;
  assign n5328 = ( ~n5079 & n5325 ) | ( ~n5079 & n5326 ) | ( n5325 & n5326 ) ;
  assign n5329 = ( n5079 & ~n5327 ) | ( n5079 & n5328 ) | ( ~n5327 & n5328 ) ;
  assign n5330 = ( x69 & n5324 ) | ( x69 & ~n5329 ) | ( n5324 & ~n5329 ) ;
  assign n5331 = ( x69 & n5080 ) | ( x69 & ~n5301 ) | ( n5080 & ~n5301 ) ;
  assign n5332 = x69 & n5080 ;
  assign n5333 = ( ~n5085 & n5331 ) | ( ~n5085 & n5332 ) | ( n5331 & n5332 ) ;
  assign n5334 = ( n5085 & n5331 ) | ( n5085 & n5332 ) | ( n5331 & n5332 ) ;
  assign n5335 = ( n5085 & n5333 ) | ( n5085 & ~n5334 ) | ( n5333 & ~n5334 ) ;
  assign n5336 = ( x70 & n5330 ) | ( x70 & ~n5335 ) | ( n5330 & ~n5335 ) ;
  assign n5337 = ( x70 & n5086 ) | ( x70 & ~n5301 ) | ( n5086 & ~n5301 ) ;
  assign n5338 = x70 & n5086 ;
  assign n5339 = ( n5091 & n5337 ) | ( n5091 & n5338 ) | ( n5337 & n5338 ) ;
  assign n5340 = ( ~n5091 & n5337 ) | ( ~n5091 & n5338 ) | ( n5337 & n5338 ) ;
  assign n5341 = ( n5091 & ~n5339 ) | ( n5091 & n5340 ) | ( ~n5339 & n5340 ) ;
  assign n5342 = ( x71 & n5336 ) | ( x71 & ~n5341 ) | ( n5336 & ~n5341 ) ;
  assign n5343 = ( x71 & n5092 ) | ( x71 & ~n5301 ) | ( n5092 & ~n5301 ) ;
  assign n5344 = x71 & n5092 ;
  assign n5345 = ( ~n5097 & n5343 ) | ( ~n5097 & n5344 ) | ( n5343 & n5344 ) ;
  assign n5346 = ( n5097 & n5343 ) | ( n5097 & n5344 ) | ( n5343 & n5344 ) ;
  assign n5347 = ( n5097 & n5345 ) | ( n5097 & ~n5346 ) | ( n5345 & ~n5346 ) ;
  assign n5348 = ( x72 & n5342 ) | ( x72 & ~n5347 ) | ( n5342 & ~n5347 ) ;
  assign n5349 = ( x72 & n5098 ) | ( x72 & ~n5301 ) | ( n5098 & ~n5301 ) ;
  assign n5350 = x72 & n5098 ;
  assign n5351 = ( n5103 & n5349 ) | ( n5103 & n5350 ) | ( n5349 & n5350 ) ;
  assign n5352 = ( ~n5103 & n5349 ) | ( ~n5103 & n5350 ) | ( n5349 & n5350 ) ;
  assign n5353 = ( n5103 & ~n5351 ) | ( n5103 & n5352 ) | ( ~n5351 & n5352 ) ;
  assign n5354 = ( x73 & n5348 ) | ( x73 & ~n5353 ) | ( n5348 & ~n5353 ) ;
  assign n5355 = ( x73 & n5104 ) | ( x73 & ~n5301 ) | ( n5104 & ~n5301 ) ;
  assign n5356 = x73 & n5104 ;
  assign n5357 = ( ~n5109 & n5355 ) | ( ~n5109 & n5356 ) | ( n5355 & n5356 ) ;
  assign n5358 = ( n5109 & n5355 ) | ( n5109 & n5356 ) | ( n5355 & n5356 ) ;
  assign n5359 = ( n5109 & n5357 ) | ( n5109 & ~n5358 ) | ( n5357 & ~n5358 ) ;
  assign n5360 = ( x74 & n5354 ) | ( x74 & ~n5359 ) | ( n5354 & ~n5359 ) ;
  assign n5361 = ( x74 & n5110 ) | ( x74 & ~n5301 ) | ( n5110 & ~n5301 ) ;
  assign n5362 = x74 & n5110 ;
  assign n5363 = ( n5115 & n5361 ) | ( n5115 & n5362 ) | ( n5361 & n5362 ) ;
  assign n5364 = ( ~n5115 & n5361 ) | ( ~n5115 & n5362 ) | ( n5361 & n5362 ) ;
  assign n5365 = ( n5115 & ~n5363 ) | ( n5115 & n5364 ) | ( ~n5363 & n5364 ) ;
  assign n5366 = ( x75 & n5360 ) | ( x75 & ~n5365 ) | ( n5360 & ~n5365 ) ;
  assign n5367 = ( x75 & n5116 ) | ( x75 & ~n5301 ) | ( n5116 & ~n5301 ) ;
  assign n5368 = x75 & n5116 ;
  assign n5369 = ( ~n5121 & n5367 ) | ( ~n5121 & n5368 ) | ( n5367 & n5368 ) ;
  assign n5370 = ( n5121 & n5367 ) | ( n5121 & n5368 ) | ( n5367 & n5368 ) ;
  assign n5371 = ( n5121 & n5369 ) | ( n5121 & ~n5370 ) | ( n5369 & ~n5370 ) ;
  assign n5372 = ( x76 & n5366 ) | ( x76 & ~n5371 ) | ( n5366 & ~n5371 ) ;
  assign n5373 = ( x76 & n5122 ) | ( x76 & ~n5301 ) | ( n5122 & ~n5301 ) ;
  assign n5374 = x76 & n5122 ;
  assign n5375 = ( n5127 & n5373 ) | ( n5127 & n5374 ) | ( n5373 & n5374 ) ;
  assign n5376 = ( ~n5127 & n5373 ) | ( ~n5127 & n5374 ) | ( n5373 & n5374 ) ;
  assign n5377 = ( n5127 & ~n5375 ) | ( n5127 & n5376 ) | ( ~n5375 & n5376 ) ;
  assign n5378 = ( x77 & n5372 ) | ( x77 & ~n5377 ) | ( n5372 & ~n5377 ) ;
  assign n5379 = ( x77 & n5128 ) | ( x77 & ~n5301 ) | ( n5128 & ~n5301 ) ;
  assign n5380 = x77 & n5128 ;
  assign n5381 = ( ~n5133 & n5379 ) | ( ~n5133 & n5380 ) | ( n5379 & n5380 ) ;
  assign n5382 = ( n5133 & n5379 ) | ( n5133 & n5380 ) | ( n5379 & n5380 ) ;
  assign n5383 = ( n5133 & n5381 ) | ( n5133 & ~n5382 ) | ( n5381 & ~n5382 ) ;
  assign n5384 = ( x78 & n5378 ) | ( x78 & ~n5383 ) | ( n5378 & ~n5383 ) ;
  assign n5385 = ( x78 & n5134 ) | ( x78 & ~n5301 ) | ( n5134 & ~n5301 ) ;
  assign n5386 = x78 & n5134 ;
  assign n5387 = ( n5139 & n5385 ) | ( n5139 & n5386 ) | ( n5385 & n5386 ) ;
  assign n5388 = ( ~n5139 & n5385 ) | ( ~n5139 & n5386 ) | ( n5385 & n5386 ) ;
  assign n5389 = ( n5139 & ~n5387 ) | ( n5139 & n5388 ) | ( ~n5387 & n5388 ) ;
  assign n5390 = ( x79 & n5384 ) | ( x79 & ~n5389 ) | ( n5384 & ~n5389 ) ;
  assign n5391 = ( x79 & n5140 ) | ( x79 & ~n5301 ) | ( n5140 & ~n5301 ) ;
  assign n5392 = x79 & n5140 ;
  assign n5393 = ( ~n5145 & n5391 ) | ( ~n5145 & n5392 ) | ( n5391 & n5392 ) ;
  assign n5394 = ( n5145 & n5391 ) | ( n5145 & n5392 ) | ( n5391 & n5392 ) ;
  assign n5395 = ( n5145 & n5393 ) | ( n5145 & ~n5394 ) | ( n5393 & ~n5394 ) ;
  assign n5396 = ( x80 & n5390 ) | ( x80 & ~n5395 ) | ( n5390 & ~n5395 ) ;
  assign n5397 = ( x80 & n5146 ) | ( x80 & ~n5301 ) | ( n5146 & ~n5301 ) ;
  assign n5398 = x80 & n5146 ;
  assign n5399 = ( n5151 & n5397 ) | ( n5151 & n5398 ) | ( n5397 & n5398 ) ;
  assign n5400 = ( ~n5151 & n5397 ) | ( ~n5151 & n5398 ) | ( n5397 & n5398 ) ;
  assign n5401 = ( n5151 & ~n5399 ) | ( n5151 & n5400 ) | ( ~n5399 & n5400 ) ;
  assign n5402 = ( x81 & n5396 ) | ( x81 & ~n5401 ) | ( n5396 & ~n5401 ) ;
  assign n5403 = ( x81 & n5152 ) | ( x81 & ~n5301 ) | ( n5152 & ~n5301 ) ;
  assign n5404 = x81 & n5152 ;
  assign n5405 = ( ~n5157 & n5403 ) | ( ~n5157 & n5404 ) | ( n5403 & n5404 ) ;
  assign n5406 = ( n5157 & n5403 ) | ( n5157 & n5404 ) | ( n5403 & n5404 ) ;
  assign n5407 = ( n5157 & n5405 ) | ( n5157 & ~n5406 ) | ( n5405 & ~n5406 ) ;
  assign n5408 = ( x82 & n5402 ) | ( x82 & ~n5407 ) | ( n5402 & ~n5407 ) ;
  assign n5409 = ( x82 & n5158 ) | ( x82 & ~n5301 ) | ( n5158 & ~n5301 ) ;
  assign n5410 = x82 & n5158 ;
  assign n5411 = ( n5163 & n5409 ) | ( n5163 & n5410 ) | ( n5409 & n5410 ) ;
  assign n5412 = ( ~n5163 & n5409 ) | ( ~n5163 & n5410 ) | ( n5409 & n5410 ) ;
  assign n5413 = ( n5163 & ~n5411 ) | ( n5163 & n5412 ) | ( ~n5411 & n5412 ) ;
  assign n5414 = ( x83 & n5408 ) | ( x83 & ~n5413 ) | ( n5408 & ~n5413 ) ;
  assign n5415 = ( x83 & n5164 ) | ( x83 & ~n5301 ) | ( n5164 & ~n5301 ) ;
  assign n5416 = x83 & n5164 ;
  assign n5417 = ( ~n5169 & n5415 ) | ( ~n5169 & n5416 ) | ( n5415 & n5416 ) ;
  assign n5418 = ( n5169 & n5415 ) | ( n5169 & n5416 ) | ( n5415 & n5416 ) ;
  assign n5419 = ( n5169 & n5417 ) | ( n5169 & ~n5418 ) | ( n5417 & ~n5418 ) ;
  assign n5420 = ( x84 & n5414 ) | ( x84 & ~n5419 ) | ( n5414 & ~n5419 ) ;
  assign n5421 = ( x84 & n5170 ) | ( x84 & ~n5301 ) | ( n5170 & ~n5301 ) ;
  assign n5422 = x84 & n5170 ;
  assign n5423 = ( n5175 & n5421 ) | ( n5175 & n5422 ) | ( n5421 & n5422 ) ;
  assign n5424 = ( ~n5175 & n5421 ) | ( ~n5175 & n5422 ) | ( n5421 & n5422 ) ;
  assign n5425 = ( n5175 & ~n5423 ) | ( n5175 & n5424 ) | ( ~n5423 & n5424 ) ;
  assign n5426 = ( x85 & n5420 ) | ( x85 & ~n5425 ) | ( n5420 & ~n5425 ) ;
  assign n5427 = ( x85 & n5176 ) | ( x85 & ~n5301 ) | ( n5176 & ~n5301 ) ;
  assign n5428 = x85 & n5176 ;
  assign n5429 = ( ~n5181 & n5427 ) | ( ~n5181 & n5428 ) | ( n5427 & n5428 ) ;
  assign n5430 = ( n5181 & n5427 ) | ( n5181 & n5428 ) | ( n5427 & n5428 ) ;
  assign n5431 = ( n5181 & n5429 ) | ( n5181 & ~n5430 ) | ( n5429 & ~n5430 ) ;
  assign n5432 = ( x86 & n5426 ) | ( x86 & ~n5431 ) | ( n5426 & ~n5431 ) ;
  assign n5433 = ( x86 & n5182 ) | ( x86 & ~n5301 ) | ( n5182 & ~n5301 ) ;
  assign n5434 = x86 & n5182 ;
  assign n5435 = ( n5187 & n5433 ) | ( n5187 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5436 = ( ~n5187 & n5433 ) | ( ~n5187 & n5434 ) | ( n5433 & n5434 ) ;
  assign n5437 = ( n5187 & ~n5435 ) | ( n5187 & n5436 ) | ( ~n5435 & n5436 ) ;
  assign n5438 = ( x87 & n5432 ) | ( x87 & ~n5437 ) | ( n5432 & ~n5437 ) ;
  assign n5439 = ( x87 & n5188 ) | ( x87 & ~n5301 ) | ( n5188 & ~n5301 ) ;
  assign n5440 = x87 & n5188 ;
  assign n5441 = ( ~n5193 & n5439 ) | ( ~n5193 & n5440 ) | ( n5439 & n5440 ) ;
  assign n5442 = ( n5193 & n5439 ) | ( n5193 & n5440 ) | ( n5439 & n5440 ) ;
  assign n5443 = ( n5193 & n5441 ) | ( n5193 & ~n5442 ) | ( n5441 & ~n5442 ) ;
  assign n5444 = ( x88 & n5438 ) | ( x88 & ~n5443 ) | ( n5438 & ~n5443 ) ;
  assign n5445 = ( x88 & n5194 ) | ( x88 & ~n5301 ) | ( n5194 & ~n5301 ) ;
  assign n5446 = x88 & n5194 ;
  assign n5447 = ( n5199 & n5445 ) | ( n5199 & n5446 ) | ( n5445 & n5446 ) ;
  assign n5448 = ( ~n5199 & n5445 ) | ( ~n5199 & n5446 ) | ( n5445 & n5446 ) ;
  assign n5449 = ( n5199 & ~n5447 ) | ( n5199 & n5448 ) | ( ~n5447 & n5448 ) ;
  assign n5450 = ( x89 & n5444 ) | ( x89 & ~n5449 ) | ( n5444 & ~n5449 ) ;
  assign n5451 = ( x89 & n5200 ) | ( x89 & ~n5301 ) | ( n5200 & ~n5301 ) ;
  assign n5452 = x89 & n5200 ;
  assign n5453 = ( ~n5205 & n5451 ) | ( ~n5205 & n5452 ) | ( n5451 & n5452 ) ;
  assign n5454 = ( n5205 & n5451 ) | ( n5205 & n5452 ) | ( n5451 & n5452 ) ;
  assign n5455 = ( n5205 & n5453 ) | ( n5205 & ~n5454 ) | ( n5453 & ~n5454 ) ;
  assign n5456 = ( x90 & n5450 ) | ( x90 & ~n5455 ) | ( n5450 & ~n5455 ) ;
  assign n5457 = ( x90 & n5206 ) | ( x90 & ~n5301 ) | ( n5206 & ~n5301 ) ;
  assign n5458 = x90 & n5206 ;
  assign n5459 = ( n5211 & n5457 ) | ( n5211 & n5458 ) | ( n5457 & n5458 ) ;
  assign n5460 = ( ~n5211 & n5457 ) | ( ~n5211 & n5458 ) | ( n5457 & n5458 ) ;
  assign n5461 = ( n5211 & ~n5459 ) | ( n5211 & n5460 ) | ( ~n5459 & n5460 ) ;
  assign n5462 = ( x91 & n5456 ) | ( x91 & ~n5461 ) | ( n5456 & ~n5461 ) ;
  assign n5463 = ( x91 & n5212 ) | ( x91 & ~n5301 ) | ( n5212 & ~n5301 ) ;
  assign n5464 = x91 & n5212 ;
  assign n5465 = ( ~n5217 & n5463 ) | ( ~n5217 & n5464 ) | ( n5463 & n5464 ) ;
  assign n5466 = ( n5217 & n5463 ) | ( n5217 & n5464 ) | ( n5463 & n5464 ) ;
  assign n5467 = ( n5217 & n5465 ) | ( n5217 & ~n5466 ) | ( n5465 & ~n5466 ) ;
  assign n5468 = ( x92 & n5462 ) | ( x92 & ~n5467 ) | ( n5462 & ~n5467 ) ;
  assign n5469 = ( x92 & n5218 ) | ( x92 & ~n5301 ) | ( n5218 & ~n5301 ) ;
  assign n5470 = x92 & n5218 ;
  assign n5471 = ( n5223 & n5469 ) | ( n5223 & n5470 ) | ( n5469 & n5470 ) ;
  assign n5472 = ( ~n5223 & n5469 ) | ( ~n5223 & n5470 ) | ( n5469 & n5470 ) ;
  assign n5473 = ( n5223 & ~n5471 ) | ( n5223 & n5472 ) | ( ~n5471 & n5472 ) ;
  assign n5474 = ( x93 & n5468 ) | ( x93 & ~n5473 ) | ( n5468 & ~n5473 ) ;
  assign n5475 = ( x93 & n5224 ) | ( x93 & ~n5301 ) | ( n5224 & ~n5301 ) ;
  assign n5476 = x93 & n5224 ;
  assign n5477 = ( ~n5229 & n5475 ) | ( ~n5229 & n5476 ) | ( n5475 & n5476 ) ;
  assign n5478 = ( n5229 & n5475 ) | ( n5229 & n5476 ) | ( n5475 & n5476 ) ;
  assign n5479 = ( n5229 & n5477 ) | ( n5229 & ~n5478 ) | ( n5477 & ~n5478 ) ;
  assign n5480 = ( x94 & n5474 ) | ( x94 & ~n5479 ) | ( n5474 & ~n5479 ) ;
  assign n5481 = ( x94 & n5230 ) | ( x94 & ~n5301 ) | ( n5230 & ~n5301 ) ;
  assign n5482 = x94 & n5230 ;
  assign n5483 = ( n5235 & n5481 ) | ( n5235 & n5482 ) | ( n5481 & n5482 ) ;
  assign n5484 = ( ~n5235 & n5481 ) | ( ~n5235 & n5482 ) | ( n5481 & n5482 ) ;
  assign n5485 = ( n5235 & ~n5483 ) | ( n5235 & n5484 ) | ( ~n5483 & n5484 ) ;
  assign n5486 = ( x95 & n5480 ) | ( x95 & ~n5485 ) | ( n5480 & ~n5485 ) ;
  assign n5487 = ( x95 & n5236 ) | ( x95 & ~n5301 ) | ( n5236 & ~n5301 ) ;
  assign n5488 = x95 & n5236 ;
  assign n5489 = ( ~n5241 & n5487 ) | ( ~n5241 & n5488 ) | ( n5487 & n5488 ) ;
  assign n5490 = ( n5241 & n5487 ) | ( n5241 & n5488 ) | ( n5487 & n5488 ) ;
  assign n5491 = ( n5241 & n5489 ) | ( n5241 & ~n5490 ) | ( n5489 & ~n5490 ) ;
  assign n5492 = ( x96 & n5486 ) | ( x96 & ~n5491 ) | ( n5486 & ~n5491 ) ;
  assign n5493 = ( x96 & n5242 ) | ( x96 & ~n5301 ) | ( n5242 & ~n5301 ) ;
  assign n5494 = x96 & n5242 ;
  assign n5495 = ( n5247 & n5493 ) | ( n5247 & n5494 ) | ( n5493 & n5494 ) ;
  assign n5496 = ( ~n5247 & n5493 ) | ( ~n5247 & n5494 ) | ( n5493 & n5494 ) ;
  assign n5497 = ( n5247 & ~n5495 ) | ( n5247 & n5496 ) | ( ~n5495 & n5496 ) ;
  assign n5498 = ( x97 & n5492 ) | ( x97 & ~n5497 ) | ( n5492 & ~n5497 ) ;
  assign n5499 = ( x97 & n5248 ) | ( x97 & ~n5301 ) | ( n5248 & ~n5301 ) ;
  assign n5500 = x97 & n5248 ;
  assign n5501 = ( ~n5253 & n5499 ) | ( ~n5253 & n5500 ) | ( n5499 & n5500 ) ;
  assign n5502 = ( n5253 & n5499 ) | ( n5253 & n5500 ) | ( n5499 & n5500 ) ;
  assign n5503 = ( n5253 & n5501 ) | ( n5253 & ~n5502 ) | ( n5501 & ~n5502 ) ;
  assign n5504 = ( x98 & n5498 ) | ( x98 & ~n5503 ) | ( n5498 & ~n5503 ) ;
  assign n5505 = ( x98 & n5254 ) | ( x98 & ~n5301 ) | ( n5254 & ~n5301 ) ;
  assign n5506 = x98 & n5254 ;
  assign n5507 = ( n5259 & n5505 ) | ( n5259 & n5506 ) | ( n5505 & n5506 ) ;
  assign n5508 = ( ~n5259 & n5505 ) | ( ~n5259 & n5506 ) | ( n5505 & n5506 ) ;
  assign n5509 = ( n5259 & ~n5507 ) | ( n5259 & n5508 ) | ( ~n5507 & n5508 ) ;
  assign n5510 = ( x99 & n5504 ) | ( x99 & ~n5509 ) | ( n5504 & ~n5509 ) ;
  assign n5511 = ( x99 & n5260 ) | ( x99 & ~n5301 ) | ( n5260 & ~n5301 ) ;
  assign n5512 = x99 & n5260 ;
  assign n5513 = ( ~n5265 & n5511 ) | ( ~n5265 & n5512 ) | ( n5511 & n5512 ) ;
  assign n5514 = ( n5265 & n5511 ) | ( n5265 & n5512 ) | ( n5511 & n5512 ) ;
  assign n5515 = ( n5265 & n5513 ) | ( n5265 & ~n5514 ) | ( n5513 & ~n5514 ) ;
  assign n5516 = ( x100 & n5510 ) | ( x100 & ~n5515 ) | ( n5510 & ~n5515 ) ;
  assign n5517 = ( x100 & n5266 ) | ( x100 & ~n5301 ) | ( n5266 & ~n5301 ) ;
  assign n5518 = x100 & n5266 ;
  assign n5519 = ( n5271 & n5517 ) | ( n5271 & n5518 ) | ( n5517 & n5518 ) ;
  assign n5520 = ( ~n5271 & n5517 ) | ( ~n5271 & n5518 ) | ( n5517 & n5518 ) ;
  assign n5521 = ( n5271 & ~n5519 ) | ( n5271 & n5520 ) | ( ~n5519 & n5520 ) ;
  assign n5522 = ( x101 & n5516 ) | ( x101 & ~n5521 ) | ( n5516 & ~n5521 ) ;
  assign n5523 = ( x101 & n5272 ) | ( x101 & ~n5301 ) | ( n5272 & ~n5301 ) ;
  assign n5524 = x101 & n5272 ;
  assign n5525 = ( ~n5277 & n5523 ) | ( ~n5277 & n5524 ) | ( n5523 & n5524 ) ;
  assign n5526 = ( n5277 & n5523 ) | ( n5277 & n5524 ) | ( n5523 & n5524 ) ;
  assign n5527 = ( n5277 & n5525 ) | ( n5277 & ~n5526 ) | ( n5525 & ~n5526 ) ;
  assign n5528 = ( x102 & n5522 ) | ( x102 & ~n5527 ) | ( n5522 & ~n5527 ) ;
  assign n5529 = ( x102 & n5278 ) | ( x102 & ~n5301 ) | ( n5278 & ~n5301 ) ;
  assign n5530 = x102 & n5278 ;
  assign n5531 = ( n5283 & n5529 ) | ( n5283 & n5530 ) | ( n5529 & n5530 ) ;
  assign n5532 = ( ~n5283 & n5529 ) | ( ~n5283 & n5530 ) | ( n5529 & n5530 ) ;
  assign n5533 = ( n5283 & ~n5531 ) | ( n5283 & n5532 ) | ( ~n5531 & n5532 ) ;
  assign n5534 = ( x103 & n5528 ) | ( x103 & ~n5533 ) | ( n5528 & ~n5533 ) ;
  assign n5535 = ( x103 & n5284 ) | ( x103 & ~n5301 ) | ( n5284 & ~n5301 ) ;
  assign n5536 = x103 & n5284 ;
  assign n5537 = ( ~n5289 & n5535 ) | ( ~n5289 & n5536 ) | ( n5535 & n5536 ) ;
  assign n5538 = ( n5289 & n5535 ) | ( n5289 & n5536 ) | ( n5535 & n5536 ) ;
  assign n5539 = ( n5289 & n5537 ) | ( n5289 & ~n5538 ) | ( n5537 & ~n5538 ) ;
  assign n5540 = ( x104 & n5534 ) | ( x104 & ~n5539 ) | ( n5534 & ~n5539 ) ;
  assign n5541 = ( x104 & n5290 ) | ( x104 & ~n5301 ) | ( n5290 & ~n5301 ) ;
  assign n5542 = x104 & n5290 ;
  assign n5543 = ( ~n5295 & n5541 ) | ( ~n5295 & n5542 ) | ( n5541 & n5542 ) ;
  assign n5544 = ( n5295 & n5541 ) | ( n5295 & n5542 ) | ( n5541 & n5542 ) ;
  assign n5545 = ( n5295 & n5543 ) | ( n5295 & ~n5544 ) | ( n5543 & ~n5544 ) ;
  assign n5546 = ( x105 & n5540 ) | ( x105 & ~n5545 ) | ( n5540 & ~n5545 ) ;
  assign n5547 = x106 | n5546 ;
  assign n5548 = ( x106 & n151 ) | ( x106 & n5546 ) | ( n151 & n5546 ) ;
  assign n5549 = ( n5299 & ~n5547 ) | ( n5299 & n5548 ) | ( ~n5547 & n5548 ) ;
  assign n5550 = ( x106 & ~n5299 ) | ( x106 & n5546 ) | ( ~n5299 & n5546 ) ;
  assign n5551 = n151 | n5550 ;
  assign n5552 = ( x21 & ~x64 ) | ( x21 & n5551 ) | ( ~x64 & n5551 ) ;
  assign n5553 = ~x21 & n5551 ;
  assign n5554 = ( n5305 & n5552 ) | ( n5305 & ~n5553 ) | ( n5552 & ~n5553 ) ;
  assign n5555 = ~x20 & x64 ;
  assign n5556 = ( x65 & ~n5554 ) | ( x65 & n5555 ) | ( ~n5554 & n5555 ) ;
  assign n5557 = ( x65 & n5305 ) | ( x65 & ~n5551 ) | ( n5305 & ~n5551 ) ;
  assign n5558 = x65 & n5305 ;
  assign n5559 = ( n5304 & n5557 ) | ( n5304 & n5558 ) | ( n5557 & n5558 ) ;
  assign n5560 = ( ~n5304 & n5557 ) | ( ~n5304 & n5558 ) | ( n5557 & n5558 ) ;
  assign n5561 = ( n5304 & ~n5559 ) | ( n5304 & n5560 ) | ( ~n5559 & n5560 ) ;
  assign n5562 = ( x66 & n5556 ) | ( x66 & ~n5561 ) | ( n5556 & ~n5561 ) ;
  assign n5563 = ( x66 & n5306 ) | ( x66 & ~n5551 ) | ( n5306 & ~n5551 ) ;
  assign n5564 = x66 & n5306 ;
  assign n5565 = ( n5311 & n5563 ) | ( n5311 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5566 = ( ~n5311 & n5563 ) | ( ~n5311 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5567 = ( n5311 & ~n5565 ) | ( n5311 & n5566 ) | ( ~n5565 & n5566 ) ;
  assign n5568 = ( x67 & n5562 ) | ( x67 & ~n5567 ) | ( n5562 & ~n5567 ) ;
  assign n5569 = ( x67 & n5312 ) | ( x67 & ~n5551 ) | ( n5312 & ~n5551 ) ;
  assign n5570 = x67 & n5312 ;
  assign n5571 = ( ~n5317 & n5569 ) | ( ~n5317 & n5570 ) | ( n5569 & n5570 ) ;
  assign n5572 = ( n5317 & n5569 ) | ( n5317 & n5570 ) | ( n5569 & n5570 ) ;
  assign n5573 = ( n5317 & n5571 ) | ( n5317 & ~n5572 ) | ( n5571 & ~n5572 ) ;
  assign n5574 = ( x68 & n5568 ) | ( x68 & ~n5573 ) | ( n5568 & ~n5573 ) ;
  assign n5575 = ( x68 & n5318 ) | ( x68 & ~n5551 ) | ( n5318 & ~n5551 ) ;
  assign n5576 = x68 & n5318 ;
  assign n5577 = ( n5323 & n5575 ) | ( n5323 & n5576 ) | ( n5575 & n5576 ) ;
  assign n5578 = ( ~n5323 & n5575 ) | ( ~n5323 & n5576 ) | ( n5575 & n5576 ) ;
  assign n5579 = ( n5323 & ~n5577 ) | ( n5323 & n5578 ) | ( ~n5577 & n5578 ) ;
  assign n5580 = ( x69 & n5574 ) | ( x69 & ~n5579 ) | ( n5574 & ~n5579 ) ;
  assign n5581 = ( x69 & n5324 ) | ( x69 & ~n5551 ) | ( n5324 & ~n5551 ) ;
  assign n5582 = x69 & n5324 ;
  assign n5583 = ( ~n5329 & n5581 ) | ( ~n5329 & n5582 ) | ( n5581 & n5582 ) ;
  assign n5584 = ( n5329 & n5581 ) | ( n5329 & n5582 ) | ( n5581 & n5582 ) ;
  assign n5585 = ( n5329 & n5583 ) | ( n5329 & ~n5584 ) | ( n5583 & ~n5584 ) ;
  assign n5586 = ( x70 & n5580 ) | ( x70 & ~n5585 ) | ( n5580 & ~n5585 ) ;
  assign n5587 = ( x70 & n5330 ) | ( x70 & ~n5551 ) | ( n5330 & ~n5551 ) ;
  assign n5588 = x70 & n5330 ;
  assign n5589 = ( n5335 & n5587 ) | ( n5335 & n5588 ) | ( n5587 & n5588 ) ;
  assign n5590 = ( ~n5335 & n5587 ) | ( ~n5335 & n5588 ) | ( n5587 & n5588 ) ;
  assign n5591 = ( n5335 & ~n5589 ) | ( n5335 & n5590 ) | ( ~n5589 & n5590 ) ;
  assign n5592 = ( x71 & n5586 ) | ( x71 & ~n5591 ) | ( n5586 & ~n5591 ) ;
  assign n5593 = ( x71 & n5336 ) | ( x71 & ~n5551 ) | ( n5336 & ~n5551 ) ;
  assign n5594 = x71 & n5336 ;
  assign n5595 = ( ~n5341 & n5593 ) | ( ~n5341 & n5594 ) | ( n5593 & n5594 ) ;
  assign n5596 = ( n5341 & n5593 ) | ( n5341 & n5594 ) | ( n5593 & n5594 ) ;
  assign n5597 = ( n5341 & n5595 ) | ( n5341 & ~n5596 ) | ( n5595 & ~n5596 ) ;
  assign n5598 = ( x72 & n5592 ) | ( x72 & ~n5597 ) | ( n5592 & ~n5597 ) ;
  assign n5599 = ( x72 & n5342 ) | ( x72 & ~n5551 ) | ( n5342 & ~n5551 ) ;
  assign n5600 = x72 & n5342 ;
  assign n5601 = ( n5347 & n5599 ) | ( n5347 & n5600 ) | ( n5599 & n5600 ) ;
  assign n5602 = ( ~n5347 & n5599 ) | ( ~n5347 & n5600 ) | ( n5599 & n5600 ) ;
  assign n5603 = ( n5347 & ~n5601 ) | ( n5347 & n5602 ) | ( ~n5601 & n5602 ) ;
  assign n5604 = ( x73 & n5598 ) | ( x73 & ~n5603 ) | ( n5598 & ~n5603 ) ;
  assign n5605 = ( x73 & n5348 ) | ( x73 & ~n5551 ) | ( n5348 & ~n5551 ) ;
  assign n5606 = x73 & n5348 ;
  assign n5607 = ( ~n5353 & n5605 ) | ( ~n5353 & n5606 ) | ( n5605 & n5606 ) ;
  assign n5608 = ( n5353 & n5605 ) | ( n5353 & n5606 ) | ( n5605 & n5606 ) ;
  assign n5609 = ( n5353 & n5607 ) | ( n5353 & ~n5608 ) | ( n5607 & ~n5608 ) ;
  assign n5610 = ( x74 & n5604 ) | ( x74 & ~n5609 ) | ( n5604 & ~n5609 ) ;
  assign n5611 = ( x74 & n5354 ) | ( x74 & ~n5551 ) | ( n5354 & ~n5551 ) ;
  assign n5612 = x74 & n5354 ;
  assign n5613 = ( n5359 & n5611 ) | ( n5359 & n5612 ) | ( n5611 & n5612 ) ;
  assign n5614 = ( ~n5359 & n5611 ) | ( ~n5359 & n5612 ) | ( n5611 & n5612 ) ;
  assign n5615 = ( n5359 & ~n5613 ) | ( n5359 & n5614 ) | ( ~n5613 & n5614 ) ;
  assign n5616 = ( x75 & n5610 ) | ( x75 & ~n5615 ) | ( n5610 & ~n5615 ) ;
  assign n5617 = ( x75 & n5360 ) | ( x75 & ~n5551 ) | ( n5360 & ~n5551 ) ;
  assign n5618 = x75 & n5360 ;
  assign n5619 = ( ~n5365 & n5617 ) | ( ~n5365 & n5618 ) | ( n5617 & n5618 ) ;
  assign n5620 = ( n5365 & n5617 ) | ( n5365 & n5618 ) | ( n5617 & n5618 ) ;
  assign n5621 = ( n5365 & n5619 ) | ( n5365 & ~n5620 ) | ( n5619 & ~n5620 ) ;
  assign n5622 = ( x76 & n5616 ) | ( x76 & ~n5621 ) | ( n5616 & ~n5621 ) ;
  assign n5623 = ( x76 & n5366 ) | ( x76 & ~n5551 ) | ( n5366 & ~n5551 ) ;
  assign n5624 = x76 & n5366 ;
  assign n5625 = ( n5371 & n5623 ) | ( n5371 & n5624 ) | ( n5623 & n5624 ) ;
  assign n5626 = ( ~n5371 & n5623 ) | ( ~n5371 & n5624 ) | ( n5623 & n5624 ) ;
  assign n5627 = ( n5371 & ~n5625 ) | ( n5371 & n5626 ) | ( ~n5625 & n5626 ) ;
  assign n5628 = ( x77 & n5622 ) | ( x77 & ~n5627 ) | ( n5622 & ~n5627 ) ;
  assign n5629 = ( x77 & n5372 ) | ( x77 & ~n5551 ) | ( n5372 & ~n5551 ) ;
  assign n5630 = x77 & n5372 ;
  assign n5631 = ( ~n5377 & n5629 ) | ( ~n5377 & n5630 ) | ( n5629 & n5630 ) ;
  assign n5632 = ( n5377 & n5629 ) | ( n5377 & n5630 ) | ( n5629 & n5630 ) ;
  assign n5633 = ( n5377 & n5631 ) | ( n5377 & ~n5632 ) | ( n5631 & ~n5632 ) ;
  assign n5634 = ( x78 & n5628 ) | ( x78 & ~n5633 ) | ( n5628 & ~n5633 ) ;
  assign n5635 = ( x78 & n5378 ) | ( x78 & ~n5551 ) | ( n5378 & ~n5551 ) ;
  assign n5636 = x78 & n5378 ;
  assign n5637 = ( n5383 & n5635 ) | ( n5383 & n5636 ) | ( n5635 & n5636 ) ;
  assign n5638 = ( ~n5383 & n5635 ) | ( ~n5383 & n5636 ) | ( n5635 & n5636 ) ;
  assign n5639 = ( n5383 & ~n5637 ) | ( n5383 & n5638 ) | ( ~n5637 & n5638 ) ;
  assign n5640 = ( x79 & n5634 ) | ( x79 & ~n5639 ) | ( n5634 & ~n5639 ) ;
  assign n5641 = ( x79 & n5384 ) | ( x79 & ~n5551 ) | ( n5384 & ~n5551 ) ;
  assign n5642 = x79 & n5384 ;
  assign n5643 = ( ~n5389 & n5641 ) | ( ~n5389 & n5642 ) | ( n5641 & n5642 ) ;
  assign n5644 = ( n5389 & n5641 ) | ( n5389 & n5642 ) | ( n5641 & n5642 ) ;
  assign n5645 = ( n5389 & n5643 ) | ( n5389 & ~n5644 ) | ( n5643 & ~n5644 ) ;
  assign n5646 = ( x80 & n5640 ) | ( x80 & ~n5645 ) | ( n5640 & ~n5645 ) ;
  assign n5647 = ( x80 & n5390 ) | ( x80 & ~n5551 ) | ( n5390 & ~n5551 ) ;
  assign n5648 = x80 & n5390 ;
  assign n5649 = ( n5395 & n5647 ) | ( n5395 & n5648 ) | ( n5647 & n5648 ) ;
  assign n5650 = ( ~n5395 & n5647 ) | ( ~n5395 & n5648 ) | ( n5647 & n5648 ) ;
  assign n5651 = ( n5395 & ~n5649 ) | ( n5395 & n5650 ) | ( ~n5649 & n5650 ) ;
  assign n5652 = ( x81 & n5646 ) | ( x81 & ~n5651 ) | ( n5646 & ~n5651 ) ;
  assign n5653 = ( x81 & n5396 ) | ( x81 & ~n5551 ) | ( n5396 & ~n5551 ) ;
  assign n5654 = x81 & n5396 ;
  assign n5655 = ( ~n5401 & n5653 ) | ( ~n5401 & n5654 ) | ( n5653 & n5654 ) ;
  assign n5656 = ( n5401 & n5653 ) | ( n5401 & n5654 ) | ( n5653 & n5654 ) ;
  assign n5657 = ( n5401 & n5655 ) | ( n5401 & ~n5656 ) | ( n5655 & ~n5656 ) ;
  assign n5658 = ( x82 & n5652 ) | ( x82 & ~n5657 ) | ( n5652 & ~n5657 ) ;
  assign n5659 = ( x82 & n5402 ) | ( x82 & ~n5551 ) | ( n5402 & ~n5551 ) ;
  assign n5660 = x82 & n5402 ;
  assign n5661 = ( n5407 & n5659 ) | ( n5407 & n5660 ) | ( n5659 & n5660 ) ;
  assign n5662 = ( ~n5407 & n5659 ) | ( ~n5407 & n5660 ) | ( n5659 & n5660 ) ;
  assign n5663 = ( n5407 & ~n5661 ) | ( n5407 & n5662 ) | ( ~n5661 & n5662 ) ;
  assign n5664 = ( x83 & n5658 ) | ( x83 & ~n5663 ) | ( n5658 & ~n5663 ) ;
  assign n5665 = ( x83 & n5408 ) | ( x83 & ~n5551 ) | ( n5408 & ~n5551 ) ;
  assign n5666 = x83 & n5408 ;
  assign n5667 = ( ~n5413 & n5665 ) | ( ~n5413 & n5666 ) | ( n5665 & n5666 ) ;
  assign n5668 = ( n5413 & n5665 ) | ( n5413 & n5666 ) | ( n5665 & n5666 ) ;
  assign n5669 = ( n5413 & n5667 ) | ( n5413 & ~n5668 ) | ( n5667 & ~n5668 ) ;
  assign n5670 = ( x84 & n5664 ) | ( x84 & ~n5669 ) | ( n5664 & ~n5669 ) ;
  assign n5671 = ( x84 & n5414 ) | ( x84 & ~n5551 ) | ( n5414 & ~n5551 ) ;
  assign n5672 = x84 & n5414 ;
  assign n5673 = ( n5419 & n5671 ) | ( n5419 & n5672 ) | ( n5671 & n5672 ) ;
  assign n5674 = ( ~n5419 & n5671 ) | ( ~n5419 & n5672 ) | ( n5671 & n5672 ) ;
  assign n5675 = ( n5419 & ~n5673 ) | ( n5419 & n5674 ) | ( ~n5673 & n5674 ) ;
  assign n5676 = ( x85 & n5670 ) | ( x85 & ~n5675 ) | ( n5670 & ~n5675 ) ;
  assign n5677 = ( x85 & n5420 ) | ( x85 & ~n5551 ) | ( n5420 & ~n5551 ) ;
  assign n5678 = x85 & n5420 ;
  assign n5679 = ( ~n5425 & n5677 ) | ( ~n5425 & n5678 ) | ( n5677 & n5678 ) ;
  assign n5680 = ( n5425 & n5677 ) | ( n5425 & n5678 ) | ( n5677 & n5678 ) ;
  assign n5681 = ( n5425 & n5679 ) | ( n5425 & ~n5680 ) | ( n5679 & ~n5680 ) ;
  assign n5682 = ( x86 & n5676 ) | ( x86 & ~n5681 ) | ( n5676 & ~n5681 ) ;
  assign n5683 = ( x86 & n5426 ) | ( x86 & ~n5551 ) | ( n5426 & ~n5551 ) ;
  assign n5684 = x86 & n5426 ;
  assign n5685 = ( n5431 & n5683 ) | ( n5431 & n5684 ) | ( n5683 & n5684 ) ;
  assign n5686 = ( ~n5431 & n5683 ) | ( ~n5431 & n5684 ) | ( n5683 & n5684 ) ;
  assign n5687 = ( n5431 & ~n5685 ) | ( n5431 & n5686 ) | ( ~n5685 & n5686 ) ;
  assign n5688 = ( x87 & n5682 ) | ( x87 & ~n5687 ) | ( n5682 & ~n5687 ) ;
  assign n5689 = ( x87 & n5432 ) | ( x87 & ~n5551 ) | ( n5432 & ~n5551 ) ;
  assign n5690 = x87 & n5432 ;
  assign n5691 = ( ~n5437 & n5689 ) | ( ~n5437 & n5690 ) | ( n5689 & n5690 ) ;
  assign n5692 = ( n5437 & n5689 ) | ( n5437 & n5690 ) | ( n5689 & n5690 ) ;
  assign n5693 = ( n5437 & n5691 ) | ( n5437 & ~n5692 ) | ( n5691 & ~n5692 ) ;
  assign n5694 = ( x88 & n5688 ) | ( x88 & ~n5693 ) | ( n5688 & ~n5693 ) ;
  assign n5695 = ( x88 & n5438 ) | ( x88 & ~n5551 ) | ( n5438 & ~n5551 ) ;
  assign n5696 = x88 & n5438 ;
  assign n5697 = ( n5443 & n5695 ) | ( n5443 & n5696 ) | ( n5695 & n5696 ) ;
  assign n5698 = ( ~n5443 & n5695 ) | ( ~n5443 & n5696 ) | ( n5695 & n5696 ) ;
  assign n5699 = ( n5443 & ~n5697 ) | ( n5443 & n5698 ) | ( ~n5697 & n5698 ) ;
  assign n5700 = ( x89 & n5694 ) | ( x89 & ~n5699 ) | ( n5694 & ~n5699 ) ;
  assign n5701 = ( x89 & n5444 ) | ( x89 & ~n5551 ) | ( n5444 & ~n5551 ) ;
  assign n5702 = x89 & n5444 ;
  assign n5703 = ( ~n5449 & n5701 ) | ( ~n5449 & n5702 ) | ( n5701 & n5702 ) ;
  assign n5704 = ( n5449 & n5701 ) | ( n5449 & n5702 ) | ( n5701 & n5702 ) ;
  assign n5705 = ( n5449 & n5703 ) | ( n5449 & ~n5704 ) | ( n5703 & ~n5704 ) ;
  assign n5706 = ( x90 & n5700 ) | ( x90 & ~n5705 ) | ( n5700 & ~n5705 ) ;
  assign n5707 = ( x90 & n5450 ) | ( x90 & ~n5551 ) | ( n5450 & ~n5551 ) ;
  assign n5708 = x90 & n5450 ;
  assign n5709 = ( n5455 & n5707 ) | ( n5455 & n5708 ) | ( n5707 & n5708 ) ;
  assign n5710 = ( ~n5455 & n5707 ) | ( ~n5455 & n5708 ) | ( n5707 & n5708 ) ;
  assign n5711 = ( n5455 & ~n5709 ) | ( n5455 & n5710 ) | ( ~n5709 & n5710 ) ;
  assign n5712 = ( x91 & n5706 ) | ( x91 & ~n5711 ) | ( n5706 & ~n5711 ) ;
  assign n5713 = ( x91 & n5456 ) | ( x91 & ~n5551 ) | ( n5456 & ~n5551 ) ;
  assign n5714 = x91 & n5456 ;
  assign n5715 = ( ~n5461 & n5713 ) | ( ~n5461 & n5714 ) | ( n5713 & n5714 ) ;
  assign n5716 = ( n5461 & n5713 ) | ( n5461 & n5714 ) | ( n5713 & n5714 ) ;
  assign n5717 = ( n5461 & n5715 ) | ( n5461 & ~n5716 ) | ( n5715 & ~n5716 ) ;
  assign n5718 = ( x92 & n5712 ) | ( x92 & ~n5717 ) | ( n5712 & ~n5717 ) ;
  assign n5719 = ( x92 & n5462 ) | ( x92 & ~n5551 ) | ( n5462 & ~n5551 ) ;
  assign n5720 = x92 & n5462 ;
  assign n5721 = ( n5467 & n5719 ) | ( n5467 & n5720 ) | ( n5719 & n5720 ) ;
  assign n5722 = ( ~n5467 & n5719 ) | ( ~n5467 & n5720 ) | ( n5719 & n5720 ) ;
  assign n5723 = ( n5467 & ~n5721 ) | ( n5467 & n5722 ) | ( ~n5721 & n5722 ) ;
  assign n5724 = ( x93 & n5718 ) | ( x93 & ~n5723 ) | ( n5718 & ~n5723 ) ;
  assign n5725 = ( x93 & n5468 ) | ( x93 & ~n5551 ) | ( n5468 & ~n5551 ) ;
  assign n5726 = x93 & n5468 ;
  assign n5727 = ( ~n5473 & n5725 ) | ( ~n5473 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5728 = ( n5473 & n5725 ) | ( n5473 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5729 = ( n5473 & n5727 ) | ( n5473 & ~n5728 ) | ( n5727 & ~n5728 ) ;
  assign n5730 = ( x94 & n5724 ) | ( x94 & ~n5729 ) | ( n5724 & ~n5729 ) ;
  assign n5731 = ( x94 & n5474 ) | ( x94 & ~n5551 ) | ( n5474 & ~n5551 ) ;
  assign n5732 = x94 & n5474 ;
  assign n5733 = ( n5479 & n5731 ) | ( n5479 & n5732 ) | ( n5731 & n5732 ) ;
  assign n5734 = ( ~n5479 & n5731 ) | ( ~n5479 & n5732 ) | ( n5731 & n5732 ) ;
  assign n5735 = ( n5479 & ~n5733 ) | ( n5479 & n5734 ) | ( ~n5733 & n5734 ) ;
  assign n5736 = ( x95 & n5730 ) | ( x95 & ~n5735 ) | ( n5730 & ~n5735 ) ;
  assign n5737 = ( x95 & n5480 ) | ( x95 & ~n5551 ) | ( n5480 & ~n5551 ) ;
  assign n5738 = x95 & n5480 ;
  assign n5739 = ( ~n5485 & n5737 ) | ( ~n5485 & n5738 ) | ( n5737 & n5738 ) ;
  assign n5740 = ( n5485 & n5737 ) | ( n5485 & n5738 ) | ( n5737 & n5738 ) ;
  assign n5741 = ( n5485 & n5739 ) | ( n5485 & ~n5740 ) | ( n5739 & ~n5740 ) ;
  assign n5742 = ( x96 & n5736 ) | ( x96 & ~n5741 ) | ( n5736 & ~n5741 ) ;
  assign n5743 = ( x96 & n5486 ) | ( x96 & ~n5551 ) | ( n5486 & ~n5551 ) ;
  assign n5744 = x96 & n5486 ;
  assign n5745 = ( n5491 & n5743 ) | ( n5491 & n5744 ) | ( n5743 & n5744 ) ;
  assign n5746 = ( ~n5491 & n5743 ) | ( ~n5491 & n5744 ) | ( n5743 & n5744 ) ;
  assign n5747 = ( n5491 & ~n5745 ) | ( n5491 & n5746 ) | ( ~n5745 & n5746 ) ;
  assign n5748 = ( x97 & n5742 ) | ( x97 & ~n5747 ) | ( n5742 & ~n5747 ) ;
  assign n5749 = ( x97 & n5492 ) | ( x97 & ~n5551 ) | ( n5492 & ~n5551 ) ;
  assign n5750 = x97 & n5492 ;
  assign n5751 = ( ~n5497 & n5749 ) | ( ~n5497 & n5750 ) | ( n5749 & n5750 ) ;
  assign n5752 = ( n5497 & n5749 ) | ( n5497 & n5750 ) | ( n5749 & n5750 ) ;
  assign n5753 = ( n5497 & n5751 ) | ( n5497 & ~n5752 ) | ( n5751 & ~n5752 ) ;
  assign n5754 = ( x98 & n5748 ) | ( x98 & ~n5753 ) | ( n5748 & ~n5753 ) ;
  assign n5755 = ( x98 & n5498 ) | ( x98 & ~n5551 ) | ( n5498 & ~n5551 ) ;
  assign n5756 = x98 & n5498 ;
  assign n5757 = ( n5503 & n5755 ) | ( n5503 & n5756 ) | ( n5755 & n5756 ) ;
  assign n5758 = ( ~n5503 & n5755 ) | ( ~n5503 & n5756 ) | ( n5755 & n5756 ) ;
  assign n5759 = ( n5503 & ~n5757 ) | ( n5503 & n5758 ) | ( ~n5757 & n5758 ) ;
  assign n5760 = ( x99 & n5754 ) | ( x99 & ~n5759 ) | ( n5754 & ~n5759 ) ;
  assign n5761 = ( x99 & n5504 ) | ( x99 & ~n5551 ) | ( n5504 & ~n5551 ) ;
  assign n5762 = x99 & n5504 ;
  assign n5763 = ( ~n5509 & n5761 ) | ( ~n5509 & n5762 ) | ( n5761 & n5762 ) ;
  assign n5764 = ( n5509 & n5761 ) | ( n5509 & n5762 ) | ( n5761 & n5762 ) ;
  assign n5765 = ( n5509 & n5763 ) | ( n5509 & ~n5764 ) | ( n5763 & ~n5764 ) ;
  assign n5766 = ( x100 & n5760 ) | ( x100 & ~n5765 ) | ( n5760 & ~n5765 ) ;
  assign n5767 = ( x100 & n5510 ) | ( x100 & ~n5551 ) | ( n5510 & ~n5551 ) ;
  assign n5768 = x100 & n5510 ;
  assign n5769 = ( n5515 & n5767 ) | ( n5515 & n5768 ) | ( n5767 & n5768 ) ;
  assign n5770 = ( ~n5515 & n5767 ) | ( ~n5515 & n5768 ) | ( n5767 & n5768 ) ;
  assign n5771 = ( n5515 & ~n5769 ) | ( n5515 & n5770 ) | ( ~n5769 & n5770 ) ;
  assign n5772 = ( x101 & n5766 ) | ( x101 & ~n5771 ) | ( n5766 & ~n5771 ) ;
  assign n5773 = ( x101 & n5516 ) | ( x101 & ~n5551 ) | ( n5516 & ~n5551 ) ;
  assign n5774 = x101 & n5516 ;
  assign n5775 = ( ~n5521 & n5773 ) | ( ~n5521 & n5774 ) | ( n5773 & n5774 ) ;
  assign n5776 = ( n5521 & n5773 ) | ( n5521 & n5774 ) | ( n5773 & n5774 ) ;
  assign n5777 = ( n5521 & n5775 ) | ( n5521 & ~n5776 ) | ( n5775 & ~n5776 ) ;
  assign n5778 = ( x102 & n5772 ) | ( x102 & ~n5777 ) | ( n5772 & ~n5777 ) ;
  assign n5779 = ( x102 & n5522 ) | ( x102 & ~n5551 ) | ( n5522 & ~n5551 ) ;
  assign n5780 = x102 & n5522 ;
  assign n5781 = ( n5527 & n5779 ) | ( n5527 & n5780 ) | ( n5779 & n5780 ) ;
  assign n5782 = ( ~n5527 & n5779 ) | ( ~n5527 & n5780 ) | ( n5779 & n5780 ) ;
  assign n5783 = ( n5527 & ~n5781 ) | ( n5527 & n5782 ) | ( ~n5781 & n5782 ) ;
  assign n5784 = ( x103 & n5778 ) | ( x103 & ~n5783 ) | ( n5778 & ~n5783 ) ;
  assign n5785 = ( x103 & n5528 ) | ( x103 & ~n5551 ) | ( n5528 & ~n5551 ) ;
  assign n5786 = x103 & n5528 ;
  assign n5787 = ( ~n5533 & n5785 ) | ( ~n5533 & n5786 ) | ( n5785 & n5786 ) ;
  assign n5788 = ( n5533 & n5785 ) | ( n5533 & n5786 ) | ( n5785 & n5786 ) ;
  assign n5789 = ( n5533 & n5787 ) | ( n5533 & ~n5788 ) | ( n5787 & ~n5788 ) ;
  assign n5790 = ( x104 & n5784 ) | ( x104 & ~n5789 ) | ( n5784 & ~n5789 ) ;
  assign n5791 = ( x104 & n5534 ) | ( x104 & ~n5551 ) | ( n5534 & ~n5551 ) ;
  assign n5792 = x104 & n5534 ;
  assign n5793 = ( n5539 & n5791 ) | ( n5539 & n5792 ) | ( n5791 & n5792 ) ;
  assign n5794 = ( ~n5539 & n5791 ) | ( ~n5539 & n5792 ) | ( n5791 & n5792 ) ;
  assign n5795 = ( n5539 & ~n5793 ) | ( n5539 & n5794 ) | ( ~n5793 & n5794 ) ;
  assign n5796 = ( x105 & n5790 ) | ( x105 & ~n5795 ) | ( n5790 & ~n5795 ) ;
  assign n5797 = ( x105 & n5540 ) | ( x105 & ~n5551 ) | ( n5540 & ~n5551 ) ;
  assign n5798 = x105 & n5540 ;
  assign n5799 = ( n5545 & n5797 ) | ( n5545 & n5798 ) | ( n5797 & n5798 ) ;
  assign n5800 = ( ~n5545 & n5797 ) | ( ~n5545 & n5798 ) | ( n5797 & n5798 ) ;
  assign n5801 = ( n5545 & ~n5799 ) | ( n5545 & n5800 ) | ( ~n5799 & n5800 ) ;
  assign n5802 = ( x106 & n5796 ) | ( x106 & ~n5801 ) | ( n5796 & ~n5801 ) ;
  assign n5803 = x107 | n5802 ;
  assign n5804 = ( x107 & n150 ) | ( x107 & n5802 ) | ( n150 & n5802 ) ;
  assign n5805 = ( n5549 & ~n5803 ) | ( n5549 & n5804 ) | ( ~n5803 & n5804 ) ;
  assign n5806 = ( x107 & ~n5549 ) | ( x107 & n5802 ) | ( ~n5549 & n5802 ) ;
  assign n5807 = n150 | n5806 ;
  assign n5808 = ( x20 & ~x64 ) | ( x20 & n5807 ) | ( ~x64 & n5807 ) ;
  assign n5809 = ~x20 & n5807 ;
  assign n5810 = ( n5555 & n5808 ) | ( n5555 & ~n5809 ) | ( n5808 & ~n5809 ) ;
  assign n5811 = ~x19 & x64 ;
  assign n5812 = ( x65 & ~n5810 ) | ( x65 & n5811 ) | ( ~n5810 & n5811 ) ;
  assign n5813 = ( x65 & n5555 ) | ( x65 & ~n5807 ) | ( n5555 & ~n5807 ) ;
  assign n5814 = x65 & n5555 ;
  assign n5815 = ( n5554 & n5813 ) | ( n5554 & n5814 ) | ( n5813 & n5814 ) ;
  assign n5816 = ( ~n5554 & n5813 ) | ( ~n5554 & n5814 ) | ( n5813 & n5814 ) ;
  assign n5817 = ( n5554 & ~n5815 ) | ( n5554 & n5816 ) | ( ~n5815 & n5816 ) ;
  assign n5818 = ( x66 & n5812 ) | ( x66 & ~n5817 ) | ( n5812 & ~n5817 ) ;
  assign n5819 = ( x66 & n5556 ) | ( x66 & ~n5807 ) | ( n5556 & ~n5807 ) ;
  assign n5820 = x66 & n5556 ;
  assign n5821 = ( n5561 & n5819 ) | ( n5561 & n5820 ) | ( n5819 & n5820 ) ;
  assign n5822 = ( ~n5561 & n5819 ) | ( ~n5561 & n5820 ) | ( n5819 & n5820 ) ;
  assign n5823 = ( n5561 & ~n5821 ) | ( n5561 & n5822 ) | ( ~n5821 & n5822 ) ;
  assign n5824 = ( x67 & n5818 ) | ( x67 & ~n5823 ) | ( n5818 & ~n5823 ) ;
  assign n5825 = ( x67 & n5562 ) | ( x67 & ~n5807 ) | ( n5562 & ~n5807 ) ;
  assign n5826 = x67 & n5562 ;
  assign n5827 = ( ~n5567 & n5825 ) | ( ~n5567 & n5826 ) | ( n5825 & n5826 ) ;
  assign n5828 = ( n5567 & n5825 ) | ( n5567 & n5826 ) | ( n5825 & n5826 ) ;
  assign n5829 = ( n5567 & n5827 ) | ( n5567 & ~n5828 ) | ( n5827 & ~n5828 ) ;
  assign n5830 = ( x68 & n5824 ) | ( x68 & ~n5829 ) | ( n5824 & ~n5829 ) ;
  assign n5831 = ( x68 & n5568 ) | ( x68 & ~n5807 ) | ( n5568 & ~n5807 ) ;
  assign n5832 = x68 & n5568 ;
  assign n5833 = ( n5573 & n5831 ) | ( n5573 & n5832 ) | ( n5831 & n5832 ) ;
  assign n5834 = ( ~n5573 & n5831 ) | ( ~n5573 & n5832 ) | ( n5831 & n5832 ) ;
  assign n5835 = ( n5573 & ~n5833 ) | ( n5573 & n5834 ) | ( ~n5833 & n5834 ) ;
  assign n5836 = ( x69 & n5830 ) | ( x69 & ~n5835 ) | ( n5830 & ~n5835 ) ;
  assign n5837 = ( x69 & n5574 ) | ( x69 & ~n5807 ) | ( n5574 & ~n5807 ) ;
  assign n5838 = x69 & n5574 ;
  assign n5839 = ( ~n5579 & n5837 ) | ( ~n5579 & n5838 ) | ( n5837 & n5838 ) ;
  assign n5840 = ( n5579 & n5837 ) | ( n5579 & n5838 ) | ( n5837 & n5838 ) ;
  assign n5841 = ( n5579 & n5839 ) | ( n5579 & ~n5840 ) | ( n5839 & ~n5840 ) ;
  assign n5842 = ( x70 & n5836 ) | ( x70 & ~n5841 ) | ( n5836 & ~n5841 ) ;
  assign n5843 = ( x70 & n5580 ) | ( x70 & ~n5807 ) | ( n5580 & ~n5807 ) ;
  assign n5844 = x70 & n5580 ;
  assign n5845 = ( n5585 & n5843 ) | ( n5585 & n5844 ) | ( n5843 & n5844 ) ;
  assign n5846 = ( ~n5585 & n5843 ) | ( ~n5585 & n5844 ) | ( n5843 & n5844 ) ;
  assign n5847 = ( n5585 & ~n5845 ) | ( n5585 & n5846 ) | ( ~n5845 & n5846 ) ;
  assign n5848 = ( x71 & n5842 ) | ( x71 & ~n5847 ) | ( n5842 & ~n5847 ) ;
  assign n5849 = ( x71 & n5586 ) | ( x71 & ~n5807 ) | ( n5586 & ~n5807 ) ;
  assign n5850 = x71 & n5586 ;
  assign n5851 = ( ~n5591 & n5849 ) | ( ~n5591 & n5850 ) | ( n5849 & n5850 ) ;
  assign n5852 = ( n5591 & n5849 ) | ( n5591 & n5850 ) | ( n5849 & n5850 ) ;
  assign n5853 = ( n5591 & n5851 ) | ( n5591 & ~n5852 ) | ( n5851 & ~n5852 ) ;
  assign n5854 = ( x72 & n5848 ) | ( x72 & ~n5853 ) | ( n5848 & ~n5853 ) ;
  assign n5855 = ( x72 & n5592 ) | ( x72 & ~n5807 ) | ( n5592 & ~n5807 ) ;
  assign n5856 = x72 & n5592 ;
  assign n5857 = ( n5597 & n5855 ) | ( n5597 & n5856 ) | ( n5855 & n5856 ) ;
  assign n5858 = ( ~n5597 & n5855 ) | ( ~n5597 & n5856 ) | ( n5855 & n5856 ) ;
  assign n5859 = ( n5597 & ~n5857 ) | ( n5597 & n5858 ) | ( ~n5857 & n5858 ) ;
  assign n5860 = ( x73 & n5854 ) | ( x73 & ~n5859 ) | ( n5854 & ~n5859 ) ;
  assign n5861 = ( x73 & n5598 ) | ( x73 & ~n5807 ) | ( n5598 & ~n5807 ) ;
  assign n5862 = x73 & n5598 ;
  assign n5863 = ( ~n5603 & n5861 ) | ( ~n5603 & n5862 ) | ( n5861 & n5862 ) ;
  assign n5864 = ( n5603 & n5861 ) | ( n5603 & n5862 ) | ( n5861 & n5862 ) ;
  assign n5865 = ( n5603 & n5863 ) | ( n5603 & ~n5864 ) | ( n5863 & ~n5864 ) ;
  assign n5866 = ( x74 & n5860 ) | ( x74 & ~n5865 ) | ( n5860 & ~n5865 ) ;
  assign n5867 = ( x74 & n5604 ) | ( x74 & ~n5807 ) | ( n5604 & ~n5807 ) ;
  assign n5868 = x74 & n5604 ;
  assign n5869 = ( n5609 & n5867 ) | ( n5609 & n5868 ) | ( n5867 & n5868 ) ;
  assign n5870 = ( ~n5609 & n5867 ) | ( ~n5609 & n5868 ) | ( n5867 & n5868 ) ;
  assign n5871 = ( n5609 & ~n5869 ) | ( n5609 & n5870 ) | ( ~n5869 & n5870 ) ;
  assign n5872 = ( x75 & n5866 ) | ( x75 & ~n5871 ) | ( n5866 & ~n5871 ) ;
  assign n5873 = ( x75 & n5610 ) | ( x75 & ~n5807 ) | ( n5610 & ~n5807 ) ;
  assign n5874 = x75 & n5610 ;
  assign n5875 = ( ~n5615 & n5873 ) | ( ~n5615 & n5874 ) | ( n5873 & n5874 ) ;
  assign n5876 = ( n5615 & n5873 ) | ( n5615 & n5874 ) | ( n5873 & n5874 ) ;
  assign n5877 = ( n5615 & n5875 ) | ( n5615 & ~n5876 ) | ( n5875 & ~n5876 ) ;
  assign n5878 = ( x76 & n5872 ) | ( x76 & ~n5877 ) | ( n5872 & ~n5877 ) ;
  assign n5879 = ( x76 & n5616 ) | ( x76 & ~n5807 ) | ( n5616 & ~n5807 ) ;
  assign n5880 = x76 & n5616 ;
  assign n5881 = ( n5621 & n5879 ) | ( n5621 & n5880 ) | ( n5879 & n5880 ) ;
  assign n5882 = ( ~n5621 & n5879 ) | ( ~n5621 & n5880 ) | ( n5879 & n5880 ) ;
  assign n5883 = ( n5621 & ~n5881 ) | ( n5621 & n5882 ) | ( ~n5881 & n5882 ) ;
  assign n5884 = ( x77 & n5878 ) | ( x77 & ~n5883 ) | ( n5878 & ~n5883 ) ;
  assign n5885 = ( x77 & n5622 ) | ( x77 & ~n5807 ) | ( n5622 & ~n5807 ) ;
  assign n5886 = x77 & n5622 ;
  assign n5887 = ( ~n5627 & n5885 ) | ( ~n5627 & n5886 ) | ( n5885 & n5886 ) ;
  assign n5888 = ( n5627 & n5885 ) | ( n5627 & n5886 ) | ( n5885 & n5886 ) ;
  assign n5889 = ( n5627 & n5887 ) | ( n5627 & ~n5888 ) | ( n5887 & ~n5888 ) ;
  assign n5890 = ( x78 & n5884 ) | ( x78 & ~n5889 ) | ( n5884 & ~n5889 ) ;
  assign n5891 = ( x78 & n5628 ) | ( x78 & ~n5807 ) | ( n5628 & ~n5807 ) ;
  assign n5892 = x78 & n5628 ;
  assign n5893 = ( n5633 & n5891 ) | ( n5633 & n5892 ) | ( n5891 & n5892 ) ;
  assign n5894 = ( ~n5633 & n5891 ) | ( ~n5633 & n5892 ) | ( n5891 & n5892 ) ;
  assign n5895 = ( n5633 & ~n5893 ) | ( n5633 & n5894 ) | ( ~n5893 & n5894 ) ;
  assign n5896 = ( x79 & n5890 ) | ( x79 & ~n5895 ) | ( n5890 & ~n5895 ) ;
  assign n5897 = ( x79 & n5634 ) | ( x79 & ~n5807 ) | ( n5634 & ~n5807 ) ;
  assign n5898 = x79 & n5634 ;
  assign n5899 = ( ~n5639 & n5897 ) | ( ~n5639 & n5898 ) | ( n5897 & n5898 ) ;
  assign n5900 = ( n5639 & n5897 ) | ( n5639 & n5898 ) | ( n5897 & n5898 ) ;
  assign n5901 = ( n5639 & n5899 ) | ( n5639 & ~n5900 ) | ( n5899 & ~n5900 ) ;
  assign n5902 = ( x80 & n5896 ) | ( x80 & ~n5901 ) | ( n5896 & ~n5901 ) ;
  assign n5903 = ( x80 & n5640 ) | ( x80 & ~n5807 ) | ( n5640 & ~n5807 ) ;
  assign n5904 = x80 & n5640 ;
  assign n5905 = ( n5645 & n5903 ) | ( n5645 & n5904 ) | ( n5903 & n5904 ) ;
  assign n5906 = ( ~n5645 & n5903 ) | ( ~n5645 & n5904 ) | ( n5903 & n5904 ) ;
  assign n5907 = ( n5645 & ~n5905 ) | ( n5645 & n5906 ) | ( ~n5905 & n5906 ) ;
  assign n5908 = ( x81 & n5902 ) | ( x81 & ~n5907 ) | ( n5902 & ~n5907 ) ;
  assign n5909 = ( x81 & n5646 ) | ( x81 & ~n5807 ) | ( n5646 & ~n5807 ) ;
  assign n5910 = x81 & n5646 ;
  assign n5911 = ( ~n5651 & n5909 ) | ( ~n5651 & n5910 ) | ( n5909 & n5910 ) ;
  assign n5912 = ( n5651 & n5909 ) | ( n5651 & n5910 ) | ( n5909 & n5910 ) ;
  assign n5913 = ( n5651 & n5911 ) | ( n5651 & ~n5912 ) | ( n5911 & ~n5912 ) ;
  assign n5914 = ( x82 & n5908 ) | ( x82 & ~n5913 ) | ( n5908 & ~n5913 ) ;
  assign n5915 = ( x82 & n5652 ) | ( x82 & ~n5807 ) | ( n5652 & ~n5807 ) ;
  assign n5916 = x82 & n5652 ;
  assign n5917 = ( n5657 & n5915 ) | ( n5657 & n5916 ) | ( n5915 & n5916 ) ;
  assign n5918 = ( ~n5657 & n5915 ) | ( ~n5657 & n5916 ) | ( n5915 & n5916 ) ;
  assign n5919 = ( n5657 & ~n5917 ) | ( n5657 & n5918 ) | ( ~n5917 & n5918 ) ;
  assign n5920 = ( x83 & n5914 ) | ( x83 & ~n5919 ) | ( n5914 & ~n5919 ) ;
  assign n5921 = ( x83 & n5658 ) | ( x83 & ~n5807 ) | ( n5658 & ~n5807 ) ;
  assign n5922 = x83 & n5658 ;
  assign n5923 = ( ~n5663 & n5921 ) | ( ~n5663 & n5922 ) | ( n5921 & n5922 ) ;
  assign n5924 = ( n5663 & n5921 ) | ( n5663 & n5922 ) | ( n5921 & n5922 ) ;
  assign n5925 = ( n5663 & n5923 ) | ( n5663 & ~n5924 ) | ( n5923 & ~n5924 ) ;
  assign n5926 = ( x84 & n5920 ) | ( x84 & ~n5925 ) | ( n5920 & ~n5925 ) ;
  assign n5927 = ( x84 & n5664 ) | ( x84 & ~n5807 ) | ( n5664 & ~n5807 ) ;
  assign n5928 = x84 & n5664 ;
  assign n5929 = ( n5669 & n5927 ) | ( n5669 & n5928 ) | ( n5927 & n5928 ) ;
  assign n5930 = ( ~n5669 & n5927 ) | ( ~n5669 & n5928 ) | ( n5927 & n5928 ) ;
  assign n5931 = ( n5669 & ~n5929 ) | ( n5669 & n5930 ) | ( ~n5929 & n5930 ) ;
  assign n5932 = ( x85 & n5926 ) | ( x85 & ~n5931 ) | ( n5926 & ~n5931 ) ;
  assign n5933 = ( x85 & n5670 ) | ( x85 & ~n5807 ) | ( n5670 & ~n5807 ) ;
  assign n5934 = x85 & n5670 ;
  assign n5935 = ( ~n5675 & n5933 ) | ( ~n5675 & n5934 ) | ( n5933 & n5934 ) ;
  assign n5936 = ( n5675 & n5933 ) | ( n5675 & n5934 ) | ( n5933 & n5934 ) ;
  assign n5937 = ( n5675 & n5935 ) | ( n5675 & ~n5936 ) | ( n5935 & ~n5936 ) ;
  assign n5938 = ( x86 & n5932 ) | ( x86 & ~n5937 ) | ( n5932 & ~n5937 ) ;
  assign n5939 = ( x86 & n5676 ) | ( x86 & ~n5807 ) | ( n5676 & ~n5807 ) ;
  assign n5940 = x86 & n5676 ;
  assign n5941 = ( n5681 & n5939 ) | ( n5681 & n5940 ) | ( n5939 & n5940 ) ;
  assign n5942 = ( ~n5681 & n5939 ) | ( ~n5681 & n5940 ) | ( n5939 & n5940 ) ;
  assign n5943 = ( n5681 & ~n5941 ) | ( n5681 & n5942 ) | ( ~n5941 & n5942 ) ;
  assign n5944 = ( x87 & n5938 ) | ( x87 & ~n5943 ) | ( n5938 & ~n5943 ) ;
  assign n5945 = ( x87 & n5682 ) | ( x87 & ~n5807 ) | ( n5682 & ~n5807 ) ;
  assign n5946 = x87 & n5682 ;
  assign n5947 = ( ~n5687 & n5945 ) | ( ~n5687 & n5946 ) | ( n5945 & n5946 ) ;
  assign n5948 = ( n5687 & n5945 ) | ( n5687 & n5946 ) | ( n5945 & n5946 ) ;
  assign n5949 = ( n5687 & n5947 ) | ( n5687 & ~n5948 ) | ( n5947 & ~n5948 ) ;
  assign n5950 = ( x88 & n5944 ) | ( x88 & ~n5949 ) | ( n5944 & ~n5949 ) ;
  assign n5951 = ( x88 & n5688 ) | ( x88 & ~n5807 ) | ( n5688 & ~n5807 ) ;
  assign n5952 = x88 & n5688 ;
  assign n5953 = ( n5693 & n5951 ) | ( n5693 & n5952 ) | ( n5951 & n5952 ) ;
  assign n5954 = ( ~n5693 & n5951 ) | ( ~n5693 & n5952 ) | ( n5951 & n5952 ) ;
  assign n5955 = ( n5693 & ~n5953 ) | ( n5693 & n5954 ) | ( ~n5953 & n5954 ) ;
  assign n5956 = ( x89 & n5950 ) | ( x89 & ~n5955 ) | ( n5950 & ~n5955 ) ;
  assign n5957 = ( x89 & n5694 ) | ( x89 & ~n5807 ) | ( n5694 & ~n5807 ) ;
  assign n5958 = x89 & n5694 ;
  assign n5959 = ( ~n5699 & n5957 ) | ( ~n5699 & n5958 ) | ( n5957 & n5958 ) ;
  assign n5960 = ( n5699 & n5957 ) | ( n5699 & n5958 ) | ( n5957 & n5958 ) ;
  assign n5961 = ( n5699 & n5959 ) | ( n5699 & ~n5960 ) | ( n5959 & ~n5960 ) ;
  assign n5962 = ( x90 & n5956 ) | ( x90 & ~n5961 ) | ( n5956 & ~n5961 ) ;
  assign n5963 = ( x90 & n5700 ) | ( x90 & ~n5807 ) | ( n5700 & ~n5807 ) ;
  assign n5964 = x90 & n5700 ;
  assign n5965 = ( n5705 & n5963 ) | ( n5705 & n5964 ) | ( n5963 & n5964 ) ;
  assign n5966 = ( ~n5705 & n5963 ) | ( ~n5705 & n5964 ) | ( n5963 & n5964 ) ;
  assign n5967 = ( n5705 & ~n5965 ) | ( n5705 & n5966 ) | ( ~n5965 & n5966 ) ;
  assign n5968 = ( x91 & n5962 ) | ( x91 & ~n5967 ) | ( n5962 & ~n5967 ) ;
  assign n5969 = ( x91 & n5706 ) | ( x91 & ~n5807 ) | ( n5706 & ~n5807 ) ;
  assign n5970 = x91 & n5706 ;
  assign n5971 = ( ~n5711 & n5969 ) | ( ~n5711 & n5970 ) | ( n5969 & n5970 ) ;
  assign n5972 = ( n5711 & n5969 ) | ( n5711 & n5970 ) | ( n5969 & n5970 ) ;
  assign n5973 = ( n5711 & n5971 ) | ( n5711 & ~n5972 ) | ( n5971 & ~n5972 ) ;
  assign n5974 = ( x92 & n5968 ) | ( x92 & ~n5973 ) | ( n5968 & ~n5973 ) ;
  assign n5975 = ( x92 & n5712 ) | ( x92 & ~n5807 ) | ( n5712 & ~n5807 ) ;
  assign n5976 = x92 & n5712 ;
  assign n5977 = ( n5717 & n5975 ) | ( n5717 & n5976 ) | ( n5975 & n5976 ) ;
  assign n5978 = ( ~n5717 & n5975 ) | ( ~n5717 & n5976 ) | ( n5975 & n5976 ) ;
  assign n5979 = ( n5717 & ~n5977 ) | ( n5717 & n5978 ) | ( ~n5977 & n5978 ) ;
  assign n5980 = ( x93 & n5974 ) | ( x93 & ~n5979 ) | ( n5974 & ~n5979 ) ;
  assign n5981 = ( x93 & n5718 ) | ( x93 & ~n5807 ) | ( n5718 & ~n5807 ) ;
  assign n5982 = x93 & n5718 ;
  assign n5983 = ( ~n5723 & n5981 ) | ( ~n5723 & n5982 ) | ( n5981 & n5982 ) ;
  assign n5984 = ( n5723 & n5981 ) | ( n5723 & n5982 ) | ( n5981 & n5982 ) ;
  assign n5985 = ( n5723 & n5983 ) | ( n5723 & ~n5984 ) | ( n5983 & ~n5984 ) ;
  assign n5986 = ( x94 & n5980 ) | ( x94 & ~n5985 ) | ( n5980 & ~n5985 ) ;
  assign n5987 = ( x94 & n5724 ) | ( x94 & ~n5807 ) | ( n5724 & ~n5807 ) ;
  assign n5988 = x94 & n5724 ;
  assign n5989 = ( n5729 & n5987 ) | ( n5729 & n5988 ) | ( n5987 & n5988 ) ;
  assign n5990 = ( ~n5729 & n5987 ) | ( ~n5729 & n5988 ) | ( n5987 & n5988 ) ;
  assign n5991 = ( n5729 & ~n5989 ) | ( n5729 & n5990 ) | ( ~n5989 & n5990 ) ;
  assign n5992 = ( x95 & n5986 ) | ( x95 & ~n5991 ) | ( n5986 & ~n5991 ) ;
  assign n5993 = ( x95 & n5730 ) | ( x95 & ~n5807 ) | ( n5730 & ~n5807 ) ;
  assign n5994 = x95 & n5730 ;
  assign n5995 = ( ~n5735 & n5993 ) | ( ~n5735 & n5994 ) | ( n5993 & n5994 ) ;
  assign n5996 = ( n5735 & n5993 ) | ( n5735 & n5994 ) | ( n5993 & n5994 ) ;
  assign n5997 = ( n5735 & n5995 ) | ( n5735 & ~n5996 ) | ( n5995 & ~n5996 ) ;
  assign n5998 = ( x96 & n5992 ) | ( x96 & ~n5997 ) | ( n5992 & ~n5997 ) ;
  assign n5999 = ( x96 & n5736 ) | ( x96 & ~n5807 ) | ( n5736 & ~n5807 ) ;
  assign n6000 = x96 & n5736 ;
  assign n6001 = ( n5741 & n5999 ) | ( n5741 & n6000 ) | ( n5999 & n6000 ) ;
  assign n6002 = ( ~n5741 & n5999 ) | ( ~n5741 & n6000 ) | ( n5999 & n6000 ) ;
  assign n6003 = ( n5741 & ~n6001 ) | ( n5741 & n6002 ) | ( ~n6001 & n6002 ) ;
  assign n6004 = ( x97 & n5998 ) | ( x97 & ~n6003 ) | ( n5998 & ~n6003 ) ;
  assign n6005 = ( x97 & n5742 ) | ( x97 & ~n5807 ) | ( n5742 & ~n5807 ) ;
  assign n6006 = x97 & n5742 ;
  assign n6007 = ( ~n5747 & n6005 ) | ( ~n5747 & n6006 ) | ( n6005 & n6006 ) ;
  assign n6008 = ( n5747 & n6005 ) | ( n5747 & n6006 ) | ( n6005 & n6006 ) ;
  assign n6009 = ( n5747 & n6007 ) | ( n5747 & ~n6008 ) | ( n6007 & ~n6008 ) ;
  assign n6010 = ( x98 & n6004 ) | ( x98 & ~n6009 ) | ( n6004 & ~n6009 ) ;
  assign n6011 = ( x98 & n5748 ) | ( x98 & ~n5807 ) | ( n5748 & ~n5807 ) ;
  assign n6012 = x98 & n5748 ;
  assign n6013 = ( n5753 & n6011 ) | ( n5753 & n6012 ) | ( n6011 & n6012 ) ;
  assign n6014 = ( ~n5753 & n6011 ) | ( ~n5753 & n6012 ) | ( n6011 & n6012 ) ;
  assign n6015 = ( n5753 & ~n6013 ) | ( n5753 & n6014 ) | ( ~n6013 & n6014 ) ;
  assign n6016 = ( x99 & n6010 ) | ( x99 & ~n6015 ) | ( n6010 & ~n6015 ) ;
  assign n6017 = ( x99 & n5754 ) | ( x99 & ~n5807 ) | ( n5754 & ~n5807 ) ;
  assign n6018 = x99 & n5754 ;
  assign n6019 = ( ~n5759 & n6017 ) | ( ~n5759 & n6018 ) | ( n6017 & n6018 ) ;
  assign n6020 = ( n5759 & n6017 ) | ( n5759 & n6018 ) | ( n6017 & n6018 ) ;
  assign n6021 = ( n5759 & n6019 ) | ( n5759 & ~n6020 ) | ( n6019 & ~n6020 ) ;
  assign n6022 = ( x100 & n6016 ) | ( x100 & ~n6021 ) | ( n6016 & ~n6021 ) ;
  assign n6023 = ( x100 & n5760 ) | ( x100 & ~n5807 ) | ( n5760 & ~n5807 ) ;
  assign n6024 = x100 & n5760 ;
  assign n6025 = ( n5765 & n6023 ) | ( n5765 & n6024 ) | ( n6023 & n6024 ) ;
  assign n6026 = ( ~n5765 & n6023 ) | ( ~n5765 & n6024 ) | ( n6023 & n6024 ) ;
  assign n6027 = ( n5765 & ~n6025 ) | ( n5765 & n6026 ) | ( ~n6025 & n6026 ) ;
  assign n6028 = ( x101 & n6022 ) | ( x101 & ~n6027 ) | ( n6022 & ~n6027 ) ;
  assign n6029 = ( x101 & n5766 ) | ( x101 & ~n5807 ) | ( n5766 & ~n5807 ) ;
  assign n6030 = x101 & n5766 ;
  assign n6031 = ( ~n5771 & n6029 ) | ( ~n5771 & n6030 ) | ( n6029 & n6030 ) ;
  assign n6032 = ( n5771 & n6029 ) | ( n5771 & n6030 ) | ( n6029 & n6030 ) ;
  assign n6033 = ( n5771 & n6031 ) | ( n5771 & ~n6032 ) | ( n6031 & ~n6032 ) ;
  assign n6034 = ( x102 & n6028 ) | ( x102 & ~n6033 ) | ( n6028 & ~n6033 ) ;
  assign n6035 = ( x102 & n5772 ) | ( x102 & ~n5807 ) | ( n5772 & ~n5807 ) ;
  assign n6036 = x102 & n5772 ;
  assign n6037 = ( n5777 & n6035 ) | ( n5777 & n6036 ) | ( n6035 & n6036 ) ;
  assign n6038 = ( ~n5777 & n6035 ) | ( ~n5777 & n6036 ) | ( n6035 & n6036 ) ;
  assign n6039 = ( n5777 & ~n6037 ) | ( n5777 & n6038 ) | ( ~n6037 & n6038 ) ;
  assign n6040 = ( x103 & n6034 ) | ( x103 & ~n6039 ) | ( n6034 & ~n6039 ) ;
  assign n6041 = ( x103 & n5778 ) | ( x103 & ~n5807 ) | ( n5778 & ~n5807 ) ;
  assign n6042 = x103 & n5778 ;
  assign n6043 = ( ~n5783 & n6041 ) | ( ~n5783 & n6042 ) | ( n6041 & n6042 ) ;
  assign n6044 = ( n5783 & n6041 ) | ( n5783 & n6042 ) | ( n6041 & n6042 ) ;
  assign n6045 = ( n5783 & n6043 ) | ( n5783 & ~n6044 ) | ( n6043 & ~n6044 ) ;
  assign n6046 = ( x104 & n6040 ) | ( x104 & ~n6045 ) | ( n6040 & ~n6045 ) ;
  assign n6047 = ( x104 & n5784 ) | ( x104 & ~n5807 ) | ( n5784 & ~n5807 ) ;
  assign n6048 = x104 & n5784 ;
  assign n6049 = ( n5789 & n6047 ) | ( n5789 & n6048 ) | ( n6047 & n6048 ) ;
  assign n6050 = ( ~n5789 & n6047 ) | ( ~n5789 & n6048 ) | ( n6047 & n6048 ) ;
  assign n6051 = ( n5789 & ~n6049 ) | ( n5789 & n6050 ) | ( ~n6049 & n6050 ) ;
  assign n6052 = ( x105 & n6046 ) | ( x105 & ~n6051 ) | ( n6046 & ~n6051 ) ;
  assign n6053 = ( x105 & n5790 ) | ( x105 & ~n5807 ) | ( n5790 & ~n5807 ) ;
  assign n6054 = x105 & n5790 ;
  assign n6055 = ( ~n5795 & n6053 ) | ( ~n5795 & n6054 ) | ( n6053 & n6054 ) ;
  assign n6056 = ( n5795 & n6053 ) | ( n5795 & n6054 ) | ( n6053 & n6054 ) ;
  assign n6057 = ( n5795 & n6055 ) | ( n5795 & ~n6056 ) | ( n6055 & ~n6056 ) ;
  assign n6058 = ( x106 & n6052 ) | ( x106 & ~n6057 ) | ( n6052 & ~n6057 ) ;
  assign n6059 = ( x106 & n5796 ) | ( x106 & ~n5807 ) | ( n5796 & ~n5807 ) ;
  assign n6060 = x106 & n5796 ;
  assign n6061 = ( ~n5801 & n6059 ) | ( ~n5801 & n6060 ) | ( n6059 & n6060 ) ;
  assign n6062 = ( n5801 & n6059 ) | ( n5801 & n6060 ) | ( n6059 & n6060 ) ;
  assign n6063 = ( n5801 & n6061 ) | ( n5801 & ~n6062 ) | ( n6061 & ~n6062 ) ;
  assign n6064 = ( x107 & n6058 ) | ( x107 & ~n6063 ) | ( n6058 & ~n6063 ) ;
  assign n6065 = x108 | n6064 ;
  assign n6066 = ( x108 & n149 ) | ( x108 & n6064 ) | ( n149 & n6064 ) ;
  assign n6067 = ( n5805 & ~n6065 ) | ( n5805 & n6066 ) | ( ~n6065 & n6066 ) ;
  assign n6068 = ( x108 & ~n5805 ) | ( x108 & n6064 ) | ( ~n5805 & n6064 ) ;
  assign n6069 = n149 | n6068 ;
  assign n6070 = ( x19 & ~x64 ) | ( x19 & n6069 ) | ( ~x64 & n6069 ) ;
  assign n6071 = ~x19 & n6069 ;
  assign n6072 = ( n5811 & n6070 ) | ( n5811 & ~n6071 ) | ( n6070 & ~n6071 ) ;
  assign n6073 = ~x18 & x64 ;
  assign n6074 = ( x65 & ~n6072 ) | ( x65 & n6073 ) | ( ~n6072 & n6073 ) ;
  assign n6075 = ( x65 & n5811 ) | ( x65 & ~n6069 ) | ( n5811 & ~n6069 ) ;
  assign n6076 = x65 & n5811 ;
  assign n6077 = ( n5810 & n6075 ) | ( n5810 & n6076 ) | ( n6075 & n6076 ) ;
  assign n6078 = ( ~n5810 & n6075 ) | ( ~n5810 & n6076 ) | ( n6075 & n6076 ) ;
  assign n6079 = ( n5810 & ~n6077 ) | ( n5810 & n6078 ) | ( ~n6077 & n6078 ) ;
  assign n6080 = ( x66 & n6074 ) | ( x66 & ~n6079 ) | ( n6074 & ~n6079 ) ;
  assign n6081 = ( x66 & n5812 ) | ( x66 & ~n6069 ) | ( n5812 & ~n6069 ) ;
  assign n6082 = x66 & n5812 ;
  assign n6083 = ( n5817 & n6081 ) | ( n5817 & n6082 ) | ( n6081 & n6082 ) ;
  assign n6084 = ( ~n5817 & n6081 ) | ( ~n5817 & n6082 ) | ( n6081 & n6082 ) ;
  assign n6085 = ( n5817 & ~n6083 ) | ( n5817 & n6084 ) | ( ~n6083 & n6084 ) ;
  assign n6086 = ( x67 & n6080 ) | ( x67 & ~n6085 ) | ( n6080 & ~n6085 ) ;
  assign n6087 = ( x67 & n5818 ) | ( x67 & ~n6069 ) | ( n5818 & ~n6069 ) ;
  assign n6088 = x67 & n5818 ;
  assign n6089 = ( ~n5823 & n6087 ) | ( ~n5823 & n6088 ) | ( n6087 & n6088 ) ;
  assign n6090 = ( n5823 & n6087 ) | ( n5823 & n6088 ) | ( n6087 & n6088 ) ;
  assign n6091 = ( n5823 & n6089 ) | ( n5823 & ~n6090 ) | ( n6089 & ~n6090 ) ;
  assign n6092 = ( x68 & n6086 ) | ( x68 & ~n6091 ) | ( n6086 & ~n6091 ) ;
  assign n6093 = ( x68 & n5824 ) | ( x68 & ~n6069 ) | ( n5824 & ~n6069 ) ;
  assign n6094 = x68 & n5824 ;
  assign n6095 = ( n5829 & n6093 ) | ( n5829 & n6094 ) | ( n6093 & n6094 ) ;
  assign n6096 = ( ~n5829 & n6093 ) | ( ~n5829 & n6094 ) | ( n6093 & n6094 ) ;
  assign n6097 = ( n5829 & ~n6095 ) | ( n5829 & n6096 ) | ( ~n6095 & n6096 ) ;
  assign n6098 = ( x69 & n6092 ) | ( x69 & ~n6097 ) | ( n6092 & ~n6097 ) ;
  assign n6099 = ( x69 & n5830 ) | ( x69 & ~n6069 ) | ( n5830 & ~n6069 ) ;
  assign n6100 = x69 & n5830 ;
  assign n6101 = ( ~n5835 & n6099 ) | ( ~n5835 & n6100 ) | ( n6099 & n6100 ) ;
  assign n6102 = ( n5835 & n6099 ) | ( n5835 & n6100 ) | ( n6099 & n6100 ) ;
  assign n6103 = ( n5835 & n6101 ) | ( n5835 & ~n6102 ) | ( n6101 & ~n6102 ) ;
  assign n6104 = ( x70 & n6098 ) | ( x70 & ~n6103 ) | ( n6098 & ~n6103 ) ;
  assign n6105 = ( x70 & n5836 ) | ( x70 & ~n6069 ) | ( n5836 & ~n6069 ) ;
  assign n6106 = x70 & n5836 ;
  assign n6107 = ( n5841 & n6105 ) | ( n5841 & n6106 ) | ( n6105 & n6106 ) ;
  assign n6108 = ( ~n5841 & n6105 ) | ( ~n5841 & n6106 ) | ( n6105 & n6106 ) ;
  assign n6109 = ( n5841 & ~n6107 ) | ( n5841 & n6108 ) | ( ~n6107 & n6108 ) ;
  assign n6110 = ( x71 & n6104 ) | ( x71 & ~n6109 ) | ( n6104 & ~n6109 ) ;
  assign n6111 = ( x71 & n5842 ) | ( x71 & ~n6069 ) | ( n5842 & ~n6069 ) ;
  assign n6112 = x71 & n5842 ;
  assign n6113 = ( ~n5847 & n6111 ) | ( ~n5847 & n6112 ) | ( n6111 & n6112 ) ;
  assign n6114 = ( n5847 & n6111 ) | ( n5847 & n6112 ) | ( n6111 & n6112 ) ;
  assign n6115 = ( n5847 & n6113 ) | ( n5847 & ~n6114 ) | ( n6113 & ~n6114 ) ;
  assign n6116 = ( x72 & n6110 ) | ( x72 & ~n6115 ) | ( n6110 & ~n6115 ) ;
  assign n6117 = ( x72 & n5848 ) | ( x72 & ~n6069 ) | ( n5848 & ~n6069 ) ;
  assign n6118 = x72 & n5848 ;
  assign n6119 = ( n5853 & n6117 ) | ( n5853 & n6118 ) | ( n6117 & n6118 ) ;
  assign n6120 = ( ~n5853 & n6117 ) | ( ~n5853 & n6118 ) | ( n6117 & n6118 ) ;
  assign n6121 = ( n5853 & ~n6119 ) | ( n5853 & n6120 ) | ( ~n6119 & n6120 ) ;
  assign n6122 = ( x73 & n6116 ) | ( x73 & ~n6121 ) | ( n6116 & ~n6121 ) ;
  assign n6123 = ( x73 & n5854 ) | ( x73 & ~n6069 ) | ( n5854 & ~n6069 ) ;
  assign n6124 = x73 & n5854 ;
  assign n6125 = ( ~n5859 & n6123 ) | ( ~n5859 & n6124 ) | ( n6123 & n6124 ) ;
  assign n6126 = ( n5859 & n6123 ) | ( n5859 & n6124 ) | ( n6123 & n6124 ) ;
  assign n6127 = ( n5859 & n6125 ) | ( n5859 & ~n6126 ) | ( n6125 & ~n6126 ) ;
  assign n6128 = ( x74 & n6122 ) | ( x74 & ~n6127 ) | ( n6122 & ~n6127 ) ;
  assign n6129 = ( x74 & n5860 ) | ( x74 & ~n6069 ) | ( n5860 & ~n6069 ) ;
  assign n6130 = x74 & n5860 ;
  assign n6131 = ( n5865 & n6129 ) | ( n5865 & n6130 ) | ( n6129 & n6130 ) ;
  assign n6132 = ( ~n5865 & n6129 ) | ( ~n5865 & n6130 ) | ( n6129 & n6130 ) ;
  assign n6133 = ( n5865 & ~n6131 ) | ( n5865 & n6132 ) | ( ~n6131 & n6132 ) ;
  assign n6134 = ( x75 & n6128 ) | ( x75 & ~n6133 ) | ( n6128 & ~n6133 ) ;
  assign n6135 = ( x75 & n5866 ) | ( x75 & ~n6069 ) | ( n5866 & ~n6069 ) ;
  assign n6136 = x75 & n5866 ;
  assign n6137 = ( ~n5871 & n6135 ) | ( ~n5871 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6138 = ( n5871 & n6135 ) | ( n5871 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6139 = ( n5871 & n6137 ) | ( n5871 & ~n6138 ) | ( n6137 & ~n6138 ) ;
  assign n6140 = ( x76 & n6134 ) | ( x76 & ~n6139 ) | ( n6134 & ~n6139 ) ;
  assign n6141 = ( x76 & n5872 ) | ( x76 & ~n6069 ) | ( n5872 & ~n6069 ) ;
  assign n6142 = x76 & n5872 ;
  assign n6143 = ( n5877 & n6141 ) | ( n5877 & n6142 ) | ( n6141 & n6142 ) ;
  assign n6144 = ( ~n5877 & n6141 ) | ( ~n5877 & n6142 ) | ( n6141 & n6142 ) ;
  assign n6145 = ( n5877 & ~n6143 ) | ( n5877 & n6144 ) | ( ~n6143 & n6144 ) ;
  assign n6146 = ( x77 & n6140 ) | ( x77 & ~n6145 ) | ( n6140 & ~n6145 ) ;
  assign n6147 = ( x77 & n5878 ) | ( x77 & ~n6069 ) | ( n5878 & ~n6069 ) ;
  assign n6148 = x77 & n5878 ;
  assign n6149 = ( ~n5883 & n6147 ) | ( ~n5883 & n6148 ) | ( n6147 & n6148 ) ;
  assign n6150 = ( n5883 & n6147 ) | ( n5883 & n6148 ) | ( n6147 & n6148 ) ;
  assign n6151 = ( n5883 & n6149 ) | ( n5883 & ~n6150 ) | ( n6149 & ~n6150 ) ;
  assign n6152 = ( x78 & n6146 ) | ( x78 & ~n6151 ) | ( n6146 & ~n6151 ) ;
  assign n6153 = ( x78 & n5884 ) | ( x78 & ~n6069 ) | ( n5884 & ~n6069 ) ;
  assign n6154 = x78 & n5884 ;
  assign n6155 = ( n5889 & n6153 ) | ( n5889 & n6154 ) | ( n6153 & n6154 ) ;
  assign n6156 = ( ~n5889 & n6153 ) | ( ~n5889 & n6154 ) | ( n6153 & n6154 ) ;
  assign n6157 = ( n5889 & ~n6155 ) | ( n5889 & n6156 ) | ( ~n6155 & n6156 ) ;
  assign n6158 = ( x79 & n6152 ) | ( x79 & ~n6157 ) | ( n6152 & ~n6157 ) ;
  assign n6159 = ( x79 & n5890 ) | ( x79 & ~n6069 ) | ( n5890 & ~n6069 ) ;
  assign n6160 = x79 & n5890 ;
  assign n6161 = ( ~n5895 & n6159 ) | ( ~n5895 & n6160 ) | ( n6159 & n6160 ) ;
  assign n6162 = ( n5895 & n6159 ) | ( n5895 & n6160 ) | ( n6159 & n6160 ) ;
  assign n6163 = ( n5895 & n6161 ) | ( n5895 & ~n6162 ) | ( n6161 & ~n6162 ) ;
  assign n6164 = ( x80 & n6158 ) | ( x80 & ~n6163 ) | ( n6158 & ~n6163 ) ;
  assign n6165 = ( x80 & n5896 ) | ( x80 & ~n6069 ) | ( n5896 & ~n6069 ) ;
  assign n6166 = x80 & n5896 ;
  assign n6167 = ( n5901 & n6165 ) | ( n5901 & n6166 ) | ( n6165 & n6166 ) ;
  assign n6168 = ( ~n5901 & n6165 ) | ( ~n5901 & n6166 ) | ( n6165 & n6166 ) ;
  assign n6169 = ( n5901 & ~n6167 ) | ( n5901 & n6168 ) | ( ~n6167 & n6168 ) ;
  assign n6170 = ( x81 & n6164 ) | ( x81 & ~n6169 ) | ( n6164 & ~n6169 ) ;
  assign n6171 = ( x81 & n5902 ) | ( x81 & ~n6069 ) | ( n5902 & ~n6069 ) ;
  assign n6172 = x81 & n5902 ;
  assign n6173 = ( ~n5907 & n6171 ) | ( ~n5907 & n6172 ) | ( n6171 & n6172 ) ;
  assign n6174 = ( n5907 & n6171 ) | ( n5907 & n6172 ) | ( n6171 & n6172 ) ;
  assign n6175 = ( n5907 & n6173 ) | ( n5907 & ~n6174 ) | ( n6173 & ~n6174 ) ;
  assign n6176 = ( x82 & n6170 ) | ( x82 & ~n6175 ) | ( n6170 & ~n6175 ) ;
  assign n6177 = ( x82 & n5908 ) | ( x82 & ~n6069 ) | ( n5908 & ~n6069 ) ;
  assign n6178 = x82 & n5908 ;
  assign n6179 = ( n5913 & n6177 ) | ( n5913 & n6178 ) | ( n6177 & n6178 ) ;
  assign n6180 = ( ~n5913 & n6177 ) | ( ~n5913 & n6178 ) | ( n6177 & n6178 ) ;
  assign n6181 = ( n5913 & ~n6179 ) | ( n5913 & n6180 ) | ( ~n6179 & n6180 ) ;
  assign n6182 = ( x83 & n6176 ) | ( x83 & ~n6181 ) | ( n6176 & ~n6181 ) ;
  assign n6183 = ( x83 & n5914 ) | ( x83 & ~n6069 ) | ( n5914 & ~n6069 ) ;
  assign n6184 = x83 & n5914 ;
  assign n6185 = ( ~n5919 & n6183 ) | ( ~n5919 & n6184 ) | ( n6183 & n6184 ) ;
  assign n6186 = ( n5919 & n6183 ) | ( n5919 & n6184 ) | ( n6183 & n6184 ) ;
  assign n6187 = ( n5919 & n6185 ) | ( n5919 & ~n6186 ) | ( n6185 & ~n6186 ) ;
  assign n6188 = ( x84 & n6182 ) | ( x84 & ~n6187 ) | ( n6182 & ~n6187 ) ;
  assign n6189 = ( x84 & n5920 ) | ( x84 & ~n6069 ) | ( n5920 & ~n6069 ) ;
  assign n6190 = x84 & n5920 ;
  assign n6191 = ( n5925 & n6189 ) | ( n5925 & n6190 ) | ( n6189 & n6190 ) ;
  assign n6192 = ( ~n5925 & n6189 ) | ( ~n5925 & n6190 ) | ( n6189 & n6190 ) ;
  assign n6193 = ( n5925 & ~n6191 ) | ( n5925 & n6192 ) | ( ~n6191 & n6192 ) ;
  assign n6194 = ( x85 & n6188 ) | ( x85 & ~n6193 ) | ( n6188 & ~n6193 ) ;
  assign n6195 = ( x85 & n5926 ) | ( x85 & ~n6069 ) | ( n5926 & ~n6069 ) ;
  assign n6196 = x85 & n5926 ;
  assign n6197 = ( ~n5931 & n6195 ) | ( ~n5931 & n6196 ) | ( n6195 & n6196 ) ;
  assign n6198 = ( n5931 & n6195 ) | ( n5931 & n6196 ) | ( n6195 & n6196 ) ;
  assign n6199 = ( n5931 & n6197 ) | ( n5931 & ~n6198 ) | ( n6197 & ~n6198 ) ;
  assign n6200 = ( x86 & n6194 ) | ( x86 & ~n6199 ) | ( n6194 & ~n6199 ) ;
  assign n6201 = ( x86 & n5932 ) | ( x86 & ~n6069 ) | ( n5932 & ~n6069 ) ;
  assign n6202 = x86 & n5932 ;
  assign n6203 = ( n5937 & n6201 ) | ( n5937 & n6202 ) | ( n6201 & n6202 ) ;
  assign n6204 = ( ~n5937 & n6201 ) | ( ~n5937 & n6202 ) | ( n6201 & n6202 ) ;
  assign n6205 = ( n5937 & ~n6203 ) | ( n5937 & n6204 ) | ( ~n6203 & n6204 ) ;
  assign n6206 = ( x87 & n6200 ) | ( x87 & ~n6205 ) | ( n6200 & ~n6205 ) ;
  assign n6207 = ( x87 & n5938 ) | ( x87 & ~n6069 ) | ( n5938 & ~n6069 ) ;
  assign n6208 = x87 & n5938 ;
  assign n6209 = ( ~n5943 & n6207 ) | ( ~n5943 & n6208 ) | ( n6207 & n6208 ) ;
  assign n6210 = ( n5943 & n6207 ) | ( n5943 & n6208 ) | ( n6207 & n6208 ) ;
  assign n6211 = ( n5943 & n6209 ) | ( n5943 & ~n6210 ) | ( n6209 & ~n6210 ) ;
  assign n6212 = ( x88 & n6206 ) | ( x88 & ~n6211 ) | ( n6206 & ~n6211 ) ;
  assign n6213 = ( x88 & n5944 ) | ( x88 & ~n6069 ) | ( n5944 & ~n6069 ) ;
  assign n6214 = x88 & n5944 ;
  assign n6215 = ( n5949 & n6213 ) | ( n5949 & n6214 ) | ( n6213 & n6214 ) ;
  assign n6216 = ( ~n5949 & n6213 ) | ( ~n5949 & n6214 ) | ( n6213 & n6214 ) ;
  assign n6217 = ( n5949 & ~n6215 ) | ( n5949 & n6216 ) | ( ~n6215 & n6216 ) ;
  assign n6218 = ( x89 & n6212 ) | ( x89 & ~n6217 ) | ( n6212 & ~n6217 ) ;
  assign n6219 = ( x89 & n5950 ) | ( x89 & ~n6069 ) | ( n5950 & ~n6069 ) ;
  assign n6220 = x89 & n5950 ;
  assign n6221 = ( ~n5955 & n6219 ) | ( ~n5955 & n6220 ) | ( n6219 & n6220 ) ;
  assign n6222 = ( n5955 & n6219 ) | ( n5955 & n6220 ) | ( n6219 & n6220 ) ;
  assign n6223 = ( n5955 & n6221 ) | ( n5955 & ~n6222 ) | ( n6221 & ~n6222 ) ;
  assign n6224 = ( x90 & n6218 ) | ( x90 & ~n6223 ) | ( n6218 & ~n6223 ) ;
  assign n6225 = ( x90 & n5956 ) | ( x90 & ~n6069 ) | ( n5956 & ~n6069 ) ;
  assign n6226 = x90 & n5956 ;
  assign n6227 = ( n5961 & n6225 ) | ( n5961 & n6226 ) | ( n6225 & n6226 ) ;
  assign n6228 = ( ~n5961 & n6225 ) | ( ~n5961 & n6226 ) | ( n6225 & n6226 ) ;
  assign n6229 = ( n5961 & ~n6227 ) | ( n5961 & n6228 ) | ( ~n6227 & n6228 ) ;
  assign n6230 = ( x91 & n6224 ) | ( x91 & ~n6229 ) | ( n6224 & ~n6229 ) ;
  assign n6231 = ( x91 & n5962 ) | ( x91 & ~n6069 ) | ( n5962 & ~n6069 ) ;
  assign n6232 = x91 & n5962 ;
  assign n6233 = ( ~n5967 & n6231 ) | ( ~n5967 & n6232 ) | ( n6231 & n6232 ) ;
  assign n6234 = ( n5967 & n6231 ) | ( n5967 & n6232 ) | ( n6231 & n6232 ) ;
  assign n6235 = ( n5967 & n6233 ) | ( n5967 & ~n6234 ) | ( n6233 & ~n6234 ) ;
  assign n6236 = ( x92 & n6230 ) | ( x92 & ~n6235 ) | ( n6230 & ~n6235 ) ;
  assign n6237 = ( x92 & n5968 ) | ( x92 & ~n6069 ) | ( n5968 & ~n6069 ) ;
  assign n6238 = x92 & n5968 ;
  assign n6239 = ( n5973 & n6237 ) | ( n5973 & n6238 ) | ( n6237 & n6238 ) ;
  assign n6240 = ( ~n5973 & n6237 ) | ( ~n5973 & n6238 ) | ( n6237 & n6238 ) ;
  assign n6241 = ( n5973 & ~n6239 ) | ( n5973 & n6240 ) | ( ~n6239 & n6240 ) ;
  assign n6242 = ( x93 & n6236 ) | ( x93 & ~n6241 ) | ( n6236 & ~n6241 ) ;
  assign n6243 = ( x93 & n5974 ) | ( x93 & ~n6069 ) | ( n5974 & ~n6069 ) ;
  assign n6244 = x93 & n5974 ;
  assign n6245 = ( ~n5979 & n6243 ) | ( ~n5979 & n6244 ) | ( n6243 & n6244 ) ;
  assign n6246 = ( n5979 & n6243 ) | ( n5979 & n6244 ) | ( n6243 & n6244 ) ;
  assign n6247 = ( n5979 & n6245 ) | ( n5979 & ~n6246 ) | ( n6245 & ~n6246 ) ;
  assign n6248 = ( x94 & n6242 ) | ( x94 & ~n6247 ) | ( n6242 & ~n6247 ) ;
  assign n6249 = ( x94 & n5980 ) | ( x94 & ~n6069 ) | ( n5980 & ~n6069 ) ;
  assign n6250 = x94 & n5980 ;
  assign n6251 = ( n5985 & n6249 ) | ( n5985 & n6250 ) | ( n6249 & n6250 ) ;
  assign n6252 = ( ~n5985 & n6249 ) | ( ~n5985 & n6250 ) | ( n6249 & n6250 ) ;
  assign n6253 = ( n5985 & ~n6251 ) | ( n5985 & n6252 ) | ( ~n6251 & n6252 ) ;
  assign n6254 = ( x95 & n6248 ) | ( x95 & ~n6253 ) | ( n6248 & ~n6253 ) ;
  assign n6255 = ( x95 & n5986 ) | ( x95 & ~n6069 ) | ( n5986 & ~n6069 ) ;
  assign n6256 = x95 & n5986 ;
  assign n6257 = ( ~n5991 & n6255 ) | ( ~n5991 & n6256 ) | ( n6255 & n6256 ) ;
  assign n6258 = ( n5991 & n6255 ) | ( n5991 & n6256 ) | ( n6255 & n6256 ) ;
  assign n6259 = ( n5991 & n6257 ) | ( n5991 & ~n6258 ) | ( n6257 & ~n6258 ) ;
  assign n6260 = ( x96 & n6254 ) | ( x96 & ~n6259 ) | ( n6254 & ~n6259 ) ;
  assign n6261 = ( x96 & n5992 ) | ( x96 & ~n6069 ) | ( n5992 & ~n6069 ) ;
  assign n6262 = x96 & n5992 ;
  assign n6263 = ( n5997 & n6261 ) | ( n5997 & n6262 ) | ( n6261 & n6262 ) ;
  assign n6264 = ( ~n5997 & n6261 ) | ( ~n5997 & n6262 ) | ( n6261 & n6262 ) ;
  assign n6265 = ( n5997 & ~n6263 ) | ( n5997 & n6264 ) | ( ~n6263 & n6264 ) ;
  assign n6266 = ( x97 & n6260 ) | ( x97 & ~n6265 ) | ( n6260 & ~n6265 ) ;
  assign n6267 = ( x97 & n5998 ) | ( x97 & ~n6069 ) | ( n5998 & ~n6069 ) ;
  assign n6268 = x97 & n5998 ;
  assign n6269 = ( ~n6003 & n6267 ) | ( ~n6003 & n6268 ) | ( n6267 & n6268 ) ;
  assign n6270 = ( n6003 & n6267 ) | ( n6003 & n6268 ) | ( n6267 & n6268 ) ;
  assign n6271 = ( n6003 & n6269 ) | ( n6003 & ~n6270 ) | ( n6269 & ~n6270 ) ;
  assign n6272 = ( x98 & n6266 ) | ( x98 & ~n6271 ) | ( n6266 & ~n6271 ) ;
  assign n6273 = ( x98 & n6004 ) | ( x98 & ~n6069 ) | ( n6004 & ~n6069 ) ;
  assign n6274 = x98 & n6004 ;
  assign n6275 = ( n6009 & n6273 ) | ( n6009 & n6274 ) | ( n6273 & n6274 ) ;
  assign n6276 = ( ~n6009 & n6273 ) | ( ~n6009 & n6274 ) | ( n6273 & n6274 ) ;
  assign n6277 = ( n6009 & ~n6275 ) | ( n6009 & n6276 ) | ( ~n6275 & n6276 ) ;
  assign n6278 = ( x99 & n6272 ) | ( x99 & ~n6277 ) | ( n6272 & ~n6277 ) ;
  assign n6279 = ( x99 & n6010 ) | ( x99 & ~n6069 ) | ( n6010 & ~n6069 ) ;
  assign n6280 = x99 & n6010 ;
  assign n6281 = ( ~n6015 & n6279 ) | ( ~n6015 & n6280 ) | ( n6279 & n6280 ) ;
  assign n6282 = ( n6015 & n6279 ) | ( n6015 & n6280 ) | ( n6279 & n6280 ) ;
  assign n6283 = ( n6015 & n6281 ) | ( n6015 & ~n6282 ) | ( n6281 & ~n6282 ) ;
  assign n6284 = ( x100 & n6278 ) | ( x100 & ~n6283 ) | ( n6278 & ~n6283 ) ;
  assign n6285 = ( x100 & n6016 ) | ( x100 & ~n6069 ) | ( n6016 & ~n6069 ) ;
  assign n6286 = x100 & n6016 ;
  assign n6287 = ( n6021 & n6285 ) | ( n6021 & n6286 ) | ( n6285 & n6286 ) ;
  assign n6288 = ( ~n6021 & n6285 ) | ( ~n6021 & n6286 ) | ( n6285 & n6286 ) ;
  assign n6289 = ( n6021 & ~n6287 ) | ( n6021 & n6288 ) | ( ~n6287 & n6288 ) ;
  assign n6290 = ( x101 & n6284 ) | ( x101 & ~n6289 ) | ( n6284 & ~n6289 ) ;
  assign n6291 = ( x101 & n6022 ) | ( x101 & ~n6069 ) | ( n6022 & ~n6069 ) ;
  assign n6292 = x101 & n6022 ;
  assign n6293 = ( ~n6027 & n6291 ) | ( ~n6027 & n6292 ) | ( n6291 & n6292 ) ;
  assign n6294 = ( n6027 & n6291 ) | ( n6027 & n6292 ) | ( n6291 & n6292 ) ;
  assign n6295 = ( n6027 & n6293 ) | ( n6027 & ~n6294 ) | ( n6293 & ~n6294 ) ;
  assign n6296 = ( x102 & n6290 ) | ( x102 & ~n6295 ) | ( n6290 & ~n6295 ) ;
  assign n6297 = ( x102 & n6028 ) | ( x102 & ~n6069 ) | ( n6028 & ~n6069 ) ;
  assign n6298 = x102 & n6028 ;
  assign n6299 = ( n6033 & n6297 ) | ( n6033 & n6298 ) | ( n6297 & n6298 ) ;
  assign n6300 = ( ~n6033 & n6297 ) | ( ~n6033 & n6298 ) | ( n6297 & n6298 ) ;
  assign n6301 = ( n6033 & ~n6299 ) | ( n6033 & n6300 ) | ( ~n6299 & n6300 ) ;
  assign n6302 = ( x103 & n6296 ) | ( x103 & ~n6301 ) | ( n6296 & ~n6301 ) ;
  assign n6303 = ( x103 & n6034 ) | ( x103 & ~n6069 ) | ( n6034 & ~n6069 ) ;
  assign n6304 = x103 & n6034 ;
  assign n6305 = ( ~n6039 & n6303 ) | ( ~n6039 & n6304 ) | ( n6303 & n6304 ) ;
  assign n6306 = ( n6039 & n6303 ) | ( n6039 & n6304 ) | ( n6303 & n6304 ) ;
  assign n6307 = ( n6039 & n6305 ) | ( n6039 & ~n6306 ) | ( n6305 & ~n6306 ) ;
  assign n6308 = ( x104 & n6302 ) | ( x104 & ~n6307 ) | ( n6302 & ~n6307 ) ;
  assign n6309 = ( x104 & n6040 ) | ( x104 & ~n6069 ) | ( n6040 & ~n6069 ) ;
  assign n6310 = x104 & n6040 ;
  assign n6311 = ( n6045 & n6309 ) | ( n6045 & n6310 ) | ( n6309 & n6310 ) ;
  assign n6312 = ( ~n6045 & n6309 ) | ( ~n6045 & n6310 ) | ( n6309 & n6310 ) ;
  assign n6313 = ( n6045 & ~n6311 ) | ( n6045 & n6312 ) | ( ~n6311 & n6312 ) ;
  assign n6314 = ( x105 & n6308 ) | ( x105 & ~n6313 ) | ( n6308 & ~n6313 ) ;
  assign n6315 = ( x105 & n6046 ) | ( x105 & ~n6069 ) | ( n6046 & ~n6069 ) ;
  assign n6316 = x105 & n6046 ;
  assign n6317 = ( ~n6051 & n6315 ) | ( ~n6051 & n6316 ) | ( n6315 & n6316 ) ;
  assign n6318 = ( n6051 & n6315 ) | ( n6051 & n6316 ) | ( n6315 & n6316 ) ;
  assign n6319 = ( n6051 & n6317 ) | ( n6051 & ~n6318 ) | ( n6317 & ~n6318 ) ;
  assign n6320 = ( x106 & n6314 ) | ( x106 & ~n6319 ) | ( n6314 & ~n6319 ) ;
  assign n6321 = ( x106 & n6052 ) | ( x106 & ~n6069 ) | ( n6052 & ~n6069 ) ;
  assign n6322 = x106 & n6052 ;
  assign n6323 = ( n6057 & n6321 ) | ( n6057 & n6322 ) | ( n6321 & n6322 ) ;
  assign n6324 = ( ~n6057 & n6321 ) | ( ~n6057 & n6322 ) | ( n6321 & n6322 ) ;
  assign n6325 = ( n6057 & ~n6323 ) | ( n6057 & n6324 ) | ( ~n6323 & n6324 ) ;
  assign n6326 = ( x107 & n6320 ) | ( x107 & ~n6325 ) | ( n6320 & ~n6325 ) ;
  assign n6327 = ( x107 & n6058 ) | ( x107 & ~n6069 ) | ( n6058 & ~n6069 ) ;
  assign n6328 = x107 & n6058 ;
  assign n6329 = ( n6063 & n6327 ) | ( n6063 & n6328 ) | ( n6327 & n6328 ) ;
  assign n6330 = ( ~n6063 & n6327 ) | ( ~n6063 & n6328 ) | ( n6327 & n6328 ) ;
  assign n6331 = ( n6063 & ~n6329 ) | ( n6063 & n6330 ) | ( ~n6329 & n6330 ) ;
  assign n6332 = ( x108 & n6326 ) | ( x108 & ~n6331 ) | ( n6326 & ~n6331 ) ;
  assign n6333 = ( x109 & ~n6067 ) | ( x109 & n6332 ) | ( ~n6067 & n6332 ) ;
  assign n6334 = n148 | n6333 ;
  assign n6335 = n6067 & n6334 ;
  assign n6336 = n280 | n6335 ;
  assign n6337 = ( x18 & ~x64 ) | ( x18 & n6334 ) | ( ~x64 & n6334 ) ;
  assign n6338 = ~x18 & n6334 ;
  assign n6339 = ( n6073 & n6337 ) | ( n6073 & ~n6338 ) | ( n6337 & ~n6338 ) ;
  assign n6340 = ~x17 & x64 ;
  assign n6341 = ( x65 & ~n6339 ) | ( x65 & n6340 ) | ( ~n6339 & n6340 ) ;
  assign n6342 = ( x65 & n6073 ) | ( x65 & ~n6334 ) | ( n6073 & ~n6334 ) ;
  assign n6343 = x65 & n6073 ;
  assign n6344 = ( n6072 & n6342 ) | ( n6072 & n6343 ) | ( n6342 & n6343 ) ;
  assign n6345 = ( ~n6072 & n6342 ) | ( ~n6072 & n6343 ) | ( n6342 & n6343 ) ;
  assign n6346 = ( n6072 & ~n6344 ) | ( n6072 & n6345 ) | ( ~n6344 & n6345 ) ;
  assign n6347 = ( x66 & n6341 ) | ( x66 & ~n6346 ) | ( n6341 & ~n6346 ) ;
  assign n6348 = ( x66 & n6074 ) | ( x66 & ~n6334 ) | ( n6074 & ~n6334 ) ;
  assign n6349 = x66 & n6074 ;
  assign n6350 = ( n6079 & n6348 ) | ( n6079 & n6349 ) | ( n6348 & n6349 ) ;
  assign n6351 = ( ~n6079 & n6348 ) | ( ~n6079 & n6349 ) | ( n6348 & n6349 ) ;
  assign n6352 = ( n6079 & ~n6350 ) | ( n6079 & n6351 ) | ( ~n6350 & n6351 ) ;
  assign n6353 = ( x67 & n6347 ) | ( x67 & ~n6352 ) | ( n6347 & ~n6352 ) ;
  assign n6354 = ( x67 & n6080 ) | ( x67 & ~n6334 ) | ( n6080 & ~n6334 ) ;
  assign n6355 = x67 & n6080 ;
  assign n6356 = ( ~n6085 & n6354 ) | ( ~n6085 & n6355 ) | ( n6354 & n6355 ) ;
  assign n6357 = ( n6085 & n6354 ) | ( n6085 & n6355 ) | ( n6354 & n6355 ) ;
  assign n6358 = ( n6085 & n6356 ) | ( n6085 & ~n6357 ) | ( n6356 & ~n6357 ) ;
  assign n6359 = ( x68 & n6353 ) | ( x68 & ~n6358 ) | ( n6353 & ~n6358 ) ;
  assign n6360 = ( x68 & n6086 ) | ( x68 & ~n6334 ) | ( n6086 & ~n6334 ) ;
  assign n6361 = x68 & n6086 ;
  assign n6362 = ( n6091 & n6360 ) | ( n6091 & n6361 ) | ( n6360 & n6361 ) ;
  assign n6363 = ( ~n6091 & n6360 ) | ( ~n6091 & n6361 ) | ( n6360 & n6361 ) ;
  assign n6364 = ( n6091 & ~n6362 ) | ( n6091 & n6363 ) | ( ~n6362 & n6363 ) ;
  assign n6365 = ( x69 & n6359 ) | ( x69 & ~n6364 ) | ( n6359 & ~n6364 ) ;
  assign n6366 = ( x69 & n6092 ) | ( x69 & ~n6334 ) | ( n6092 & ~n6334 ) ;
  assign n6367 = x69 & n6092 ;
  assign n6368 = ( ~n6097 & n6366 ) | ( ~n6097 & n6367 ) | ( n6366 & n6367 ) ;
  assign n6369 = ( n6097 & n6366 ) | ( n6097 & n6367 ) | ( n6366 & n6367 ) ;
  assign n6370 = ( n6097 & n6368 ) | ( n6097 & ~n6369 ) | ( n6368 & ~n6369 ) ;
  assign n6371 = ( x70 & n6365 ) | ( x70 & ~n6370 ) | ( n6365 & ~n6370 ) ;
  assign n6372 = ( x70 & n6098 ) | ( x70 & ~n6334 ) | ( n6098 & ~n6334 ) ;
  assign n6373 = x70 & n6098 ;
  assign n6374 = ( n6103 & n6372 ) | ( n6103 & n6373 ) | ( n6372 & n6373 ) ;
  assign n6375 = ( ~n6103 & n6372 ) | ( ~n6103 & n6373 ) | ( n6372 & n6373 ) ;
  assign n6376 = ( n6103 & ~n6374 ) | ( n6103 & n6375 ) | ( ~n6374 & n6375 ) ;
  assign n6377 = ( x71 & n6371 ) | ( x71 & ~n6376 ) | ( n6371 & ~n6376 ) ;
  assign n6378 = ( x71 & n6104 ) | ( x71 & ~n6334 ) | ( n6104 & ~n6334 ) ;
  assign n6379 = x71 & n6104 ;
  assign n6380 = ( ~n6109 & n6378 ) | ( ~n6109 & n6379 ) | ( n6378 & n6379 ) ;
  assign n6381 = ( n6109 & n6378 ) | ( n6109 & n6379 ) | ( n6378 & n6379 ) ;
  assign n6382 = ( n6109 & n6380 ) | ( n6109 & ~n6381 ) | ( n6380 & ~n6381 ) ;
  assign n6383 = ( x72 & n6377 ) | ( x72 & ~n6382 ) | ( n6377 & ~n6382 ) ;
  assign n6384 = ( x72 & n6110 ) | ( x72 & ~n6334 ) | ( n6110 & ~n6334 ) ;
  assign n6385 = x72 & n6110 ;
  assign n6386 = ( n6115 & n6384 ) | ( n6115 & n6385 ) | ( n6384 & n6385 ) ;
  assign n6387 = ( ~n6115 & n6384 ) | ( ~n6115 & n6385 ) | ( n6384 & n6385 ) ;
  assign n6388 = ( n6115 & ~n6386 ) | ( n6115 & n6387 ) | ( ~n6386 & n6387 ) ;
  assign n6389 = ( x73 & n6383 ) | ( x73 & ~n6388 ) | ( n6383 & ~n6388 ) ;
  assign n6390 = ( x73 & n6116 ) | ( x73 & ~n6334 ) | ( n6116 & ~n6334 ) ;
  assign n6391 = x73 & n6116 ;
  assign n6392 = ( ~n6121 & n6390 ) | ( ~n6121 & n6391 ) | ( n6390 & n6391 ) ;
  assign n6393 = ( n6121 & n6390 ) | ( n6121 & n6391 ) | ( n6390 & n6391 ) ;
  assign n6394 = ( n6121 & n6392 ) | ( n6121 & ~n6393 ) | ( n6392 & ~n6393 ) ;
  assign n6395 = ( x74 & n6389 ) | ( x74 & ~n6394 ) | ( n6389 & ~n6394 ) ;
  assign n6396 = ( x74 & n6122 ) | ( x74 & ~n6334 ) | ( n6122 & ~n6334 ) ;
  assign n6397 = x74 & n6122 ;
  assign n6398 = ( n6127 & n6396 ) | ( n6127 & n6397 ) | ( n6396 & n6397 ) ;
  assign n6399 = ( ~n6127 & n6396 ) | ( ~n6127 & n6397 ) | ( n6396 & n6397 ) ;
  assign n6400 = ( n6127 & ~n6398 ) | ( n6127 & n6399 ) | ( ~n6398 & n6399 ) ;
  assign n6401 = ( x75 & n6395 ) | ( x75 & ~n6400 ) | ( n6395 & ~n6400 ) ;
  assign n6402 = ( x75 & n6128 ) | ( x75 & ~n6334 ) | ( n6128 & ~n6334 ) ;
  assign n6403 = x75 & n6128 ;
  assign n6404 = ( ~n6133 & n6402 ) | ( ~n6133 & n6403 ) | ( n6402 & n6403 ) ;
  assign n6405 = ( n6133 & n6402 ) | ( n6133 & n6403 ) | ( n6402 & n6403 ) ;
  assign n6406 = ( n6133 & n6404 ) | ( n6133 & ~n6405 ) | ( n6404 & ~n6405 ) ;
  assign n6407 = ( x76 & n6401 ) | ( x76 & ~n6406 ) | ( n6401 & ~n6406 ) ;
  assign n6408 = ( x76 & n6134 ) | ( x76 & ~n6334 ) | ( n6134 & ~n6334 ) ;
  assign n6409 = x76 & n6134 ;
  assign n6410 = ( n6139 & n6408 ) | ( n6139 & n6409 ) | ( n6408 & n6409 ) ;
  assign n6411 = ( ~n6139 & n6408 ) | ( ~n6139 & n6409 ) | ( n6408 & n6409 ) ;
  assign n6412 = ( n6139 & ~n6410 ) | ( n6139 & n6411 ) | ( ~n6410 & n6411 ) ;
  assign n6413 = ( x77 & n6407 ) | ( x77 & ~n6412 ) | ( n6407 & ~n6412 ) ;
  assign n6414 = ( x77 & n6140 ) | ( x77 & ~n6334 ) | ( n6140 & ~n6334 ) ;
  assign n6415 = x77 & n6140 ;
  assign n6416 = ( ~n6145 & n6414 ) | ( ~n6145 & n6415 ) | ( n6414 & n6415 ) ;
  assign n6417 = ( n6145 & n6414 ) | ( n6145 & n6415 ) | ( n6414 & n6415 ) ;
  assign n6418 = ( n6145 & n6416 ) | ( n6145 & ~n6417 ) | ( n6416 & ~n6417 ) ;
  assign n6419 = ( x78 & n6413 ) | ( x78 & ~n6418 ) | ( n6413 & ~n6418 ) ;
  assign n6420 = ( x78 & n6146 ) | ( x78 & ~n6334 ) | ( n6146 & ~n6334 ) ;
  assign n6421 = x78 & n6146 ;
  assign n6422 = ( n6151 & n6420 ) | ( n6151 & n6421 ) | ( n6420 & n6421 ) ;
  assign n6423 = ( ~n6151 & n6420 ) | ( ~n6151 & n6421 ) | ( n6420 & n6421 ) ;
  assign n6424 = ( n6151 & ~n6422 ) | ( n6151 & n6423 ) | ( ~n6422 & n6423 ) ;
  assign n6425 = ( x79 & n6419 ) | ( x79 & ~n6424 ) | ( n6419 & ~n6424 ) ;
  assign n6426 = ( x79 & n6152 ) | ( x79 & ~n6334 ) | ( n6152 & ~n6334 ) ;
  assign n6427 = x79 & n6152 ;
  assign n6428 = ( ~n6157 & n6426 ) | ( ~n6157 & n6427 ) | ( n6426 & n6427 ) ;
  assign n6429 = ( n6157 & n6426 ) | ( n6157 & n6427 ) | ( n6426 & n6427 ) ;
  assign n6430 = ( n6157 & n6428 ) | ( n6157 & ~n6429 ) | ( n6428 & ~n6429 ) ;
  assign n6431 = ( x80 & n6425 ) | ( x80 & ~n6430 ) | ( n6425 & ~n6430 ) ;
  assign n6432 = ( x80 & n6158 ) | ( x80 & ~n6334 ) | ( n6158 & ~n6334 ) ;
  assign n6433 = x80 & n6158 ;
  assign n6434 = ( n6163 & n6432 ) | ( n6163 & n6433 ) | ( n6432 & n6433 ) ;
  assign n6435 = ( ~n6163 & n6432 ) | ( ~n6163 & n6433 ) | ( n6432 & n6433 ) ;
  assign n6436 = ( n6163 & ~n6434 ) | ( n6163 & n6435 ) | ( ~n6434 & n6435 ) ;
  assign n6437 = ( x81 & n6431 ) | ( x81 & ~n6436 ) | ( n6431 & ~n6436 ) ;
  assign n6438 = ( x81 & n6164 ) | ( x81 & ~n6334 ) | ( n6164 & ~n6334 ) ;
  assign n6439 = x81 & n6164 ;
  assign n6440 = ( ~n6169 & n6438 ) | ( ~n6169 & n6439 ) | ( n6438 & n6439 ) ;
  assign n6441 = ( n6169 & n6438 ) | ( n6169 & n6439 ) | ( n6438 & n6439 ) ;
  assign n6442 = ( n6169 & n6440 ) | ( n6169 & ~n6441 ) | ( n6440 & ~n6441 ) ;
  assign n6443 = ( x82 & n6437 ) | ( x82 & ~n6442 ) | ( n6437 & ~n6442 ) ;
  assign n6444 = ( x82 & n6170 ) | ( x82 & ~n6334 ) | ( n6170 & ~n6334 ) ;
  assign n6445 = x82 & n6170 ;
  assign n6446 = ( n6175 & n6444 ) | ( n6175 & n6445 ) | ( n6444 & n6445 ) ;
  assign n6447 = ( ~n6175 & n6444 ) | ( ~n6175 & n6445 ) | ( n6444 & n6445 ) ;
  assign n6448 = ( n6175 & ~n6446 ) | ( n6175 & n6447 ) | ( ~n6446 & n6447 ) ;
  assign n6449 = ( x83 & n6443 ) | ( x83 & ~n6448 ) | ( n6443 & ~n6448 ) ;
  assign n6450 = ( x83 & n6176 ) | ( x83 & ~n6334 ) | ( n6176 & ~n6334 ) ;
  assign n6451 = x83 & n6176 ;
  assign n6452 = ( ~n6181 & n6450 ) | ( ~n6181 & n6451 ) | ( n6450 & n6451 ) ;
  assign n6453 = ( n6181 & n6450 ) | ( n6181 & n6451 ) | ( n6450 & n6451 ) ;
  assign n6454 = ( n6181 & n6452 ) | ( n6181 & ~n6453 ) | ( n6452 & ~n6453 ) ;
  assign n6455 = ( x84 & n6449 ) | ( x84 & ~n6454 ) | ( n6449 & ~n6454 ) ;
  assign n6456 = ( x84 & n6182 ) | ( x84 & ~n6334 ) | ( n6182 & ~n6334 ) ;
  assign n6457 = x84 & n6182 ;
  assign n6458 = ( n6187 & n6456 ) | ( n6187 & n6457 ) | ( n6456 & n6457 ) ;
  assign n6459 = ( ~n6187 & n6456 ) | ( ~n6187 & n6457 ) | ( n6456 & n6457 ) ;
  assign n6460 = ( n6187 & ~n6458 ) | ( n6187 & n6459 ) | ( ~n6458 & n6459 ) ;
  assign n6461 = ( x85 & n6455 ) | ( x85 & ~n6460 ) | ( n6455 & ~n6460 ) ;
  assign n6462 = ( x85 & n6188 ) | ( x85 & ~n6334 ) | ( n6188 & ~n6334 ) ;
  assign n6463 = x85 & n6188 ;
  assign n6464 = ( ~n6193 & n6462 ) | ( ~n6193 & n6463 ) | ( n6462 & n6463 ) ;
  assign n6465 = ( n6193 & n6462 ) | ( n6193 & n6463 ) | ( n6462 & n6463 ) ;
  assign n6466 = ( n6193 & n6464 ) | ( n6193 & ~n6465 ) | ( n6464 & ~n6465 ) ;
  assign n6467 = ( x86 & n6461 ) | ( x86 & ~n6466 ) | ( n6461 & ~n6466 ) ;
  assign n6468 = ( x86 & n6194 ) | ( x86 & ~n6334 ) | ( n6194 & ~n6334 ) ;
  assign n6469 = x86 & n6194 ;
  assign n6470 = ( n6199 & n6468 ) | ( n6199 & n6469 ) | ( n6468 & n6469 ) ;
  assign n6471 = ( ~n6199 & n6468 ) | ( ~n6199 & n6469 ) | ( n6468 & n6469 ) ;
  assign n6472 = ( n6199 & ~n6470 ) | ( n6199 & n6471 ) | ( ~n6470 & n6471 ) ;
  assign n6473 = ( x87 & n6467 ) | ( x87 & ~n6472 ) | ( n6467 & ~n6472 ) ;
  assign n6474 = ( x87 & n6200 ) | ( x87 & ~n6334 ) | ( n6200 & ~n6334 ) ;
  assign n6475 = x87 & n6200 ;
  assign n6476 = ( ~n6205 & n6474 ) | ( ~n6205 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6477 = ( n6205 & n6474 ) | ( n6205 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6478 = ( n6205 & n6476 ) | ( n6205 & ~n6477 ) | ( n6476 & ~n6477 ) ;
  assign n6479 = ( x88 & n6473 ) | ( x88 & ~n6478 ) | ( n6473 & ~n6478 ) ;
  assign n6480 = ( x88 & n6206 ) | ( x88 & ~n6334 ) | ( n6206 & ~n6334 ) ;
  assign n6481 = x88 & n6206 ;
  assign n6482 = ( n6211 & n6480 ) | ( n6211 & n6481 ) | ( n6480 & n6481 ) ;
  assign n6483 = ( ~n6211 & n6480 ) | ( ~n6211 & n6481 ) | ( n6480 & n6481 ) ;
  assign n6484 = ( n6211 & ~n6482 ) | ( n6211 & n6483 ) | ( ~n6482 & n6483 ) ;
  assign n6485 = ( x89 & n6479 ) | ( x89 & ~n6484 ) | ( n6479 & ~n6484 ) ;
  assign n6486 = ( x89 & n6212 ) | ( x89 & ~n6334 ) | ( n6212 & ~n6334 ) ;
  assign n6487 = x89 & n6212 ;
  assign n6488 = ( ~n6217 & n6486 ) | ( ~n6217 & n6487 ) | ( n6486 & n6487 ) ;
  assign n6489 = ( n6217 & n6486 ) | ( n6217 & n6487 ) | ( n6486 & n6487 ) ;
  assign n6490 = ( n6217 & n6488 ) | ( n6217 & ~n6489 ) | ( n6488 & ~n6489 ) ;
  assign n6491 = ( x90 & n6485 ) | ( x90 & ~n6490 ) | ( n6485 & ~n6490 ) ;
  assign n6492 = ( x90 & n6218 ) | ( x90 & ~n6334 ) | ( n6218 & ~n6334 ) ;
  assign n6493 = x90 & n6218 ;
  assign n6494 = ( n6223 & n6492 ) | ( n6223 & n6493 ) | ( n6492 & n6493 ) ;
  assign n6495 = ( ~n6223 & n6492 ) | ( ~n6223 & n6493 ) | ( n6492 & n6493 ) ;
  assign n6496 = ( n6223 & ~n6494 ) | ( n6223 & n6495 ) | ( ~n6494 & n6495 ) ;
  assign n6497 = ( x91 & n6491 ) | ( x91 & ~n6496 ) | ( n6491 & ~n6496 ) ;
  assign n6498 = ( x91 & n6224 ) | ( x91 & ~n6334 ) | ( n6224 & ~n6334 ) ;
  assign n6499 = x91 & n6224 ;
  assign n6500 = ( ~n6229 & n6498 ) | ( ~n6229 & n6499 ) | ( n6498 & n6499 ) ;
  assign n6501 = ( n6229 & n6498 ) | ( n6229 & n6499 ) | ( n6498 & n6499 ) ;
  assign n6502 = ( n6229 & n6500 ) | ( n6229 & ~n6501 ) | ( n6500 & ~n6501 ) ;
  assign n6503 = ( x92 & n6497 ) | ( x92 & ~n6502 ) | ( n6497 & ~n6502 ) ;
  assign n6504 = ( x92 & n6230 ) | ( x92 & ~n6334 ) | ( n6230 & ~n6334 ) ;
  assign n6505 = x92 & n6230 ;
  assign n6506 = ( n6235 & n6504 ) | ( n6235 & n6505 ) | ( n6504 & n6505 ) ;
  assign n6507 = ( ~n6235 & n6504 ) | ( ~n6235 & n6505 ) | ( n6504 & n6505 ) ;
  assign n6508 = ( n6235 & ~n6506 ) | ( n6235 & n6507 ) | ( ~n6506 & n6507 ) ;
  assign n6509 = ( x93 & n6503 ) | ( x93 & ~n6508 ) | ( n6503 & ~n6508 ) ;
  assign n6510 = ( x93 & n6236 ) | ( x93 & ~n6334 ) | ( n6236 & ~n6334 ) ;
  assign n6511 = x93 & n6236 ;
  assign n6512 = ( ~n6241 & n6510 ) | ( ~n6241 & n6511 ) | ( n6510 & n6511 ) ;
  assign n6513 = ( n6241 & n6510 ) | ( n6241 & n6511 ) | ( n6510 & n6511 ) ;
  assign n6514 = ( n6241 & n6512 ) | ( n6241 & ~n6513 ) | ( n6512 & ~n6513 ) ;
  assign n6515 = ( x94 & n6509 ) | ( x94 & ~n6514 ) | ( n6509 & ~n6514 ) ;
  assign n6516 = ( x94 & n6242 ) | ( x94 & ~n6334 ) | ( n6242 & ~n6334 ) ;
  assign n6517 = x94 & n6242 ;
  assign n6518 = ( n6247 & n6516 ) | ( n6247 & n6517 ) | ( n6516 & n6517 ) ;
  assign n6519 = ( ~n6247 & n6516 ) | ( ~n6247 & n6517 ) | ( n6516 & n6517 ) ;
  assign n6520 = ( n6247 & ~n6518 ) | ( n6247 & n6519 ) | ( ~n6518 & n6519 ) ;
  assign n6521 = ( x95 & n6515 ) | ( x95 & ~n6520 ) | ( n6515 & ~n6520 ) ;
  assign n6522 = ( x95 & n6248 ) | ( x95 & ~n6334 ) | ( n6248 & ~n6334 ) ;
  assign n6523 = x95 & n6248 ;
  assign n6524 = ( ~n6253 & n6522 ) | ( ~n6253 & n6523 ) | ( n6522 & n6523 ) ;
  assign n6525 = ( n6253 & n6522 ) | ( n6253 & n6523 ) | ( n6522 & n6523 ) ;
  assign n6526 = ( n6253 & n6524 ) | ( n6253 & ~n6525 ) | ( n6524 & ~n6525 ) ;
  assign n6527 = ( x96 & n6521 ) | ( x96 & ~n6526 ) | ( n6521 & ~n6526 ) ;
  assign n6528 = ( x96 & n6254 ) | ( x96 & ~n6334 ) | ( n6254 & ~n6334 ) ;
  assign n6529 = x96 & n6254 ;
  assign n6530 = ( n6259 & n6528 ) | ( n6259 & n6529 ) | ( n6528 & n6529 ) ;
  assign n6531 = ( ~n6259 & n6528 ) | ( ~n6259 & n6529 ) | ( n6528 & n6529 ) ;
  assign n6532 = ( n6259 & ~n6530 ) | ( n6259 & n6531 ) | ( ~n6530 & n6531 ) ;
  assign n6533 = ( x97 & n6527 ) | ( x97 & ~n6532 ) | ( n6527 & ~n6532 ) ;
  assign n6534 = ( x97 & n6260 ) | ( x97 & ~n6334 ) | ( n6260 & ~n6334 ) ;
  assign n6535 = x97 & n6260 ;
  assign n6536 = ( ~n6265 & n6534 ) | ( ~n6265 & n6535 ) | ( n6534 & n6535 ) ;
  assign n6537 = ( n6265 & n6534 ) | ( n6265 & n6535 ) | ( n6534 & n6535 ) ;
  assign n6538 = ( n6265 & n6536 ) | ( n6265 & ~n6537 ) | ( n6536 & ~n6537 ) ;
  assign n6539 = ( x98 & n6533 ) | ( x98 & ~n6538 ) | ( n6533 & ~n6538 ) ;
  assign n6540 = ( x98 & n6266 ) | ( x98 & ~n6334 ) | ( n6266 & ~n6334 ) ;
  assign n6541 = x98 & n6266 ;
  assign n6542 = ( n6271 & n6540 ) | ( n6271 & n6541 ) | ( n6540 & n6541 ) ;
  assign n6543 = ( ~n6271 & n6540 ) | ( ~n6271 & n6541 ) | ( n6540 & n6541 ) ;
  assign n6544 = ( n6271 & ~n6542 ) | ( n6271 & n6543 ) | ( ~n6542 & n6543 ) ;
  assign n6545 = ( x99 & n6539 ) | ( x99 & ~n6544 ) | ( n6539 & ~n6544 ) ;
  assign n6546 = ( x99 & n6272 ) | ( x99 & ~n6334 ) | ( n6272 & ~n6334 ) ;
  assign n6547 = x99 & n6272 ;
  assign n6548 = ( ~n6277 & n6546 ) | ( ~n6277 & n6547 ) | ( n6546 & n6547 ) ;
  assign n6549 = ( n6277 & n6546 ) | ( n6277 & n6547 ) | ( n6546 & n6547 ) ;
  assign n6550 = ( n6277 & n6548 ) | ( n6277 & ~n6549 ) | ( n6548 & ~n6549 ) ;
  assign n6551 = ( x100 & n6545 ) | ( x100 & ~n6550 ) | ( n6545 & ~n6550 ) ;
  assign n6552 = ( x100 & n6278 ) | ( x100 & ~n6334 ) | ( n6278 & ~n6334 ) ;
  assign n6553 = x100 & n6278 ;
  assign n6554 = ( n6283 & n6552 ) | ( n6283 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6555 = ( ~n6283 & n6552 ) | ( ~n6283 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6556 = ( n6283 & ~n6554 ) | ( n6283 & n6555 ) | ( ~n6554 & n6555 ) ;
  assign n6557 = ( x101 & n6551 ) | ( x101 & ~n6556 ) | ( n6551 & ~n6556 ) ;
  assign n6558 = ( x101 & n6284 ) | ( x101 & ~n6334 ) | ( n6284 & ~n6334 ) ;
  assign n6559 = x101 & n6284 ;
  assign n6560 = ( ~n6289 & n6558 ) | ( ~n6289 & n6559 ) | ( n6558 & n6559 ) ;
  assign n6561 = ( n6289 & n6558 ) | ( n6289 & n6559 ) | ( n6558 & n6559 ) ;
  assign n6562 = ( n6289 & n6560 ) | ( n6289 & ~n6561 ) | ( n6560 & ~n6561 ) ;
  assign n6563 = ( x102 & n6557 ) | ( x102 & ~n6562 ) | ( n6557 & ~n6562 ) ;
  assign n6564 = ( x102 & n6290 ) | ( x102 & ~n6334 ) | ( n6290 & ~n6334 ) ;
  assign n6565 = x102 & n6290 ;
  assign n6566 = ( n6295 & n6564 ) | ( n6295 & n6565 ) | ( n6564 & n6565 ) ;
  assign n6567 = ( ~n6295 & n6564 ) | ( ~n6295 & n6565 ) | ( n6564 & n6565 ) ;
  assign n6568 = ( n6295 & ~n6566 ) | ( n6295 & n6567 ) | ( ~n6566 & n6567 ) ;
  assign n6569 = ( x103 & n6563 ) | ( x103 & ~n6568 ) | ( n6563 & ~n6568 ) ;
  assign n6570 = ( x103 & n6296 ) | ( x103 & ~n6334 ) | ( n6296 & ~n6334 ) ;
  assign n6571 = x103 & n6296 ;
  assign n6572 = ( ~n6301 & n6570 ) | ( ~n6301 & n6571 ) | ( n6570 & n6571 ) ;
  assign n6573 = ( n6301 & n6570 ) | ( n6301 & n6571 ) | ( n6570 & n6571 ) ;
  assign n6574 = ( n6301 & n6572 ) | ( n6301 & ~n6573 ) | ( n6572 & ~n6573 ) ;
  assign n6575 = ( x104 & n6569 ) | ( x104 & ~n6574 ) | ( n6569 & ~n6574 ) ;
  assign n6576 = ( x104 & n6302 ) | ( x104 & ~n6334 ) | ( n6302 & ~n6334 ) ;
  assign n6577 = x104 & n6302 ;
  assign n6578 = ( n6307 & n6576 ) | ( n6307 & n6577 ) | ( n6576 & n6577 ) ;
  assign n6579 = ( ~n6307 & n6576 ) | ( ~n6307 & n6577 ) | ( n6576 & n6577 ) ;
  assign n6580 = ( n6307 & ~n6578 ) | ( n6307 & n6579 ) | ( ~n6578 & n6579 ) ;
  assign n6581 = ( x105 & n6575 ) | ( x105 & ~n6580 ) | ( n6575 & ~n6580 ) ;
  assign n6582 = ( x105 & n6308 ) | ( x105 & ~n6334 ) | ( n6308 & ~n6334 ) ;
  assign n6583 = x105 & n6308 ;
  assign n6584 = ( ~n6313 & n6582 ) | ( ~n6313 & n6583 ) | ( n6582 & n6583 ) ;
  assign n6585 = ( n6313 & n6582 ) | ( n6313 & n6583 ) | ( n6582 & n6583 ) ;
  assign n6586 = ( n6313 & n6584 ) | ( n6313 & ~n6585 ) | ( n6584 & ~n6585 ) ;
  assign n6587 = ( x106 & n6581 ) | ( x106 & ~n6586 ) | ( n6581 & ~n6586 ) ;
  assign n6588 = ( x106 & n6314 ) | ( x106 & ~n6334 ) | ( n6314 & ~n6334 ) ;
  assign n6589 = x106 & n6314 ;
  assign n6590 = ( n6319 & n6588 ) | ( n6319 & n6589 ) | ( n6588 & n6589 ) ;
  assign n6591 = ( ~n6319 & n6588 ) | ( ~n6319 & n6589 ) | ( n6588 & n6589 ) ;
  assign n6592 = ( n6319 & ~n6590 ) | ( n6319 & n6591 ) | ( ~n6590 & n6591 ) ;
  assign n6593 = ( x107 & n6587 ) | ( x107 & ~n6592 ) | ( n6587 & ~n6592 ) ;
  assign n6594 = ( x107 & n6320 ) | ( x107 & ~n6334 ) | ( n6320 & ~n6334 ) ;
  assign n6595 = x107 & n6320 ;
  assign n6596 = ( ~n6325 & n6594 ) | ( ~n6325 & n6595 ) | ( n6594 & n6595 ) ;
  assign n6597 = ( n6325 & n6594 ) | ( n6325 & n6595 ) | ( n6594 & n6595 ) ;
  assign n6598 = ( n6325 & n6596 ) | ( n6325 & ~n6597 ) | ( n6596 & ~n6597 ) ;
  assign n6599 = ( x108 & n6593 ) | ( x108 & ~n6598 ) | ( n6593 & ~n6598 ) ;
  assign n6600 = ( x108 & n6326 ) | ( x108 & ~n6334 ) | ( n6326 & ~n6334 ) ;
  assign n6601 = x108 & n6326 ;
  assign n6602 = ( ~n6331 & n6600 ) | ( ~n6331 & n6601 ) | ( n6600 & n6601 ) ;
  assign n6603 = ( n6331 & n6600 ) | ( n6331 & n6601 ) | ( n6600 & n6601 ) ;
  assign n6604 = ( n6331 & n6602 ) | ( n6331 & ~n6603 ) | ( n6602 & ~n6603 ) ;
  assign n6605 = ( x109 & n6599 ) | ( x109 & ~n6604 ) | ( n6599 & ~n6604 ) ;
  assign n6606 = x110 | n6605 ;
  assign n6607 = ( x110 & n147 ) | ( x110 & n6605 ) | ( n147 & n6605 ) ;
  assign n6608 = ( n6336 & ~n6606 ) | ( n6336 & n6607 ) | ( ~n6606 & n6607 ) ;
  assign n6609 = ( x110 & ~n6336 ) | ( x110 & n6605 ) | ( ~n6336 & n6605 ) ;
  assign n6610 = n147 | n6609 ;
  assign n6611 = ( x17 & ~x64 ) | ( x17 & n6610 ) | ( ~x64 & n6610 ) ;
  assign n6612 = ~x17 & n6610 ;
  assign n6613 = ( n6340 & n6611 ) | ( n6340 & ~n6612 ) | ( n6611 & ~n6612 ) ;
  assign n6614 = ~x16 & x64 ;
  assign n6615 = ( x65 & ~n6613 ) | ( x65 & n6614 ) | ( ~n6613 & n6614 ) ;
  assign n6616 = ( x65 & n6340 ) | ( x65 & ~n6610 ) | ( n6340 & ~n6610 ) ;
  assign n6617 = x65 & n6340 ;
  assign n6618 = ( n6339 & n6616 ) | ( n6339 & n6617 ) | ( n6616 & n6617 ) ;
  assign n6619 = ( ~n6339 & n6616 ) | ( ~n6339 & n6617 ) | ( n6616 & n6617 ) ;
  assign n6620 = ( n6339 & ~n6618 ) | ( n6339 & n6619 ) | ( ~n6618 & n6619 ) ;
  assign n6621 = ( x66 & n6615 ) | ( x66 & ~n6620 ) | ( n6615 & ~n6620 ) ;
  assign n6622 = ( x66 & n6341 ) | ( x66 & ~n6610 ) | ( n6341 & ~n6610 ) ;
  assign n6623 = x66 & n6341 ;
  assign n6624 = ( n6346 & n6622 ) | ( n6346 & n6623 ) | ( n6622 & n6623 ) ;
  assign n6625 = ( ~n6346 & n6622 ) | ( ~n6346 & n6623 ) | ( n6622 & n6623 ) ;
  assign n6626 = ( n6346 & ~n6624 ) | ( n6346 & n6625 ) | ( ~n6624 & n6625 ) ;
  assign n6627 = ( x67 & n6621 ) | ( x67 & ~n6626 ) | ( n6621 & ~n6626 ) ;
  assign n6628 = ( x67 & n6347 ) | ( x67 & ~n6610 ) | ( n6347 & ~n6610 ) ;
  assign n6629 = x67 & n6347 ;
  assign n6630 = ( ~n6352 & n6628 ) | ( ~n6352 & n6629 ) | ( n6628 & n6629 ) ;
  assign n6631 = ( n6352 & n6628 ) | ( n6352 & n6629 ) | ( n6628 & n6629 ) ;
  assign n6632 = ( n6352 & n6630 ) | ( n6352 & ~n6631 ) | ( n6630 & ~n6631 ) ;
  assign n6633 = ( x68 & n6627 ) | ( x68 & ~n6632 ) | ( n6627 & ~n6632 ) ;
  assign n6634 = ( x68 & n6353 ) | ( x68 & ~n6610 ) | ( n6353 & ~n6610 ) ;
  assign n6635 = x68 & n6353 ;
  assign n6636 = ( n6358 & n6634 ) | ( n6358 & n6635 ) | ( n6634 & n6635 ) ;
  assign n6637 = ( ~n6358 & n6634 ) | ( ~n6358 & n6635 ) | ( n6634 & n6635 ) ;
  assign n6638 = ( n6358 & ~n6636 ) | ( n6358 & n6637 ) | ( ~n6636 & n6637 ) ;
  assign n6639 = ( x69 & n6633 ) | ( x69 & ~n6638 ) | ( n6633 & ~n6638 ) ;
  assign n6640 = ( x69 & n6359 ) | ( x69 & ~n6610 ) | ( n6359 & ~n6610 ) ;
  assign n6641 = x69 & n6359 ;
  assign n6642 = ( ~n6364 & n6640 ) | ( ~n6364 & n6641 ) | ( n6640 & n6641 ) ;
  assign n6643 = ( n6364 & n6640 ) | ( n6364 & n6641 ) | ( n6640 & n6641 ) ;
  assign n6644 = ( n6364 & n6642 ) | ( n6364 & ~n6643 ) | ( n6642 & ~n6643 ) ;
  assign n6645 = ( x70 & n6639 ) | ( x70 & ~n6644 ) | ( n6639 & ~n6644 ) ;
  assign n6646 = ( x70 & n6365 ) | ( x70 & ~n6610 ) | ( n6365 & ~n6610 ) ;
  assign n6647 = x70 & n6365 ;
  assign n6648 = ( n6370 & n6646 ) | ( n6370 & n6647 ) | ( n6646 & n6647 ) ;
  assign n6649 = ( ~n6370 & n6646 ) | ( ~n6370 & n6647 ) | ( n6646 & n6647 ) ;
  assign n6650 = ( n6370 & ~n6648 ) | ( n6370 & n6649 ) | ( ~n6648 & n6649 ) ;
  assign n6651 = ( x71 & n6645 ) | ( x71 & ~n6650 ) | ( n6645 & ~n6650 ) ;
  assign n6652 = ( x71 & n6371 ) | ( x71 & ~n6610 ) | ( n6371 & ~n6610 ) ;
  assign n6653 = x71 & n6371 ;
  assign n6654 = ( ~n6376 & n6652 ) | ( ~n6376 & n6653 ) | ( n6652 & n6653 ) ;
  assign n6655 = ( n6376 & n6652 ) | ( n6376 & n6653 ) | ( n6652 & n6653 ) ;
  assign n6656 = ( n6376 & n6654 ) | ( n6376 & ~n6655 ) | ( n6654 & ~n6655 ) ;
  assign n6657 = ( x72 & n6651 ) | ( x72 & ~n6656 ) | ( n6651 & ~n6656 ) ;
  assign n6658 = ( x72 & n6377 ) | ( x72 & ~n6610 ) | ( n6377 & ~n6610 ) ;
  assign n6659 = x72 & n6377 ;
  assign n6660 = ( n6382 & n6658 ) | ( n6382 & n6659 ) | ( n6658 & n6659 ) ;
  assign n6661 = ( ~n6382 & n6658 ) | ( ~n6382 & n6659 ) | ( n6658 & n6659 ) ;
  assign n6662 = ( n6382 & ~n6660 ) | ( n6382 & n6661 ) | ( ~n6660 & n6661 ) ;
  assign n6663 = ( x73 & n6657 ) | ( x73 & ~n6662 ) | ( n6657 & ~n6662 ) ;
  assign n6664 = ( x73 & n6383 ) | ( x73 & ~n6610 ) | ( n6383 & ~n6610 ) ;
  assign n6665 = x73 & n6383 ;
  assign n6666 = ( ~n6388 & n6664 ) | ( ~n6388 & n6665 ) | ( n6664 & n6665 ) ;
  assign n6667 = ( n6388 & n6664 ) | ( n6388 & n6665 ) | ( n6664 & n6665 ) ;
  assign n6668 = ( n6388 & n6666 ) | ( n6388 & ~n6667 ) | ( n6666 & ~n6667 ) ;
  assign n6669 = ( x74 & n6663 ) | ( x74 & ~n6668 ) | ( n6663 & ~n6668 ) ;
  assign n6670 = ( x74 & n6389 ) | ( x74 & ~n6610 ) | ( n6389 & ~n6610 ) ;
  assign n6671 = x74 & n6389 ;
  assign n6672 = ( n6394 & n6670 ) | ( n6394 & n6671 ) | ( n6670 & n6671 ) ;
  assign n6673 = ( ~n6394 & n6670 ) | ( ~n6394 & n6671 ) | ( n6670 & n6671 ) ;
  assign n6674 = ( n6394 & ~n6672 ) | ( n6394 & n6673 ) | ( ~n6672 & n6673 ) ;
  assign n6675 = ( x75 & n6669 ) | ( x75 & ~n6674 ) | ( n6669 & ~n6674 ) ;
  assign n6676 = ( x75 & n6395 ) | ( x75 & ~n6610 ) | ( n6395 & ~n6610 ) ;
  assign n6677 = x75 & n6395 ;
  assign n6678 = ( ~n6400 & n6676 ) | ( ~n6400 & n6677 ) | ( n6676 & n6677 ) ;
  assign n6679 = ( n6400 & n6676 ) | ( n6400 & n6677 ) | ( n6676 & n6677 ) ;
  assign n6680 = ( n6400 & n6678 ) | ( n6400 & ~n6679 ) | ( n6678 & ~n6679 ) ;
  assign n6681 = ( x76 & n6675 ) | ( x76 & ~n6680 ) | ( n6675 & ~n6680 ) ;
  assign n6682 = ( x76 & n6401 ) | ( x76 & ~n6610 ) | ( n6401 & ~n6610 ) ;
  assign n6683 = x76 & n6401 ;
  assign n6684 = ( n6406 & n6682 ) | ( n6406 & n6683 ) | ( n6682 & n6683 ) ;
  assign n6685 = ( ~n6406 & n6682 ) | ( ~n6406 & n6683 ) | ( n6682 & n6683 ) ;
  assign n6686 = ( n6406 & ~n6684 ) | ( n6406 & n6685 ) | ( ~n6684 & n6685 ) ;
  assign n6687 = ( x77 & n6681 ) | ( x77 & ~n6686 ) | ( n6681 & ~n6686 ) ;
  assign n6688 = ( x77 & n6407 ) | ( x77 & ~n6610 ) | ( n6407 & ~n6610 ) ;
  assign n6689 = x77 & n6407 ;
  assign n6690 = ( ~n6412 & n6688 ) | ( ~n6412 & n6689 ) | ( n6688 & n6689 ) ;
  assign n6691 = ( n6412 & n6688 ) | ( n6412 & n6689 ) | ( n6688 & n6689 ) ;
  assign n6692 = ( n6412 & n6690 ) | ( n6412 & ~n6691 ) | ( n6690 & ~n6691 ) ;
  assign n6693 = ( x78 & n6687 ) | ( x78 & ~n6692 ) | ( n6687 & ~n6692 ) ;
  assign n6694 = ( x78 & n6413 ) | ( x78 & ~n6610 ) | ( n6413 & ~n6610 ) ;
  assign n6695 = x78 & n6413 ;
  assign n6696 = ( n6418 & n6694 ) | ( n6418 & n6695 ) | ( n6694 & n6695 ) ;
  assign n6697 = ( ~n6418 & n6694 ) | ( ~n6418 & n6695 ) | ( n6694 & n6695 ) ;
  assign n6698 = ( n6418 & ~n6696 ) | ( n6418 & n6697 ) | ( ~n6696 & n6697 ) ;
  assign n6699 = ( x79 & n6693 ) | ( x79 & ~n6698 ) | ( n6693 & ~n6698 ) ;
  assign n6700 = ( x79 & n6419 ) | ( x79 & ~n6610 ) | ( n6419 & ~n6610 ) ;
  assign n6701 = x79 & n6419 ;
  assign n6702 = ( ~n6424 & n6700 ) | ( ~n6424 & n6701 ) | ( n6700 & n6701 ) ;
  assign n6703 = ( n6424 & n6700 ) | ( n6424 & n6701 ) | ( n6700 & n6701 ) ;
  assign n6704 = ( n6424 & n6702 ) | ( n6424 & ~n6703 ) | ( n6702 & ~n6703 ) ;
  assign n6705 = ( x80 & n6699 ) | ( x80 & ~n6704 ) | ( n6699 & ~n6704 ) ;
  assign n6706 = ( x80 & n6425 ) | ( x80 & ~n6610 ) | ( n6425 & ~n6610 ) ;
  assign n6707 = x80 & n6425 ;
  assign n6708 = ( n6430 & n6706 ) | ( n6430 & n6707 ) | ( n6706 & n6707 ) ;
  assign n6709 = ( ~n6430 & n6706 ) | ( ~n6430 & n6707 ) | ( n6706 & n6707 ) ;
  assign n6710 = ( n6430 & ~n6708 ) | ( n6430 & n6709 ) | ( ~n6708 & n6709 ) ;
  assign n6711 = ( x81 & n6705 ) | ( x81 & ~n6710 ) | ( n6705 & ~n6710 ) ;
  assign n6712 = ( x81 & n6431 ) | ( x81 & ~n6610 ) | ( n6431 & ~n6610 ) ;
  assign n6713 = x81 & n6431 ;
  assign n6714 = ( ~n6436 & n6712 ) | ( ~n6436 & n6713 ) | ( n6712 & n6713 ) ;
  assign n6715 = ( n6436 & n6712 ) | ( n6436 & n6713 ) | ( n6712 & n6713 ) ;
  assign n6716 = ( n6436 & n6714 ) | ( n6436 & ~n6715 ) | ( n6714 & ~n6715 ) ;
  assign n6717 = ( x82 & n6711 ) | ( x82 & ~n6716 ) | ( n6711 & ~n6716 ) ;
  assign n6718 = ( x82 & n6437 ) | ( x82 & ~n6610 ) | ( n6437 & ~n6610 ) ;
  assign n6719 = x82 & n6437 ;
  assign n6720 = ( n6442 & n6718 ) | ( n6442 & n6719 ) | ( n6718 & n6719 ) ;
  assign n6721 = ( ~n6442 & n6718 ) | ( ~n6442 & n6719 ) | ( n6718 & n6719 ) ;
  assign n6722 = ( n6442 & ~n6720 ) | ( n6442 & n6721 ) | ( ~n6720 & n6721 ) ;
  assign n6723 = ( x83 & n6717 ) | ( x83 & ~n6722 ) | ( n6717 & ~n6722 ) ;
  assign n6724 = ( x83 & n6443 ) | ( x83 & ~n6610 ) | ( n6443 & ~n6610 ) ;
  assign n6725 = x83 & n6443 ;
  assign n6726 = ( ~n6448 & n6724 ) | ( ~n6448 & n6725 ) | ( n6724 & n6725 ) ;
  assign n6727 = ( n6448 & n6724 ) | ( n6448 & n6725 ) | ( n6724 & n6725 ) ;
  assign n6728 = ( n6448 & n6726 ) | ( n6448 & ~n6727 ) | ( n6726 & ~n6727 ) ;
  assign n6729 = ( x84 & n6723 ) | ( x84 & ~n6728 ) | ( n6723 & ~n6728 ) ;
  assign n6730 = ( x84 & n6449 ) | ( x84 & ~n6610 ) | ( n6449 & ~n6610 ) ;
  assign n6731 = x84 & n6449 ;
  assign n6732 = ( n6454 & n6730 ) | ( n6454 & n6731 ) | ( n6730 & n6731 ) ;
  assign n6733 = ( ~n6454 & n6730 ) | ( ~n6454 & n6731 ) | ( n6730 & n6731 ) ;
  assign n6734 = ( n6454 & ~n6732 ) | ( n6454 & n6733 ) | ( ~n6732 & n6733 ) ;
  assign n6735 = ( x85 & n6729 ) | ( x85 & ~n6734 ) | ( n6729 & ~n6734 ) ;
  assign n6736 = ( x85 & n6455 ) | ( x85 & ~n6610 ) | ( n6455 & ~n6610 ) ;
  assign n6737 = x85 & n6455 ;
  assign n6738 = ( ~n6460 & n6736 ) | ( ~n6460 & n6737 ) | ( n6736 & n6737 ) ;
  assign n6739 = ( n6460 & n6736 ) | ( n6460 & n6737 ) | ( n6736 & n6737 ) ;
  assign n6740 = ( n6460 & n6738 ) | ( n6460 & ~n6739 ) | ( n6738 & ~n6739 ) ;
  assign n6741 = ( x86 & n6735 ) | ( x86 & ~n6740 ) | ( n6735 & ~n6740 ) ;
  assign n6742 = ( x86 & n6461 ) | ( x86 & ~n6610 ) | ( n6461 & ~n6610 ) ;
  assign n6743 = x86 & n6461 ;
  assign n6744 = ( n6466 & n6742 ) | ( n6466 & n6743 ) | ( n6742 & n6743 ) ;
  assign n6745 = ( ~n6466 & n6742 ) | ( ~n6466 & n6743 ) | ( n6742 & n6743 ) ;
  assign n6746 = ( n6466 & ~n6744 ) | ( n6466 & n6745 ) | ( ~n6744 & n6745 ) ;
  assign n6747 = ( x87 & n6741 ) | ( x87 & ~n6746 ) | ( n6741 & ~n6746 ) ;
  assign n6748 = ( x87 & n6467 ) | ( x87 & ~n6610 ) | ( n6467 & ~n6610 ) ;
  assign n6749 = x87 & n6467 ;
  assign n6750 = ( ~n6472 & n6748 ) | ( ~n6472 & n6749 ) | ( n6748 & n6749 ) ;
  assign n6751 = ( n6472 & n6748 ) | ( n6472 & n6749 ) | ( n6748 & n6749 ) ;
  assign n6752 = ( n6472 & n6750 ) | ( n6472 & ~n6751 ) | ( n6750 & ~n6751 ) ;
  assign n6753 = ( x88 & n6747 ) | ( x88 & ~n6752 ) | ( n6747 & ~n6752 ) ;
  assign n6754 = ( x88 & n6473 ) | ( x88 & ~n6610 ) | ( n6473 & ~n6610 ) ;
  assign n6755 = x88 & n6473 ;
  assign n6756 = ( n6478 & n6754 ) | ( n6478 & n6755 ) | ( n6754 & n6755 ) ;
  assign n6757 = ( ~n6478 & n6754 ) | ( ~n6478 & n6755 ) | ( n6754 & n6755 ) ;
  assign n6758 = ( n6478 & ~n6756 ) | ( n6478 & n6757 ) | ( ~n6756 & n6757 ) ;
  assign n6759 = ( x89 & n6753 ) | ( x89 & ~n6758 ) | ( n6753 & ~n6758 ) ;
  assign n6760 = ( x89 & n6479 ) | ( x89 & ~n6610 ) | ( n6479 & ~n6610 ) ;
  assign n6761 = x89 & n6479 ;
  assign n6762 = ( ~n6484 & n6760 ) | ( ~n6484 & n6761 ) | ( n6760 & n6761 ) ;
  assign n6763 = ( n6484 & n6760 ) | ( n6484 & n6761 ) | ( n6760 & n6761 ) ;
  assign n6764 = ( n6484 & n6762 ) | ( n6484 & ~n6763 ) | ( n6762 & ~n6763 ) ;
  assign n6765 = ( x90 & n6759 ) | ( x90 & ~n6764 ) | ( n6759 & ~n6764 ) ;
  assign n6766 = ( x90 & n6485 ) | ( x90 & ~n6610 ) | ( n6485 & ~n6610 ) ;
  assign n6767 = x90 & n6485 ;
  assign n6768 = ( n6490 & n6766 ) | ( n6490 & n6767 ) | ( n6766 & n6767 ) ;
  assign n6769 = ( ~n6490 & n6766 ) | ( ~n6490 & n6767 ) | ( n6766 & n6767 ) ;
  assign n6770 = ( n6490 & ~n6768 ) | ( n6490 & n6769 ) | ( ~n6768 & n6769 ) ;
  assign n6771 = ( x91 & n6765 ) | ( x91 & ~n6770 ) | ( n6765 & ~n6770 ) ;
  assign n6772 = ( x91 & n6491 ) | ( x91 & ~n6610 ) | ( n6491 & ~n6610 ) ;
  assign n6773 = x91 & n6491 ;
  assign n6774 = ( ~n6496 & n6772 ) | ( ~n6496 & n6773 ) | ( n6772 & n6773 ) ;
  assign n6775 = ( n6496 & n6772 ) | ( n6496 & n6773 ) | ( n6772 & n6773 ) ;
  assign n6776 = ( n6496 & n6774 ) | ( n6496 & ~n6775 ) | ( n6774 & ~n6775 ) ;
  assign n6777 = ( x92 & n6771 ) | ( x92 & ~n6776 ) | ( n6771 & ~n6776 ) ;
  assign n6778 = ( x92 & n6497 ) | ( x92 & ~n6610 ) | ( n6497 & ~n6610 ) ;
  assign n6779 = x92 & n6497 ;
  assign n6780 = ( n6502 & n6778 ) | ( n6502 & n6779 ) | ( n6778 & n6779 ) ;
  assign n6781 = ( ~n6502 & n6778 ) | ( ~n6502 & n6779 ) | ( n6778 & n6779 ) ;
  assign n6782 = ( n6502 & ~n6780 ) | ( n6502 & n6781 ) | ( ~n6780 & n6781 ) ;
  assign n6783 = ( x93 & n6777 ) | ( x93 & ~n6782 ) | ( n6777 & ~n6782 ) ;
  assign n6784 = ( x93 & n6503 ) | ( x93 & ~n6610 ) | ( n6503 & ~n6610 ) ;
  assign n6785 = x93 & n6503 ;
  assign n6786 = ( ~n6508 & n6784 ) | ( ~n6508 & n6785 ) | ( n6784 & n6785 ) ;
  assign n6787 = ( n6508 & n6784 ) | ( n6508 & n6785 ) | ( n6784 & n6785 ) ;
  assign n6788 = ( n6508 & n6786 ) | ( n6508 & ~n6787 ) | ( n6786 & ~n6787 ) ;
  assign n6789 = ( x94 & n6783 ) | ( x94 & ~n6788 ) | ( n6783 & ~n6788 ) ;
  assign n6790 = ( x94 & n6509 ) | ( x94 & ~n6610 ) | ( n6509 & ~n6610 ) ;
  assign n6791 = x94 & n6509 ;
  assign n6792 = ( n6514 & n6790 ) | ( n6514 & n6791 ) | ( n6790 & n6791 ) ;
  assign n6793 = ( ~n6514 & n6790 ) | ( ~n6514 & n6791 ) | ( n6790 & n6791 ) ;
  assign n6794 = ( n6514 & ~n6792 ) | ( n6514 & n6793 ) | ( ~n6792 & n6793 ) ;
  assign n6795 = ( x95 & n6789 ) | ( x95 & ~n6794 ) | ( n6789 & ~n6794 ) ;
  assign n6796 = ( x95 & n6515 ) | ( x95 & ~n6610 ) | ( n6515 & ~n6610 ) ;
  assign n6797 = x95 & n6515 ;
  assign n6798 = ( ~n6520 & n6796 ) | ( ~n6520 & n6797 ) | ( n6796 & n6797 ) ;
  assign n6799 = ( n6520 & n6796 ) | ( n6520 & n6797 ) | ( n6796 & n6797 ) ;
  assign n6800 = ( n6520 & n6798 ) | ( n6520 & ~n6799 ) | ( n6798 & ~n6799 ) ;
  assign n6801 = ( x96 & n6795 ) | ( x96 & ~n6800 ) | ( n6795 & ~n6800 ) ;
  assign n6802 = ( x96 & n6521 ) | ( x96 & ~n6610 ) | ( n6521 & ~n6610 ) ;
  assign n6803 = x96 & n6521 ;
  assign n6804 = ( n6526 & n6802 ) | ( n6526 & n6803 ) | ( n6802 & n6803 ) ;
  assign n6805 = ( ~n6526 & n6802 ) | ( ~n6526 & n6803 ) | ( n6802 & n6803 ) ;
  assign n6806 = ( n6526 & ~n6804 ) | ( n6526 & n6805 ) | ( ~n6804 & n6805 ) ;
  assign n6807 = ( x97 & n6801 ) | ( x97 & ~n6806 ) | ( n6801 & ~n6806 ) ;
  assign n6808 = ( x97 & n6527 ) | ( x97 & ~n6610 ) | ( n6527 & ~n6610 ) ;
  assign n6809 = x97 & n6527 ;
  assign n6810 = ( ~n6532 & n6808 ) | ( ~n6532 & n6809 ) | ( n6808 & n6809 ) ;
  assign n6811 = ( n6532 & n6808 ) | ( n6532 & n6809 ) | ( n6808 & n6809 ) ;
  assign n6812 = ( n6532 & n6810 ) | ( n6532 & ~n6811 ) | ( n6810 & ~n6811 ) ;
  assign n6813 = ( x98 & n6807 ) | ( x98 & ~n6812 ) | ( n6807 & ~n6812 ) ;
  assign n6814 = ( x98 & n6533 ) | ( x98 & ~n6610 ) | ( n6533 & ~n6610 ) ;
  assign n6815 = x98 & n6533 ;
  assign n6816 = ( n6538 & n6814 ) | ( n6538 & n6815 ) | ( n6814 & n6815 ) ;
  assign n6817 = ( ~n6538 & n6814 ) | ( ~n6538 & n6815 ) | ( n6814 & n6815 ) ;
  assign n6818 = ( n6538 & ~n6816 ) | ( n6538 & n6817 ) | ( ~n6816 & n6817 ) ;
  assign n6819 = ( x99 & n6813 ) | ( x99 & ~n6818 ) | ( n6813 & ~n6818 ) ;
  assign n6820 = ( x99 & n6539 ) | ( x99 & ~n6610 ) | ( n6539 & ~n6610 ) ;
  assign n6821 = x99 & n6539 ;
  assign n6822 = ( ~n6544 & n6820 ) | ( ~n6544 & n6821 ) | ( n6820 & n6821 ) ;
  assign n6823 = ( n6544 & n6820 ) | ( n6544 & n6821 ) | ( n6820 & n6821 ) ;
  assign n6824 = ( n6544 & n6822 ) | ( n6544 & ~n6823 ) | ( n6822 & ~n6823 ) ;
  assign n6825 = ( x100 & n6819 ) | ( x100 & ~n6824 ) | ( n6819 & ~n6824 ) ;
  assign n6826 = ( x100 & n6545 ) | ( x100 & ~n6610 ) | ( n6545 & ~n6610 ) ;
  assign n6827 = x100 & n6545 ;
  assign n6828 = ( n6550 & n6826 ) | ( n6550 & n6827 ) | ( n6826 & n6827 ) ;
  assign n6829 = ( ~n6550 & n6826 ) | ( ~n6550 & n6827 ) | ( n6826 & n6827 ) ;
  assign n6830 = ( n6550 & ~n6828 ) | ( n6550 & n6829 ) | ( ~n6828 & n6829 ) ;
  assign n6831 = ( x101 & n6825 ) | ( x101 & ~n6830 ) | ( n6825 & ~n6830 ) ;
  assign n6832 = ( x101 & n6551 ) | ( x101 & ~n6610 ) | ( n6551 & ~n6610 ) ;
  assign n6833 = x101 & n6551 ;
  assign n6834 = ( ~n6556 & n6832 ) | ( ~n6556 & n6833 ) | ( n6832 & n6833 ) ;
  assign n6835 = ( n6556 & n6832 ) | ( n6556 & n6833 ) | ( n6832 & n6833 ) ;
  assign n6836 = ( n6556 & n6834 ) | ( n6556 & ~n6835 ) | ( n6834 & ~n6835 ) ;
  assign n6837 = ( x102 & n6831 ) | ( x102 & ~n6836 ) | ( n6831 & ~n6836 ) ;
  assign n6838 = ( x102 & n6557 ) | ( x102 & ~n6610 ) | ( n6557 & ~n6610 ) ;
  assign n6839 = x102 & n6557 ;
  assign n6840 = ( n6562 & n6838 ) | ( n6562 & n6839 ) | ( n6838 & n6839 ) ;
  assign n6841 = ( ~n6562 & n6838 ) | ( ~n6562 & n6839 ) | ( n6838 & n6839 ) ;
  assign n6842 = ( n6562 & ~n6840 ) | ( n6562 & n6841 ) | ( ~n6840 & n6841 ) ;
  assign n6843 = ( x103 & n6837 ) | ( x103 & ~n6842 ) | ( n6837 & ~n6842 ) ;
  assign n6844 = ( x103 & n6563 ) | ( x103 & ~n6610 ) | ( n6563 & ~n6610 ) ;
  assign n6845 = x103 & n6563 ;
  assign n6846 = ( ~n6568 & n6844 ) | ( ~n6568 & n6845 ) | ( n6844 & n6845 ) ;
  assign n6847 = ( n6568 & n6844 ) | ( n6568 & n6845 ) | ( n6844 & n6845 ) ;
  assign n6848 = ( n6568 & n6846 ) | ( n6568 & ~n6847 ) | ( n6846 & ~n6847 ) ;
  assign n6849 = ( x104 & n6843 ) | ( x104 & ~n6848 ) | ( n6843 & ~n6848 ) ;
  assign n6850 = ( x104 & n6569 ) | ( x104 & ~n6610 ) | ( n6569 & ~n6610 ) ;
  assign n6851 = x104 & n6569 ;
  assign n6852 = ( n6574 & n6850 ) | ( n6574 & n6851 ) | ( n6850 & n6851 ) ;
  assign n6853 = ( ~n6574 & n6850 ) | ( ~n6574 & n6851 ) | ( n6850 & n6851 ) ;
  assign n6854 = ( n6574 & ~n6852 ) | ( n6574 & n6853 ) | ( ~n6852 & n6853 ) ;
  assign n6855 = ( x105 & n6849 ) | ( x105 & ~n6854 ) | ( n6849 & ~n6854 ) ;
  assign n6856 = ( x105 & n6575 ) | ( x105 & ~n6610 ) | ( n6575 & ~n6610 ) ;
  assign n6857 = x105 & n6575 ;
  assign n6858 = ( ~n6580 & n6856 ) | ( ~n6580 & n6857 ) | ( n6856 & n6857 ) ;
  assign n6859 = ( n6580 & n6856 ) | ( n6580 & n6857 ) | ( n6856 & n6857 ) ;
  assign n6860 = ( n6580 & n6858 ) | ( n6580 & ~n6859 ) | ( n6858 & ~n6859 ) ;
  assign n6861 = ( x106 & n6855 ) | ( x106 & ~n6860 ) | ( n6855 & ~n6860 ) ;
  assign n6862 = ( x106 & n6581 ) | ( x106 & ~n6610 ) | ( n6581 & ~n6610 ) ;
  assign n6863 = x106 & n6581 ;
  assign n6864 = ( n6586 & n6862 ) | ( n6586 & n6863 ) | ( n6862 & n6863 ) ;
  assign n6865 = ( ~n6586 & n6862 ) | ( ~n6586 & n6863 ) | ( n6862 & n6863 ) ;
  assign n6866 = ( n6586 & ~n6864 ) | ( n6586 & n6865 ) | ( ~n6864 & n6865 ) ;
  assign n6867 = ( x107 & n6861 ) | ( x107 & ~n6866 ) | ( n6861 & ~n6866 ) ;
  assign n6868 = ( x107 & n6587 ) | ( x107 & ~n6610 ) | ( n6587 & ~n6610 ) ;
  assign n6869 = x107 & n6587 ;
  assign n6870 = ( ~n6592 & n6868 ) | ( ~n6592 & n6869 ) | ( n6868 & n6869 ) ;
  assign n6871 = ( n6592 & n6868 ) | ( n6592 & n6869 ) | ( n6868 & n6869 ) ;
  assign n6872 = ( n6592 & n6870 ) | ( n6592 & ~n6871 ) | ( n6870 & ~n6871 ) ;
  assign n6873 = ( x108 & n6867 ) | ( x108 & ~n6872 ) | ( n6867 & ~n6872 ) ;
  assign n6874 = ( x108 & n6593 ) | ( x108 & ~n6610 ) | ( n6593 & ~n6610 ) ;
  assign n6875 = x108 & n6593 ;
  assign n6876 = ( n6598 & n6874 ) | ( n6598 & n6875 ) | ( n6874 & n6875 ) ;
  assign n6877 = ( ~n6598 & n6874 ) | ( ~n6598 & n6875 ) | ( n6874 & n6875 ) ;
  assign n6878 = ( n6598 & ~n6876 ) | ( n6598 & n6877 ) | ( ~n6876 & n6877 ) ;
  assign n6879 = ( x109 & n6873 ) | ( x109 & ~n6878 ) | ( n6873 & ~n6878 ) ;
  assign n6880 = ( x109 & n6599 ) | ( x109 & ~n6610 ) | ( n6599 & ~n6610 ) ;
  assign n6881 = x109 & n6599 ;
  assign n6882 = ( n6604 & n6880 ) | ( n6604 & n6881 ) | ( n6880 & n6881 ) ;
  assign n6883 = ( ~n6604 & n6880 ) | ( ~n6604 & n6881 ) | ( n6880 & n6881 ) ;
  assign n6884 = ( n6604 & ~n6882 ) | ( n6604 & n6883 ) | ( ~n6882 & n6883 ) ;
  assign n6885 = ( x110 & n6879 ) | ( x110 & ~n6884 ) | ( n6879 & ~n6884 ) ;
  assign n6886 = x111 | n6885 ;
  assign n6887 = ( x111 & n146 ) | ( x111 & n6885 ) | ( n146 & n6885 ) ;
  assign n6888 = ( n6608 & ~n6886 ) | ( n6608 & n6887 ) | ( ~n6886 & n6887 ) ;
  assign n6889 = ( x111 & ~n6608 ) | ( x111 & n6885 ) | ( ~n6608 & n6885 ) ;
  assign n6890 = n146 | n6889 ;
  assign n6891 = ( x16 & ~x64 ) | ( x16 & n6890 ) | ( ~x64 & n6890 ) ;
  assign n6892 = ~x16 & n6890 ;
  assign n6893 = ( n6614 & n6891 ) | ( n6614 & ~n6892 ) | ( n6891 & ~n6892 ) ;
  assign n6894 = ~x15 & x64 ;
  assign n6895 = ( x65 & ~n6893 ) | ( x65 & n6894 ) | ( ~n6893 & n6894 ) ;
  assign n6896 = ( x65 & n6614 ) | ( x65 & ~n6890 ) | ( n6614 & ~n6890 ) ;
  assign n6897 = x65 & n6614 ;
  assign n6898 = ( n6613 & n6896 ) | ( n6613 & n6897 ) | ( n6896 & n6897 ) ;
  assign n6899 = ( ~n6613 & n6896 ) | ( ~n6613 & n6897 ) | ( n6896 & n6897 ) ;
  assign n6900 = ( n6613 & ~n6898 ) | ( n6613 & n6899 ) | ( ~n6898 & n6899 ) ;
  assign n6901 = ( x66 & n6895 ) | ( x66 & ~n6900 ) | ( n6895 & ~n6900 ) ;
  assign n6902 = ( x66 & n6615 ) | ( x66 & ~n6890 ) | ( n6615 & ~n6890 ) ;
  assign n6903 = x66 & n6615 ;
  assign n6904 = ( n6620 & n6902 ) | ( n6620 & n6903 ) | ( n6902 & n6903 ) ;
  assign n6905 = ( ~n6620 & n6902 ) | ( ~n6620 & n6903 ) | ( n6902 & n6903 ) ;
  assign n6906 = ( n6620 & ~n6904 ) | ( n6620 & n6905 ) | ( ~n6904 & n6905 ) ;
  assign n6907 = ( x67 & n6901 ) | ( x67 & ~n6906 ) | ( n6901 & ~n6906 ) ;
  assign n6908 = ( x67 & n6621 ) | ( x67 & ~n6890 ) | ( n6621 & ~n6890 ) ;
  assign n6909 = x67 & n6621 ;
  assign n6910 = ( ~n6626 & n6908 ) | ( ~n6626 & n6909 ) | ( n6908 & n6909 ) ;
  assign n6911 = ( n6626 & n6908 ) | ( n6626 & n6909 ) | ( n6908 & n6909 ) ;
  assign n6912 = ( n6626 & n6910 ) | ( n6626 & ~n6911 ) | ( n6910 & ~n6911 ) ;
  assign n6913 = ( x68 & n6907 ) | ( x68 & ~n6912 ) | ( n6907 & ~n6912 ) ;
  assign n6914 = ( x68 & n6627 ) | ( x68 & ~n6890 ) | ( n6627 & ~n6890 ) ;
  assign n6915 = x68 & n6627 ;
  assign n6916 = ( n6632 & n6914 ) | ( n6632 & n6915 ) | ( n6914 & n6915 ) ;
  assign n6917 = ( ~n6632 & n6914 ) | ( ~n6632 & n6915 ) | ( n6914 & n6915 ) ;
  assign n6918 = ( n6632 & ~n6916 ) | ( n6632 & n6917 ) | ( ~n6916 & n6917 ) ;
  assign n6919 = ( x69 & n6913 ) | ( x69 & ~n6918 ) | ( n6913 & ~n6918 ) ;
  assign n6920 = ( x69 & n6633 ) | ( x69 & ~n6890 ) | ( n6633 & ~n6890 ) ;
  assign n6921 = x69 & n6633 ;
  assign n6922 = ( ~n6638 & n6920 ) | ( ~n6638 & n6921 ) | ( n6920 & n6921 ) ;
  assign n6923 = ( n6638 & n6920 ) | ( n6638 & n6921 ) | ( n6920 & n6921 ) ;
  assign n6924 = ( n6638 & n6922 ) | ( n6638 & ~n6923 ) | ( n6922 & ~n6923 ) ;
  assign n6925 = ( x70 & n6919 ) | ( x70 & ~n6924 ) | ( n6919 & ~n6924 ) ;
  assign n6926 = ( x70 & n6639 ) | ( x70 & ~n6890 ) | ( n6639 & ~n6890 ) ;
  assign n6927 = x70 & n6639 ;
  assign n6928 = ( n6644 & n6926 ) | ( n6644 & n6927 ) | ( n6926 & n6927 ) ;
  assign n6929 = ( ~n6644 & n6926 ) | ( ~n6644 & n6927 ) | ( n6926 & n6927 ) ;
  assign n6930 = ( n6644 & ~n6928 ) | ( n6644 & n6929 ) | ( ~n6928 & n6929 ) ;
  assign n6931 = ( x71 & n6925 ) | ( x71 & ~n6930 ) | ( n6925 & ~n6930 ) ;
  assign n6932 = ( x71 & n6645 ) | ( x71 & ~n6890 ) | ( n6645 & ~n6890 ) ;
  assign n6933 = x71 & n6645 ;
  assign n6934 = ( ~n6650 & n6932 ) | ( ~n6650 & n6933 ) | ( n6932 & n6933 ) ;
  assign n6935 = ( n6650 & n6932 ) | ( n6650 & n6933 ) | ( n6932 & n6933 ) ;
  assign n6936 = ( n6650 & n6934 ) | ( n6650 & ~n6935 ) | ( n6934 & ~n6935 ) ;
  assign n6937 = ( x72 & n6931 ) | ( x72 & ~n6936 ) | ( n6931 & ~n6936 ) ;
  assign n6938 = ( x72 & n6651 ) | ( x72 & ~n6890 ) | ( n6651 & ~n6890 ) ;
  assign n6939 = x72 & n6651 ;
  assign n6940 = ( n6656 & n6938 ) | ( n6656 & n6939 ) | ( n6938 & n6939 ) ;
  assign n6941 = ( ~n6656 & n6938 ) | ( ~n6656 & n6939 ) | ( n6938 & n6939 ) ;
  assign n6942 = ( n6656 & ~n6940 ) | ( n6656 & n6941 ) | ( ~n6940 & n6941 ) ;
  assign n6943 = ( x73 & n6937 ) | ( x73 & ~n6942 ) | ( n6937 & ~n6942 ) ;
  assign n6944 = ( x73 & n6657 ) | ( x73 & ~n6890 ) | ( n6657 & ~n6890 ) ;
  assign n6945 = x73 & n6657 ;
  assign n6946 = ( ~n6662 & n6944 ) | ( ~n6662 & n6945 ) | ( n6944 & n6945 ) ;
  assign n6947 = ( n6662 & n6944 ) | ( n6662 & n6945 ) | ( n6944 & n6945 ) ;
  assign n6948 = ( n6662 & n6946 ) | ( n6662 & ~n6947 ) | ( n6946 & ~n6947 ) ;
  assign n6949 = ( x74 & n6943 ) | ( x74 & ~n6948 ) | ( n6943 & ~n6948 ) ;
  assign n6950 = ( x74 & n6663 ) | ( x74 & ~n6890 ) | ( n6663 & ~n6890 ) ;
  assign n6951 = x74 & n6663 ;
  assign n6952 = ( n6668 & n6950 ) | ( n6668 & n6951 ) | ( n6950 & n6951 ) ;
  assign n6953 = ( ~n6668 & n6950 ) | ( ~n6668 & n6951 ) | ( n6950 & n6951 ) ;
  assign n6954 = ( n6668 & ~n6952 ) | ( n6668 & n6953 ) | ( ~n6952 & n6953 ) ;
  assign n6955 = ( x75 & n6949 ) | ( x75 & ~n6954 ) | ( n6949 & ~n6954 ) ;
  assign n6956 = ( x75 & n6669 ) | ( x75 & ~n6890 ) | ( n6669 & ~n6890 ) ;
  assign n6957 = x75 & n6669 ;
  assign n6958 = ( ~n6674 & n6956 ) | ( ~n6674 & n6957 ) | ( n6956 & n6957 ) ;
  assign n6959 = ( n6674 & n6956 ) | ( n6674 & n6957 ) | ( n6956 & n6957 ) ;
  assign n6960 = ( n6674 & n6958 ) | ( n6674 & ~n6959 ) | ( n6958 & ~n6959 ) ;
  assign n6961 = ( x76 & n6955 ) | ( x76 & ~n6960 ) | ( n6955 & ~n6960 ) ;
  assign n6962 = ( x76 & n6675 ) | ( x76 & ~n6890 ) | ( n6675 & ~n6890 ) ;
  assign n6963 = x76 & n6675 ;
  assign n6964 = ( n6680 & n6962 ) | ( n6680 & n6963 ) | ( n6962 & n6963 ) ;
  assign n6965 = ( ~n6680 & n6962 ) | ( ~n6680 & n6963 ) | ( n6962 & n6963 ) ;
  assign n6966 = ( n6680 & ~n6964 ) | ( n6680 & n6965 ) | ( ~n6964 & n6965 ) ;
  assign n6967 = ( x77 & n6961 ) | ( x77 & ~n6966 ) | ( n6961 & ~n6966 ) ;
  assign n6968 = ( x77 & n6681 ) | ( x77 & ~n6890 ) | ( n6681 & ~n6890 ) ;
  assign n6969 = x77 & n6681 ;
  assign n6970 = ( ~n6686 & n6968 ) | ( ~n6686 & n6969 ) | ( n6968 & n6969 ) ;
  assign n6971 = ( n6686 & n6968 ) | ( n6686 & n6969 ) | ( n6968 & n6969 ) ;
  assign n6972 = ( n6686 & n6970 ) | ( n6686 & ~n6971 ) | ( n6970 & ~n6971 ) ;
  assign n6973 = ( x78 & n6967 ) | ( x78 & ~n6972 ) | ( n6967 & ~n6972 ) ;
  assign n6974 = ( x78 & n6687 ) | ( x78 & ~n6890 ) | ( n6687 & ~n6890 ) ;
  assign n6975 = x78 & n6687 ;
  assign n6976 = ( n6692 & n6974 ) | ( n6692 & n6975 ) | ( n6974 & n6975 ) ;
  assign n6977 = ( ~n6692 & n6974 ) | ( ~n6692 & n6975 ) | ( n6974 & n6975 ) ;
  assign n6978 = ( n6692 & ~n6976 ) | ( n6692 & n6977 ) | ( ~n6976 & n6977 ) ;
  assign n6979 = ( x79 & n6973 ) | ( x79 & ~n6978 ) | ( n6973 & ~n6978 ) ;
  assign n6980 = ( x79 & n6693 ) | ( x79 & ~n6890 ) | ( n6693 & ~n6890 ) ;
  assign n6981 = x79 & n6693 ;
  assign n6982 = ( ~n6698 & n6980 ) | ( ~n6698 & n6981 ) | ( n6980 & n6981 ) ;
  assign n6983 = ( n6698 & n6980 ) | ( n6698 & n6981 ) | ( n6980 & n6981 ) ;
  assign n6984 = ( n6698 & n6982 ) | ( n6698 & ~n6983 ) | ( n6982 & ~n6983 ) ;
  assign n6985 = ( x80 & n6979 ) | ( x80 & ~n6984 ) | ( n6979 & ~n6984 ) ;
  assign n6986 = ( x80 & n6699 ) | ( x80 & ~n6890 ) | ( n6699 & ~n6890 ) ;
  assign n6987 = x80 & n6699 ;
  assign n6988 = ( n6704 & n6986 ) | ( n6704 & n6987 ) | ( n6986 & n6987 ) ;
  assign n6989 = ( ~n6704 & n6986 ) | ( ~n6704 & n6987 ) | ( n6986 & n6987 ) ;
  assign n6990 = ( n6704 & ~n6988 ) | ( n6704 & n6989 ) | ( ~n6988 & n6989 ) ;
  assign n6991 = ( x81 & n6985 ) | ( x81 & ~n6990 ) | ( n6985 & ~n6990 ) ;
  assign n6992 = ( x81 & n6705 ) | ( x81 & ~n6890 ) | ( n6705 & ~n6890 ) ;
  assign n6993 = x81 & n6705 ;
  assign n6994 = ( ~n6710 & n6992 ) | ( ~n6710 & n6993 ) | ( n6992 & n6993 ) ;
  assign n6995 = ( n6710 & n6992 ) | ( n6710 & n6993 ) | ( n6992 & n6993 ) ;
  assign n6996 = ( n6710 & n6994 ) | ( n6710 & ~n6995 ) | ( n6994 & ~n6995 ) ;
  assign n6997 = ( x82 & n6991 ) | ( x82 & ~n6996 ) | ( n6991 & ~n6996 ) ;
  assign n6998 = ( x82 & n6711 ) | ( x82 & ~n6890 ) | ( n6711 & ~n6890 ) ;
  assign n6999 = x82 & n6711 ;
  assign n7000 = ( n6716 & n6998 ) | ( n6716 & n6999 ) | ( n6998 & n6999 ) ;
  assign n7001 = ( ~n6716 & n6998 ) | ( ~n6716 & n6999 ) | ( n6998 & n6999 ) ;
  assign n7002 = ( n6716 & ~n7000 ) | ( n6716 & n7001 ) | ( ~n7000 & n7001 ) ;
  assign n7003 = ( x83 & n6997 ) | ( x83 & ~n7002 ) | ( n6997 & ~n7002 ) ;
  assign n7004 = ( x83 & n6717 ) | ( x83 & ~n6890 ) | ( n6717 & ~n6890 ) ;
  assign n7005 = x83 & n6717 ;
  assign n7006 = ( ~n6722 & n7004 ) | ( ~n6722 & n7005 ) | ( n7004 & n7005 ) ;
  assign n7007 = ( n6722 & n7004 ) | ( n6722 & n7005 ) | ( n7004 & n7005 ) ;
  assign n7008 = ( n6722 & n7006 ) | ( n6722 & ~n7007 ) | ( n7006 & ~n7007 ) ;
  assign n7009 = ( x84 & n7003 ) | ( x84 & ~n7008 ) | ( n7003 & ~n7008 ) ;
  assign n7010 = ( x84 & n6723 ) | ( x84 & ~n6890 ) | ( n6723 & ~n6890 ) ;
  assign n7011 = x84 & n6723 ;
  assign n7012 = ( n6728 & n7010 ) | ( n6728 & n7011 ) | ( n7010 & n7011 ) ;
  assign n7013 = ( ~n6728 & n7010 ) | ( ~n6728 & n7011 ) | ( n7010 & n7011 ) ;
  assign n7014 = ( n6728 & ~n7012 ) | ( n6728 & n7013 ) | ( ~n7012 & n7013 ) ;
  assign n7015 = ( x85 & n7009 ) | ( x85 & ~n7014 ) | ( n7009 & ~n7014 ) ;
  assign n7016 = ( x85 & n6729 ) | ( x85 & ~n6890 ) | ( n6729 & ~n6890 ) ;
  assign n7017 = x85 & n6729 ;
  assign n7018 = ( ~n6734 & n7016 ) | ( ~n6734 & n7017 ) | ( n7016 & n7017 ) ;
  assign n7019 = ( n6734 & n7016 ) | ( n6734 & n7017 ) | ( n7016 & n7017 ) ;
  assign n7020 = ( n6734 & n7018 ) | ( n6734 & ~n7019 ) | ( n7018 & ~n7019 ) ;
  assign n7021 = ( x86 & n7015 ) | ( x86 & ~n7020 ) | ( n7015 & ~n7020 ) ;
  assign n7022 = ( x86 & n6735 ) | ( x86 & ~n6890 ) | ( n6735 & ~n6890 ) ;
  assign n7023 = x86 & n6735 ;
  assign n7024 = ( n6740 & n7022 ) | ( n6740 & n7023 ) | ( n7022 & n7023 ) ;
  assign n7025 = ( ~n6740 & n7022 ) | ( ~n6740 & n7023 ) | ( n7022 & n7023 ) ;
  assign n7026 = ( n6740 & ~n7024 ) | ( n6740 & n7025 ) | ( ~n7024 & n7025 ) ;
  assign n7027 = ( x87 & n7021 ) | ( x87 & ~n7026 ) | ( n7021 & ~n7026 ) ;
  assign n7028 = ( x87 & n6741 ) | ( x87 & ~n6890 ) | ( n6741 & ~n6890 ) ;
  assign n7029 = x87 & n6741 ;
  assign n7030 = ( ~n6746 & n7028 ) | ( ~n6746 & n7029 ) | ( n7028 & n7029 ) ;
  assign n7031 = ( n6746 & n7028 ) | ( n6746 & n7029 ) | ( n7028 & n7029 ) ;
  assign n7032 = ( n6746 & n7030 ) | ( n6746 & ~n7031 ) | ( n7030 & ~n7031 ) ;
  assign n7033 = ( x88 & n7027 ) | ( x88 & ~n7032 ) | ( n7027 & ~n7032 ) ;
  assign n7034 = ( x88 & n6747 ) | ( x88 & ~n6890 ) | ( n6747 & ~n6890 ) ;
  assign n7035 = x88 & n6747 ;
  assign n7036 = ( n6752 & n7034 ) | ( n6752 & n7035 ) | ( n7034 & n7035 ) ;
  assign n7037 = ( ~n6752 & n7034 ) | ( ~n6752 & n7035 ) | ( n7034 & n7035 ) ;
  assign n7038 = ( n6752 & ~n7036 ) | ( n6752 & n7037 ) | ( ~n7036 & n7037 ) ;
  assign n7039 = ( x89 & n7033 ) | ( x89 & ~n7038 ) | ( n7033 & ~n7038 ) ;
  assign n7040 = ( x89 & n6753 ) | ( x89 & ~n6890 ) | ( n6753 & ~n6890 ) ;
  assign n7041 = x89 & n6753 ;
  assign n7042 = ( ~n6758 & n7040 ) | ( ~n6758 & n7041 ) | ( n7040 & n7041 ) ;
  assign n7043 = ( n6758 & n7040 ) | ( n6758 & n7041 ) | ( n7040 & n7041 ) ;
  assign n7044 = ( n6758 & n7042 ) | ( n6758 & ~n7043 ) | ( n7042 & ~n7043 ) ;
  assign n7045 = ( x90 & n7039 ) | ( x90 & ~n7044 ) | ( n7039 & ~n7044 ) ;
  assign n7046 = ( x90 & n6759 ) | ( x90 & ~n6890 ) | ( n6759 & ~n6890 ) ;
  assign n7047 = x90 & n6759 ;
  assign n7048 = ( n6764 & n7046 ) | ( n6764 & n7047 ) | ( n7046 & n7047 ) ;
  assign n7049 = ( ~n6764 & n7046 ) | ( ~n6764 & n7047 ) | ( n7046 & n7047 ) ;
  assign n7050 = ( n6764 & ~n7048 ) | ( n6764 & n7049 ) | ( ~n7048 & n7049 ) ;
  assign n7051 = ( x91 & n7045 ) | ( x91 & ~n7050 ) | ( n7045 & ~n7050 ) ;
  assign n7052 = ( x91 & n6765 ) | ( x91 & ~n6890 ) | ( n6765 & ~n6890 ) ;
  assign n7053 = x91 & n6765 ;
  assign n7054 = ( ~n6770 & n7052 ) | ( ~n6770 & n7053 ) | ( n7052 & n7053 ) ;
  assign n7055 = ( n6770 & n7052 ) | ( n6770 & n7053 ) | ( n7052 & n7053 ) ;
  assign n7056 = ( n6770 & n7054 ) | ( n6770 & ~n7055 ) | ( n7054 & ~n7055 ) ;
  assign n7057 = ( x92 & n7051 ) | ( x92 & ~n7056 ) | ( n7051 & ~n7056 ) ;
  assign n7058 = ( x92 & n6771 ) | ( x92 & ~n6890 ) | ( n6771 & ~n6890 ) ;
  assign n7059 = x92 & n6771 ;
  assign n7060 = ( n6776 & n7058 ) | ( n6776 & n7059 ) | ( n7058 & n7059 ) ;
  assign n7061 = ( ~n6776 & n7058 ) | ( ~n6776 & n7059 ) | ( n7058 & n7059 ) ;
  assign n7062 = ( n6776 & ~n7060 ) | ( n6776 & n7061 ) | ( ~n7060 & n7061 ) ;
  assign n7063 = ( x93 & n7057 ) | ( x93 & ~n7062 ) | ( n7057 & ~n7062 ) ;
  assign n7064 = ( x93 & n6777 ) | ( x93 & ~n6890 ) | ( n6777 & ~n6890 ) ;
  assign n7065 = x93 & n6777 ;
  assign n7066 = ( ~n6782 & n7064 ) | ( ~n6782 & n7065 ) | ( n7064 & n7065 ) ;
  assign n7067 = ( n6782 & n7064 ) | ( n6782 & n7065 ) | ( n7064 & n7065 ) ;
  assign n7068 = ( n6782 & n7066 ) | ( n6782 & ~n7067 ) | ( n7066 & ~n7067 ) ;
  assign n7069 = ( x94 & n7063 ) | ( x94 & ~n7068 ) | ( n7063 & ~n7068 ) ;
  assign n7070 = ( x94 & n6783 ) | ( x94 & ~n6890 ) | ( n6783 & ~n6890 ) ;
  assign n7071 = x94 & n6783 ;
  assign n7072 = ( n6788 & n7070 ) | ( n6788 & n7071 ) | ( n7070 & n7071 ) ;
  assign n7073 = ( ~n6788 & n7070 ) | ( ~n6788 & n7071 ) | ( n7070 & n7071 ) ;
  assign n7074 = ( n6788 & ~n7072 ) | ( n6788 & n7073 ) | ( ~n7072 & n7073 ) ;
  assign n7075 = ( x95 & n7069 ) | ( x95 & ~n7074 ) | ( n7069 & ~n7074 ) ;
  assign n7076 = ( x95 & n6789 ) | ( x95 & ~n6890 ) | ( n6789 & ~n6890 ) ;
  assign n7077 = x95 & n6789 ;
  assign n7078 = ( ~n6794 & n7076 ) | ( ~n6794 & n7077 ) | ( n7076 & n7077 ) ;
  assign n7079 = ( n6794 & n7076 ) | ( n6794 & n7077 ) | ( n7076 & n7077 ) ;
  assign n7080 = ( n6794 & n7078 ) | ( n6794 & ~n7079 ) | ( n7078 & ~n7079 ) ;
  assign n7081 = ( x96 & n7075 ) | ( x96 & ~n7080 ) | ( n7075 & ~n7080 ) ;
  assign n7082 = ( x96 & n6795 ) | ( x96 & ~n6890 ) | ( n6795 & ~n6890 ) ;
  assign n7083 = x96 & n6795 ;
  assign n7084 = ( n6800 & n7082 ) | ( n6800 & n7083 ) | ( n7082 & n7083 ) ;
  assign n7085 = ( ~n6800 & n7082 ) | ( ~n6800 & n7083 ) | ( n7082 & n7083 ) ;
  assign n7086 = ( n6800 & ~n7084 ) | ( n6800 & n7085 ) | ( ~n7084 & n7085 ) ;
  assign n7087 = ( x97 & n7081 ) | ( x97 & ~n7086 ) | ( n7081 & ~n7086 ) ;
  assign n7088 = ( x97 & n6801 ) | ( x97 & ~n6890 ) | ( n6801 & ~n6890 ) ;
  assign n7089 = x97 & n6801 ;
  assign n7090 = ( ~n6806 & n7088 ) | ( ~n6806 & n7089 ) | ( n7088 & n7089 ) ;
  assign n7091 = ( n6806 & n7088 ) | ( n6806 & n7089 ) | ( n7088 & n7089 ) ;
  assign n7092 = ( n6806 & n7090 ) | ( n6806 & ~n7091 ) | ( n7090 & ~n7091 ) ;
  assign n7093 = ( x98 & n7087 ) | ( x98 & ~n7092 ) | ( n7087 & ~n7092 ) ;
  assign n7094 = ( x98 & n6807 ) | ( x98 & ~n6890 ) | ( n6807 & ~n6890 ) ;
  assign n7095 = x98 & n6807 ;
  assign n7096 = ( n6812 & n7094 ) | ( n6812 & n7095 ) | ( n7094 & n7095 ) ;
  assign n7097 = ( ~n6812 & n7094 ) | ( ~n6812 & n7095 ) | ( n7094 & n7095 ) ;
  assign n7098 = ( n6812 & ~n7096 ) | ( n6812 & n7097 ) | ( ~n7096 & n7097 ) ;
  assign n7099 = ( x99 & n7093 ) | ( x99 & ~n7098 ) | ( n7093 & ~n7098 ) ;
  assign n7100 = ( x99 & n6813 ) | ( x99 & ~n6890 ) | ( n6813 & ~n6890 ) ;
  assign n7101 = x99 & n6813 ;
  assign n7102 = ( ~n6818 & n7100 ) | ( ~n6818 & n7101 ) | ( n7100 & n7101 ) ;
  assign n7103 = ( n6818 & n7100 ) | ( n6818 & n7101 ) | ( n7100 & n7101 ) ;
  assign n7104 = ( n6818 & n7102 ) | ( n6818 & ~n7103 ) | ( n7102 & ~n7103 ) ;
  assign n7105 = ( x100 & n7099 ) | ( x100 & ~n7104 ) | ( n7099 & ~n7104 ) ;
  assign n7106 = ( x100 & n6819 ) | ( x100 & ~n6890 ) | ( n6819 & ~n6890 ) ;
  assign n7107 = x100 & n6819 ;
  assign n7108 = ( n6824 & n7106 ) | ( n6824 & n7107 ) | ( n7106 & n7107 ) ;
  assign n7109 = ( ~n6824 & n7106 ) | ( ~n6824 & n7107 ) | ( n7106 & n7107 ) ;
  assign n7110 = ( n6824 & ~n7108 ) | ( n6824 & n7109 ) | ( ~n7108 & n7109 ) ;
  assign n7111 = ( x101 & n7105 ) | ( x101 & ~n7110 ) | ( n7105 & ~n7110 ) ;
  assign n7112 = ( x101 & n6825 ) | ( x101 & ~n6890 ) | ( n6825 & ~n6890 ) ;
  assign n7113 = x101 & n6825 ;
  assign n7114 = ( ~n6830 & n7112 ) | ( ~n6830 & n7113 ) | ( n7112 & n7113 ) ;
  assign n7115 = ( n6830 & n7112 ) | ( n6830 & n7113 ) | ( n7112 & n7113 ) ;
  assign n7116 = ( n6830 & n7114 ) | ( n6830 & ~n7115 ) | ( n7114 & ~n7115 ) ;
  assign n7117 = ( x102 & n7111 ) | ( x102 & ~n7116 ) | ( n7111 & ~n7116 ) ;
  assign n7118 = ( x102 & n6831 ) | ( x102 & ~n6890 ) | ( n6831 & ~n6890 ) ;
  assign n7119 = x102 & n6831 ;
  assign n7120 = ( n6836 & n7118 ) | ( n6836 & n7119 ) | ( n7118 & n7119 ) ;
  assign n7121 = ( ~n6836 & n7118 ) | ( ~n6836 & n7119 ) | ( n7118 & n7119 ) ;
  assign n7122 = ( n6836 & ~n7120 ) | ( n6836 & n7121 ) | ( ~n7120 & n7121 ) ;
  assign n7123 = ( x103 & n7117 ) | ( x103 & ~n7122 ) | ( n7117 & ~n7122 ) ;
  assign n7124 = ( x103 & n6837 ) | ( x103 & ~n6890 ) | ( n6837 & ~n6890 ) ;
  assign n7125 = x103 & n6837 ;
  assign n7126 = ( ~n6842 & n7124 ) | ( ~n6842 & n7125 ) | ( n7124 & n7125 ) ;
  assign n7127 = ( n6842 & n7124 ) | ( n6842 & n7125 ) | ( n7124 & n7125 ) ;
  assign n7128 = ( n6842 & n7126 ) | ( n6842 & ~n7127 ) | ( n7126 & ~n7127 ) ;
  assign n7129 = ( x104 & n7123 ) | ( x104 & ~n7128 ) | ( n7123 & ~n7128 ) ;
  assign n7130 = ( x104 & n6843 ) | ( x104 & ~n6890 ) | ( n6843 & ~n6890 ) ;
  assign n7131 = x104 & n6843 ;
  assign n7132 = ( n6848 & n7130 ) | ( n6848 & n7131 ) | ( n7130 & n7131 ) ;
  assign n7133 = ( ~n6848 & n7130 ) | ( ~n6848 & n7131 ) | ( n7130 & n7131 ) ;
  assign n7134 = ( n6848 & ~n7132 ) | ( n6848 & n7133 ) | ( ~n7132 & n7133 ) ;
  assign n7135 = ( x105 & n7129 ) | ( x105 & ~n7134 ) | ( n7129 & ~n7134 ) ;
  assign n7136 = ( x105 & n6849 ) | ( x105 & ~n6890 ) | ( n6849 & ~n6890 ) ;
  assign n7137 = x105 & n6849 ;
  assign n7138 = ( ~n6854 & n7136 ) | ( ~n6854 & n7137 ) | ( n7136 & n7137 ) ;
  assign n7139 = ( n6854 & n7136 ) | ( n6854 & n7137 ) | ( n7136 & n7137 ) ;
  assign n7140 = ( n6854 & n7138 ) | ( n6854 & ~n7139 ) | ( n7138 & ~n7139 ) ;
  assign n7141 = ( x106 & n7135 ) | ( x106 & ~n7140 ) | ( n7135 & ~n7140 ) ;
  assign n7142 = ( x106 & n6855 ) | ( x106 & ~n6890 ) | ( n6855 & ~n6890 ) ;
  assign n7143 = x106 & n6855 ;
  assign n7144 = ( n6860 & n7142 ) | ( n6860 & n7143 ) | ( n7142 & n7143 ) ;
  assign n7145 = ( ~n6860 & n7142 ) | ( ~n6860 & n7143 ) | ( n7142 & n7143 ) ;
  assign n7146 = ( n6860 & ~n7144 ) | ( n6860 & n7145 ) | ( ~n7144 & n7145 ) ;
  assign n7147 = ( x107 & n7141 ) | ( x107 & ~n7146 ) | ( n7141 & ~n7146 ) ;
  assign n7148 = ( x107 & n6861 ) | ( x107 & ~n6890 ) | ( n6861 & ~n6890 ) ;
  assign n7149 = x107 & n6861 ;
  assign n7150 = ( ~n6866 & n7148 ) | ( ~n6866 & n7149 ) | ( n7148 & n7149 ) ;
  assign n7151 = ( n6866 & n7148 ) | ( n6866 & n7149 ) | ( n7148 & n7149 ) ;
  assign n7152 = ( n6866 & n7150 ) | ( n6866 & ~n7151 ) | ( n7150 & ~n7151 ) ;
  assign n7153 = ( x108 & n7147 ) | ( x108 & ~n7152 ) | ( n7147 & ~n7152 ) ;
  assign n7154 = ( x108 & n6867 ) | ( x108 & ~n6890 ) | ( n6867 & ~n6890 ) ;
  assign n7155 = x108 & n6867 ;
  assign n7156 = ( n6872 & n7154 ) | ( n6872 & n7155 ) | ( n7154 & n7155 ) ;
  assign n7157 = ( ~n6872 & n7154 ) | ( ~n6872 & n7155 ) | ( n7154 & n7155 ) ;
  assign n7158 = ( n6872 & ~n7156 ) | ( n6872 & n7157 ) | ( ~n7156 & n7157 ) ;
  assign n7159 = ( x109 & n7153 ) | ( x109 & ~n7158 ) | ( n7153 & ~n7158 ) ;
  assign n7160 = ( x109 & n6873 ) | ( x109 & ~n6890 ) | ( n6873 & ~n6890 ) ;
  assign n7161 = x109 & n6873 ;
  assign n7162 = ( ~n6878 & n7160 ) | ( ~n6878 & n7161 ) | ( n7160 & n7161 ) ;
  assign n7163 = ( n6878 & n7160 ) | ( n6878 & n7161 ) | ( n7160 & n7161 ) ;
  assign n7164 = ( n6878 & n7162 ) | ( n6878 & ~n7163 ) | ( n7162 & ~n7163 ) ;
  assign n7165 = ( x110 & n7159 ) | ( x110 & ~n7164 ) | ( n7159 & ~n7164 ) ;
  assign n7166 = ( x110 & n6879 ) | ( x110 & ~n6890 ) | ( n6879 & ~n6890 ) ;
  assign n7167 = x110 & n6879 ;
  assign n7168 = ( ~n6884 & n7166 ) | ( ~n6884 & n7167 ) | ( n7166 & n7167 ) ;
  assign n7169 = ( n6884 & n7166 ) | ( n6884 & n7167 ) | ( n7166 & n7167 ) ;
  assign n7170 = ( n6884 & n7168 ) | ( n6884 & ~n7169 ) | ( n7168 & ~n7169 ) ;
  assign n7171 = ( x111 & n7165 ) | ( x111 & ~n7170 ) | ( n7165 & ~n7170 ) ;
  assign n7172 = ( x112 & ~n6888 ) | ( x112 & n7171 ) | ( ~n6888 & n7171 ) ;
  assign n7173 = n145 | n7172 ;
  assign n7174 = n6888 & n7173 ;
  assign n7175 = n280 | n7174 ;
  assign n7176 = ( x15 & ~x64 ) | ( x15 & n7173 ) | ( ~x64 & n7173 ) ;
  assign n7177 = ~x15 & n7173 ;
  assign n7178 = ( n6894 & n7176 ) | ( n6894 & ~n7177 ) | ( n7176 & ~n7177 ) ;
  assign n7179 = ~x14 & x64 ;
  assign n7180 = ( x65 & ~n7178 ) | ( x65 & n7179 ) | ( ~n7178 & n7179 ) ;
  assign n7181 = ( x65 & n6894 ) | ( x65 & ~n7173 ) | ( n6894 & ~n7173 ) ;
  assign n7182 = x65 & n6894 ;
  assign n7183 = ( n6893 & n7181 ) | ( n6893 & n7182 ) | ( n7181 & n7182 ) ;
  assign n7184 = ( ~n6893 & n7181 ) | ( ~n6893 & n7182 ) | ( n7181 & n7182 ) ;
  assign n7185 = ( n6893 & ~n7183 ) | ( n6893 & n7184 ) | ( ~n7183 & n7184 ) ;
  assign n7186 = ( x66 & n7180 ) | ( x66 & ~n7185 ) | ( n7180 & ~n7185 ) ;
  assign n7187 = ( x66 & n6895 ) | ( x66 & ~n7173 ) | ( n6895 & ~n7173 ) ;
  assign n7188 = x66 & n6895 ;
  assign n7189 = ( n6900 & n7187 ) | ( n6900 & n7188 ) | ( n7187 & n7188 ) ;
  assign n7190 = ( ~n6900 & n7187 ) | ( ~n6900 & n7188 ) | ( n7187 & n7188 ) ;
  assign n7191 = ( n6900 & ~n7189 ) | ( n6900 & n7190 ) | ( ~n7189 & n7190 ) ;
  assign n7192 = ( x67 & n7186 ) | ( x67 & ~n7191 ) | ( n7186 & ~n7191 ) ;
  assign n7193 = ( x67 & n6901 ) | ( x67 & ~n7173 ) | ( n6901 & ~n7173 ) ;
  assign n7194 = x67 & n6901 ;
  assign n7195 = ( ~n6906 & n7193 ) | ( ~n6906 & n7194 ) | ( n7193 & n7194 ) ;
  assign n7196 = ( n6906 & n7193 ) | ( n6906 & n7194 ) | ( n7193 & n7194 ) ;
  assign n7197 = ( n6906 & n7195 ) | ( n6906 & ~n7196 ) | ( n7195 & ~n7196 ) ;
  assign n7198 = ( x68 & n7192 ) | ( x68 & ~n7197 ) | ( n7192 & ~n7197 ) ;
  assign n7199 = ( x68 & n6907 ) | ( x68 & ~n7173 ) | ( n6907 & ~n7173 ) ;
  assign n7200 = x68 & n6907 ;
  assign n7201 = ( n6912 & n7199 ) | ( n6912 & n7200 ) | ( n7199 & n7200 ) ;
  assign n7202 = ( ~n6912 & n7199 ) | ( ~n6912 & n7200 ) | ( n7199 & n7200 ) ;
  assign n7203 = ( n6912 & ~n7201 ) | ( n6912 & n7202 ) | ( ~n7201 & n7202 ) ;
  assign n7204 = ( x69 & n7198 ) | ( x69 & ~n7203 ) | ( n7198 & ~n7203 ) ;
  assign n7205 = ( x69 & n6913 ) | ( x69 & ~n7173 ) | ( n6913 & ~n7173 ) ;
  assign n7206 = x69 & n6913 ;
  assign n7207 = ( ~n6918 & n7205 ) | ( ~n6918 & n7206 ) | ( n7205 & n7206 ) ;
  assign n7208 = ( n6918 & n7205 ) | ( n6918 & n7206 ) | ( n7205 & n7206 ) ;
  assign n7209 = ( n6918 & n7207 ) | ( n6918 & ~n7208 ) | ( n7207 & ~n7208 ) ;
  assign n7210 = ( x70 & n7204 ) | ( x70 & ~n7209 ) | ( n7204 & ~n7209 ) ;
  assign n7211 = ( x70 & n6919 ) | ( x70 & ~n7173 ) | ( n6919 & ~n7173 ) ;
  assign n7212 = x70 & n6919 ;
  assign n7213 = ( n6924 & n7211 ) | ( n6924 & n7212 ) | ( n7211 & n7212 ) ;
  assign n7214 = ( ~n6924 & n7211 ) | ( ~n6924 & n7212 ) | ( n7211 & n7212 ) ;
  assign n7215 = ( n6924 & ~n7213 ) | ( n6924 & n7214 ) | ( ~n7213 & n7214 ) ;
  assign n7216 = ( x71 & n7210 ) | ( x71 & ~n7215 ) | ( n7210 & ~n7215 ) ;
  assign n7217 = ( x71 & n6925 ) | ( x71 & ~n7173 ) | ( n6925 & ~n7173 ) ;
  assign n7218 = x71 & n6925 ;
  assign n7219 = ( ~n6930 & n7217 ) | ( ~n6930 & n7218 ) | ( n7217 & n7218 ) ;
  assign n7220 = ( n6930 & n7217 ) | ( n6930 & n7218 ) | ( n7217 & n7218 ) ;
  assign n7221 = ( n6930 & n7219 ) | ( n6930 & ~n7220 ) | ( n7219 & ~n7220 ) ;
  assign n7222 = ( x72 & n7216 ) | ( x72 & ~n7221 ) | ( n7216 & ~n7221 ) ;
  assign n7223 = ( x72 & n6931 ) | ( x72 & ~n7173 ) | ( n6931 & ~n7173 ) ;
  assign n7224 = x72 & n6931 ;
  assign n7225 = ( n6936 & n7223 ) | ( n6936 & n7224 ) | ( n7223 & n7224 ) ;
  assign n7226 = ( ~n6936 & n7223 ) | ( ~n6936 & n7224 ) | ( n7223 & n7224 ) ;
  assign n7227 = ( n6936 & ~n7225 ) | ( n6936 & n7226 ) | ( ~n7225 & n7226 ) ;
  assign n7228 = ( x73 & n7222 ) | ( x73 & ~n7227 ) | ( n7222 & ~n7227 ) ;
  assign n7229 = ( x73 & n6937 ) | ( x73 & ~n7173 ) | ( n6937 & ~n7173 ) ;
  assign n7230 = x73 & n6937 ;
  assign n7231 = ( ~n6942 & n7229 ) | ( ~n6942 & n7230 ) | ( n7229 & n7230 ) ;
  assign n7232 = ( n6942 & n7229 ) | ( n6942 & n7230 ) | ( n7229 & n7230 ) ;
  assign n7233 = ( n6942 & n7231 ) | ( n6942 & ~n7232 ) | ( n7231 & ~n7232 ) ;
  assign n7234 = ( x74 & n7228 ) | ( x74 & ~n7233 ) | ( n7228 & ~n7233 ) ;
  assign n7235 = ( x74 & n6943 ) | ( x74 & ~n7173 ) | ( n6943 & ~n7173 ) ;
  assign n7236 = x74 & n6943 ;
  assign n7237 = ( n6948 & n7235 ) | ( n6948 & n7236 ) | ( n7235 & n7236 ) ;
  assign n7238 = ( ~n6948 & n7235 ) | ( ~n6948 & n7236 ) | ( n7235 & n7236 ) ;
  assign n7239 = ( n6948 & ~n7237 ) | ( n6948 & n7238 ) | ( ~n7237 & n7238 ) ;
  assign n7240 = ( x75 & n7234 ) | ( x75 & ~n7239 ) | ( n7234 & ~n7239 ) ;
  assign n7241 = ( x75 & n6949 ) | ( x75 & ~n7173 ) | ( n6949 & ~n7173 ) ;
  assign n7242 = x75 & n6949 ;
  assign n7243 = ( ~n6954 & n7241 ) | ( ~n6954 & n7242 ) | ( n7241 & n7242 ) ;
  assign n7244 = ( n6954 & n7241 ) | ( n6954 & n7242 ) | ( n7241 & n7242 ) ;
  assign n7245 = ( n6954 & n7243 ) | ( n6954 & ~n7244 ) | ( n7243 & ~n7244 ) ;
  assign n7246 = ( x76 & n7240 ) | ( x76 & ~n7245 ) | ( n7240 & ~n7245 ) ;
  assign n7247 = ( x76 & n6955 ) | ( x76 & ~n7173 ) | ( n6955 & ~n7173 ) ;
  assign n7248 = x76 & n6955 ;
  assign n7249 = ( n6960 & n7247 ) | ( n6960 & n7248 ) | ( n7247 & n7248 ) ;
  assign n7250 = ( ~n6960 & n7247 ) | ( ~n6960 & n7248 ) | ( n7247 & n7248 ) ;
  assign n7251 = ( n6960 & ~n7249 ) | ( n6960 & n7250 ) | ( ~n7249 & n7250 ) ;
  assign n7252 = ( x77 & n7246 ) | ( x77 & ~n7251 ) | ( n7246 & ~n7251 ) ;
  assign n7253 = ( x77 & n6961 ) | ( x77 & ~n7173 ) | ( n6961 & ~n7173 ) ;
  assign n7254 = x77 & n6961 ;
  assign n7255 = ( ~n6966 & n7253 ) | ( ~n6966 & n7254 ) | ( n7253 & n7254 ) ;
  assign n7256 = ( n6966 & n7253 ) | ( n6966 & n7254 ) | ( n7253 & n7254 ) ;
  assign n7257 = ( n6966 & n7255 ) | ( n6966 & ~n7256 ) | ( n7255 & ~n7256 ) ;
  assign n7258 = ( x78 & n7252 ) | ( x78 & ~n7257 ) | ( n7252 & ~n7257 ) ;
  assign n7259 = ( x78 & n6967 ) | ( x78 & ~n7173 ) | ( n6967 & ~n7173 ) ;
  assign n7260 = x78 & n6967 ;
  assign n7261 = ( n6972 & n7259 ) | ( n6972 & n7260 ) | ( n7259 & n7260 ) ;
  assign n7262 = ( ~n6972 & n7259 ) | ( ~n6972 & n7260 ) | ( n7259 & n7260 ) ;
  assign n7263 = ( n6972 & ~n7261 ) | ( n6972 & n7262 ) | ( ~n7261 & n7262 ) ;
  assign n7264 = ( x79 & n7258 ) | ( x79 & ~n7263 ) | ( n7258 & ~n7263 ) ;
  assign n7265 = ( x79 & n6973 ) | ( x79 & ~n7173 ) | ( n6973 & ~n7173 ) ;
  assign n7266 = x79 & n6973 ;
  assign n7267 = ( ~n6978 & n7265 ) | ( ~n6978 & n7266 ) | ( n7265 & n7266 ) ;
  assign n7268 = ( n6978 & n7265 ) | ( n6978 & n7266 ) | ( n7265 & n7266 ) ;
  assign n7269 = ( n6978 & n7267 ) | ( n6978 & ~n7268 ) | ( n7267 & ~n7268 ) ;
  assign n7270 = ( x80 & n7264 ) | ( x80 & ~n7269 ) | ( n7264 & ~n7269 ) ;
  assign n7271 = ( x80 & n6979 ) | ( x80 & ~n7173 ) | ( n6979 & ~n7173 ) ;
  assign n7272 = x80 & n6979 ;
  assign n7273 = ( n6984 & n7271 ) | ( n6984 & n7272 ) | ( n7271 & n7272 ) ;
  assign n7274 = ( ~n6984 & n7271 ) | ( ~n6984 & n7272 ) | ( n7271 & n7272 ) ;
  assign n7275 = ( n6984 & ~n7273 ) | ( n6984 & n7274 ) | ( ~n7273 & n7274 ) ;
  assign n7276 = ( x81 & n7270 ) | ( x81 & ~n7275 ) | ( n7270 & ~n7275 ) ;
  assign n7277 = ( x81 & n6985 ) | ( x81 & ~n7173 ) | ( n6985 & ~n7173 ) ;
  assign n7278 = x81 & n6985 ;
  assign n7279 = ( ~n6990 & n7277 ) | ( ~n6990 & n7278 ) | ( n7277 & n7278 ) ;
  assign n7280 = ( n6990 & n7277 ) | ( n6990 & n7278 ) | ( n7277 & n7278 ) ;
  assign n7281 = ( n6990 & n7279 ) | ( n6990 & ~n7280 ) | ( n7279 & ~n7280 ) ;
  assign n7282 = ( x82 & n7276 ) | ( x82 & ~n7281 ) | ( n7276 & ~n7281 ) ;
  assign n7283 = ( x82 & n6991 ) | ( x82 & ~n7173 ) | ( n6991 & ~n7173 ) ;
  assign n7284 = x82 & n6991 ;
  assign n7285 = ( n6996 & n7283 ) | ( n6996 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7286 = ( ~n6996 & n7283 ) | ( ~n6996 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7287 = ( n6996 & ~n7285 ) | ( n6996 & n7286 ) | ( ~n7285 & n7286 ) ;
  assign n7288 = ( x83 & n7282 ) | ( x83 & ~n7287 ) | ( n7282 & ~n7287 ) ;
  assign n7289 = ( x83 & n6997 ) | ( x83 & ~n7173 ) | ( n6997 & ~n7173 ) ;
  assign n7290 = x83 & n6997 ;
  assign n7291 = ( ~n7002 & n7289 ) | ( ~n7002 & n7290 ) | ( n7289 & n7290 ) ;
  assign n7292 = ( n7002 & n7289 ) | ( n7002 & n7290 ) | ( n7289 & n7290 ) ;
  assign n7293 = ( n7002 & n7291 ) | ( n7002 & ~n7292 ) | ( n7291 & ~n7292 ) ;
  assign n7294 = ( x84 & n7288 ) | ( x84 & ~n7293 ) | ( n7288 & ~n7293 ) ;
  assign n7295 = ( x84 & n7003 ) | ( x84 & ~n7173 ) | ( n7003 & ~n7173 ) ;
  assign n7296 = x84 & n7003 ;
  assign n7297 = ( n7008 & n7295 ) | ( n7008 & n7296 ) | ( n7295 & n7296 ) ;
  assign n7298 = ( ~n7008 & n7295 ) | ( ~n7008 & n7296 ) | ( n7295 & n7296 ) ;
  assign n7299 = ( n7008 & ~n7297 ) | ( n7008 & n7298 ) | ( ~n7297 & n7298 ) ;
  assign n7300 = ( x85 & n7294 ) | ( x85 & ~n7299 ) | ( n7294 & ~n7299 ) ;
  assign n7301 = ( x85 & n7009 ) | ( x85 & ~n7173 ) | ( n7009 & ~n7173 ) ;
  assign n7302 = x85 & n7009 ;
  assign n7303 = ( ~n7014 & n7301 ) | ( ~n7014 & n7302 ) | ( n7301 & n7302 ) ;
  assign n7304 = ( n7014 & n7301 ) | ( n7014 & n7302 ) | ( n7301 & n7302 ) ;
  assign n7305 = ( n7014 & n7303 ) | ( n7014 & ~n7304 ) | ( n7303 & ~n7304 ) ;
  assign n7306 = ( x86 & n7300 ) | ( x86 & ~n7305 ) | ( n7300 & ~n7305 ) ;
  assign n7307 = ( x86 & n7015 ) | ( x86 & ~n7173 ) | ( n7015 & ~n7173 ) ;
  assign n7308 = x86 & n7015 ;
  assign n7309 = ( n7020 & n7307 ) | ( n7020 & n7308 ) | ( n7307 & n7308 ) ;
  assign n7310 = ( ~n7020 & n7307 ) | ( ~n7020 & n7308 ) | ( n7307 & n7308 ) ;
  assign n7311 = ( n7020 & ~n7309 ) | ( n7020 & n7310 ) | ( ~n7309 & n7310 ) ;
  assign n7312 = ( x87 & n7306 ) | ( x87 & ~n7311 ) | ( n7306 & ~n7311 ) ;
  assign n7313 = ( x87 & n7021 ) | ( x87 & ~n7173 ) | ( n7021 & ~n7173 ) ;
  assign n7314 = x87 & n7021 ;
  assign n7315 = ( ~n7026 & n7313 ) | ( ~n7026 & n7314 ) | ( n7313 & n7314 ) ;
  assign n7316 = ( n7026 & n7313 ) | ( n7026 & n7314 ) | ( n7313 & n7314 ) ;
  assign n7317 = ( n7026 & n7315 ) | ( n7026 & ~n7316 ) | ( n7315 & ~n7316 ) ;
  assign n7318 = ( x88 & n7312 ) | ( x88 & ~n7317 ) | ( n7312 & ~n7317 ) ;
  assign n7319 = ( x88 & n7027 ) | ( x88 & ~n7173 ) | ( n7027 & ~n7173 ) ;
  assign n7320 = x88 & n7027 ;
  assign n7321 = ( n7032 & n7319 ) | ( n7032 & n7320 ) | ( n7319 & n7320 ) ;
  assign n7322 = ( ~n7032 & n7319 ) | ( ~n7032 & n7320 ) | ( n7319 & n7320 ) ;
  assign n7323 = ( n7032 & ~n7321 ) | ( n7032 & n7322 ) | ( ~n7321 & n7322 ) ;
  assign n7324 = ( x89 & n7318 ) | ( x89 & ~n7323 ) | ( n7318 & ~n7323 ) ;
  assign n7325 = ( x89 & n7033 ) | ( x89 & ~n7173 ) | ( n7033 & ~n7173 ) ;
  assign n7326 = x89 & n7033 ;
  assign n7327 = ( ~n7038 & n7325 ) | ( ~n7038 & n7326 ) | ( n7325 & n7326 ) ;
  assign n7328 = ( n7038 & n7325 ) | ( n7038 & n7326 ) | ( n7325 & n7326 ) ;
  assign n7329 = ( n7038 & n7327 ) | ( n7038 & ~n7328 ) | ( n7327 & ~n7328 ) ;
  assign n7330 = ( x90 & n7324 ) | ( x90 & ~n7329 ) | ( n7324 & ~n7329 ) ;
  assign n7331 = ( x90 & n7039 ) | ( x90 & ~n7173 ) | ( n7039 & ~n7173 ) ;
  assign n7332 = x90 & n7039 ;
  assign n7333 = ( n7044 & n7331 ) | ( n7044 & n7332 ) | ( n7331 & n7332 ) ;
  assign n7334 = ( ~n7044 & n7331 ) | ( ~n7044 & n7332 ) | ( n7331 & n7332 ) ;
  assign n7335 = ( n7044 & ~n7333 ) | ( n7044 & n7334 ) | ( ~n7333 & n7334 ) ;
  assign n7336 = ( x91 & n7330 ) | ( x91 & ~n7335 ) | ( n7330 & ~n7335 ) ;
  assign n7337 = ( x91 & n7045 ) | ( x91 & ~n7173 ) | ( n7045 & ~n7173 ) ;
  assign n7338 = x91 & n7045 ;
  assign n7339 = ( ~n7050 & n7337 ) | ( ~n7050 & n7338 ) | ( n7337 & n7338 ) ;
  assign n7340 = ( n7050 & n7337 ) | ( n7050 & n7338 ) | ( n7337 & n7338 ) ;
  assign n7341 = ( n7050 & n7339 ) | ( n7050 & ~n7340 ) | ( n7339 & ~n7340 ) ;
  assign n7342 = ( x92 & n7336 ) | ( x92 & ~n7341 ) | ( n7336 & ~n7341 ) ;
  assign n7343 = ( x92 & n7051 ) | ( x92 & ~n7173 ) | ( n7051 & ~n7173 ) ;
  assign n7344 = x92 & n7051 ;
  assign n7345 = ( n7056 & n7343 ) | ( n7056 & n7344 ) | ( n7343 & n7344 ) ;
  assign n7346 = ( ~n7056 & n7343 ) | ( ~n7056 & n7344 ) | ( n7343 & n7344 ) ;
  assign n7347 = ( n7056 & ~n7345 ) | ( n7056 & n7346 ) | ( ~n7345 & n7346 ) ;
  assign n7348 = ( x93 & n7342 ) | ( x93 & ~n7347 ) | ( n7342 & ~n7347 ) ;
  assign n7349 = ( x93 & n7057 ) | ( x93 & ~n7173 ) | ( n7057 & ~n7173 ) ;
  assign n7350 = x93 & n7057 ;
  assign n7351 = ( ~n7062 & n7349 ) | ( ~n7062 & n7350 ) | ( n7349 & n7350 ) ;
  assign n7352 = ( n7062 & n7349 ) | ( n7062 & n7350 ) | ( n7349 & n7350 ) ;
  assign n7353 = ( n7062 & n7351 ) | ( n7062 & ~n7352 ) | ( n7351 & ~n7352 ) ;
  assign n7354 = ( x94 & n7348 ) | ( x94 & ~n7353 ) | ( n7348 & ~n7353 ) ;
  assign n7355 = ( x94 & n7063 ) | ( x94 & ~n7173 ) | ( n7063 & ~n7173 ) ;
  assign n7356 = x94 & n7063 ;
  assign n7357 = ( n7068 & n7355 ) | ( n7068 & n7356 ) | ( n7355 & n7356 ) ;
  assign n7358 = ( ~n7068 & n7355 ) | ( ~n7068 & n7356 ) | ( n7355 & n7356 ) ;
  assign n7359 = ( n7068 & ~n7357 ) | ( n7068 & n7358 ) | ( ~n7357 & n7358 ) ;
  assign n7360 = ( x95 & n7354 ) | ( x95 & ~n7359 ) | ( n7354 & ~n7359 ) ;
  assign n7361 = ( x95 & n7069 ) | ( x95 & ~n7173 ) | ( n7069 & ~n7173 ) ;
  assign n7362 = x95 & n7069 ;
  assign n7363 = ( ~n7074 & n7361 ) | ( ~n7074 & n7362 ) | ( n7361 & n7362 ) ;
  assign n7364 = ( n7074 & n7361 ) | ( n7074 & n7362 ) | ( n7361 & n7362 ) ;
  assign n7365 = ( n7074 & n7363 ) | ( n7074 & ~n7364 ) | ( n7363 & ~n7364 ) ;
  assign n7366 = ( x96 & n7360 ) | ( x96 & ~n7365 ) | ( n7360 & ~n7365 ) ;
  assign n7367 = ( x96 & n7075 ) | ( x96 & ~n7173 ) | ( n7075 & ~n7173 ) ;
  assign n7368 = x96 & n7075 ;
  assign n7369 = ( n7080 & n7367 ) | ( n7080 & n7368 ) | ( n7367 & n7368 ) ;
  assign n7370 = ( ~n7080 & n7367 ) | ( ~n7080 & n7368 ) | ( n7367 & n7368 ) ;
  assign n7371 = ( n7080 & ~n7369 ) | ( n7080 & n7370 ) | ( ~n7369 & n7370 ) ;
  assign n7372 = ( x97 & n7366 ) | ( x97 & ~n7371 ) | ( n7366 & ~n7371 ) ;
  assign n7373 = ( x97 & n7081 ) | ( x97 & ~n7173 ) | ( n7081 & ~n7173 ) ;
  assign n7374 = x97 & n7081 ;
  assign n7375 = ( ~n7086 & n7373 ) | ( ~n7086 & n7374 ) | ( n7373 & n7374 ) ;
  assign n7376 = ( n7086 & n7373 ) | ( n7086 & n7374 ) | ( n7373 & n7374 ) ;
  assign n7377 = ( n7086 & n7375 ) | ( n7086 & ~n7376 ) | ( n7375 & ~n7376 ) ;
  assign n7378 = ( x98 & n7372 ) | ( x98 & ~n7377 ) | ( n7372 & ~n7377 ) ;
  assign n7379 = ( x98 & n7087 ) | ( x98 & ~n7173 ) | ( n7087 & ~n7173 ) ;
  assign n7380 = x98 & n7087 ;
  assign n7381 = ( n7092 & n7379 ) | ( n7092 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7382 = ( ~n7092 & n7379 ) | ( ~n7092 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7383 = ( n7092 & ~n7381 ) | ( n7092 & n7382 ) | ( ~n7381 & n7382 ) ;
  assign n7384 = ( x99 & n7378 ) | ( x99 & ~n7383 ) | ( n7378 & ~n7383 ) ;
  assign n7385 = ( x99 & n7093 ) | ( x99 & ~n7173 ) | ( n7093 & ~n7173 ) ;
  assign n7386 = x99 & n7093 ;
  assign n7387 = ( ~n7098 & n7385 ) | ( ~n7098 & n7386 ) | ( n7385 & n7386 ) ;
  assign n7388 = ( n7098 & n7385 ) | ( n7098 & n7386 ) | ( n7385 & n7386 ) ;
  assign n7389 = ( n7098 & n7387 ) | ( n7098 & ~n7388 ) | ( n7387 & ~n7388 ) ;
  assign n7390 = ( x100 & n7384 ) | ( x100 & ~n7389 ) | ( n7384 & ~n7389 ) ;
  assign n7391 = ( x100 & n7099 ) | ( x100 & ~n7173 ) | ( n7099 & ~n7173 ) ;
  assign n7392 = x100 & n7099 ;
  assign n7393 = ( n7104 & n7391 ) | ( n7104 & n7392 ) | ( n7391 & n7392 ) ;
  assign n7394 = ( ~n7104 & n7391 ) | ( ~n7104 & n7392 ) | ( n7391 & n7392 ) ;
  assign n7395 = ( n7104 & ~n7393 ) | ( n7104 & n7394 ) | ( ~n7393 & n7394 ) ;
  assign n7396 = ( x101 & n7390 ) | ( x101 & ~n7395 ) | ( n7390 & ~n7395 ) ;
  assign n7397 = ( x101 & n7105 ) | ( x101 & ~n7173 ) | ( n7105 & ~n7173 ) ;
  assign n7398 = x101 & n7105 ;
  assign n7399 = ( ~n7110 & n7397 ) | ( ~n7110 & n7398 ) | ( n7397 & n7398 ) ;
  assign n7400 = ( n7110 & n7397 ) | ( n7110 & n7398 ) | ( n7397 & n7398 ) ;
  assign n7401 = ( n7110 & n7399 ) | ( n7110 & ~n7400 ) | ( n7399 & ~n7400 ) ;
  assign n7402 = ( x102 & n7396 ) | ( x102 & ~n7401 ) | ( n7396 & ~n7401 ) ;
  assign n7403 = ( x102 & n7111 ) | ( x102 & ~n7173 ) | ( n7111 & ~n7173 ) ;
  assign n7404 = x102 & n7111 ;
  assign n7405 = ( n7116 & n7403 ) | ( n7116 & n7404 ) | ( n7403 & n7404 ) ;
  assign n7406 = ( ~n7116 & n7403 ) | ( ~n7116 & n7404 ) | ( n7403 & n7404 ) ;
  assign n7407 = ( n7116 & ~n7405 ) | ( n7116 & n7406 ) | ( ~n7405 & n7406 ) ;
  assign n7408 = ( x103 & n7402 ) | ( x103 & ~n7407 ) | ( n7402 & ~n7407 ) ;
  assign n7409 = ( x103 & n7117 ) | ( x103 & ~n7173 ) | ( n7117 & ~n7173 ) ;
  assign n7410 = x103 & n7117 ;
  assign n7411 = ( ~n7122 & n7409 ) | ( ~n7122 & n7410 ) | ( n7409 & n7410 ) ;
  assign n7412 = ( n7122 & n7409 ) | ( n7122 & n7410 ) | ( n7409 & n7410 ) ;
  assign n7413 = ( n7122 & n7411 ) | ( n7122 & ~n7412 ) | ( n7411 & ~n7412 ) ;
  assign n7414 = ( x104 & n7408 ) | ( x104 & ~n7413 ) | ( n7408 & ~n7413 ) ;
  assign n7415 = ( x104 & n7123 ) | ( x104 & ~n7173 ) | ( n7123 & ~n7173 ) ;
  assign n7416 = x104 & n7123 ;
  assign n7417 = ( n7128 & n7415 ) | ( n7128 & n7416 ) | ( n7415 & n7416 ) ;
  assign n7418 = ( ~n7128 & n7415 ) | ( ~n7128 & n7416 ) | ( n7415 & n7416 ) ;
  assign n7419 = ( n7128 & ~n7417 ) | ( n7128 & n7418 ) | ( ~n7417 & n7418 ) ;
  assign n7420 = ( x105 & n7414 ) | ( x105 & ~n7419 ) | ( n7414 & ~n7419 ) ;
  assign n7421 = ( x105 & n7129 ) | ( x105 & ~n7173 ) | ( n7129 & ~n7173 ) ;
  assign n7422 = x105 & n7129 ;
  assign n7423 = ( ~n7134 & n7421 ) | ( ~n7134 & n7422 ) | ( n7421 & n7422 ) ;
  assign n7424 = ( n7134 & n7421 ) | ( n7134 & n7422 ) | ( n7421 & n7422 ) ;
  assign n7425 = ( n7134 & n7423 ) | ( n7134 & ~n7424 ) | ( n7423 & ~n7424 ) ;
  assign n7426 = ( x106 & n7420 ) | ( x106 & ~n7425 ) | ( n7420 & ~n7425 ) ;
  assign n7427 = ( x106 & n7135 ) | ( x106 & ~n7173 ) | ( n7135 & ~n7173 ) ;
  assign n7428 = x106 & n7135 ;
  assign n7429 = ( n7140 & n7427 ) | ( n7140 & n7428 ) | ( n7427 & n7428 ) ;
  assign n7430 = ( ~n7140 & n7427 ) | ( ~n7140 & n7428 ) | ( n7427 & n7428 ) ;
  assign n7431 = ( n7140 & ~n7429 ) | ( n7140 & n7430 ) | ( ~n7429 & n7430 ) ;
  assign n7432 = ( x107 & n7426 ) | ( x107 & ~n7431 ) | ( n7426 & ~n7431 ) ;
  assign n7433 = ( x107 & n7141 ) | ( x107 & ~n7173 ) | ( n7141 & ~n7173 ) ;
  assign n7434 = x107 & n7141 ;
  assign n7435 = ( ~n7146 & n7433 ) | ( ~n7146 & n7434 ) | ( n7433 & n7434 ) ;
  assign n7436 = ( n7146 & n7433 ) | ( n7146 & n7434 ) | ( n7433 & n7434 ) ;
  assign n7437 = ( n7146 & n7435 ) | ( n7146 & ~n7436 ) | ( n7435 & ~n7436 ) ;
  assign n7438 = ( x108 & n7432 ) | ( x108 & ~n7437 ) | ( n7432 & ~n7437 ) ;
  assign n7439 = ( x108 & n7147 ) | ( x108 & ~n7173 ) | ( n7147 & ~n7173 ) ;
  assign n7440 = x108 & n7147 ;
  assign n7441 = ( n7152 & n7439 ) | ( n7152 & n7440 ) | ( n7439 & n7440 ) ;
  assign n7442 = ( ~n7152 & n7439 ) | ( ~n7152 & n7440 ) | ( n7439 & n7440 ) ;
  assign n7443 = ( n7152 & ~n7441 ) | ( n7152 & n7442 ) | ( ~n7441 & n7442 ) ;
  assign n7444 = ( x109 & n7438 ) | ( x109 & ~n7443 ) | ( n7438 & ~n7443 ) ;
  assign n7445 = ( x109 & n7153 ) | ( x109 & ~n7173 ) | ( n7153 & ~n7173 ) ;
  assign n7446 = x109 & n7153 ;
  assign n7447 = ( ~n7158 & n7445 ) | ( ~n7158 & n7446 ) | ( n7445 & n7446 ) ;
  assign n7448 = ( n7158 & n7445 ) | ( n7158 & n7446 ) | ( n7445 & n7446 ) ;
  assign n7449 = ( n7158 & n7447 ) | ( n7158 & ~n7448 ) | ( n7447 & ~n7448 ) ;
  assign n7450 = ( x110 & n7444 ) | ( x110 & ~n7449 ) | ( n7444 & ~n7449 ) ;
  assign n7451 = ( x110 & n7159 ) | ( x110 & ~n7173 ) | ( n7159 & ~n7173 ) ;
  assign n7452 = x110 & n7159 ;
  assign n7453 = ( n7164 & n7451 ) | ( n7164 & n7452 ) | ( n7451 & n7452 ) ;
  assign n7454 = ( ~n7164 & n7451 ) | ( ~n7164 & n7452 ) | ( n7451 & n7452 ) ;
  assign n7455 = ( n7164 & ~n7453 ) | ( n7164 & n7454 ) | ( ~n7453 & n7454 ) ;
  assign n7456 = ( x111 & n7450 ) | ( x111 & ~n7455 ) | ( n7450 & ~n7455 ) ;
  assign n7457 = ( x111 & n7165 ) | ( x111 & ~n7173 ) | ( n7165 & ~n7173 ) ;
  assign n7458 = x111 & n7165 ;
  assign n7459 = ( n7170 & n7457 ) | ( n7170 & n7458 ) | ( n7457 & n7458 ) ;
  assign n7460 = ( ~n7170 & n7457 ) | ( ~n7170 & n7458 ) | ( n7457 & n7458 ) ;
  assign n7461 = ( n7170 & ~n7459 ) | ( n7170 & n7460 ) | ( ~n7459 & n7460 ) ;
  assign n7462 = ( x112 & n7456 ) | ( x112 & ~n7461 ) | ( n7456 & ~n7461 ) ;
  assign n7463 = ( x113 & ~n7175 ) | ( x113 & n7462 ) | ( ~n7175 & n7462 ) ;
  assign n7464 = n144 | n7463 ;
  assign n7465 = ( n280 & n7175 ) | ( n280 & n7464 ) | ( n7175 & n7464 ) ;
  assign n7466 = ( x14 & ~x64 ) | ( x14 & n7464 ) | ( ~x64 & n7464 ) ;
  assign n7467 = ~x14 & n7464 ;
  assign n7468 = ( n7179 & n7466 ) | ( n7179 & ~n7467 ) | ( n7466 & ~n7467 ) ;
  assign n7469 = ~x13 & x64 ;
  assign n7470 = ( x65 & ~n7468 ) | ( x65 & n7469 ) | ( ~n7468 & n7469 ) ;
  assign n7471 = ( x65 & n7179 ) | ( x65 & ~n7464 ) | ( n7179 & ~n7464 ) ;
  assign n7472 = x65 & n7179 ;
  assign n7473 = ( n7178 & n7471 ) | ( n7178 & n7472 ) | ( n7471 & n7472 ) ;
  assign n7474 = ( ~n7178 & n7471 ) | ( ~n7178 & n7472 ) | ( n7471 & n7472 ) ;
  assign n7475 = ( n7178 & ~n7473 ) | ( n7178 & n7474 ) | ( ~n7473 & n7474 ) ;
  assign n7476 = ( x66 & n7470 ) | ( x66 & ~n7475 ) | ( n7470 & ~n7475 ) ;
  assign n7477 = ( x66 & n7180 ) | ( x66 & ~n7464 ) | ( n7180 & ~n7464 ) ;
  assign n7478 = x66 & n7180 ;
  assign n7479 = ( n7185 & n7477 ) | ( n7185 & n7478 ) | ( n7477 & n7478 ) ;
  assign n7480 = ( ~n7185 & n7477 ) | ( ~n7185 & n7478 ) | ( n7477 & n7478 ) ;
  assign n7481 = ( n7185 & ~n7479 ) | ( n7185 & n7480 ) | ( ~n7479 & n7480 ) ;
  assign n7482 = ( x67 & n7476 ) | ( x67 & ~n7481 ) | ( n7476 & ~n7481 ) ;
  assign n7483 = ( x67 & n7186 ) | ( x67 & ~n7464 ) | ( n7186 & ~n7464 ) ;
  assign n7484 = x67 & n7186 ;
  assign n7485 = ( ~n7191 & n7483 ) | ( ~n7191 & n7484 ) | ( n7483 & n7484 ) ;
  assign n7486 = ( n7191 & n7483 ) | ( n7191 & n7484 ) | ( n7483 & n7484 ) ;
  assign n7487 = ( n7191 & n7485 ) | ( n7191 & ~n7486 ) | ( n7485 & ~n7486 ) ;
  assign n7488 = ( x68 & n7482 ) | ( x68 & ~n7487 ) | ( n7482 & ~n7487 ) ;
  assign n7489 = ( x68 & n7192 ) | ( x68 & ~n7464 ) | ( n7192 & ~n7464 ) ;
  assign n7490 = x68 & n7192 ;
  assign n7491 = ( n7197 & n7489 ) | ( n7197 & n7490 ) | ( n7489 & n7490 ) ;
  assign n7492 = ( ~n7197 & n7489 ) | ( ~n7197 & n7490 ) | ( n7489 & n7490 ) ;
  assign n7493 = ( n7197 & ~n7491 ) | ( n7197 & n7492 ) | ( ~n7491 & n7492 ) ;
  assign n7494 = ( x69 & n7488 ) | ( x69 & ~n7493 ) | ( n7488 & ~n7493 ) ;
  assign n7495 = ( x69 & n7198 ) | ( x69 & ~n7464 ) | ( n7198 & ~n7464 ) ;
  assign n7496 = x69 & n7198 ;
  assign n7497 = ( ~n7203 & n7495 ) | ( ~n7203 & n7496 ) | ( n7495 & n7496 ) ;
  assign n7498 = ( n7203 & n7495 ) | ( n7203 & n7496 ) | ( n7495 & n7496 ) ;
  assign n7499 = ( n7203 & n7497 ) | ( n7203 & ~n7498 ) | ( n7497 & ~n7498 ) ;
  assign n7500 = ( x70 & n7494 ) | ( x70 & ~n7499 ) | ( n7494 & ~n7499 ) ;
  assign n7501 = ( x70 & n7204 ) | ( x70 & ~n7464 ) | ( n7204 & ~n7464 ) ;
  assign n7502 = x70 & n7204 ;
  assign n7503 = ( n7209 & n7501 ) | ( n7209 & n7502 ) | ( n7501 & n7502 ) ;
  assign n7504 = ( ~n7209 & n7501 ) | ( ~n7209 & n7502 ) | ( n7501 & n7502 ) ;
  assign n7505 = ( n7209 & ~n7503 ) | ( n7209 & n7504 ) | ( ~n7503 & n7504 ) ;
  assign n7506 = ( x71 & n7500 ) | ( x71 & ~n7505 ) | ( n7500 & ~n7505 ) ;
  assign n7507 = ( x71 & n7210 ) | ( x71 & ~n7464 ) | ( n7210 & ~n7464 ) ;
  assign n7508 = x71 & n7210 ;
  assign n7509 = ( ~n7215 & n7507 ) | ( ~n7215 & n7508 ) | ( n7507 & n7508 ) ;
  assign n7510 = ( n7215 & n7507 ) | ( n7215 & n7508 ) | ( n7507 & n7508 ) ;
  assign n7511 = ( n7215 & n7509 ) | ( n7215 & ~n7510 ) | ( n7509 & ~n7510 ) ;
  assign n7512 = ( x72 & n7506 ) | ( x72 & ~n7511 ) | ( n7506 & ~n7511 ) ;
  assign n7513 = ( x72 & n7216 ) | ( x72 & ~n7464 ) | ( n7216 & ~n7464 ) ;
  assign n7514 = x72 & n7216 ;
  assign n7515 = ( n7221 & n7513 ) | ( n7221 & n7514 ) | ( n7513 & n7514 ) ;
  assign n7516 = ( ~n7221 & n7513 ) | ( ~n7221 & n7514 ) | ( n7513 & n7514 ) ;
  assign n7517 = ( n7221 & ~n7515 ) | ( n7221 & n7516 ) | ( ~n7515 & n7516 ) ;
  assign n7518 = ( x73 & n7512 ) | ( x73 & ~n7517 ) | ( n7512 & ~n7517 ) ;
  assign n7519 = ( x73 & n7222 ) | ( x73 & ~n7464 ) | ( n7222 & ~n7464 ) ;
  assign n7520 = x73 & n7222 ;
  assign n7521 = ( ~n7227 & n7519 ) | ( ~n7227 & n7520 ) | ( n7519 & n7520 ) ;
  assign n7522 = ( n7227 & n7519 ) | ( n7227 & n7520 ) | ( n7519 & n7520 ) ;
  assign n7523 = ( n7227 & n7521 ) | ( n7227 & ~n7522 ) | ( n7521 & ~n7522 ) ;
  assign n7524 = ( x74 & n7518 ) | ( x74 & ~n7523 ) | ( n7518 & ~n7523 ) ;
  assign n7525 = ( x74 & n7228 ) | ( x74 & ~n7464 ) | ( n7228 & ~n7464 ) ;
  assign n7526 = x74 & n7228 ;
  assign n7527 = ( n7233 & n7525 ) | ( n7233 & n7526 ) | ( n7525 & n7526 ) ;
  assign n7528 = ( ~n7233 & n7525 ) | ( ~n7233 & n7526 ) | ( n7525 & n7526 ) ;
  assign n7529 = ( n7233 & ~n7527 ) | ( n7233 & n7528 ) | ( ~n7527 & n7528 ) ;
  assign n7530 = ( x75 & n7524 ) | ( x75 & ~n7529 ) | ( n7524 & ~n7529 ) ;
  assign n7531 = ( x75 & n7234 ) | ( x75 & ~n7464 ) | ( n7234 & ~n7464 ) ;
  assign n7532 = x75 & n7234 ;
  assign n7533 = ( ~n7239 & n7531 ) | ( ~n7239 & n7532 ) | ( n7531 & n7532 ) ;
  assign n7534 = ( n7239 & n7531 ) | ( n7239 & n7532 ) | ( n7531 & n7532 ) ;
  assign n7535 = ( n7239 & n7533 ) | ( n7239 & ~n7534 ) | ( n7533 & ~n7534 ) ;
  assign n7536 = ( x76 & n7530 ) | ( x76 & ~n7535 ) | ( n7530 & ~n7535 ) ;
  assign n7537 = ( x76 & n7240 ) | ( x76 & ~n7464 ) | ( n7240 & ~n7464 ) ;
  assign n7538 = x76 & n7240 ;
  assign n7539 = ( n7245 & n7537 ) | ( n7245 & n7538 ) | ( n7537 & n7538 ) ;
  assign n7540 = ( ~n7245 & n7537 ) | ( ~n7245 & n7538 ) | ( n7537 & n7538 ) ;
  assign n7541 = ( n7245 & ~n7539 ) | ( n7245 & n7540 ) | ( ~n7539 & n7540 ) ;
  assign n7542 = ( x77 & n7536 ) | ( x77 & ~n7541 ) | ( n7536 & ~n7541 ) ;
  assign n7543 = ( x77 & n7246 ) | ( x77 & ~n7464 ) | ( n7246 & ~n7464 ) ;
  assign n7544 = x77 & n7246 ;
  assign n7545 = ( ~n7251 & n7543 ) | ( ~n7251 & n7544 ) | ( n7543 & n7544 ) ;
  assign n7546 = ( n7251 & n7543 ) | ( n7251 & n7544 ) | ( n7543 & n7544 ) ;
  assign n7547 = ( n7251 & n7545 ) | ( n7251 & ~n7546 ) | ( n7545 & ~n7546 ) ;
  assign n7548 = ( x78 & n7542 ) | ( x78 & ~n7547 ) | ( n7542 & ~n7547 ) ;
  assign n7549 = ( x78 & n7252 ) | ( x78 & ~n7464 ) | ( n7252 & ~n7464 ) ;
  assign n7550 = x78 & n7252 ;
  assign n7551 = ( n7257 & n7549 ) | ( n7257 & n7550 ) | ( n7549 & n7550 ) ;
  assign n7552 = ( ~n7257 & n7549 ) | ( ~n7257 & n7550 ) | ( n7549 & n7550 ) ;
  assign n7553 = ( n7257 & ~n7551 ) | ( n7257 & n7552 ) | ( ~n7551 & n7552 ) ;
  assign n7554 = ( x79 & n7548 ) | ( x79 & ~n7553 ) | ( n7548 & ~n7553 ) ;
  assign n7555 = ( x79 & n7258 ) | ( x79 & ~n7464 ) | ( n7258 & ~n7464 ) ;
  assign n7556 = x79 & n7258 ;
  assign n7557 = ( ~n7263 & n7555 ) | ( ~n7263 & n7556 ) | ( n7555 & n7556 ) ;
  assign n7558 = ( n7263 & n7555 ) | ( n7263 & n7556 ) | ( n7555 & n7556 ) ;
  assign n7559 = ( n7263 & n7557 ) | ( n7263 & ~n7558 ) | ( n7557 & ~n7558 ) ;
  assign n7560 = ( x80 & n7554 ) | ( x80 & ~n7559 ) | ( n7554 & ~n7559 ) ;
  assign n7561 = ( x80 & n7264 ) | ( x80 & ~n7464 ) | ( n7264 & ~n7464 ) ;
  assign n7562 = x80 & n7264 ;
  assign n7563 = ( n7269 & n7561 ) | ( n7269 & n7562 ) | ( n7561 & n7562 ) ;
  assign n7564 = ( ~n7269 & n7561 ) | ( ~n7269 & n7562 ) | ( n7561 & n7562 ) ;
  assign n7565 = ( n7269 & ~n7563 ) | ( n7269 & n7564 ) | ( ~n7563 & n7564 ) ;
  assign n7566 = ( x81 & n7560 ) | ( x81 & ~n7565 ) | ( n7560 & ~n7565 ) ;
  assign n7567 = ( x81 & n7270 ) | ( x81 & ~n7464 ) | ( n7270 & ~n7464 ) ;
  assign n7568 = x81 & n7270 ;
  assign n7569 = ( ~n7275 & n7567 ) | ( ~n7275 & n7568 ) | ( n7567 & n7568 ) ;
  assign n7570 = ( n7275 & n7567 ) | ( n7275 & n7568 ) | ( n7567 & n7568 ) ;
  assign n7571 = ( n7275 & n7569 ) | ( n7275 & ~n7570 ) | ( n7569 & ~n7570 ) ;
  assign n7572 = ( x82 & n7566 ) | ( x82 & ~n7571 ) | ( n7566 & ~n7571 ) ;
  assign n7573 = ( x82 & n7276 ) | ( x82 & ~n7464 ) | ( n7276 & ~n7464 ) ;
  assign n7574 = x82 & n7276 ;
  assign n7575 = ( n7281 & n7573 ) | ( n7281 & n7574 ) | ( n7573 & n7574 ) ;
  assign n7576 = ( ~n7281 & n7573 ) | ( ~n7281 & n7574 ) | ( n7573 & n7574 ) ;
  assign n7577 = ( n7281 & ~n7575 ) | ( n7281 & n7576 ) | ( ~n7575 & n7576 ) ;
  assign n7578 = ( x83 & n7572 ) | ( x83 & ~n7577 ) | ( n7572 & ~n7577 ) ;
  assign n7579 = ( x83 & n7282 ) | ( x83 & ~n7464 ) | ( n7282 & ~n7464 ) ;
  assign n7580 = x83 & n7282 ;
  assign n7581 = ( ~n7287 & n7579 ) | ( ~n7287 & n7580 ) | ( n7579 & n7580 ) ;
  assign n7582 = ( n7287 & n7579 ) | ( n7287 & n7580 ) | ( n7579 & n7580 ) ;
  assign n7583 = ( n7287 & n7581 ) | ( n7287 & ~n7582 ) | ( n7581 & ~n7582 ) ;
  assign n7584 = ( x84 & n7578 ) | ( x84 & ~n7583 ) | ( n7578 & ~n7583 ) ;
  assign n7585 = ( x84 & n7288 ) | ( x84 & ~n7464 ) | ( n7288 & ~n7464 ) ;
  assign n7586 = x84 & n7288 ;
  assign n7587 = ( n7293 & n7585 ) | ( n7293 & n7586 ) | ( n7585 & n7586 ) ;
  assign n7588 = ( ~n7293 & n7585 ) | ( ~n7293 & n7586 ) | ( n7585 & n7586 ) ;
  assign n7589 = ( n7293 & ~n7587 ) | ( n7293 & n7588 ) | ( ~n7587 & n7588 ) ;
  assign n7590 = ( x85 & n7584 ) | ( x85 & ~n7589 ) | ( n7584 & ~n7589 ) ;
  assign n7591 = ( x85 & n7294 ) | ( x85 & ~n7464 ) | ( n7294 & ~n7464 ) ;
  assign n7592 = x85 & n7294 ;
  assign n7593 = ( ~n7299 & n7591 ) | ( ~n7299 & n7592 ) | ( n7591 & n7592 ) ;
  assign n7594 = ( n7299 & n7591 ) | ( n7299 & n7592 ) | ( n7591 & n7592 ) ;
  assign n7595 = ( n7299 & n7593 ) | ( n7299 & ~n7594 ) | ( n7593 & ~n7594 ) ;
  assign n7596 = ( x86 & n7590 ) | ( x86 & ~n7595 ) | ( n7590 & ~n7595 ) ;
  assign n7597 = ( x86 & n7300 ) | ( x86 & ~n7464 ) | ( n7300 & ~n7464 ) ;
  assign n7598 = x86 & n7300 ;
  assign n7599 = ( n7305 & n7597 ) | ( n7305 & n7598 ) | ( n7597 & n7598 ) ;
  assign n7600 = ( ~n7305 & n7597 ) | ( ~n7305 & n7598 ) | ( n7597 & n7598 ) ;
  assign n7601 = ( n7305 & ~n7599 ) | ( n7305 & n7600 ) | ( ~n7599 & n7600 ) ;
  assign n7602 = ( x87 & n7596 ) | ( x87 & ~n7601 ) | ( n7596 & ~n7601 ) ;
  assign n7603 = ( x87 & n7306 ) | ( x87 & ~n7464 ) | ( n7306 & ~n7464 ) ;
  assign n7604 = x87 & n7306 ;
  assign n7605 = ( ~n7311 & n7603 ) | ( ~n7311 & n7604 ) | ( n7603 & n7604 ) ;
  assign n7606 = ( n7311 & n7603 ) | ( n7311 & n7604 ) | ( n7603 & n7604 ) ;
  assign n7607 = ( n7311 & n7605 ) | ( n7311 & ~n7606 ) | ( n7605 & ~n7606 ) ;
  assign n7608 = ( x88 & n7602 ) | ( x88 & ~n7607 ) | ( n7602 & ~n7607 ) ;
  assign n7609 = ( x88 & n7312 ) | ( x88 & ~n7464 ) | ( n7312 & ~n7464 ) ;
  assign n7610 = x88 & n7312 ;
  assign n7611 = ( n7317 & n7609 ) | ( n7317 & n7610 ) | ( n7609 & n7610 ) ;
  assign n7612 = ( ~n7317 & n7609 ) | ( ~n7317 & n7610 ) | ( n7609 & n7610 ) ;
  assign n7613 = ( n7317 & ~n7611 ) | ( n7317 & n7612 ) | ( ~n7611 & n7612 ) ;
  assign n7614 = ( x89 & n7608 ) | ( x89 & ~n7613 ) | ( n7608 & ~n7613 ) ;
  assign n7615 = ( x89 & n7318 ) | ( x89 & ~n7464 ) | ( n7318 & ~n7464 ) ;
  assign n7616 = x89 & n7318 ;
  assign n7617 = ( ~n7323 & n7615 ) | ( ~n7323 & n7616 ) | ( n7615 & n7616 ) ;
  assign n7618 = ( n7323 & n7615 ) | ( n7323 & n7616 ) | ( n7615 & n7616 ) ;
  assign n7619 = ( n7323 & n7617 ) | ( n7323 & ~n7618 ) | ( n7617 & ~n7618 ) ;
  assign n7620 = ( x90 & n7614 ) | ( x90 & ~n7619 ) | ( n7614 & ~n7619 ) ;
  assign n7621 = ( x90 & n7324 ) | ( x90 & ~n7464 ) | ( n7324 & ~n7464 ) ;
  assign n7622 = x90 & n7324 ;
  assign n7623 = ( n7329 & n7621 ) | ( n7329 & n7622 ) | ( n7621 & n7622 ) ;
  assign n7624 = ( ~n7329 & n7621 ) | ( ~n7329 & n7622 ) | ( n7621 & n7622 ) ;
  assign n7625 = ( n7329 & ~n7623 ) | ( n7329 & n7624 ) | ( ~n7623 & n7624 ) ;
  assign n7626 = ( x91 & n7620 ) | ( x91 & ~n7625 ) | ( n7620 & ~n7625 ) ;
  assign n7627 = ( x91 & n7330 ) | ( x91 & ~n7464 ) | ( n7330 & ~n7464 ) ;
  assign n7628 = x91 & n7330 ;
  assign n7629 = ( ~n7335 & n7627 ) | ( ~n7335 & n7628 ) | ( n7627 & n7628 ) ;
  assign n7630 = ( n7335 & n7627 ) | ( n7335 & n7628 ) | ( n7627 & n7628 ) ;
  assign n7631 = ( n7335 & n7629 ) | ( n7335 & ~n7630 ) | ( n7629 & ~n7630 ) ;
  assign n7632 = ( x92 & n7626 ) | ( x92 & ~n7631 ) | ( n7626 & ~n7631 ) ;
  assign n7633 = ( x92 & n7336 ) | ( x92 & ~n7464 ) | ( n7336 & ~n7464 ) ;
  assign n7634 = x92 & n7336 ;
  assign n7635 = ( n7341 & n7633 ) | ( n7341 & n7634 ) | ( n7633 & n7634 ) ;
  assign n7636 = ( ~n7341 & n7633 ) | ( ~n7341 & n7634 ) | ( n7633 & n7634 ) ;
  assign n7637 = ( n7341 & ~n7635 ) | ( n7341 & n7636 ) | ( ~n7635 & n7636 ) ;
  assign n7638 = ( x93 & n7632 ) | ( x93 & ~n7637 ) | ( n7632 & ~n7637 ) ;
  assign n7639 = ( x93 & n7342 ) | ( x93 & ~n7464 ) | ( n7342 & ~n7464 ) ;
  assign n7640 = x93 & n7342 ;
  assign n7641 = ( ~n7347 & n7639 ) | ( ~n7347 & n7640 ) | ( n7639 & n7640 ) ;
  assign n7642 = ( n7347 & n7639 ) | ( n7347 & n7640 ) | ( n7639 & n7640 ) ;
  assign n7643 = ( n7347 & n7641 ) | ( n7347 & ~n7642 ) | ( n7641 & ~n7642 ) ;
  assign n7644 = ( x94 & n7638 ) | ( x94 & ~n7643 ) | ( n7638 & ~n7643 ) ;
  assign n7645 = ( x94 & n7348 ) | ( x94 & ~n7464 ) | ( n7348 & ~n7464 ) ;
  assign n7646 = x94 & n7348 ;
  assign n7647 = ( n7353 & n7645 ) | ( n7353 & n7646 ) | ( n7645 & n7646 ) ;
  assign n7648 = ( ~n7353 & n7645 ) | ( ~n7353 & n7646 ) | ( n7645 & n7646 ) ;
  assign n7649 = ( n7353 & ~n7647 ) | ( n7353 & n7648 ) | ( ~n7647 & n7648 ) ;
  assign n7650 = ( x95 & n7644 ) | ( x95 & ~n7649 ) | ( n7644 & ~n7649 ) ;
  assign n7651 = ( x95 & n7354 ) | ( x95 & ~n7464 ) | ( n7354 & ~n7464 ) ;
  assign n7652 = x95 & n7354 ;
  assign n7653 = ( ~n7359 & n7651 ) | ( ~n7359 & n7652 ) | ( n7651 & n7652 ) ;
  assign n7654 = ( n7359 & n7651 ) | ( n7359 & n7652 ) | ( n7651 & n7652 ) ;
  assign n7655 = ( n7359 & n7653 ) | ( n7359 & ~n7654 ) | ( n7653 & ~n7654 ) ;
  assign n7656 = ( x96 & n7650 ) | ( x96 & ~n7655 ) | ( n7650 & ~n7655 ) ;
  assign n7657 = ( x96 & n7360 ) | ( x96 & ~n7464 ) | ( n7360 & ~n7464 ) ;
  assign n7658 = x96 & n7360 ;
  assign n7659 = ( n7365 & n7657 ) | ( n7365 & n7658 ) | ( n7657 & n7658 ) ;
  assign n7660 = ( ~n7365 & n7657 ) | ( ~n7365 & n7658 ) | ( n7657 & n7658 ) ;
  assign n7661 = ( n7365 & ~n7659 ) | ( n7365 & n7660 ) | ( ~n7659 & n7660 ) ;
  assign n7662 = ( x97 & n7656 ) | ( x97 & ~n7661 ) | ( n7656 & ~n7661 ) ;
  assign n7663 = ( x97 & n7366 ) | ( x97 & ~n7464 ) | ( n7366 & ~n7464 ) ;
  assign n7664 = x97 & n7366 ;
  assign n7665 = ( ~n7371 & n7663 ) | ( ~n7371 & n7664 ) | ( n7663 & n7664 ) ;
  assign n7666 = ( n7371 & n7663 ) | ( n7371 & n7664 ) | ( n7663 & n7664 ) ;
  assign n7667 = ( n7371 & n7665 ) | ( n7371 & ~n7666 ) | ( n7665 & ~n7666 ) ;
  assign n7668 = ( x98 & n7662 ) | ( x98 & ~n7667 ) | ( n7662 & ~n7667 ) ;
  assign n7669 = ( x98 & n7372 ) | ( x98 & ~n7464 ) | ( n7372 & ~n7464 ) ;
  assign n7670 = x98 & n7372 ;
  assign n7671 = ( n7377 & n7669 ) | ( n7377 & n7670 ) | ( n7669 & n7670 ) ;
  assign n7672 = ( ~n7377 & n7669 ) | ( ~n7377 & n7670 ) | ( n7669 & n7670 ) ;
  assign n7673 = ( n7377 & ~n7671 ) | ( n7377 & n7672 ) | ( ~n7671 & n7672 ) ;
  assign n7674 = ( x99 & n7668 ) | ( x99 & ~n7673 ) | ( n7668 & ~n7673 ) ;
  assign n7675 = ( x99 & n7378 ) | ( x99 & ~n7464 ) | ( n7378 & ~n7464 ) ;
  assign n7676 = x99 & n7378 ;
  assign n7677 = ( ~n7383 & n7675 ) | ( ~n7383 & n7676 ) | ( n7675 & n7676 ) ;
  assign n7678 = ( n7383 & n7675 ) | ( n7383 & n7676 ) | ( n7675 & n7676 ) ;
  assign n7679 = ( n7383 & n7677 ) | ( n7383 & ~n7678 ) | ( n7677 & ~n7678 ) ;
  assign n7680 = ( x100 & n7674 ) | ( x100 & ~n7679 ) | ( n7674 & ~n7679 ) ;
  assign n7681 = ( x100 & n7384 ) | ( x100 & ~n7464 ) | ( n7384 & ~n7464 ) ;
  assign n7682 = x100 & n7384 ;
  assign n7683 = ( n7389 & n7681 ) | ( n7389 & n7682 ) | ( n7681 & n7682 ) ;
  assign n7684 = ( ~n7389 & n7681 ) | ( ~n7389 & n7682 ) | ( n7681 & n7682 ) ;
  assign n7685 = ( n7389 & ~n7683 ) | ( n7389 & n7684 ) | ( ~n7683 & n7684 ) ;
  assign n7686 = ( x101 & n7680 ) | ( x101 & ~n7685 ) | ( n7680 & ~n7685 ) ;
  assign n7687 = ( x101 & n7390 ) | ( x101 & ~n7464 ) | ( n7390 & ~n7464 ) ;
  assign n7688 = x101 & n7390 ;
  assign n7689 = ( ~n7395 & n7687 ) | ( ~n7395 & n7688 ) | ( n7687 & n7688 ) ;
  assign n7690 = ( n7395 & n7687 ) | ( n7395 & n7688 ) | ( n7687 & n7688 ) ;
  assign n7691 = ( n7395 & n7689 ) | ( n7395 & ~n7690 ) | ( n7689 & ~n7690 ) ;
  assign n7692 = ( x102 & n7686 ) | ( x102 & ~n7691 ) | ( n7686 & ~n7691 ) ;
  assign n7693 = ( x102 & n7396 ) | ( x102 & ~n7464 ) | ( n7396 & ~n7464 ) ;
  assign n7694 = x102 & n7396 ;
  assign n7695 = ( n7401 & n7693 ) | ( n7401 & n7694 ) | ( n7693 & n7694 ) ;
  assign n7696 = ( ~n7401 & n7693 ) | ( ~n7401 & n7694 ) | ( n7693 & n7694 ) ;
  assign n7697 = ( n7401 & ~n7695 ) | ( n7401 & n7696 ) | ( ~n7695 & n7696 ) ;
  assign n7698 = ( x103 & n7692 ) | ( x103 & ~n7697 ) | ( n7692 & ~n7697 ) ;
  assign n7699 = ( x103 & n7402 ) | ( x103 & ~n7464 ) | ( n7402 & ~n7464 ) ;
  assign n7700 = x103 & n7402 ;
  assign n7701 = ( ~n7407 & n7699 ) | ( ~n7407 & n7700 ) | ( n7699 & n7700 ) ;
  assign n7702 = ( n7407 & n7699 ) | ( n7407 & n7700 ) | ( n7699 & n7700 ) ;
  assign n7703 = ( n7407 & n7701 ) | ( n7407 & ~n7702 ) | ( n7701 & ~n7702 ) ;
  assign n7704 = ( x104 & n7698 ) | ( x104 & ~n7703 ) | ( n7698 & ~n7703 ) ;
  assign n7705 = ( x104 & n7408 ) | ( x104 & ~n7464 ) | ( n7408 & ~n7464 ) ;
  assign n7706 = x104 & n7408 ;
  assign n7707 = ( n7413 & n7705 ) | ( n7413 & n7706 ) | ( n7705 & n7706 ) ;
  assign n7708 = ( ~n7413 & n7705 ) | ( ~n7413 & n7706 ) | ( n7705 & n7706 ) ;
  assign n7709 = ( n7413 & ~n7707 ) | ( n7413 & n7708 ) | ( ~n7707 & n7708 ) ;
  assign n7710 = ( x105 & n7704 ) | ( x105 & ~n7709 ) | ( n7704 & ~n7709 ) ;
  assign n7711 = ( x105 & n7414 ) | ( x105 & ~n7464 ) | ( n7414 & ~n7464 ) ;
  assign n7712 = x105 & n7414 ;
  assign n7713 = ( ~n7419 & n7711 ) | ( ~n7419 & n7712 ) | ( n7711 & n7712 ) ;
  assign n7714 = ( n7419 & n7711 ) | ( n7419 & n7712 ) | ( n7711 & n7712 ) ;
  assign n7715 = ( n7419 & n7713 ) | ( n7419 & ~n7714 ) | ( n7713 & ~n7714 ) ;
  assign n7716 = ( x106 & n7710 ) | ( x106 & ~n7715 ) | ( n7710 & ~n7715 ) ;
  assign n7717 = ( x106 & n7420 ) | ( x106 & ~n7464 ) | ( n7420 & ~n7464 ) ;
  assign n7718 = x106 & n7420 ;
  assign n7719 = ( n7425 & n7717 ) | ( n7425 & n7718 ) | ( n7717 & n7718 ) ;
  assign n7720 = ( ~n7425 & n7717 ) | ( ~n7425 & n7718 ) | ( n7717 & n7718 ) ;
  assign n7721 = ( n7425 & ~n7719 ) | ( n7425 & n7720 ) | ( ~n7719 & n7720 ) ;
  assign n7722 = ( x107 & n7716 ) | ( x107 & ~n7721 ) | ( n7716 & ~n7721 ) ;
  assign n7723 = ( x107 & n7426 ) | ( x107 & ~n7464 ) | ( n7426 & ~n7464 ) ;
  assign n7724 = x107 & n7426 ;
  assign n7725 = ( ~n7431 & n7723 ) | ( ~n7431 & n7724 ) | ( n7723 & n7724 ) ;
  assign n7726 = ( n7431 & n7723 ) | ( n7431 & n7724 ) | ( n7723 & n7724 ) ;
  assign n7727 = ( n7431 & n7725 ) | ( n7431 & ~n7726 ) | ( n7725 & ~n7726 ) ;
  assign n7728 = ( x108 & n7722 ) | ( x108 & ~n7727 ) | ( n7722 & ~n7727 ) ;
  assign n7729 = ( x108 & n7432 ) | ( x108 & ~n7464 ) | ( n7432 & ~n7464 ) ;
  assign n7730 = x108 & n7432 ;
  assign n7731 = ( n7437 & n7729 ) | ( n7437 & n7730 ) | ( n7729 & n7730 ) ;
  assign n7732 = ( ~n7437 & n7729 ) | ( ~n7437 & n7730 ) | ( n7729 & n7730 ) ;
  assign n7733 = ( n7437 & ~n7731 ) | ( n7437 & n7732 ) | ( ~n7731 & n7732 ) ;
  assign n7734 = ( x109 & n7728 ) | ( x109 & ~n7733 ) | ( n7728 & ~n7733 ) ;
  assign n7735 = ( x109 & n7438 ) | ( x109 & ~n7464 ) | ( n7438 & ~n7464 ) ;
  assign n7736 = x109 & n7438 ;
  assign n7737 = ( ~n7443 & n7735 ) | ( ~n7443 & n7736 ) | ( n7735 & n7736 ) ;
  assign n7738 = ( n7443 & n7735 ) | ( n7443 & n7736 ) | ( n7735 & n7736 ) ;
  assign n7739 = ( n7443 & n7737 ) | ( n7443 & ~n7738 ) | ( n7737 & ~n7738 ) ;
  assign n7740 = ( x110 & n7734 ) | ( x110 & ~n7739 ) | ( n7734 & ~n7739 ) ;
  assign n7741 = ( x110 & n7444 ) | ( x110 & ~n7464 ) | ( n7444 & ~n7464 ) ;
  assign n7742 = x110 & n7444 ;
  assign n7743 = ( n7449 & n7741 ) | ( n7449 & n7742 ) | ( n7741 & n7742 ) ;
  assign n7744 = ( ~n7449 & n7741 ) | ( ~n7449 & n7742 ) | ( n7741 & n7742 ) ;
  assign n7745 = ( n7449 & ~n7743 ) | ( n7449 & n7744 ) | ( ~n7743 & n7744 ) ;
  assign n7746 = ( x111 & n7740 ) | ( x111 & ~n7745 ) | ( n7740 & ~n7745 ) ;
  assign n7747 = ( x111 & n7450 ) | ( x111 & ~n7464 ) | ( n7450 & ~n7464 ) ;
  assign n7748 = x111 & n7450 ;
  assign n7749 = ( ~n7455 & n7747 ) | ( ~n7455 & n7748 ) | ( n7747 & n7748 ) ;
  assign n7750 = ( n7455 & n7747 ) | ( n7455 & n7748 ) | ( n7747 & n7748 ) ;
  assign n7751 = ( n7455 & n7749 ) | ( n7455 & ~n7750 ) | ( n7749 & ~n7750 ) ;
  assign n7752 = ( x112 & n7746 ) | ( x112 & ~n7751 ) | ( n7746 & ~n7751 ) ;
  assign n7753 = ( x112 & n7456 ) | ( x112 & ~n7464 ) | ( n7456 & ~n7464 ) ;
  assign n7754 = x112 & n7456 ;
  assign n7755 = ( ~n7461 & n7753 ) | ( ~n7461 & n7754 ) | ( n7753 & n7754 ) ;
  assign n7756 = ( n7461 & n7753 ) | ( n7461 & n7754 ) | ( n7753 & n7754 ) ;
  assign n7757 = ( n7461 & n7755 ) | ( n7461 & ~n7756 ) | ( n7755 & ~n7756 ) ;
  assign n7758 = ( x113 & n7752 ) | ( x113 & ~n7757 ) | ( n7752 & ~n7757 ) ;
  assign n7759 = x114 | n7758 ;
  assign n7760 = ( x114 & n143 ) | ( x114 & n7758 ) | ( n143 & n7758 ) ;
  assign n7761 = ( n7465 & ~n7759 ) | ( n7465 & n7760 ) | ( ~n7759 & n7760 ) ;
  assign n7762 = ( x114 & ~n7465 ) | ( x114 & n7758 ) | ( ~n7465 & n7758 ) ;
  assign n7763 = n143 | n7762 ;
  assign n7764 = ( x13 & ~x64 ) | ( x13 & n7763 ) | ( ~x64 & n7763 ) ;
  assign n7765 = ~x13 & n7763 ;
  assign n7766 = ( n7469 & n7764 ) | ( n7469 & ~n7765 ) | ( n7764 & ~n7765 ) ;
  assign n7767 = ~x12 & x64 ;
  assign n7768 = ( x65 & ~n7766 ) | ( x65 & n7767 ) | ( ~n7766 & n7767 ) ;
  assign n7769 = ( x65 & n7469 ) | ( x65 & ~n7763 ) | ( n7469 & ~n7763 ) ;
  assign n7770 = x65 & n7469 ;
  assign n7771 = ( n7468 & n7769 ) | ( n7468 & n7770 ) | ( n7769 & n7770 ) ;
  assign n7772 = ( ~n7468 & n7769 ) | ( ~n7468 & n7770 ) | ( n7769 & n7770 ) ;
  assign n7773 = ( n7468 & ~n7771 ) | ( n7468 & n7772 ) | ( ~n7771 & n7772 ) ;
  assign n7774 = ( x66 & n7768 ) | ( x66 & ~n7773 ) | ( n7768 & ~n7773 ) ;
  assign n7775 = ( x66 & n7470 ) | ( x66 & ~n7763 ) | ( n7470 & ~n7763 ) ;
  assign n7776 = x66 & n7470 ;
  assign n7777 = ( n7475 & n7775 ) | ( n7475 & n7776 ) | ( n7775 & n7776 ) ;
  assign n7778 = ( ~n7475 & n7775 ) | ( ~n7475 & n7776 ) | ( n7775 & n7776 ) ;
  assign n7779 = ( n7475 & ~n7777 ) | ( n7475 & n7778 ) | ( ~n7777 & n7778 ) ;
  assign n7780 = ( x67 & n7774 ) | ( x67 & ~n7779 ) | ( n7774 & ~n7779 ) ;
  assign n7781 = ( x67 & n7476 ) | ( x67 & ~n7763 ) | ( n7476 & ~n7763 ) ;
  assign n7782 = x67 & n7476 ;
  assign n7783 = ( ~n7481 & n7781 ) | ( ~n7481 & n7782 ) | ( n7781 & n7782 ) ;
  assign n7784 = ( n7481 & n7781 ) | ( n7481 & n7782 ) | ( n7781 & n7782 ) ;
  assign n7785 = ( n7481 & n7783 ) | ( n7481 & ~n7784 ) | ( n7783 & ~n7784 ) ;
  assign n7786 = ( x68 & n7780 ) | ( x68 & ~n7785 ) | ( n7780 & ~n7785 ) ;
  assign n7787 = ( x68 & n7482 ) | ( x68 & ~n7763 ) | ( n7482 & ~n7763 ) ;
  assign n7788 = x68 & n7482 ;
  assign n7789 = ( n7487 & n7787 ) | ( n7487 & n7788 ) | ( n7787 & n7788 ) ;
  assign n7790 = ( ~n7487 & n7787 ) | ( ~n7487 & n7788 ) | ( n7787 & n7788 ) ;
  assign n7791 = ( n7487 & ~n7789 ) | ( n7487 & n7790 ) | ( ~n7789 & n7790 ) ;
  assign n7792 = ( x69 & n7786 ) | ( x69 & ~n7791 ) | ( n7786 & ~n7791 ) ;
  assign n7793 = ( x69 & n7488 ) | ( x69 & ~n7763 ) | ( n7488 & ~n7763 ) ;
  assign n7794 = x69 & n7488 ;
  assign n7795 = ( ~n7493 & n7793 ) | ( ~n7493 & n7794 ) | ( n7793 & n7794 ) ;
  assign n7796 = ( n7493 & n7793 ) | ( n7493 & n7794 ) | ( n7793 & n7794 ) ;
  assign n7797 = ( n7493 & n7795 ) | ( n7493 & ~n7796 ) | ( n7795 & ~n7796 ) ;
  assign n7798 = ( x70 & n7792 ) | ( x70 & ~n7797 ) | ( n7792 & ~n7797 ) ;
  assign n7799 = ( x70 & n7494 ) | ( x70 & ~n7763 ) | ( n7494 & ~n7763 ) ;
  assign n7800 = x70 & n7494 ;
  assign n7801 = ( n7499 & n7799 ) | ( n7499 & n7800 ) | ( n7799 & n7800 ) ;
  assign n7802 = ( ~n7499 & n7799 ) | ( ~n7499 & n7800 ) | ( n7799 & n7800 ) ;
  assign n7803 = ( n7499 & ~n7801 ) | ( n7499 & n7802 ) | ( ~n7801 & n7802 ) ;
  assign n7804 = ( x71 & n7798 ) | ( x71 & ~n7803 ) | ( n7798 & ~n7803 ) ;
  assign n7805 = ( x71 & n7500 ) | ( x71 & ~n7763 ) | ( n7500 & ~n7763 ) ;
  assign n7806 = x71 & n7500 ;
  assign n7807 = ( ~n7505 & n7805 ) | ( ~n7505 & n7806 ) | ( n7805 & n7806 ) ;
  assign n7808 = ( n7505 & n7805 ) | ( n7505 & n7806 ) | ( n7805 & n7806 ) ;
  assign n7809 = ( n7505 & n7807 ) | ( n7505 & ~n7808 ) | ( n7807 & ~n7808 ) ;
  assign n7810 = ( x72 & n7804 ) | ( x72 & ~n7809 ) | ( n7804 & ~n7809 ) ;
  assign n7811 = ( x72 & n7506 ) | ( x72 & ~n7763 ) | ( n7506 & ~n7763 ) ;
  assign n7812 = x72 & n7506 ;
  assign n7813 = ( n7511 & n7811 ) | ( n7511 & n7812 ) | ( n7811 & n7812 ) ;
  assign n7814 = ( ~n7511 & n7811 ) | ( ~n7511 & n7812 ) | ( n7811 & n7812 ) ;
  assign n7815 = ( n7511 & ~n7813 ) | ( n7511 & n7814 ) | ( ~n7813 & n7814 ) ;
  assign n7816 = ( x73 & n7810 ) | ( x73 & ~n7815 ) | ( n7810 & ~n7815 ) ;
  assign n7817 = ( x73 & n7512 ) | ( x73 & ~n7763 ) | ( n7512 & ~n7763 ) ;
  assign n7818 = x73 & n7512 ;
  assign n7819 = ( ~n7517 & n7817 ) | ( ~n7517 & n7818 ) | ( n7817 & n7818 ) ;
  assign n7820 = ( n7517 & n7817 ) | ( n7517 & n7818 ) | ( n7817 & n7818 ) ;
  assign n7821 = ( n7517 & n7819 ) | ( n7517 & ~n7820 ) | ( n7819 & ~n7820 ) ;
  assign n7822 = ( x74 & n7816 ) | ( x74 & ~n7821 ) | ( n7816 & ~n7821 ) ;
  assign n7823 = ( x74 & n7518 ) | ( x74 & ~n7763 ) | ( n7518 & ~n7763 ) ;
  assign n7824 = x74 & n7518 ;
  assign n7825 = ( n7523 & n7823 ) | ( n7523 & n7824 ) | ( n7823 & n7824 ) ;
  assign n7826 = ( ~n7523 & n7823 ) | ( ~n7523 & n7824 ) | ( n7823 & n7824 ) ;
  assign n7827 = ( n7523 & ~n7825 ) | ( n7523 & n7826 ) | ( ~n7825 & n7826 ) ;
  assign n7828 = ( x75 & n7822 ) | ( x75 & ~n7827 ) | ( n7822 & ~n7827 ) ;
  assign n7829 = ( x75 & n7524 ) | ( x75 & ~n7763 ) | ( n7524 & ~n7763 ) ;
  assign n7830 = x75 & n7524 ;
  assign n7831 = ( ~n7529 & n7829 ) | ( ~n7529 & n7830 ) | ( n7829 & n7830 ) ;
  assign n7832 = ( n7529 & n7829 ) | ( n7529 & n7830 ) | ( n7829 & n7830 ) ;
  assign n7833 = ( n7529 & n7831 ) | ( n7529 & ~n7832 ) | ( n7831 & ~n7832 ) ;
  assign n7834 = ( x76 & n7828 ) | ( x76 & ~n7833 ) | ( n7828 & ~n7833 ) ;
  assign n7835 = ( x76 & n7530 ) | ( x76 & ~n7763 ) | ( n7530 & ~n7763 ) ;
  assign n7836 = x76 & n7530 ;
  assign n7837 = ( n7535 & n7835 ) | ( n7535 & n7836 ) | ( n7835 & n7836 ) ;
  assign n7838 = ( ~n7535 & n7835 ) | ( ~n7535 & n7836 ) | ( n7835 & n7836 ) ;
  assign n7839 = ( n7535 & ~n7837 ) | ( n7535 & n7838 ) | ( ~n7837 & n7838 ) ;
  assign n7840 = ( x77 & n7834 ) | ( x77 & ~n7839 ) | ( n7834 & ~n7839 ) ;
  assign n7841 = ( x77 & n7536 ) | ( x77 & ~n7763 ) | ( n7536 & ~n7763 ) ;
  assign n7842 = x77 & n7536 ;
  assign n7843 = ( ~n7541 & n7841 ) | ( ~n7541 & n7842 ) | ( n7841 & n7842 ) ;
  assign n7844 = ( n7541 & n7841 ) | ( n7541 & n7842 ) | ( n7841 & n7842 ) ;
  assign n7845 = ( n7541 & n7843 ) | ( n7541 & ~n7844 ) | ( n7843 & ~n7844 ) ;
  assign n7846 = ( x78 & n7840 ) | ( x78 & ~n7845 ) | ( n7840 & ~n7845 ) ;
  assign n7847 = ( x78 & n7542 ) | ( x78 & ~n7763 ) | ( n7542 & ~n7763 ) ;
  assign n7848 = x78 & n7542 ;
  assign n7849 = ( n7547 & n7847 ) | ( n7547 & n7848 ) | ( n7847 & n7848 ) ;
  assign n7850 = ( ~n7547 & n7847 ) | ( ~n7547 & n7848 ) | ( n7847 & n7848 ) ;
  assign n7851 = ( n7547 & ~n7849 ) | ( n7547 & n7850 ) | ( ~n7849 & n7850 ) ;
  assign n7852 = ( x79 & n7846 ) | ( x79 & ~n7851 ) | ( n7846 & ~n7851 ) ;
  assign n7853 = ( x79 & n7548 ) | ( x79 & ~n7763 ) | ( n7548 & ~n7763 ) ;
  assign n7854 = x79 & n7548 ;
  assign n7855 = ( ~n7553 & n7853 ) | ( ~n7553 & n7854 ) | ( n7853 & n7854 ) ;
  assign n7856 = ( n7553 & n7853 ) | ( n7553 & n7854 ) | ( n7853 & n7854 ) ;
  assign n7857 = ( n7553 & n7855 ) | ( n7553 & ~n7856 ) | ( n7855 & ~n7856 ) ;
  assign n7858 = ( x80 & n7852 ) | ( x80 & ~n7857 ) | ( n7852 & ~n7857 ) ;
  assign n7859 = ( x80 & n7554 ) | ( x80 & ~n7763 ) | ( n7554 & ~n7763 ) ;
  assign n7860 = x80 & n7554 ;
  assign n7861 = ( n7559 & n7859 ) | ( n7559 & n7860 ) | ( n7859 & n7860 ) ;
  assign n7862 = ( ~n7559 & n7859 ) | ( ~n7559 & n7860 ) | ( n7859 & n7860 ) ;
  assign n7863 = ( n7559 & ~n7861 ) | ( n7559 & n7862 ) | ( ~n7861 & n7862 ) ;
  assign n7864 = ( x81 & n7858 ) | ( x81 & ~n7863 ) | ( n7858 & ~n7863 ) ;
  assign n7865 = ( x81 & n7560 ) | ( x81 & ~n7763 ) | ( n7560 & ~n7763 ) ;
  assign n7866 = x81 & n7560 ;
  assign n7867 = ( ~n7565 & n7865 ) | ( ~n7565 & n7866 ) | ( n7865 & n7866 ) ;
  assign n7868 = ( n7565 & n7865 ) | ( n7565 & n7866 ) | ( n7865 & n7866 ) ;
  assign n7869 = ( n7565 & n7867 ) | ( n7565 & ~n7868 ) | ( n7867 & ~n7868 ) ;
  assign n7870 = ( x82 & n7864 ) | ( x82 & ~n7869 ) | ( n7864 & ~n7869 ) ;
  assign n7871 = ( x82 & n7566 ) | ( x82 & ~n7763 ) | ( n7566 & ~n7763 ) ;
  assign n7872 = x82 & n7566 ;
  assign n7873 = ( n7571 & n7871 ) | ( n7571 & n7872 ) | ( n7871 & n7872 ) ;
  assign n7874 = ( ~n7571 & n7871 ) | ( ~n7571 & n7872 ) | ( n7871 & n7872 ) ;
  assign n7875 = ( n7571 & ~n7873 ) | ( n7571 & n7874 ) | ( ~n7873 & n7874 ) ;
  assign n7876 = ( x83 & n7870 ) | ( x83 & ~n7875 ) | ( n7870 & ~n7875 ) ;
  assign n7877 = ( x83 & n7572 ) | ( x83 & ~n7763 ) | ( n7572 & ~n7763 ) ;
  assign n7878 = x83 & n7572 ;
  assign n7879 = ( ~n7577 & n7877 ) | ( ~n7577 & n7878 ) | ( n7877 & n7878 ) ;
  assign n7880 = ( n7577 & n7877 ) | ( n7577 & n7878 ) | ( n7877 & n7878 ) ;
  assign n7881 = ( n7577 & n7879 ) | ( n7577 & ~n7880 ) | ( n7879 & ~n7880 ) ;
  assign n7882 = ( x84 & n7876 ) | ( x84 & ~n7881 ) | ( n7876 & ~n7881 ) ;
  assign n7883 = ( x84 & n7578 ) | ( x84 & ~n7763 ) | ( n7578 & ~n7763 ) ;
  assign n7884 = x84 & n7578 ;
  assign n7885 = ( n7583 & n7883 ) | ( n7583 & n7884 ) | ( n7883 & n7884 ) ;
  assign n7886 = ( ~n7583 & n7883 ) | ( ~n7583 & n7884 ) | ( n7883 & n7884 ) ;
  assign n7887 = ( n7583 & ~n7885 ) | ( n7583 & n7886 ) | ( ~n7885 & n7886 ) ;
  assign n7888 = ( x85 & n7882 ) | ( x85 & ~n7887 ) | ( n7882 & ~n7887 ) ;
  assign n7889 = ( x85 & n7584 ) | ( x85 & ~n7763 ) | ( n7584 & ~n7763 ) ;
  assign n7890 = x85 & n7584 ;
  assign n7891 = ( ~n7589 & n7889 ) | ( ~n7589 & n7890 ) | ( n7889 & n7890 ) ;
  assign n7892 = ( n7589 & n7889 ) | ( n7589 & n7890 ) | ( n7889 & n7890 ) ;
  assign n7893 = ( n7589 & n7891 ) | ( n7589 & ~n7892 ) | ( n7891 & ~n7892 ) ;
  assign n7894 = ( x86 & n7888 ) | ( x86 & ~n7893 ) | ( n7888 & ~n7893 ) ;
  assign n7895 = ( x86 & n7590 ) | ( x86 & ~n7763 ) | ( n7590 & ~n7763 ) ;
  assign n7896 = x86 & n7590 ;
  assign n7897 = ( n7595 & n7895 ) | ( n7595 & n7896 ) | ( n7895 & n7896 ) ;
  assign n7898 = ( ~n7595 & n7895 ) | ( ~n7595 & n7896 ) | ( n7895 & n7896 ) ;
  assign n7899 = ( n7595 & ~n7897 ) | ( n7595 & n7898 ) | ( ~n7897 & n7898 ) ;
  assign n7900 = ( x87 & n7894 ) | ( x87 & ~n7899 ) | ( n7894 & ~n7899 ) ;
  assign n7901 = ( x87 & n7596 ) | ( x87 & ~n7763 ) | ( n7596 & ~n7763 ) ;
  assign n7902 = x87 & n7596 ;
  assign n7903 = ( ~n7601 & n7901 ) | ( ~n7601 & n7902 ) | ( n7901 & n7902 ) ;
  assign n7904 = ( n7601 & n7901 ) | ( n7601 & n7902 ) | ( n7901 & n7902 ) ;
  assign n7905 = ( n7601 & n7903 ) | ( n7601 & ~n7904 ) | ( n7903 & ~n7904 ) ;
  assign n7906 = ( x88 & n7900 ) | ( x88 & ~n7905 ) | ( n7900 & ~n7905 ) ;
  assign n7907 = ( x88 & n7602 ) | ( x88 & ~n7763 ) | ( n7602 & ~n7763 ) ;
  assign n7908 = x88 & n7602 ;
  assign n7909 = ( n7607 & n7907 ) | ( n7607 & n7908 ) | ( n7907 & n7908 ) ;
  assign n7910 = ( ~n7607 & n7907 ) | ( ~n7607 & n7908 ) | ( n7907 & n7908 ) ;
  assign n7911 = ( n7607 & ~n7909 ) | ( n7607 & n7910 ) | ( ~n7909 & n7910 ) ;
  assign n7912 = ( x89 & n7906 ) | ( x89 & ~n7911 ) | ( n7906 & ~n7911 ) ;
  assign n7913 = ( x89 & n7608 ) | ( x89 & ~n7763 ) | ( n7608 & ~n7763 ) ;
  assign n7914 = x89 & n7608 ;
  assign n7915 = ( ~n7613 & n7913 ) | ( ~n7613 & n7914 ) | ( n7913 & n7914 ) ;
  assign n7916 = ( n7613 & n7913 ) | ( n7613 & n7914 ) | ( n7913 & n7914 ) ;
  assign n7917 = ( n7613 & n7915 ) | ( n7613 & ~n7916 ) | ( n7915 & ~n7916 ) ;
  assign n7918 = ( x90 & n7912 ) | ( x90 & ~n7917 ) | ( n7912 & ~n7917 ) ;
  assign n7919 = ( x90 & n7614 ) | ( x90 & ~n7763 ) | ( n7614 & ~n7763 ) ;
  assign n7920 = x90 & n7614 ;
  assign n7921 = ( n7619 & n7919 ) | ( n7619 & n7920 ) | ( n7919 & n7920 ) ;
  assign n7922 = ( ~n7619 & n7919 ) | ( ~n7619 & n7920 ) | ( n7919 & n7920 ) ;
  assign n7923 = ( n7619 & ~n7921 ) | ( n7619 & n7922 ) | ( ~n7921 & n7922 ) ;
  assign n7924 = ( x91 & n7918 ) | ( x91 & ~n7923 ) | ( n7918 & ~n7923 ) ;
  assign n7925 = ( x91 & n7620 ) | ( x91 & ~n7763 ) | ( n7620 & ~n7763 ) ;
  assign n7926 = x91 & n7620 ;
  assign n7927 = ( ~n7625 & n7925 ) | ( ~n7625 & n7926 ) | ( n7925 & n7926 ) ;
  assign n7928 = ( n7625 & n7925 ) | ( n7625 & n7926 ) | ( n7925 & n7926 ) ;
  assign n7929 = ( n7625 & n7927 ) | ( n7625 & ~n7928 ) | ( n7927 & ~n7928 ) ;
  assign n7930 = ( x92 & n7924 ) | ( x92 & ~n7929 ) | ( n7924 & ~n7929 ) ;
  assign n7931 = ( x92 & n7626 ) | ( x92 & ~n7763 ) | ( n7626 & ~n7763 ) ;
  assign n7932 = x92 & n7626 ;
  assign n7933 = ( n7631 & n7931 ) | ( n7631 & n7932 ) | ( n7931 & n7932 ) ;
  assign n7934 = ( ~n7631 & n7931 ) | ( ~n7631 & n7932 ) | ( n7931 & n7932 ) ;
  assign n7935 = ( n7631 & ~n7933 ) | ( n7631 & n7934 ) | ( ~n7933 & n7934 ) ;
  assign n7936 = ( x93 & n7930 ) | ( x93 & ~n7935 ) | ( n7930 & ~n7935 ) ;
  assign n7937 = ( x93 & n7632 ) | ( x93 & ~n7763 ) | ( n7632 & ~n7763 ) ;
  assign n7938 = x93 & n7632 ;
  assign n7939 = ( ~n7637 & n7937 ) | ( ~n7637 & n7938 ) | ( n7937 & n7938 ) ;
  assign n7940 = ( n7637 & n7937 ) | ( n7637 & n7938 ) | ( n7937 & n7938 ) ;
  assign n7941 = ( n7637 & n7939 ) | ( n7637 & ~n7940 ) | ( n7939 & ~n7940 ) ;
  assign n7942 = ( x94 & n7936 ) | ( x94 & ~n7941 ) | ( n7936 & ~n7941 ) ;
  assign n7943 = ( x94 & n7638 ) | ( x94 & ~n7763 ) | ( n7638 & ~n7763 ) ;
  assign n7944 = x94 & n7638 ;
  assign n7945 = ( n7643 & n7943 ) | ( n7643 & n7944 ) | ( n7943 & n7944 ) ;
  assign n7946 = ( ~n7643 & n7943 ) | ( ~n7643 & n7944 ) | ( n7943 & n7944 ) ;
  assign n7947 = ( n7643 & ~n7945 ) | ( n7643 & n7946 ) | ( ~n7945 & n7946 ) ;
  assign n7948 = ( x95 & n7942 ) | ( x95 & ~n7947 ) | ( n7942 & ~n7947 ) ;
  assign n7949 = ( x95 & n7644 ) | ( x95 & ~n7763 ) | ( n7644 & ~n7763 ) ;
  assign n7950 = x95 & n7644 ;
  assign n7951 = ( ~n7649 & n7949 ) | ( ~n7649 & n7950 ) | ( n7949 & n7950 ) ;
  assign n7952 = ( n7649 & n7949 ) | ( n7649 & n7950 ) | ( n7949 & n7950 ) ;
  assign n7953 = ( n7649 & n7951 ) | ( n7649 & ~n7952 ) | ( n7951 & ~n7952 ) ;
  assign n7954 = ( x96 & n7948 ) | ( x96 & ~n7953 ) | ( n7948 & ~n7953 ) ;
  assign n7955 = ( x96 & n7650 ) | ( x96 & ~n7763 ) | ( n7650 & ~n7763 ) ;
  assign n7956 = x96 & n7650 ;
  assign n7957 = ( n7655 & n7955 ) | ( n7655 & n7956 ) | ( n7955 & n7956 ) ;
  assign n7958 = ( ~n7655 & n7955 ) | ( ~n7655 & n7956 ) | ( n7955 & n7956 ) ;
  assign n7959 = ( n7655 & ~n7957 ) | ( n7655 & n7958 ) | ( ~n7957 & n7958 ) ;
  assign n7960 = ( x97 & n7954 ) | ( x97 & ~n7959 ) | ( n7954 & ~n7959 ) ;
  assign n7961 = ( x97 & n7656 ) | ( x97 & ~n7763 ) | ( n7656 & ~n7763 ) ;
  assign n7962 = x97 & n7656 ;
  assign n7963 = ( ~n7661 & n7961 ) | ( ~n7661 & n7962 ) | ( n7961 & n7962 ) ;
  assign n7964 = ( n7661 & n7961 ) | ( n7661 & n7962 ) | ( n7961 & n7962 ) ;
  assign n7965 = ( n7661 & n7963 ) | ( n7661 & ~n7964 ) | ( n7963 & ~n7964 ) ;
  assign n7966 = ( x98 & n7960 ) | ( x98 & ~n7965 ) | ( n7960 & ~n7965 ) ;
  assign n7967 = ( x98 & n7662 ) | ( x98 & ~n7763 ) | ( n7662 & ~n7763 ) ;
  assign n7968 = x98 & n7662 ;
  assign n7969 = ( n7667 & n7967 ) | ( n7667 & n7968 ) | ( n7967 & n7968 ) ;
  assign n7970 = ( ~n7667 & n7967 ) | ( ~n7667 & n7968 ) | ( n7967 & n7968 ) ;
  assign n7971 = ( n7667 & ~n7969 ) | ( n7667 & n7970 ) | ( ~n7969 & n7970 ) ;
  assign n7972 = ( x99 & n7966 ) | ( x99 & ~n7971 ) | ( n7966 & ~n7971 ) ;
  assign n7973 = ( x99 & n7668 ) | ( x99 & ~n7763 ) | ( n7668 & ~n7763 ) ;
  assign n7974 = x99 & n7668 ;
  assign n7975 = ( ~n7673 & n7973 ) | ( ~n7673 & n7974 ) | ( n7973 & n7974 ) ;
  assign n7976 = ( n7673 & n7973 ) | ( n7673 & n7974 ) | ( n7973 & n7974 ) ;
  assign n7977 = ( n7673 & n7975 ) | ( n7673 & ~n7976 ) | ( n7975 & ~n7976 ) ;
  assign n7978 = ( x100 & n7972 ) | ( x100 & ~n7977 ) | ( n7972 & ~n7977 ) ;
  assign n7979 = ( x100 & n7674 ) | ( x100 & ~n7763 ) | ( n7674 & ~n7763 ) ;
  assign n7980 = x100 & n7674 ;
  assign n7981 = ( n7679 & n7979 ) | ( n7679 & n7980 ) | ( n7979 & n7980 ) ;
  assign n7982 = ( ~n7679 & n7979 ) | ( ~n7679 & n7980 ) | ( n7979 & n7980 ) ;
  assign n7983 = ( n7679 & ~n7981 ) | ( n7679 & n7982 ) | ( ~n7981 & n7982 ) ;
  assign n7984 = ( x101 & n7978 ) | ( x101 & ~n7983 ) | ( n7978 & ~n7983 ) ;
  assign n7985 = ( x101 & n7680 ) | ( x101 & ~n7763 ) | ( n7680 & ~n7763 ) ;
  assign n7986 = x101 & n7680 ;
  assign n7987 = ( ~n7685 & n7985 ) | ( ~n7685 & n7986 ) | ( n7985 & n7986 ) ;
  assign n7988 = ( n7685 & n7985 ) | ( n7685 & n7986 ) | ( n7985 & n7986 ) ;
  assign n7989 = ( n7685 & n7987 ) | ( n7685 & ~n7988 ) | ( n7987 & ~n7988 ) ;
  assign n7990 = ( x102 & n7984 ) | ( x102 & ~n7989 ) | ( n7984 & ~n7989 ) ;
  assign n7991 = ( x102 & n7686 ) | ( x102 & ~n7763 ) | ( n7686 & ~n7763 ) ;
  assign n7992 = x102 & n7686 ;
  assign n7993 = ( n7691 & n7991 ) | ( n7691 & n7992 ) | ( n7991 & n7992 ) ;
  assign n7994 = ( ~n7691 & n7991 ) | ( ~n7691 & n7992 ) | ( n7991 & n7992 ) ;
  assign n7995 = ( n7691 & ~n7993 ) | ( n7691 & n7994 ) | ( ~n7993 & n7994 ) ;
  assign n7996 = ( x103 & n7990 ) | ( x103 & ~n7995 ) | ( n7990 & ~n7995 ) ;
  assign n7997 = ( x103 & n7692 ) | ( x103 & ~n7763 ) | ( n7692 & ~n7763 ) ;
  assign n7998 = x103 & n7692 ;
  assign n7999 = ( ~n7697 & n7997 ) | ( ~n7697 & n7998 ) | ( n7997 & n7998 ) ;
  assign n8000 = ( n7697 & n7997 ) | ( n7697 & n7998 ) | ( n7997 & n7998 ) ;
  assign n8001 = ( n7697 & n7999 ) | ( n7697 & ~n8000 ) | ( n7999 & ~n8000 ) ;
  assign n8002 = ( x104 & n7996 ) | ( x104 & ~n8001 ) | ( n7996 & ~n8001 ) ;
  assign n8003 = ( x104 & n7698 ) | ( x104 & ~n7763 ) | ( n7698 & ~n7763 ) ;
  assign n8004 = x104 & n7698 ;
  assign n8005 = ( n7703 & n8003 ) | ( n7703 & n8004 ) | ( n8003 & n8004 ) ;
  assign n8006 = ( ~n7703 & n8003 ) | ( ~n7703 & n8004 ) | ( n8003 & n8004 ) ;
  assign n8007 = ( n7703 & ~n8005 ) | ( n7703 & n8006 ) | ( ~n8005 & n8006 ) ;
  assign n8008 = ( x105 & n8002 ) | ( x105 & ~n8007 ) | ( n8002 & ~n8007 ) ;
  assign n8009 = ( x105 & n7704 ) | ( x105 & ~n7763 ) | ( n7704 & ~n7763 ) ;
  assign n8010 = x105 & n7704 ;
  assign n8011 = ( ~n7709 & n8009 ) | ( ~n7709 & n8010 ) | ( n8009 & n8010 ) ;
  assign n8012 = ( n7709 & n8009 ) | ( n7709 & n8010 ) | ( n8009 & n8010 ) ;
  assign n8013 = ( n7709 & n8011 ) | ( n7709 & ~n8012 ) | ( n8011 & ~n8012 ) ;
  assign n8014 = ( x106 & n8008 ) | ( x106 & ~n8013 ) | ( n8008 & ~n8013 ) ;
  assign n8015 = ( x106 & n7710 ) | ( x106 & ~n7763 ) | ( n7710 & ~n7763 ) ;
  assign n8016 = x106 & n7710 ;
  assign n8017 = ( n7715 & n8015 ) | ( n7715 & n8016 ) | ( n8015 & n8016 ) ;
  assign n8018 = ( ~n7715 & n8015 ) | ( ~n7715 & n8016 ) | ( n8015 & n8016 ) ;
  assign n8019 = ( n7715 & ~n8017 ) | ( n7715 & n8018 ) | ( ~n8017 & n8018 ) ;
  assign n8020 = ( x107 & n8014 ) | ( x107 & ~n8019 ) | ( n8014 & ~n8019 ) ;
  assign n8021 = ( x107 & n7716 ) | ( x107 & ~n7763 ) | ( n7716 & ~n7763 ) ;
  assign n8022 = x107 & n7716 ;
  assign n8023 = ( ~n7721 & n8021 ) | ( ~n7721 & n8022 ) | ( n8021 & n8022 ) ;
  assign n8024 = ( n7721 & n8021 ) | ( n7721 & n8022 ) | ( n8021 & n8022 ) ;
  assign n8025 = ( n7721 & n8023 ) | ( n7721 & ~n8024 ) | ( n8023 & ~n8024 ) ;
  assign n8026 = ( x108 & n8020 ) | ( x108 & ~n8025 ) | ( n8020 & ~n8025 ) ;
  assign n8027 = ( x108 & n7722 ) | ( x108 & ~n7763 ) | ( n7722 & ~n7763 ) ;
  assign n8028 = x108 & n7722 ;
  assign n8029 = ( n7727 & n8027 ) | ( n7727 & n8028 ) | ( n8027 & n8028 ) ;
  assign n8030 = ( ~n7727 & n8027 ) | ( ~n7727 & n8028 ) | ( n8027 & n8028 ) ;
  assign n8031 = ( n7727 & ~n8029 ) | ( n7727 & n8030 ) | ( ~n8029 & n8030 ) ;
  assign n8032 = ( x109 & n8026 ) | ( x109 & ~n8031 ) | ( n8026 & ~n8031 ) ;
  assign n8033 = ( x109 & n7728 ) | ( x109 & ~n7763 ) | ( n7728 & ~n7763 ) ;
  assign n8034 = x109 & n7728 ;
  assign n8035 = ( ~n7733 & n8033 ) | ( ~n7733 & n8034 ) | ( n8033 & n8034 ) ;
  assign n8036 = ( n7733 & n8033 ) | ( n7733 & n8034 ) | ( n8033 & n8034 ) ;
  assign n8037 = ( n7733 & n8035 ) | ( n7733 & ~n8036 ) | ( n8035 & ~n8036 ) ;
  assign n8038 = ( x110 & n8032 ) | ( x110 & ~n8037 ) | ( n8032 & ~n8037 ) ;
  assign n8039 = ( x110 & n7734 ) | ( x110 & ~n7763 ) | ( n7734 & ~n7763 ) ;
  assign n8040 = x110 & n7734 ;
  assign n8041 = ( n7739 & n8039 ) | ( n7739 & n8040 ) | ( n8039 & n8040 ) ;
  assign n8042 = ( ~n7739 & n8039 ) | ( ~n7739 & n8040 ) | ( n8039 & n8040 ) ;
  assign n8043 = ( n7739 & ~n8041 ) | ( n7739 & n8042 ) | ( ~n8041 & n8042 ) ;
  assign n8044 = ( x111 & n8038 ) | ( x111 & ~n8043 ) | ( n8038 & ~n8043 ) ;
  assign n8045 = ( x111 & n7740 ) | ( x111 & ~n7763 ) | ( n7740 & ~n7763 ) ;
  assign n8046 = x111 & n7740 ;
  assign n8047 = ( ~n7745 & n8045 ) | ( ~n7745 & n8046 ) | ( n8045 & n8046 ) ;
  assign n8048 = ( n7745 & n8045 ) | ( n7745 & n8046 ) | ( n8045 & n8046 ) ;
  assign n8049 = ( n7745 & n8047 ) | ( n7745 & ~n8048 ) | ( n8047 & ~n8048 ) ;
  assign n8050 = ( x112 & n8044 ) | ( x112 & ~n8049 ) | ( n8044 & ~n8049 ) ;
  assign n8051 = ( x112 & n7746 ) | ( x112 & ~n7763 ) | ( n7746 & ~n7763 ) ;
  assign n8052 = x112 & n7746 ;
  assign n8053 = ( n7751 & n8051 ) | ( n7751 & n8052 ) | ( n8051 & n8052 ) ;
  assign n8054 = ( ~n7751 & n8051 ) | ( ~n7751 & n8052 ) | ( n8051 & n8052 ) ;
  assign n8055 = ( n7751 & ~n8053 ) | ( n7751 & n8054 ) | ( ~n8053 & n8054 ) ;
  assign n8056 = ( x113 & n8050 ) | ( x113 & ~n8055 ) | ( n8050 & ~n8055 ) ;
  assign n8057 = ( x113 & n7752 ) | ( x113 & ~n7763 ) | ( n7752 & ~n7763 ) ;
  assign n8058 = x113 & n7752 ;
  assign n8059 = ( n7757 & n8057 ) | ( n7757 & n8058 ) | ( n8057 & n8058 ) ;
  assign n8060 = ( ~n7757 & n8057 ) | ( ~n7757 & n8058 ) | ( n8057 & n8058 ) ;
  assign n8061 = ( n7757 & ~n8059 ) | ( n7757 & n8060 ) | ( ~n8059 & n8060 ) ;
  assign n8062 = ( x114 & n8056 ) | ( x114 & ~n8061 ) | ( n8056 & ~n8061 ) ;
  assign n8063 = x115 | n8062 ;
  assign n8064 = ( x115 & n142 ) | ( x115 & n8062 ) | ( n142 & n8062 ) ;
  assign n8065 = ( n7761 & ~n8063 ) | ( n7761 & n8064 ) | ( ~n8063 & n8064 ) ;
  assign n8066 = ( x115 & ~n7761 ) | ( x115 & n8062 ) | ( ~n7761 & n8062 ) ;
  assign n8067 = n142 | n8066 ;
  assign n8068 = ( x12 & ~x64 ) | ( x12 & n8067 ) | ( ~x64 & n8067 ) ;
  assign n8069 = ~x12 & n8067 ;
  assign n8070 = ( n7767 & n8068 ) | ( n7767 & ~n8069 ) | ( n8068 & ~n8069 ) ;
  assign n8071 = ~x11 & x64 ;
  assign n8072 = ( x65 & ~n8070 ) | ( x65 & n8071 ) | ( ~n8070 & n8071 ) ;
  assign n8073 = ( x65 & n7767 ) | ( x65 & ~n8067 ) | ( n7767 & ~n8067 ) ;
  assign n8074 = x65 & n7767 ;
  assign n8075 = ( n7766 & n8073 ) | ( n7766 & n8074 ) | ( n8073 & n8074 ) ;
  assign n8076 = ( ~n7766 & n8073 ) | ( ~n7766 & n8074 ) | ( n8073 & n8074 ) ;
  assign n8077 = ( n7766 & ~n8075 ) | ( n7766 & n8076 ) | ( ~n8075 & n8076 ) ;
  assign n8078 = ( x66 & n8072 ) | ( x66 & ~n8077 ) | ( n8072 & ~n8077 ) ;
  assign n8079 = ( x66 & n7768 ) | ( x66 & ~n8067 ) | ( n7768 & ~n8067 ) ;
  assign n8080 = x66 & n7768 ;
  assign n8081 = ( n7773 & n8079 ) | ( n7773 & n8080 ) | ( n8079 & n8080 ) ;
  assign n8082 = ( ~n7773 & n8079 ) | ( ~n7773 & n8080 ) | ( n8079 & n8080 ) ;
  assign n8083 = ( n7773 & ~n8081 ) | ( n7773 & n8082 ) | ( ~n8081 & n8082 ) ;
  assign n8084 = ( x67 & n8078 ) | ( x67 & ~n8083 ) | ( n8078 & ~n8083 ) ;
  assign n8085 = ( x67 & n7774 ) | ( x67 & ~n8067 ) | ( n7774 & ~n8067 ) ;
  assign n8086 = x67 & n7774 ;
  assign n8087 = ( ~n7779 & n8085 ) | ( ~n7779 & n8086 ) | ( n8085 & n8086 ) ;
  assign n8088 = ( n7779 & n8085 ) | ( n7779 & n8086 ) | ( n8085 & n8086 ) ;
  assign n8089 = ( n7779 & n8087 ) | ( n7779 & ~n8088 ) | ( n8087 & ~n8088 ) ;
  assign n8090 = ( x68 & n8084 ) | ( x68 & ~n8089 ) | ( n8084 & ~n8089 ) ;
  assign n8091 = ( x68 & n7780 ) | ( x68 & ~n8067 ) | ( n7780 & ~n8067 ) ;
  assign n8092 = x68 & n7780 ;
  assign n8093 = ( n7785 & n8091 ) | ( n7785 & n8092 ) | ( n8091 & n8092 ) ;
  assign n8094 = ( ~n7785 & n8091 ) | ( ~n7785 & n8092 ) | ( n8091 & n8092 ) ;
  assign n8095 = ( n7785 & ~n8093 ) | ( n7785 & n8094 ) | ( ~n8093 & n8094 ) ;
  assign n8096 = ( x69 & n8090 ) | ( x69 & ~n8095 ) | ( n8090 & ~n8095 ) ;
  assign n8097 = ( x69 & n7786 ) | ( x69 & ~n8067 ) | ( n7786 & ~n8067 ) ;
  assign n8098 = x69 & n7786 ;
  assign n8099 = ( ~n7791 & n8097 ) | ( ~n7791 & n8098 ) | ( n8097 & n8098 ) ;
  assign n8100 = ( n7791 & n8097 ) | ( n7791 & n8098 ) | ( n8097 & n8098 ) ;
  assign n8101 = ( n7791 & n8099 ) | ( n7791 & ~n8100 ) | ( n8099 & ~n8100 ) ;
  assign n8102 = ( x70 & n8096 ) | ( x70 & ~n8101 ) | ( n8096 & ~n8101 ) ;
  assign n8103 = ( x70 & n7792 ) | ( x70 & ~n8067 ) | ( n7792 & ~n8067 ) ;
  assign n8104 = x70 & n7792 ;
  assign n8105 = ( n7797 & n8103 ) | ( n7797 & n8104 ) | ( n8103 & n8104 ) ;
  assign n8106 = ( ~n7797 & n8103 ) | ( ~n7797 & n8104 ) | ( n8103 & n8104 ) ;
  assign n8107 = ( n7797 & ~n8105 ) | ( n7797 & n8106 ) | ( ~n8105 & n8106 ) ;
  assign n8108 = ( x71 & n8102 ) | ( x71 & ~n8107 ) | ( n8102 & ~n8107 ) ;
  assign n8109 = ( x71 & n7798 ) | ( x71 & ~n8067 ) | ( n7798 & ~n8067 ) ;
  assign n8110 = x71 & n7798 ;
  assign n8111 = ( ~n7803 & n8109 ) | ( ~n7803 & n8110 ) | ( n8109 & n8110 ) ;
  assign n8112 = ( n7803 & n8109 ) | ( n7803 & n8110 ) | ( n8109 & n8110 ) ;
  assign n8113 = ( n7803 & n8111 ) | ( n7803 & ~n8112 ) | ( n8111 & ~n8112 ) ;
  assign n8114 = ( x72 & n8108 ) | ( x72 & ~n8113 ) | ( n8108 & ~n8113 ) ;
  assign n8115 = ( x72 & n7804 ) | ( x72 & ~n8067 ) | ( n7804 & ~n8067 ) ;
  assign n8116 = x72 & n7804 ;
  assign n8117 = ( n7809 & n8115 ) | ( n7809 & n8116 ) | ( n8115 & n8116 ) ;
  assign n8118 = ( ~n7809 & n8115 ) | ( ~n7809 & n8116 ) | ( n8115 & n8116 ) ;
  assign n8119 = ( n7809 & ~n8117 ) | ( n7809 & n8118 ) | ( ~n8117 & n8118 ) ;
  assign n8120 = ( x73 & n8114 ) | ( x73 & ~n8119 ) | ( n8114 & ~n8119 ) ;
  assign n8121 = ( x73 & n7810 ) | ( x73 & ~n8067 ) | ( n7810 & ~n8067 ) ;
  assign n8122 = x73 & n7810 ;
  assign n8123 = ( ~n7815 & n8121 ) | ( ~n7815 & n8122 ) | ( n8121 & n8122 ) ;
  assign n8124 = ( n7815 & n8121 ) | ( n7815 & n8122 ) | ( n8121 & n8122 ) ;
  assign n8125 = ( n7815 & n8123 ) | ( n7815 & ~n8124 ) | ( n8123 & ~n8124 ) ;
  assign n8126 = ( x74 & n8120 ) | ( x74 & ~n8125 ) | ( n8120 & ~n8125 ) ;
  assign n8127 = ( x74 & n7816 ) | ( x74 & ~n8067 ) | ( n7816 & ~n8067 ) ;
  assign n8128 = x74 & n7816 ;
  assign n8129 = ( n7821 & n8127 ) | ( n7821 & n8128 ) | ( n8127 & n8128 ) ;
  assign n8130 = ( ~n7821 & n8127 ) | ( ~n7821 & n8128 ) | ( n8127 & n8128 ) ;
  assign n8131 = ( n7821 & ~n8129 ) | ( n7821 & n8130 ) | ( ~n8129 & n8130 ) ;
  assign n8132 = ( x75 & n8126 ) | ( x75 & ~n8131 ) | ( n8126 & ~n8131 ) ;
  assign n8133 = ( x75 & n7822 ) | ( x75 & ~n8067 ) | ( n7822 & ~n8067 ) ;
  assign n8134 = x75 & n7822 ;
  assign n8135 = ( ~n7827 & n8133 ) | ( ~n7827 & n8134 ) | ( n8133 & n8134 ) ;
  assign n8136 = ( n7827 & n8133 ) | ( n7827 & n8134 ) | ( n8133 & n8134 ) ;
  assign n8137 = ( n7827 & n8135 ) | ( n7827 & ~n8136 ) | ( n8135 & ~n8136 ) ;
  assign n8138 = ( x76 & n8132 ) | ( x76 & ~n8137 ) | ( n8132 & ~n8137 ) ;
  assign n8139 = ( x76 & n7828 ) | ( x76 & ~n8067 ) | ( n7828 & ~n8067 ) ;
  assign n8140 = x76 & n7828 ;
  assign n8141 = ( n7833 & n8139 ) | ( n7833 & n8140 ) | ( n8139 & n8140 ) ;
  assign n8142 = ( ~n7833 & n8139 ) | ( ~n7833 & n8140 ) | ( n8139 & n8140 ) ;
  assign n8143 = ( n7833 & ~n8141 ) | ( n7833 & n8142 ) | ( ~n8141 & n8142 ) ;
  assign n8144 = ( x77 & n8138 ) | ( x77 & ~n8143 ) | ( n8138 & ~n8143 ) ;
  assign n8145 = ( x77 & n7834 ) | ( x77 & ~n8067 ) | ( n7834 & ~n8067 ) ;
  assign n8146 = x77 & n7834 ;
  assign n8147 = ( ~n7839 & n8145 ) | ( ~n7839 & n8146 ) | ( n8145 & n8146 ) ;
  assign n8148 = ( n7839 & n8145 ) | ( n7839 & n8146 ) | ( n8145 & n8146 ) ;
  assign n8149 = ( n7839 & n8147 ) | ( n7839 & ~n8148 ) | ( n8147 & ~n8148 ) ;
  assign n8150 = ( x78 & n8144 ) | ( x78 & ~n8149 ) | ( n8144 & ~n8149 ) ;
  assign n8151 = ( x78 & n7840 ) | ( x78 & ~n8067 ) | ( n7840 & ~n8067 ) ;
  assign n8152 = x78 & n7840 ;
  assign n8153 = ( n7845 & n8151 ) | ( n7845 & n8152 ) | ( n8151 & n8152 ) ;
  assign n8154 = ( ~n7845 & n8151 ) | ( ~n7845 & n8152 ) | ( n8151 & n8152 ) ;
  assign n8155 = ( n7845 & ~n8153 ) | ( n7845 & n8154 ) | ( ~n8153 & n8154 ) ;
  assign n8156 = ( x79 & n8150 ) | ( x79 & ~n8155 ) | ( n8150 & ~n8155 ) ;
  assign n8157 = ( x79 & n7846 ) | ( x79 & ~n8067 ) | ( n7846 & ~n8067 ) ;
  assign n8158 = x79 & n7846 ;
  assign n8159 = ( ~n7851 & n8157 ) | ( ~n7851 & n8158 ) | ( n8157 & n8158 ) ;
  assign n8160 = ( n7851 & n8157 ) | ( n7851 & n8158 ) | ( n8157 & n8158 ) ;
  assign n8161 = ( n7851 & n8159 ) | ( n7851 & ~n8160 ) | ( n8159 & ~n8160 ) ;
  assign n8162 = ( x80 & n8156 ) | ( x80 & ~n8161 ) | ( n8156 & ~n8161 ) ;
  assign n8163 = ( x80 & n7852 ) | ( x80 & ~n8067 ) | ( n7852 & ~n8067 ) ;
  assign n8164 = x80 & n7852 ;
  assign n8165 = ( n7857 & n8163 ) | ( n7857 & n8164 ) | ( n8163 & n8164 ) ;
  assign n8166 = ( ~n7857 & n8163 ) | ( ~n7857 & n8164 ) | ( n8163 & n8164 ) ;
  assign n8167 = ( n7857 & ~n8165 ) | ( n7857 & n8166 ) | ( ~n8165 & n8166 ) ;
  assign n8168 = ( x81 & n8162 ) | ( x81 & ~n8167 ) | ( n8162 & ~n8167 ) ;
  assign n8169 = ( x81 & n7858 ) | ( x81 & ~n8067 ) | ( n7858 & ~n8067 ) ;
  assign n8170 = x81 & n7858 ;
  assign n8171 = ( ~n7863 & n8169 ) | ( ~n7863 & n8170 ) | ( n8169 & n8170 ) ;
  assign n8172 = ( n7863 & n8169 ) | ( n7863 & n8170 ) | ( n8169 & n8170 ) ;
  assign n8173 = ( n7863 & n8171 ) | ( n7863 & ~n8172 ) | ( n8171 & ~n8172 ) ;
  assign n8174 = ( x82 & n8168 ) | ( x82 & ~n8173 ) | ( n8168 & ~n8173 ) ;
  assign n8175 = ( x82 & n7864 ) | ( x82 & ~n8067 ) | ( n7864 & ~n8067 ) ;
  assign n8176 = x82 & n7864 ;
  assign n8177 = ( n7869 & n8175 ) | ( n7869 & n8176 ) | ( n8175 & n8176 ) ;
  assign n8178 = ( ~n7869 & n8175 ) | ( ~n7869 & n8176 ) | ( n8175 & n8176 ) ;
  assign n8179 = ( n7869 & ~n8177 ) | ( n7869 & n8178 ) | ( ~n8177 & n8178 ) ;
  assign n8180 = ( x83 & n8174 ) | ( x83 & ~n8179 ) | ( n8174 & ~n8179 ) ;
  assign n8181 = ( x83 & n7870 ) | ( x83 & ~n8067 ) | ( n7870 & ~n8067 ) ;
  assign n8182 = x83 & n7870 ;
  assign n8183 = ( ~n7875 & n8181 ) | ( ~n7875 & n8182 ) | ( n8181 & n8182 ) ;
  assign n8184 = ( n7875 & n8181 ) | ( n7875 & n8182 ) | ( n8181 & n8182 ) ;
  assign n8185 = ( n7875 & n8183 ) | ( n7875 & ~n8184 ) | ( n8183 & ~n8184 ) ;
  assign n8186 = ( x84 & n8180 ) | ( x84 & ~n8185 ) | ( n8180 & ~n8185 ) ;
  assign n8187 = ( x84 & n7876 ) | ( x84 & ~n8067 ) | ( n7876 & ~n8067 ) ;
  assign n8188 = x84 & n7876 ;
  assign n8189 = ( n7881 & n8187 ) | ( n7881 & n8188 ) | ( n8187 & n8188 ) ;
  assign n8190 = ( ~n7881 & n8187 ) | ( ~n7881 & n8188 ) | ( n8187 & n8188 ) ;
  assign n8191 = ( n7881 & ~n8189 ) | ( n7881 & n8190 ) | ( ~n8189 & n8190 ) ;
  assign n8192 = ( x85 & n8186 ) | ( x85 & ~n8191 ) | ( n8186 & ~n8191 ) ;
  assign n8193 = ( x85 & n7882 ) | ( x85 & ~n8067 ) | ( n7882 & ~n8067 ) ;
  assign n8194 = x85 & n7882 ;
  assign n8195 = ( ~n7887 & n8193 ) | ( ~n7887 & n8194 ) | ( n8193 & n8194 ) ;
  assign n8196 = ( n7887 & n8193 ) | ( n7887 & n8194 ) | ( n8193 & n8194 ) ;
  assign n8197 = ( n7887 & n8195 ) | ( n7887 & ~n8196 ) | ( n8195 & ~n8196 ) ;
  assign n8198 = ( x86 & n8192 ) | ( x86 & ~n8197 ) | ( n8192 & ~n8197 ) ;
  assign n8199 = ( x86 & n7888 ) | ( x86 & ~n8067 ) | ( n7888 & ~n8067 ) ;
  assign n8200 = x86 & n7888 ;
  assign n8201 = ( n7893 & n8199 ) | ( n7893 & n8200 ) | ( n8199 & n8200 ) ;
  assign n8202 = ( ~n7893 & n8199 ) | ( ~n7893 & n8200 ) | ( n8199 & n8200 ) ;
  assign n8203 = ( n7893 & ~n8201 ) | ( n7893 & n8202 ) | ( ~n8201 & n8202 ) ;
  assign n8204 = ( x87 & n8198 ) | ( x87 & ~n8203 ) | ( n8198 & ~n8203 ) ;
  assign n8205 = ( x87 & n7894 ) | ( x87 & ~n8067 ) | ( n7894 & ~n8067 ) ;
  assign n8206 = x87 & n7894 ;
  assign n8207 = ( ~n7899 & n8205 ) | ( ~n7899 & n8206 ) | ( n8205 & n8206 ) ;
  assign n8208 = ( n7899 & n8205 ) | ( n7899 & n8206 ) | ( n8205 & n8206 ) ;
  assign n8209 = ( n7899 & n8207 ) | ( n7899 & ~n8208 ) | ( n8207 & ~n8208 ) ;
  assign n8210 = ( x88 & n8204 ) | ( x88 & ~n8209 ) | ( n8204 & ~n8209 ) ;
  assign n8211 = ( x88 & n7900 ) | ( x88 & ~n8067 ) | ( n7900 & ~n8067 ) ;
  assign n8212 = x88 & n7900 ;
  assign n8213 = ( n7905 & n8211 ) | ( n7905 & n8212 ) | ( n8211 & n8212 ) ;
  assign n8214 = ( ~n7905 & n8211 ) | ( ~n7905 & n8212 ) | ( n8211 & n8212 ) ;
  assign n8215 = ( n7905 & ~n8213 ) | ( n7905 & n8214 ) | ( ~n8213 & n8214 ) ;
  assign n8216 = ( x89 & n8210 ) | ( x89 & ~n8215 ) | ( n8210 & ~n8215 ) ;
  assign n8217 = ( x89 & n7906 ) | ( x89 & ~n8067 ) | ( n7906 & ~n8067 ) ;
  assign n8218 = x89 & n7906 ;
  assign n8219 = ( ~n7911 & n8217 ) | ( ~n7911 & n8218 ) | ( n8217 & n8218 ) ;
  assign n8220 = ( n7911 & n8217 ) | ( n7911 & n8218 ) | ( n8217 & n8218 ) ;
  assign n8221 = ( n7911 & n8219 ) | ( n7911 & ~n8220 ) | ( n8219 & ~n8220 ) ;
  assign n8222 = ( x90 & n8216 ) | ( x90 & ~n8221 ) | ( n8216 & ~n8221 ) ;
  assign n8223 = ( x90 & n7912 ) | ( x90 & ~n8067 ) | ( n7912 & ~n8067 ) ;
  assign n8224 = x90 & n7912 ;
  assign n8225 = ( n7917 & n8223 ) | ( n7917 & n8224 ) | ( n8223 & n8224 ) ;
  assign n8226 = ( ~n7917 & n8223 ) | ( ~n7917 & n8224 ) | ( n8223 & n8224 ) ;
  assign n8227 = ( n7917 & ~n8225 ) | ( n7917 & n8226 ) | ( ~n8225 & n8226 ) ;
  assign n8228 = ( x91 & n8222 ) | ( x91 & ~n8227 ) | ( n8222 & ~n8227 ) ;
  assign n8229 = ( x91 & n7918 ) | ( x91 & ~n8067 ) | ( n7918 & ~n8067 ) ;
  assign n8230 = x91 & n7918 ;
  assign n8231 = ( ~n7923 & n8229 ) | ( ~n7923 & n8230 ) | ( n8229 & n8230 ) ;
  assign n8232 = ( n7923 & n8229 ) | ( n7923 & n8230 ) | ( n8229 & n8230 ) ;
  assign n8233 = ( n7923 & n8231 ) | ( n7923 & ~n8232 ) | ( n8231 & ~n8232 ) ;
  assign n8234 = ( x92 & n8228 ) | ( x92 & ~n8233 ) | ( n8228 & ~n8233 ) ;
  assign n8235 = ( x92 & n7924 ) | ( x92 & ~n8067 ) | ( n7924 & ~n8067 ) ;
  assign n8236 = x92 & n7924 ;
  assign n8237 = ( n7929 & n8235 ) | ( n7929 & n8236 ) | ( n8235 & n8236 ) ;
  assign n8238 = ( ~n7929 & n8235 ) | ( ~n7929 & n8236 ) | ( n8235 & n8236 ) ;
  assign n8239 = ( n7929 & ~n8237 ) | ( n7929 & n8238 ) | ( ~n8237 & n8238 ) ;
  assign n8240 = ( x93 & n8234 ) | ( x93 & ~n8239 ) | ( n8234 & ~n8239 ) ;
  assign n8241 = ( x93 & n7930 ) | ( x93 & ~n8067 ) | ( n7930 & ~n8067 ) ;
  assign n8242 = x93 & n7930 ;
  assign n8243 = ( ~n7935 & n8241 ) | ( ~n7935 & n8242 ) | ( n8241 & n8242 ) ;
  assign n8244 = ( n7935 & n8241 ) | ( n7935 & n8242 ) | ( n8241 & n8242 ) ;
  assign n8245 = ( n7935 & n8243 ) | ( n7935 & ~n8244 ) | ( n8243 & ~n8244 ) ;
  assign n8246 = ( x94 & n8240 ) | ( x94 & ~n8245 ) | ( n8240 & ~n8245 ) ;
  assign n8247 = ( x94 & n7936 ) | ( x94 & ~n8067 ) | ( n7936 & ~n8067 ) ;
  assign n8248 = x94 & n7936 ;
  assign n8249 = ( n7941 & n8247 ) | ( n7941 & n8248 ) | ( n8247 & n8248 ) ;
  assign n8250 = ( ~n7941 & n8247 ) | ( ~n7941 & n8248 ) | ( n8247 & n8248 ) ;
  assign n8251 = ( n7941 & ~n8249 ) | ( n7941 & n8250 ) | ( ~n8249 & n8250 ) ;
  assign n8252 = ( x95 & n8246 ) | ( x95 & ~n8251 ) | ( n8246 & ~n8251 ) ;
  assign n8253 = ( x95 & n7942 ) | ( x95 & ~n8067 ) | ( n7942 & ~n8067 ) ;
  assign n8254 = x95 & n7942 ;
  assign n8255 = ( ~n7947 & n8253 ) | ( ~n7947 & n8254 ) | ( n8253 & n8254 ) ;
  assign n8256 = ( n7947 & n8253 ) | ( n7947 & n8254 ) | ( n8253 & n8254 ) ;
  assign n8257 = ( n7947 & n8255 ) | ( n7947 & ~n8256 ) | ( n8255 & ~n8256 ) ;
  assign n8258 = ( x96 & n8252 ) | ( x96 & ~n8257 ) | ( n8252 & ~n8257 ) ;
  assign n8259 = ( x96 & n7948 ) | ( x96 & ~n8067 ) | ( n7948 & ~n8067 ) ;
  assign n8260 = x96 & n7948 ;
  assign n8261 = ( n7953 & n8259 ) | ( n7953 & n8260 ) | ( n8259 & n8260 ) ;
  assign n8262 = ( ~n7953 & n8259 ) | ( ~n7953 & n8260 ) | ( n8259 & n8260 ) ;
  assign n8263 = ( n7953 & ~n8261 ) | ( n7953 & n8262 ) | ( ~n8261 & n8262 ) ;
  assign n8264 = ( x97 & n8258 ) | ( x97 & ~n8263 ) | ( n8258 & ~n8263 ) ;
  assign n8265 = ( x97 & n7954 ) | ( x97 & ~n8067 ) | ( n7954 & ~n8067 ) ;
  assign n8266 = x97 & n7954 ;
  assign n8267 = ( ~n7959 & n8265 ) | ( ~n7959 & n8266 ) | ( n8265 & n8266 ) ;
  assign n8268 = ( n7959 & n8265 ) | ( n7959 & n8266 ) | ( n8265 & n8266 ) ;
  assign n8269 = ( n7959 & n8267 ) | ( n7959 & ~n8268 ) | ( n8267 & ~n8268 ) ;
  assign n8270 = ( x98 & n8264 ) | ( x98 & ~n8269 ) | ( n8264 & ~n8269 ) ;
  assign n8271 = ( x98 & n7960 ) | ( x98 & ~n8067 ) | ( n7960 & ~n8067 ) ;
  assign n8272 = x98 & n7960 ;
  assign n8273 = ( n7965 & n8271 ) | ( n7965 & n8272 ) | ( n8271 & n8272 ) ;
  assign n8274 = ( ~n7965 & n8271 ) | ( ~n7965 & n8272 ) | ( n8271 & n8272 ) ;
  assign n8275 = ( n7965 & ~n8273 ) | ( n7965 & n8274 ) | ( ~n8273 & n8274 ) ;
  assign n8276 = ( x99 & n8270 ) | ( x99 & ~n8275 ) | ( n8270 & ~n8275 ) ;
  assign n8277 = ( x99 & n7966 ) | ( x99 & ~n8067 ) | ( n7966 & ~n8067 ) ;
  assign n8278 = x99 & n7966 ;
  assign n8279 = ( ~n7971 & n8277 ) | ( ~n7971 & n8278 ) | ( n8277 & n8278 ) ;
  assign n8280 = ( n7971 & n8277 ) | ( n7971 & n8278 ) | ( n8277 & n8278 ) ;
  assign n8281 = ( n7971 & n8279 ) | ( n7971 & ~n8280 ) | ( n8279 & ~n8280 ) ;
  assign n8282 = ( x100 & n8276 ) | ( x100 & ~n8281 ) | ( n8276 & ~n8281 ) ;
  assign n8283 = ( x100 & n7972 ) | ( x100 & ~n8067 ) | ( n7972 & ~n8067 ) ;
  assign n8284 = x100 & n7972 ;
  assign n8285 = ( n7977 & n8283 ) | ( n7977 & n8284 ) | ( n8283 & n8284 ) ;
  assign n8286 = ( ~n7977 & n8283 ) | ( ~n7977 & n8284 ) | ( n8283 & n8284 ) ;
  assign n8287 = ( n7977 & ~n8285 ) | ( n7977 & n8286 ) | ( ~n8285 & n8286 ) ;
  assign n8288 = ( x101 & n8282 ) | ( x101 & ~n8287 ) | ( n8282 & ~n8287 ) ;
  assign n8289 = ( x101 & n7978 ) | ( x101 & ~n8067 ) | ( n7978 & ~n8067 ) ;
  assign n8290 = x101 & n7978 ;
  assign n8291 = ( ~n7983 & n8289 ) | ( ~n7983 & n8290 ) | ( n8289 & n8290 ) ;
  assign n8292 = ( n7983 & n8289 ) | ( n7983 & n8290 ) | ( n8289 & n8290 ) ;
  assign n8293 = ( n7983 & n8291 ) | ( n7983 & ~n8292 ) | ( n8291 & ~n8292 ) ;
  assign n8294 = ( x102 & n8288 ) | ( x102 & ~n8293 ) | ( n8288 & ~n8293 ) ;
  assign n8295 = ( x102 & n7984 ) | ( x102 & ~n8067 ) | ( n7984 & ~n8067 ) ;
  assign n8296 = x102 & n7984 ;
  assign n8297 = ( n7989 & n8295 ) | ( n7989 & n8296 ) | ( n8295 & n8296 ) ;
  assign n8298 = ( ~n7989 & n8295 ) | ( ~n7989 & n8296 ) | ( n8295 & n8296 ) ;
  assign n8299 = ( n7989 & ~n8297 ) | ( n7989 & n8298 ) | ( ~n8297 & n8298 ) ;
  assign n8300 = ( x103 & n8294 ) | ( x103 & ~n8299 ) | ( n8294 & ~n8299 ) ;
  assign n8301 = ( x103 & n7990 ) | ( x103 & ~n8067 ) | ( n7990 & ~n8067 ) ;
  assign n8302 = x103 & n7990 ;
  assign n8303 = ( ~n7995 & n8301 ) | ( ~n7995 & n8302 ) | ( n8301 & n8302 ) ;
  assign n8304 = ( n7995 & n8301 ) | ( n7995 & n8302 ) | ( n8301 & n8302 ) ;
  assign n8305 = ( n7995 & n8303 ) | ( n7995 & ~n8304 ) | ( n8303 & ~n8304 ) ;
  assign n8306 = ( x104 & n8300 ) | ( x104 & ~n8305 ) | ( n8300 & ~n8305 ) ;
  assign n8307 = ( x104 & n7996 ) | ( x104 & ~n8067 ) | ( n7996 & ~n8067 ) ;
  assign n8308 = x104 & n7996 ;
  assign n8309 = ( n8001 & n8307 ) | ( n8001 & n8308 ) | ( n8307 & n8308 ) ;
  assign n8310 = ( ~n8001 & n8307 ) | ( ~n8001 & n8308 ) | ( n8307 & n8308 ) ;
  assign n8311 = ( n8001 & ~n8309 ) | ( n8001 & n8310 ) | ( ~n8309 & n8310 ) ;
  assign n8312 = ( x105 & n8306 ) | ( x105 & ~n8311 ) | ( n8306 & ~n8311 ) ;
  assign n8313 = ( x105 & n8002 ) | ( x105 & ~n8067 ) | ( n8002 & ~n8067 ) ;
  assign n8314 = x105 & n8002 ;
  assign n8315 = ( ~n8007 & n8313 ) | ( ~n8007 & n8314 ) | ( n8313 & n8314 ) ;
  assign n8316 = ( n8007 & n8313 ) | ( n8007 & n8314 ) | ( n8313 & n8314 ) ;
  assign n8317 = ( n8007 & n8315 ) | ( n8007 & ~n8316 ) | ( n8315 & ~n8316 ) ;
  assign n8318 = ( x106 & n8312 ) | ( x106 & ~n8317 ) | ( n8312 & ~n8317 ) ;
  assign n8319 = ( x106 & n8008 ) | ( x106 & ~n8067 ) | ( n8008 & ~n8067 ) ;
  assign n8320 = x106 & n8008 ;
  assign n8321 = ( n8013 & n8319 ) | ( n8013 & n8320 ) | ( n8319 & n8320 ) ;
  assign n8322 = ( ~n8013 & n8319 ) | ( ~n8013 & n8320 ) | ( n8319 & n8320 ) ;
  assign n8323 = ( n8013 & ~n8321 ) | ( n8013 & n8322 ) | ( ~n8321 & n8322 ) ;
  assign n8324 = ( x107 & n8318 ) | ( x107 & ~n8323 ) | ( n8318 & ~n8323 ) ;
  assign n8325 = ( x107 & n8014 ) | ( x107 & ~n8067 ) | ( n8014 & ~n8067 ) ;
  assign n8326 = x107 & n8014 ;
  assign n8327 = ( ~n8019 & n8325 ) | ( ~n8019 & n8326 ) | ( n8325 & n8326 ) ;
  assign n8328 = ( n8019 & n8325 ) | ( n8019 & n8326 ) | ( n8325 & n8326 ) ;
  assign n8329 = ( n8019 & n8327 ) | ( n8019 & ~n8328 ) | ( n8327 & ~n8328 ) ;
  assign n8330 = ( x108 & n8324 ) | ( x108 & ~n8329 ) | ( n8324 & ~n8329 ) ;
  assign n8331 = ( x108 & n8020 ) | ( x108 & ~n8067 ) | ( n8020 & ~n8067 ) ;
  assign n8332 = x108 & n8020 ;
  assign n8333 = ( n8025 & n8331 ) | ( n8025 & n8332 ) | ( n8331 & n8332 ) ;
  assign n8334 = ( ~n8025 & n8331 ) | ( ~n8025 & n8332 ) | ( n8331 & n8332 ) ;
  assign n8335 = ( n8025 & ~n8333 ) | ( n8025 & n8334 ) | ( ~n8333 & n8334 ) ;
  assign n8336 = ( x109 & n8330 ) | ( x109 & ~n8335 ) | ( n8330 & ~n8335 ) ;
  assign n8337 = ( x109 & n8026 ) | ( x109 & ~n8067 ) | ( n8026 & ~n8067 ) ;
  assign n8338 = x109 & n8026 ;
  assign n8339 = ( ~n8031 & n8337 ) | ( ~n8031 & n8338 ) | ( n8337 & n8338 ) ;
  assign n8340 = ( n8031 & n8337 ) | ( n8031 & n8338 ) | ( n8337 & n8338 ) ;
  assign n8341 = ( n8031 & n8339 ) | ( n8031 & ~n8340 ) | ( n8339 & ~n8340 ) ;
  assign n8342 = ( x110 & n8336 ) | ( x110 & ~n8341 ) | ( n8336 & ~n8341 ) ;
  assign n8343 = ( x110 & n8032 ) | ( x110 & ~n8067 ) | ( n8032 & ~n8067 ) ;
  assign n8344 = x110 & n8032 ;
  assign n8345 = ( n8037 & n8343 ) | ( n8037 & n8344 ) | ( n8343 & n8344 ) ;
  assign n8346 = ( ~n8037 & n8343 ) | ( ~n8037 & n8344 ) | ( n8343 & n8344 ) ;
  assign n8347 = ( n8037 & ~n8345 ) | ( n8037 & n8346 ) | ( ~n8345 & n8346 ) ;
  assign n8348 = ( x111 & n8342 ) | ( x111 & ~n8347 ) | ( n8342 & ~n8347 ) ;
  assign n8349 = ( x111 & n8038 ) | ( x111 & ~n8067 ) | ( n8038 & ~n8067 ) ;
  assign n8350 = x111 & n8038 ;
  assign n8351 = ( ~n8043 & n8349 ) | ( ~n8043 & n8350 ) | ( n8349 & n8350 ) ;
  assign n8352 = ( n8043 & n8349 ) | ( n8043 & n8350 ) | ( n8349 & n8350 ) ;
  assign n8353 = ( n8043 & n8351 ) | ( n8043 & ~n8352 ) | ( n8351 & ~n8352 ) ;
  assign n8354 = ( x112 & n8348 ) | ( x112 & ~n8353 ) | ( n8348 & ~n8353 ) ;
  assign n8355 = ( x112 & n8044 ) | ( x112 & ~n8067 ) | ( n8044 & ~n8067 ) ;
  assign n8356 = x112 & n8044 ;
  assign n8357 = ( n8049 & n8355 ) | ( n8049 & n8356 ) | ( n8355 & n8356 ) ;
  assign n8358 = ( ~n8049 & n8355 ) | ( ~n8049 & n8356 ) | ( n8355 & n8356 ) ;
  assign n8359 = ( n8049 & ~n8357 ) | ( n8049 & n8358 ) | ( ~n8357 & n8358 ) ;
  assign n8360 = ( x113 & n8354 ) | ( x113 & ~n8359 ) | ( n8354 & ~n8359 ) ;
  assign n8361 = ( x113 & n8050 ) | ( x113 & ~n8067 ) | ( n8050 & ~n8067 ) ;
  assign n8362 = x113 & n8050 ;
  assign n8363 = ( ~n8055 & n8361 ) | ( ~n8055 & n8362 ) | ( n8361 & n8362 ) ;
  assign n8364 = ( n8055 & n8361 ) | ( n8055 & n8362 ) | ( n8361 & n8362 ) ;
  assign n8365 = ( n8055 & n8363 ) | ( n8055 & ~n8364 ) | ( n8363 & ~n8364 ) ;
  assign n8366 = ( x114 & n8360 ) | ( x114 & ~n8365 ) | ( n8360 & ~n8365 ) ;
  assign n8367 = ( x114 & n8056 ) | ( x114 & ~n8067 ) | ( n8056 & ~n8067 ) ;
  assign n8368 = x114 & n8056 ;
  assign n8369 = ( ~n8061 & n8367 ) | ( ~n8061 & n8368 ) | ( n8367 & n8368 ) ;
  assign n8370 = ( n8061 & n8367 ) | ( n8061 & n8368 ) | ( n8367 & n8368 ) ;
  assign n8371 = ( n8061 & n8369 ) | ( n8061 & ~n8370 ) | ( n8369 & ~n8370 ) ;
  assign n8372 = ( x115 & n8366 ) | ( x115 & ~n8371 ) | ( n8366 & ~n8371 ) ;
  assign n8373 = x116 | n8372 ;
  assign n8374 = ( x116 & n141 ) | ( x116 & n8372 ) | ( n141 & n8372 ) ;
  assign n8375 = ( n8065 & ~n8373 ) | ( n8065 & n8374 ) | ( ~n8373 & n8374 ) ;
  assign n8376 = ( x116 & ~n8065 ) | ( x116 & n8372 ) | ( ~n8065 & n8372 ) ;
  assign n8377 = n141 | n8376 ;
  assign n8378 = ( x11 & ~x64 ) | ( x11 & n8377 ) | ( ~x64 & n8377 ) ;
  assign n8379 = ~x11 & n8377 ;
  assign n8380 = ( n8071 & n8378 ) | ( n8071 & ~n8379 ) | ( n8378 & ~n8379 ) ;
  assign n8381 = ~x10 & x64 ;
  assign n8382 = ( x65 & ~n8380 ) | ( x65 & n8381 ) | ( ~n8380 & n8381 ) ;
  assign n8383 = ( x65 & n8071 ) | ( x65 & ~n8377 ) | ( n8071 & ~n8377 ) ;
  assign n8384 = x65 & n8071 ;
  assign n8385 = ( n8070 & n8383 ) | ( n8070 & n8384 ) | ( n8383 & n8384 ) ;
  assign n8386 = ( ~n8070 & n8383 ) | ( ~n8070 & n8384 ) | ( n8383 & n8384 ) ;
  assign n8387 = ( n8070 & ~n8385 ) | ( n8070 & n8386 ) | ( ~n8385 & n8386 ) ;
  assign n8388 = ( x66 & n8382 ) | ( x66 & ~n8387 ) | ( n8382 & ~n8387 ) ;
  assign n8389 = ( x66 & n8072 ) | ( x66 & ~n8377 ) | ( n8072 & ~n8377 ) ;
  assign n8390 = x66 & n8072 ;
  assign n8391 = ( n8077 & n8389 ) | ( n8077 & n8390 ) | ( n8389 & n8390 ) ;
  assign n8392 = ( ~n8077 & n8389 ) | ( ~n8077 & n8390 ) | ( n8389 & n8390 ) ;
  assign n8393 = ( n8077 & ~n8391 ) | ( n8077 & n8392 ) | ( ~n8391 & n8392 ) ;
  assign n8394 = ( x67 & n8388 ) | ( x67 & ~n8393 ) | ( n8388 & ~n8393 ) ;
  assign n8395 = ( x67 & n8078 ) | ( x67 & ~n8377 ) | ( n8078 & ~n8377 ) ;
  assign n8396 = x67 & n8078 ;
  assign n8397 = ( ~n8083 & n8395 ) | ( ~n8083 & n8396 ) | ( n8395 & n8396 ) ;
  assign n8398 = ( n8083 & n8395 ) | ( n8083 & n8396 ) | ( n8395 & n8396 ) ;
  assign n8399 = ( n8083 & n8397 ) | ( n8083 & ~n8398 ) | ( n8397 & ~n8398 ) ;
  assign n8400 = ( x68 & n8394 ) | ( x68 & ~n8399 ) | ( n8394 & ~n8399 ) ;
  assign n8401 = ( x68 & n8084 ) | ( x68 & ~n8377 ) | ( n8084 & ~n8377 ) ;
  assign n8402 = x68 & n8084 ;
  assign n8403 = ( n8089 & n8401 ) | ( n8089 & n8402 ) | ( n8401 & n8402 ) ;
  assign n8404 = ( ~n8089 & n8401 ) | ( ~n8089 & n8402 ) | ( n8401 & n8402 ) ;
  assign n8405 = ( n8089 & ~n8403 ) | ( n8089 & n8404 ) | ( ~n8403 & n8404 ) ;
  assign n8406 = ( x69 & n8400 ) | ( x69 & ~n8405 ) | ( n8400 & ~n8405 ) ;
  assign n8407 = ( x69 & n8090 ) | ( x69 & ~n8377 ) | ( n8090 & ~n8377 ) ;
  assign n8408 = x69 & n8090 ;
  assign n8409 = ( ~n8095 & n8407 ) | ( ~n8095 & n8408 ) | ( n8407 & n8408 ) ;
  assign n8410 = ( n8095 & n8407 ) | ( n8095 & n8408 ) | ( n8407 & n8408 ) ;
  assign n8411 = ( n8095 & n8409 ) | ( n8095 & ~n8410 ) | ( n8409 & ~n8410 ) ;
  assign n8412 = ( x70 & n8406 ) | ( x70 & ~n8411 ) | ( n8406 & ~n8411 ) ;
  assign n8413 = ( x70 & n8096 ) | ( x70 & ~n8377 ) | ( n8096 & ~n8377 ) ;
  assign n8414 = x70 & n8096 ;
  assign n8415 = ( n8101 & n8413 ) | ( n8101 & n8414 ) | ( n8413 & n8414 ) ;
  assign n8416 = ( ~n8101 & n8413 ) | ( ~n8101 & n8414 ) | ( n8413 & n8414 ) ;
  assign n8417 = ( n8101 & ~n8415 ) | ( n8101 & n8416 ) | ( ~n8415 & n8416 ) ;
  assign n8418 = ( x71 & n8412 ) | ( x71 & ~n8417 ) | ( n8412 & ~n8417 ) ;
  assign n8419 = ( x71 & n8102 ) | ( x71 & ~n8377 ) | ( n8102 & ~n8377 ) ;
  assign n8420 = x71 & n8102 ;
  assign n8421 = ( ~n8107 & n8419 ) | ( ~n8107 & n8420 ) | ( n8419 & n8420 ) ;
  assign n8422 = ( n8107 & n8419 ) | ( n8107 & n8420 ) | ( n8419 & n8420 ) ;
  assign n8423 = ( n8107 & n8421 ) | ( n8107 & ~n8422 ) | ( n8421 & ~n8422 ) ;
  assign n8424 = ( x72 & n8418 ) | ( x72 & ~n8423 ) | ( n8418 & ~n8423 ) ;
  assign n8425 = ( x72 & n8108 ) | ( x72 & ~n8377 ) | ( n8108 & ~n8377 ) ;
  assign n8426 = x72 & n8108 ;
  assign n8427 = ( n8113 & n8425 ) | ( n8113 & n8426 ) | ( n8425 & n8426 ) ;
  assign n8428 = ( ~n8113 & n8425 ) | ( ~n8113 & n8426 ) | ( n8425 & n8426 ) ;
  assign n8429 = ( n8113 & ~n8427 ) | ( n8113 & n8428 ) | ( ~n8427 & n8428 ) ;
  assign n8430 = ( x73 & n8424 ) | ( x73 & ~n8429 ) | ( n8424 & ~n8429 ) ;
  assign n8431 = ( x73 & n8114 ) | ( x73 & ~n8377 ) | ( n8114 & ~n8377 ) ;
  assign n8432 = x73 & n8114 ;
  assign n8433 = ( ~n8119 & n8431 ) | ( ~n8119 & n8432 ) | ( n8431 & n8432 ) ;
  assign n8434 = ( n8119 & n8431 ) | ( n8119 & n8432 ) | ( n8431 & n8432 ) ;
  assign n8435 = ( n8119 & n8433 ) | ( n8119 & ~n8434 ) | ( n8433 & ~n8434 ) ;
  assign n8436 = ( x74 & n8430 ) | ( x74 & ~n8435 ) | ( n8430 & ~n8435 ) ;
  assign n8437 = ( x74 & n8120 ) | ( x74 & ~n8377 ) | ( n8120 & ~n8377 ) ;
  assign n8438 = x74 & n8120 ;
  assign n8439 = ( n8125 & n8437 ) | ( n8125 & n8438 ) | ( n8437 & n8438 ) ;
  assign n8440 = ( ~n8125 & n8437 ) | ( ~n8125 & n8438 ) | ( n8437 & n8438 ) ;
  assign n8441 = ( n8125 & ~n8439 ) | ( n8125 & n8440 ) | ( ~n8439 & n8440 ) ;
  assign n8442 = ( x75 & n8436 ) | ( x75 & ~n8441 ) | ( n8436 & ~n8441 ) ;
  assign n8443 = ( x75 & n8126 ) | ( x75 & ~n8377 ) | ( n8126 & ~n8377 ) ;
  assign n8444 = x75 & n8126 ;
  assign n8445 = ( ~n8131 & n8443 ) | ( ~n8131 & n8444 ) | ( n8443 & n8444 ) ;
  assign n8446 = ( n8131 & n8443 ) | ( n8131 & n8444 ) | ( n8443 & n8444 ) ;
  assign n8447 = ( n8131 & n8445 ) | ( n8131 & ~n8446 ) | ( n8445 & ~n8446 ) ;
  assign n8448 = ( x76 & n8442 ) | ( x76 & ~n8447 ) | ( n8442 & ~n8447 ) ;
  assign n8449 = ( x76 & n8132 ) | ( x76 & ~n8377 ) | ( n8132 & ~n8377 ) ;
  assign n8450 = x76 & n8132 ;
  assign n8451 = ( n8137 & n8449 ) | ( n8137 & n8450 ) | ( n8449 & n8450 ) ;
  assign n8452 = ( ~n8137 & n8449 ) | ( ~n8137 & n8450 ) | ( n8449 & n8450 ) ;
  assign n8453 = ( n8137 & ~n8451 ) | ( n8137 & n8452 ) | ( ~n8451 & n8452 ) ;
  assign n8454 = ( x77 & n8448 ) | ( x77 & ~n8453 ) | ( n8448 & ~n8453 ) ;
  assign n8455 = ( x77 & n8138 ) | ( x77 & ~n8377 ) | ( n8138 & ~n8377 ) ;
  assign n8456 = x77 & n8138 ;
  assign n8457 = ( ~n8143 & n8455 ) | ( ~n8143 & n8456 ) | ( n8455 & n8456 ) ;
  assign n8458 = ( n8143 & n8455 ) | ( n8143 & n8456 ) | ( n8455 & n8456 ) ;
  assign n8459 = ( n8143 & n8457 ) | ( n8143 & ~n8458 ) | ( n8457 & ~n8458 ) ;
  assign n8460 = ( x78 & n8454 ) | ( x78 & ~n8459 ) | ( n8454 & ~n8459 ) ;
  assign n8461 = ( x78 & n8144 ) | ( x78 & ~n8377 ) | ( n8144 & ~n8377 ) ;
  assign n8462 = x78 & n8144 ;
  assign n8463 = ( n8149 & n8461 ) | ( n8149 & n8462 ) | ( n8461 & n8462 ) ;
  assign n8464 = ( ~n8149 & n8461 ) | ( ~n8149 & n8462 ) | ( n8461 & n8462 ) ;
  assign n8465 = ( n8149 & ~n8463 ) | ( n8149 & n8464 ) | ( ~n8463 & n8464 ) ;
  assign n8466 = ( x79 & n8460 ) | ( x79 & ~n8465 ) | ( n8460 & ~n8465 ) ;
  assign n8467 = ( x79 & n8150 ) | ( x79 & ~n8377 ) | ( n8150 & ~n8377 ) ;
  assign n8468 = x79 & n8150 ;
  assign n8469 = ( ~n8155 & n8467 ) | ( ~n8155 & n8468 ) | ( n8467 & n8468 ) ;
  assign n8470 = ( n8155 & n8467 ) | ( n8155 & n8468 ) | ( n8467 & n8468 ) ;
  assign n8471 = ( n8155 & n8469 ) | ( n8155 & ~n8470 ) | ( n8469 & ~n8470 ) ;
  assign n8472 = ( x80 & n8466 ) | ( x80 & ~n8471 ) | ( n8466 & ~n8471 ) ;
  assign n8473 = ( x80 & n8156 ) | ( x80 & ~n8377 ) | ( n8156 & ~n8377 ) ;
  assign n8474 = x80 & n8156 ;
  assign n8475 = ( n8161 & n8473 ) | ( n8161 & n8474 ) | ( n8473 & n8474 ) ;
  assign n8476 = ( ~n8161 & n8473 ) | ( ~n8161 & n8474 ) | ( n8473 & n8474 ) ;
  assign n8477 = ( n8161 & ~n8475 ) | ( n8161 & n8476 ) | ( ~n8475 & n8476 ) ;
  assign n8478 = ( x81 & n8472 ) | ( x81 & ~n8477 ) | ( n8472 & ~n8477 ) ;
  assign n8479 = ( x81 & n8162 ) | ( x81 & ~n8377 ) | ( n8162 & ~n8377 ) ;
  assign n8480 = x81 & n8162 ;
  assign n8481 = ( ~n8167 & n8479 ) | ( ~n8167 & n8480 ) | ( n8479 & n8480 ) ;
  assign n8482 = ( n8167 & n8479 ) | ( n8167 & n8480 ) | ( n8479 & n8480 ) ;
  assign n8483 = ( n8167 & n8481 ) | ( n8167 & ~n8482 ) | ( n8481 & ~n8482 ) ;
  assign n8484 = ( x82 & n8478 ) | ( x82 & ~n8483 ) | ( n8478 & ~n8483 ) ;
  assign n8485 = ( x82 & n8168 ) | ( x82 & ~n8377 ) | ( n8168 & ~n8377 ) ;
  assign n8486 = x82 & n8168 ;
  assign n8487 = ( n8173 & n8485 ) | ( n8173 & n8486 ) | ( n8485 & n8486 ) ;
  assign n8488 = ( ~n8173 & n8485 ) | ( ~n8173 & n8486 ) | ( n8485 & n8486 ) ;
  assign n8489 = ( n8173 & ~n8487 ) | ( n8173 & n8488 ) | ( ~n8487 & n8488 ) ;
  assign n8490 = ( x83 & n8484 ) | ( x83 & ~n8489 ) | ( n8484 & ~n8489 ) ;
  assign n8491 = ( x83 & n8174 ) | ( x83 & ~n8377 ) | ( n8174 & ~n8377 ) ;
  assign n8492 = x83 & n8174 ;
  assign n8493 = ( ~n8179 & n8491 ) | ( ~n8179 & n8492 ) | ( n8491 & n8492 ) ;
  assign n8494 = ( n8179 & n8491 ) | ( n8179 & n8492 ) | ( n8491 & n8492 ) ;
  assign n8495 = ( n8179 & n8493 ) | ( n8179 & ~n8494 ) | ( n8493 & ~n8494 ) ;
  assign n8496 = ( x84 & n8490 ) | ( x84 & ~n8495 ) | ( n8490 & ~n8495 ) ;
  assign n8497 = ( x84 & n8180 ) | ( x84 & ~n8377 ) | ( n8180 & ~n8377 ) ;
  assign n8498 = x84 & n8180 ;
  assign n8499 = ( n8185 & n8497 ) | ( n8185 & n8498 ) | ( n8497 & n8498 ) ;
  assign n8500 = ( ~n8185 & n8497 ) | ( ~n8185 & n8498 ) | ( n8497 & n8498 ) ;
  assign n8501 = ( n8185 & ~n8499 ) | ( n8185 & n8500 ) | ( ~n8499 & n8500 ) ;
  assign n8502 = ( x85 & n8496 ) | ( x85 & ~n8501 ) | ( n8496 & ~n8501 ) ;
  assign n8503 = ( x85 & n8186 ) | ( x85 & ~n8377 ) | ( n8186 & ~n8377 ) ;
  assign n8504 = x85 & n8186 ;
  assign n8505 = ( ~n8191 & n8503 ) | ( ~n8191 & n8504 ) | ( n8503 & n8504 ) ;
  assign n8506 = ( n8191 & n8503 ) | ( n8191 & n8504 ) | ( n8503 & n8504 ) ;
  assign n8507 = ( n8191 & n8505 ) | ( n8191 & ~n8506 ) | ( n8505 & ~n8506 ) ;
  assign n8508 = ( x86 & n8502 ) | ( x86 & ~n8507 ) | ( n8502 & ~n8507 ) ;
  assign n8509 = ( x86 & n8192 ) | ( x86 & ~n8377 ) | ( n8192 & ~n8377 ) ;
  assign n8510 = x86 & n8192 ;
  assign n8511 = ( n8197 & n8509 ) | ( n8197 & n8510 ) | ( n8509 & n8510 ) ;
  assign n8512 = ( ~n8197 & n8509 ) | ( ~n8197 & n8510 ) | ( n8509 & n8510 ) ;
  assign n8513 = ( n8197 & ~n8511 ) | ( n8197 & n8512 ) | ( ~n8511 & n8512 ) ;
  assign n8514 = ( x87 & n8508 ) | ( x87 & ~n8513 ) | ( n8508 & ~n8513 ) ;
  assign n8515 = ( x87 & n8198 ) | ( x87 & ~n8377 ) | ( n8198 & ~n8377 ) ;
  assign n8516 = x87 & n8198 ;
  assign n8517 = ( ~n8203 & n8515 ) | ( ~n8203 & n8516 ) | ( n8515 & n8516 ) ;
  assign n8518 = ( n8203 & n8515 ) | ( n8203 & n8516 ) | ( n8515 & n8516 ) ;
  assign n8519 = ( n8203 & n8517 ) | ( n8203 & ~n8518 ) | ( n8517 & ~n8518 ) ;
  assign n8520 = ( x88 & n8514 ) | ( x88 & ~n8519 ) | ( n8514 & ~n8519 ) ;
  assign n8521 = ( x88 & n8204 ) | ( x88 & ~n8377 ) | ( n8204 & ~n8377 ) ;
  assign n8522 = x88 & n8204 ;
  assign n8523 = ( n8209 & n8521 ) | ( n8209 & n8522 ) | ( n8521 & n8522 ) ;
  assign n8524 = ( ~n8209 & n8521 ) | ( ~n8209 & n8522 ) | ( n8521 & n8522 ) ;
  assign n8525 = ( n8209 & ~n8523 ) | ( n8209 & n8524 ) | ( ~n8523 & n8524 ) ;
  assign n8526 = ( x89 & n8520 ) | ( x89 & ~n8525 ) | ( n8520 & ~n8525 ) ;
  assign n8527 = ( x89 & n8210 ) | ( x89 & ~n8377 ) | ( n8210 & ~n8377 ) ;
  assign n8528 = x89 & n8210 ;
  assign n8529 = ( ~n8215 & n8527 ) | ( ~n8215 & n8528 ) | ( n8527 & n8528 ) ;
  assign n8530 = ( n8215 & n8527 ) | ( n8215 & n8528 ) | ( n8527 & n8528 ) ;
  assign n8531 = ( n8215 & n8529 ) | ( n8215 & ~n8530 ) | ( n8529 & ~n8530 ) ;
  assign n8532 = ( x90 & n8526 ) | ( x90 & ~n8531 ) | ( n8526 & ~n8531 ) ;
  assign n8533 = ( x90 & n8216 ) | ( x90 & ~n8377 ) | ( n8216 & ~n8377 ) ;
  assign n8534 = x90 & n8216 ;
  assign n8535 = ( n8221 & n8533 ) | ( n8221 & n8534 ) | ( n8533 & n8534 ) ;
  assign n8536 = ( ~n8221 & n8533 ) | ( ~n8221 & n8534 ) | ( n8533 & n8534 ) ;
  assign n8537 = ( n8221 & ~n8535 ) | ( n8221 & n8536 ) | ( ~n8535 & n8536 ) ;
  assign n8538 = ( x91 & n8532 ) | ( x91 & ~n8537 ) | ( n8532 & ~n8537 ) ;
  assign n8539 = ( x91 & n8222 ) | ( x91 & ~n8377 ) | ( n8222 & ~n8377 ) ;
  assign n8540 = x91 & n8222 ;
  assign n8541 = ( ~n8227 & n8539 ) | ( ~n8227 & n8540 ) | ( n8539 & n8540 ) ;
  assign n8542 = ( n8227 & n8539 ) | ( n8227 & n8540 ) | ( n8539 & n8540 ) ;
  assign n8543 = ( n8227 & n8541 ) | ( n8227 & ~n8542 ) | ( n8541 & ~n8542 ) ;
  assign n8544 = ( x92 & n8538 ) | ( x92 & ~n8543 ) | ( n8538 & ~n8543 ) ;
  assign n8545 = ( x92 & n8228 ) | ( x92 & ~n8377 ) | ( n8228 & ~n8377 ) ;
  assign n8546 = x92 & n8228 ;
  assign n8547 = ( n8233 & n8545 ) | ( n8233 & n8546 ) | ( n8545 & n8546 ) ;
  assign n8548 = ( ~n8233 & n8545 ) | ( ~n8233 & n8546 ) | ( n8545 & n8546 ) ;
  assign n8549 = ( n8233 & ~n8547 ) | ( n8233 & n8548 ) | ( ~n8547 & n8548 ) ;
  assign n8550 = ( x93 & n8544 ) | ( x93 & ~n8549 ) | ( n8544 & ~n8549 ) ;
  assign n8551 = ( x93 & n8234 ) | ( x93 & ~n8377 ) | ( n8234 & ~n8377 ) ;
  assign n8552 = x93 & n8234 ;
  assign n8553 = ( ~n8239 & n8551 ) | ( ~n8239 & n8552 ) | ( n8551 & n8552 ) ;
  assign n8554 = ( n8239 & n8551 ) | ( n8239 & n8552 ) | ( n8551 & n8552 ) ;
  assign n8555 = ( n8239 & n8553 ) | ( n8239 & ~n8554 ) | ( n8553 & ~n8554 ) ;
  assign n8556 = ( x94 & n8550 ) | ( x94 & ~n8555 ) | ( n8550 & ~n8555 ) ;
  assign n8557 = ( x94 & n8240 ) | ( x94 & ~n8377 ) | ( n8240 & ~n8377 ) ;
  assign n8558 = x94 & n8240 ;
  assign n8559 = ( n8245 & n8557 ) | ( n8245 & n8558 ) | ( n8557 & n8558 ) ;
  assign n8560 = ( ~n8245 & n8557 ) | ( ~n8245 & n8558 ) | ( n8557 & n8558 ) ;
  assign n8561 = ( n8245 & ~n8559 ) | ( n8245 & n8560 ) | ( ~n8559 & n8560 ) ;
  assign n8562 = ( x95 & n8556 ) | ( x95 & ~n8561 ) | ( n8556 & ~n8561 ) ;
  assign n8563 = ( x95 & n8246 ) | ( x95 & ~n8377 ) | ( n8246 & ~n8377 ) ;
  assign n8564 = x95 & n8246 ;
  assign n8565 = ( ~n8251 & n8563 ) | ( ~n8251 & n8564 ) | ( n8563 & n8564 ) ;
  assign n8566 = ( n8251 & n8563 ) | ( n8251 & n8564 ) | ( n8563 & n8564 ) ;
  assign n8567 = ( n8251 & n8565 ) | ( n8251 & ~n8566 ) | ( n8565 & ~n8566 ) ;
  assign n8568 = ( x96 & n8562 ) | ( x96 & ~n8567 ) | ( n8562 & ~n8567 ) ;
  assign n8569 = ( x96 & n8252 ) | ( x96 & ~n8377 ) | ( n8252 & ~n8377 ) ;
  assign n8570 = x96 & n8252 ;
  assign n8571 = ( n8257 & n8569 ) | ( n8257 & n8570 ) | ( n8569 & n8570 ) ;
  assign n8572 = ( ~n8257 & n8569 ) | ( ~n8257 & n8570 ) | ( n8569 & n8570 ) ;
  assign n8573 = ( n8257 & ~n8571 ) | ( n8257 & n8572 ) | ( ~n8571 & n8572 ) ;
  assign n8574 = ( x97 & n8568 ) | ( x97 & ~n8573 ) | ( n8568 & ~n8573 ) ;
  assign n8575 = ( x97 & n8258 ) | ( x97 & ~n8377 ) | ( n8258 & ~n8377 ) ;
  assign n8576 = x97 & n8258 ;
  assign n8577 = ( ~n8263 & n8575 ) | ( ~n8263 & n8576 ) | ( n8575 & n8576 ) ;
  assign n8578 = ( n8263 & n8575 ) | ( n8263 & n8576 ) | ( n8575 & n8576 ) ;
  assign n8579 = ( n8263 & n8577 ) | ( n8263 & ~n8578 ) | ( n8577 & ~n8578 ) ;
  assign n8580 = ( x98 & n8574 ) | ( x98 & ~n8579 ) | ( n8574 & ~n8579 ) ;
  assign n8581 = ( x98 & n8264 ) | ( x98 & ~n8377 ) | ( n8264 & ~n8377 ) ;
  assign n8582 = x98 & n8264 ;
  assign n8583 = ( n8269 & n8581 ) | ( n8269 & n8582 ) | ( n8581 & n8582 ) ;
  assign n8584 = ( ~n8269 & n8581 ) | ( ~n8269 & n8582 ) | ( n8581 & n8582 ) ;
  assign n8585 = ( n8269 & ~n8583 ) | ( n8269 & n8584 ) | ( ~n8583 & n8584 ) ;
  assign n8586 = ( x99 & n8580 ) | ( x99 & ~n8585 ) | ( n8580 & ~n8585 ) ;
  assign n8587 = ( x99 & n8270 ) | ( x99 & ~n8377 ) | ( n8270 & ~n8377 ) ;
  assign n8588 = x99 & n8270 ;
  assign n8589 = ( ~n8275 & n8587 ) | ( ~n8275 & n8588 ) | ( n8587 & n8588 ) ;
  assign n8590 = ( n8275 & n8587 ) | ( n8275 & n8588 ) | ( n8587 & n8588 ) ;
  assign n8591 = ( n8275 & n8589 ) | ( n8275 & ~n8590 ) | ( n8589 & ~n8590 ) ;
  assign n8592 = ( x100 & n8586 ) | ( x100 & ~n8591 ) | ( n8586 & ~n8591 ) ;
  assign n8593 = ( x100 & n8276 ) | ( x100 & ~n8377 ) | ( n8276 & ~n8377 ) ;
  assign n8594 = x100 & n8276 ;
  assign n8595 = ( n8281 & n8593 ) | ( n8281 & n8594 ) | ( n8593 & n8594 ) ;
  assign n8596 = ( ~n8281 & n8593 ) | ( ~n8281 & n8594 ) | ( n8593 & n8594 ) ;
  assign n8597 = ( n8281 & ~n8595 ) | ( n8281 & n8596 ) | ( ~n8595 & n8596 ) ;
  assign n8598 = ( x101 & n8592 ) | ( x101 & ~n8597 ) | ( n8592 & ~n8597 ) ;
  assign n8599 = ( x101 & n8282 ) | ( x101 & ~n8377 ) | ( n8282 & ~n8377 ) ;
  assign n8600 = x101 & n8282 ;
  assign n8601 = ( ~n8287 & n8599 ) | ( ~n8287 & n8600 ) | ( n8599 & n8600 ) ;
  assign n8602 = ( n8287 & n8599 ) | ( n8287 & n8600 ) | ( n8599 & n8600 ) ;
  assign n8603 = ( n8287 & n8601 ) | ( n8287 & ~n8602 ) | ( n8601 & ~n8602 ) ;
  assign n8604 = ( x102 & n8598 ) | ( x102 & ~n8603 ) | ( n8598 & ~n8603 ) ;
  assign n8605 = ( x102 & n8288 ) | ( x102 & ~n8377 ) | ( n8288 & ~n8377 ) ;
  assign n8606 = x102 & n8288 ;
  assign n8607 = ( n8293 & n8605 ) | ( n8293 & n8606 ) | ( n8605 & n8606 ) ;
  assign n8608 = ( ~n8293 & n8605 ) | ( ~n8293 & n8606 ) | ( n8605 & n8606 ) ;
  assign n8609 = ( n8293 & ~n8607 ) | ( n8293 & n8608 ) | ( ~n8607 & n8608 ) ;
  assign n8610 = ( x103 & n8604 ) | ( x103 & ~n8609 ) | ( n8604 & ~n8609 ) ;
  assign n8611 = ( x103 & n8294 ) | ( x103 & ~n8377 ) | ( n8294 & ~n8377 ) ;
  assign n8612 = x103 & n8294 ;
  assign n8613 = ( ~n8299 & n8611 ) | ( ~n8299 & n8612 ) | ( n8611 & n8612 ) ;
  assign n8614 = ( n8299 & n8611 ) | ( n8299 & n8612 ) | ( n8611 & n8612 ) ;
  assign n8615 = ( n8299 & n8613 ) | ( n8299 & ~n8614 ) | ( n8613 & ~n8614 ) ;
  assign n8616 = ( x104 & n8610 ) | ( x104 & ~n8615 ) | ( n8610 & ~n8615 ) ;
  assign n8617 = ( x104 & n8300 ) | ( x104 & ~n8377 ) | ( n8300 & ~n8377 ) ;
  assign n8618 = x104 & n8300 ;
  assign n8619 = ( n8305 & n8617 ) | ( n8305 & n8618 ) | ( n8617 & n8618 ) ;
  assign n8620 = ( ~n8305 & n8617 ) | ( ~n8305 & n8618 ) | ( n8617 & n8618 ) ;
  assign n8621 = ( n8305 & ~n8619 ) | ( n8305 & n8620 ) | ( ~n8619 & n8620 ) ;
  assign n8622 = ( x105 & n8616 ) | ( x105 & ~n8621 ) | ( n8616 & ~n8621 ) ;
  assign n8623 = ( x105 & n8306 ) | ( x105 & ~n8377 ) | ( n8306 & ~n8377 ) ;
  assign n8624 = x105 & n8306 ;
  assign n8625 = ( ~n8311 & n8623 ) | ( ~n8311 & n8624 ) | ( n8623 & n8624 ) ;
  assign n8626 = ( n8311 & n8623 ) | ( n8311 & n8624 ) | ( n8623 & n8624 ) ;
  assign n8627 = ( n8311 & n8625 ) | ( n8311 & ~n8626 ) | ( n8625 & ~n8626 ) ;
  assign n8628 = ( x106 & n8622 ) | ( x106 & ~n8627 ) | ( n8622 & ~n8627 ) ;
  assign n8629 = ( x106 & n8312 ) | ( x106 & ~n8377 ) | ( n8312 & ~n8377 ) ;
  assign n8630 = x106 & n8312 ;
  assign n8631 = ( n8317 & n8629 ) | ( n8317 & n8630 ) | ( n8629 & n8630 ) ;
  assign n8632 = ( ~n8317 & n8629 ) | ( ~n8317 & n8630 ) | ( n8629 & n8630 ) ;
  assign n8633 = ( n8317 & ~n8631 ) | ( n8317 & n8632 ) | ( ~n8631 & n8632 ) ;
  assign n8634 = ( x107 & n8628 ) | ( x107 & ~n8633 ) | ( n8628 & ~n8633 ) ;
  assign n8635 = ( x107 & n8318 ) | ( x107 & ~n8377 ) | ( n8318 & ~n8377 ) ;
  assign n8636 = x107 & n8318 ;
  assign n8637 = ( ~n8323 & n8635 ) | ( ~n8323 & n8636 ) | ( n8635 & n8636 ) ;
  assign n8638 = ( n8323 & n8635 ) | ( n8323 & n8636 ) | ( n8635 & n8636 ) ;
  assign n8639 = ( n8323 & n8637 ) | ( n8323 & ~n8638 ) | ( n8637 & ~n8638 ) ;
  assign n8640 = ( x108 & n8634 ) | ( x108 & ~n8639 ) | ( n8634 & ~n8639 ) ;
  assign n8641 = ( x108 & n8324 ) | ( x108 & ~n8377 ) | ( n8324 & ~n8377 ) ;
  assign n8642 = x108 & n8324 ;
  assign n8643 = ( n8329 & n8641 ) | ( n8329 & n8642 ) | ( n8641 & n8642 ) ;
  assign n8644 = ( ~n8329 & n8641 ) | ( ~n8329 & n8642 ) | ( n8641 & n8642 ) ;
  assign n8645 = ( n8329 & ~n8643 ) | ( n8329 & n8644 ) | ( ~n8643 & n8644 ) ;
  assign n8646 = ( x109 & n8640 ) | ( x109 & ~n8645 ) | ( n8640 & ~n8645 ) ;
  assign n8647 = ( x109 & n8330 ) | ( x109 & ~n8377 ) | ( n8330 & ~n8377 ) ;
  assign n8648 = x109 & n8330 ;
  assign n8649 = ( ~n8335 & n8647 ) | ( ~n8335 & n8648 ) | ( n8647 & n8648 ) ;
  assign n8650 = ( n8335 & n8647 ) | ( n8335 & n8648 ) | ( n8647 & n8648 ) ;
  assign n8651 = ( n8335 & n8649 ) | ( n8335 & ~n8650 ) | ( n8649 & ~n8650 ) ;
  assign n8652 = ( x110 & n8646 ) | ( x110 & ~n8651 ) | ( n8646 & ~n8651 ) ;
  assign n8653 = ( x110 & n8336 ) | ( x110 & ~n8377 ) | ( n8336 & ~n8377 ) ;
  assign n8654 = x110 & n8336 ;
  assign n8655 = ( n8341 & n8653 ) | ( n8341 & n8654 ) | ( n8653 & n8654 ) ;
  assign n8656 = ( ~n8341 & n8653 ) | ( ~n8341 & n8654 ) | ( n8653 & n8654 ) ;
  assign n8657 = ( n8341 & ~n8655 ) | ( n8341 & n8656 ) | ( ~n8655 & n8656 ) ;
  assign n8658 = ( x111 & n8652 ) | ( x111 & ~n8657 ) | ( n8652 & ~n8657 ) ;
  assign n8659 = ( x111 & n8342 ) | ( x111 & ~n8377 ) | ( n8342 & ~n8377 ) ;
  assign n8660 = x111 & n8342 ;
  assign n8661 = ( ~n8347 & n8659 ) | ( ~n8347 & n8660 ) | ( n8659 & n8660 ) ;
  assign n8662 = ( n8347 & n8659 ) | ( n8347 & n8660 ) | ( n8659 & n8660 ) ;
  assign n8663 = ( n8347 & n8661 ) | ( n8347 & ~n8662 ) | ( n8661 & ~n8662 ) ;
  assign n8664 = ( x112 & n8658 ) | ( x112 & ~n8663 ) | ( n8658 & ~n8663 ) ;
  assign n8665 = ( x112 & n8348 ) | ( x112 & ~n8377 ) | ( n8348 & ~n8377 ) ;
  assign n8666 = x112 & n8348 ;
  assign n8667 = ( n8353 & n8665 ) | ( n8353 & n8666 ) | ( n8665 & n8666 ) ;
  assign n8668 = ( ~n8353 & n8665 ) | ( ~n8353 & n8666 ) | ( n8665 & n8666 ) ;
  assign n8669 = ( n8353 & ~n8667 ) | ( n8353 & n8668 ) | ( ~n8667 & n8668 ) ;
  assign n8670 = ( x113 & n8664 ) | ( x113 & ~n8669 ) | ( n8664 & ~n8669 ) ;
  assign n8671 = ( x113 & n8354 ) | ( x113 & ~n8377 ) | ( n8354 & ~n8377 ) ;
  assign n8672 = x113 & n8354 ;
  assign n8673 = ( ~n8359 & n8671 ) | ( ~n8359 & n8672 ) | ( n8671 & n8672 ) ;
  assign n8674 = ( n8359 & n8671 ) | ( n8359 & n8672 ) | ( n8671 & n8672 ) ;
  assign n8675 = ( n8359 & n8673 ) | ( n8359 & ~n8674 ) | ( n8673 & ~n8674 ) ;
  assign n8676 = ( x114 & n8670 ) | ( x114 & ~n8675 ) | ( n8670 & ~n8675 ) ;
  assign n8677 = ( x114 & n8360 ) | ( x114 & ~n8377 ) | ( n8360 & ~n8377 ) ;
  assign n8678 = x114 & n8360 ;
  assign n8679 = ( n8365 & n8677 ) | ( n8365 & n8678 ) | ( n8677 & n8678 ) ;
  assign n8680 = ( ~n8365 & n8677 ) | ( ~n8365 & n8678 ) | ( n8677 & n8678 ) ;
  assign n8681 = ( n8365 & ~n8679 ) | ( n8365 & n8680 ) | ( ~n8679 & n8680 ) ;
  assign n8682 = ( x115 & n8676 ) | ( x115 & ~n8681 ) | ( n8676 & ~n8681 ) ;
  assign n8683 = ( x115 & n8366 ) | ( x115 & ~n8377 ) | ( n8366 & ~n8377 ) ;
  assign n8684 = x115 & n8366 ;
  assign n8685 = ( n8371 & n8683 ) | ( n8371 & n8684 ) | ( n8683 & n8684 ) ;
  assign n8686 = ( ~n8371 & n8683 ) | ( ~n8371 & n8684 ) | ( n8683 & n8684 ) ;
  assign n8687 = ( n8371 & ~n8685 ) | ( n8371 & n8686 ) | ( ~n8685 & n8686 ) ;
  assign n8688 = ( x116 & n8682 ) | ( x116 & ~n8687 ) | ( n8682 & ~n8687 ) ;
  assign n8689 = x117 | n8688 ;
  assign n8690 = ( x117 & n140 ) | ( x117 & n8688 ) | ( n140 & n8688 ) ;
  assign n8691 = ( n8375 & ~n8689 ) | ( n8375 & n8690 ) | ( ~n8689 & n8690 ) ;
  assign n8692 = ( x117 & ~n8375 ) | ( x117 & n8688 ) | ( ~n8375 & n8688 ) ;
  assign n8693 = n140 | n8692 ;
  assign n8694 = ( x10 & ~x64 ) | ( x10 & n8693 ) | ( ~x64 & n8693 ) ;
  assign n8695 = ~x10 & n8693 ;
  assign n8696 = ( n8381 & n8694 ) | ( n8381 & ~n8695 ) | ( n8694 & ~n8695 ) ;
  assign n8697 = ~x9 & x64 ;
  assign n8698 = ( x65 & ~n8696 ) | ( x65 & n8697 ) | ( ~n8696 & n8697 ) ;
  assign n8699 = ( x65 & n8381 ) | ( x65 & ~n8693 ) | ( n8381 & ~n8693 ) ;
  assign n8700 = x65 & n8381 ;
  assign n8701 = ( n8380 & n8699 ) | ( n8380 & n8700 ) | ( n8699 & n8700 ) ;
  assign n8702 = ( ~n8380 & n8699 ) | ( ~n8380 & n8700 ) | ( n8699 & n8700 ) ;
  assign n8703 = ( n8380 & ~n8701 ) | ( n8380 & n8702 ) | ( ~n8701 & n8702 ) ;
  assign n8704 = ( x66 & n8698 ) | ( x66 & ~n8703 ) | ( n8698 & ~n8703 ) ;
  assign n8705 = ( x66 & n8382 ) | ( x66 & ~n8693 ) | ( n8382 & ~n8693 ) ;
  assign n8706 = x66 & n8382 ;
  assign n8707 = ( n8387 & n8705 ) | ( n8387 & n8706 ) | ( n8705 & n8706 ) ;
  assign n8708 = ( ~n8387 & n8705 ) | ( ~n8387 & n8706 ) | ( n8705 & n8706 ) ;
  assign n8709 = ( n8387 & ~n8707 ) | ( n8387 & n8708 ) | ( ~n8707 & n8708 ) ;
  assign n8710 = ( x67 & n8704 ) | ( x67 & ~n8709 ) | ( n8704 & ~n8709 ) ;
  assign n8711 = ( x67 & n8388 ) | ( x67 & ~n8693 ) | ( n8388 & ~n8693 ) ;
  assign n8712 = x67 & n8388 ;
  assign n8713 = ( ~n8393 & n8711 ) | ( ~n8393 & n8712 ) | ( n8711 & n8712 ) ;
  assign n8714 = ( n8393 & n8711 ) | ( n8393 & n8712 ) | ( n8711 & n8712 ) ;
  assign n8715 = ( n8393 & n8713 ) | ( n8393 & ~n8714 ) | ( n8713 & ~n8714 ) ;
  assign n8716 = ( x68 & n8710 ) | ( x68 & ~n8715 ) | ( n8710 & ~n8715 ) ;
  assign n8717 = ( x68 & n8394 ) | ( x68 & ~n8693 ) | ( n8394 & ~n8693 ) ;
  assign n8718 = x68 & n8394 ;
  assign n8719 = ( n8399 & n8717 ) | ( n8399 & n8718 ) | ( n8717 & n8718 ) ;
  assign n8720 = ( ~n8399 & n8717 ) | ( ~n8399 & n8718 ) | ( n8717 & n8718 ) ;
  assign n8721 = ( n8399 & ~n8719 ) | ( n8399 & n8720 ) | ( ~n8719 & n8720 ) ;
  assign n8722 = ( x69 & n8716 ) | ( x69 & ~n8721 ) | ( n8716 & ~n8721 ) ;
  assign n8723 = ( x69 & n8400 ) | ( x69 & ~n8693 ) | ( n8400 & ~n8693 ) ;
  assign n8724 = x69 & n8400 ;
  assign n8725 = ( ~n8405 & n8723 ) | ( ~n8405 & n8724 ) | ( n8723 & n8724 ) ;
  assign n8726 = ( n8405 & n8723 ) | ( n8405 & n8724 ) | ( n8723 & n8724 ) ;
  assign n8727 = ( n8405 & n8725 ) | ( n8405 & ~n8726 ) | ( n8725 & ~n8726 ) ;
  assign n8728 = ( x70 & n8722 ) | ( x70 & ~n8727 ) | ( n8722 & ~n8727 ) ;
  assign n8729 = ( x70 & n8406 ) | ( x70 & ~n8693 ) | ( n8406 & ~n8693 ) ;
  assign n8730 = x70 & n8406 ;
  assign n8731 = ( n8411 & n8729 ) | ( n8411 & n8730 ) | ( n8729 & n8730 ) ;
  assign n8732 = ( ~n8411 & n8729 ) | ( ~n8411 & n8730 ) | ( n8729 & n8730 ) ;
  assign n8733 = ( n8411 & ~n8731 ) | ( n8411 & n8732 ) | ( ~n8731 & n8732 ) ;
  assign n8734 = ( x71 & n8728 ) | ( x71 & ~n8733 ) | ( n8728 & ~n8733 ) ;
  assign n8735 = ( x71 & n8412 ) | ( x71 & ~n8693 ) | ( n8412 & ~n8693 ) ;
  assign n8736 = x71 & n8412 ;
  assign n8737 = ( ~n8417 & n8735 ) | ( ~n8417 & n8736 ) | ( n8735 & n8736 ) ;
  assign n8738 = ( n8417 & n8735 ) | ( n8417 & n8736 ) | ( n8735 & n8736 ) ;
  assign n8739 = ( n8417 & n8737 ) | ( n8417 & ~n8738 ) | ( n8737 & ~n8738 ) ;
  assign n8740 = ( x72 & n8734 ) | ( x72 & ~n8739 ) | ( n8734 & ~n8739 ) ;
  assign n8741 = ( x72 & n8418 ) | ( x72 & ~n8693 ) | ( n8418 & ~n8693 ) ;
  assign n8742 = x72 & n8418 ;
  assign n8743 = ( n8423 & n8741 ) | ( n8423 & n8742 ) | ( n8741 & n8742 ) ;
  assign n8744 = ( ~n8423 & n8741 ) | ( ~n8423 & n8742 ) | ( n8741 & n8742 ) ;
  assign n8745 = ( n8423 & ~n8743 ) | ( n8423 & n8744 ) | ( ~n8743 & n8744 ) ;
  assign n8746 = ( x73 & n8740 ) | ( x73 & ~n8745 ) | ( n8740 & ~n8745 ) ;
  assign n8747 = ( x73 & n8424 ) | ( x73 & ~n8693 ) | ( n8424 & ~n8693 ) ;
  assign n8748 = x73 & n8424 ;
  assign n8749 = ( ~n8429 & n8747 ) | ( ~n8429 & n8748 ) | ( n8747 & n8748 ) ;
  assign n8750 = ( n8429 & n8747 ) | ( n8429 & n8748 ) | ( n8747 & n8748 ) ;
  assign n8751 = ( n8429 & n8749 ) | ( n8429 & ~n8750 ) | ( n8749 & ~n8750 ) ;
  assign n8752 = ( x74 & n8746 ) | ( x74 & ~n8751 ) | ( n8746 & ~n8751 ) ;
  assign n8753 = ( x74 & n8430 ) | ( x74 & ~n8693 ) | ( n8430 & ~n8693 ) ;
  assign n8754 = x74 & n8430 ;
  assign n8755 = ( n8435 & n8753 ) | ( n8435 & n8754 ) | ( n8753 & n8754 ) ;
  assign n8756 = ( ~n8435 & n8753 ) | ( ~n8435 & n8754 ) | ( n8753 & n8754 ) ;
  assign n8757 = ( n8435 & ~n8755 ) | ( n8435 & n8756 ) | ( ~n8755 & n8756 ) ;
  assign n8758 = ( x75 & n8752 ) | ( x75 & ~n8757 ) | ( n8752 & ~n8757 ) ;
  assign n8759 = ( x75 & n8436 ) | ( x75 & ~n8693 ) | ( n8436 & ~n8693 ) ;
  assign n8760 = x75 & n8436 ;
  assign n8761 = ( ~n8441 & n8759 ) | ( ~n8441 & n8760 ) | ( n8759 & n8760 ) ;
  assign n8762 = ( n8441 & n8759 ) | ( n8441 & n8760 ) | ( n8759 & n8760 ) ;
  assign n8763 = ( n8441 & n8761 ) | ( n8441 & ~n8762 ) | ( n8761 & ~n8762 ) ;
  assign n8764 = ( x76 & n8758 ) | ( x76 & ~n8763 ) | ( n8758 & ~n8763 ) ;
  assign n8765 = ( x76 & n8442 ) | ( x76 & ~n8693 ) | ( n8442 & ~n8693 ) ;
  assign n8766 = x76 & n8442 ;
  assign n8767 = ( n8447 & n8765 ) | ( n8447 & n8766 ) | ( n8765 & n8766 ) ;
  assign n8768 = ( ~n8447 & n8765 ) | ( ~n8447 & n8766 ) | ( n8765 & n8766 ) ;
  assign n8769 = ( n8447 & ~n8767 ) | ( n8447 & n8768 ) | ( ~n8767 & n8768 ) ;
  assign n8770 = ( x77 & n8764 ) | ( x77 & ~n8769 ) | ( n8764 & ~n8769 ) ;
  assign n8771 = ( x77 & n8448 ) | ( x77 & ~n8693 ) | ( n8448 & ~n8693 ) ;
  assign n8772 = x77 & n8448 ;
  assign n8773 = ( ~n8453 & n8771 ) | ( ~n8453 & n8772 ) | ( n8771 & n8772 ) ;
  assign n8774 = ( n8453 & n8771 ) | ( n8453 & n8772 ) | ( n8771 & n8772 ) ;
  assign n8775 = ( n8453 & n8773 ) | ( n8453 & ~n8774 ) | ( n8773 & ~n8774 ) ;
  assign n8776 = ( x78 & n8770 ) | ( x78 & ~n8775 ) | ( n8770 & ~n8775 ) ;
  assign n8777 = ( x78 & n8454 ) | ( x78 & ~n8693 ) | ( n8454 & ~n8693 ) ;
  assign n8778 = x78 & n8454 ;
  assign n8779 = ( n8459 & n8777 ) | ( n8459 & n8778 ) | ( n8777 & n8778 ) ;
  assign n8780 = ( ~n8459 & n8777 ) | ( ~n8459 & n8778 ) | ( n8777 & n8778 ) ;
  assign n8781 = ( n8459 & ~n8779 ) | ( n8459 & n8780 ) | ( ~n8779 & n8780 ) ;
  assign n8782 = ( x79 & n8776 ) | ( x79 & ~n8781 ) | ( n8776 & ~n8781 ) ;
  assign n8783 = ( x79 & n8460 ) | ( x79 & ~n8693 ) | ( n8460 & ~n8693 ) ;
  assign n8784 = x79 & n8460 ;
  assign n8785 = ( ~n8465 & n8783 ) | ( ~n8465 & n8784 ) | ( n8783 & n8784 ) ;
  assign n8786 = ( n8465 & n8783 ) | ( n8465 & n8784 ) | ( n8783 & n8784 ) ;
  assign n8787 = ( n8465 & n8785 ) | ( n8465 & ~n8786 ) | ( n8785 & ~n8786 ) ;
  assign n8788 = ( x80 & n8782 ) | ( x80 & ~n8787 ) | ( n8782 & ~n8787 ) ;
  assign n8789 = ( x80 & n8466 ) | ( x80 & ~n8693 ) | ( n8466 & ~n8693 ) ;
  assign n8790 = x80 & n8466 ;
  assign n8791 = ( n8471 & n8789 ) | ( n8471 & n8790 ) | ( n8789 & n8790 ) ;
  assign n8792 = ( ~n8471 & n8789 ) | ( ~n8471 & n8790 ) | ( n8789 & n8790 ) ;
  assign n8793 = ( n8471 & ~n8791 ) | ( n8471 & n8792 ) | ( ~n8791 & n8792 ) ;
  assign n8794 = ( x81 & n8788 ) | ( x81 & ~n8793 ) | ( n8788 & ~n8793 ) ;
  assign n8795 = ( x81 & n8472 ) | ( x81 & ~n8693 ) | ( n8472 & ~n8693 ) ;
  assign n8796 = x81 & n8472 ;
  assign n8797 = ( ~n8477 & n8795 ) | ( ~n8477 & n8796 ) | ( n8795 & n8796 ) ;
  assign n8798 = ( n8477 & n8795 ) | ( n8477 & n8796 ) | ( n8795 & n8796 ) ;
  assign n8799 = ( n8477 & n8797 ) | ( n8477 & ~n8798 ) | ( n8797 & ~n8798 ) ;
  assign n8800 = ( x82 & n8794 ) | ( x82 & ~n8799 ) | ( n8794 & ~n8799 ) ;
  assign n8801 = ( x82 & n8478 ) | ( x82 & ~n8693 ) | ( n8478 & ~n8693 ) ;
  assign n8802 = x82 & n8478 ;
  assign n8803 = ( n8483 & n8801 ) | ( n8483 & n8802 ) | ( n8801 & n8802 ) ;
  assign n8804 = ( ~n8483 & n8801 ) | ( ~n8483 & n8802 ) | ( n8801 & n8802 ) ;
  assign n8805 = ( n8483 & ~n8803 ) | ( n8483 & n8804 ) | ( ~n8803 & n8804 ) ;
  assign n8806 = ( x83 & n8800 ) | ( x83 & ~n8805 ) | ( n8800 & ~n8805 ) ;
  assign n8807 = ( x83 & n8484 ) | ( x83 & ~n8693 ) | ( n8484 & ~n8693 ) ;
  assign n8808 = x83 & n8484 ;
  assign n8809 = ( ~n8489 & n8807 ) | ( ~n8489 & n8808 ) | ( n8807 & n8808 ) ;
  assign n8810 = ( n8489 & n8807 ) | ( n8489 & n8808 ) | ( n8807 & n8808 ) ;
  assign n8811 = ( n8489 & n8809 ) | ( n8489 & ~n8810 ) | ( n8809 & ~n8810 ) ;
  assign n8812 = ( x84 & n8806 ) | ( x84 & ~n8811 ) | ( n8806 & ~n8811 ) ;
  assign n8813 = ( x84 & n8490 ) | ( x84 & ~n8693 ) | ( n8490 & ~n8693 ) ;
  assign n8814 = x84 & n8490 ;
  assign n8815 = ( n8495 & n8813 ) | ( n8495 & n8814 ) | ( n8813 & n8814 ) ;
  assign n8816 = ( ~n8495 & n8813 ) | ( ~n8495 & n8814 ) | ( n8813 & n8814 ) ;
  assign n8817 = ( n8495 & ~n8815 ) | ( n8495 & n8816 ) | ( ~n8815 & n8816 ) ;
  assign n8818 = ( x85 & n8812 ) | ( x85 & ~n8817 ) | ( n8812 & ~n8817 ) ;
  assign n8819 = ( x85 & n8496 ) | ( x85 & ~n8693 ) | ( n8496 & ~n8693 ) ;
  assign n8820 = x85 & n8496 ;
  assign n8821 = ( ~n8501 & n8819 ) | ( ~n8501 & n8820 ) | ( n8819 & n8820 ) ;
  assign n8822 = ( n8501 & n8819 ) | ( n8501 & n8820 ) | ( n8819 & n8820 ) ;
  assign n8823 = ( n8501 & n8821 ) | ( n8501 & ~n8822 ) | ( n8821 & ~n8822 ) ;
  assign n8824 = ( x86 & n8818 ) | ( x86 & ~n8823 ) | ( n8818 & ~n8823 ) ;
  assign n8825 = ( x86 & n8502 ) | ( x86 & ~n8693 ) | ( n8502 & ~n8693 ) ;
  assign n8826 = x86 & n8502 ;
  assign n8827 = ( n8507 & n8825 ) | ( n8507 & n8826 ) | ( n8825 & n8826 ) ;
  assign n8828 = ( ~n8507 & n8825 ) | ( ~n8507 & n8826 ) | ( n8825 & n8826 ) ;
  assign n8829 = ( n8507 & ~n8827 ) | ( n8507 & n8828 ) | ( ~n8827 & n8828 ) ;
  assign n8830 = ( x87 & n8824 ) | ( x87 & ~n8829 ) | ( n8824 & ~n8829 ) ;
  assign n8831 = ( x87 & n8508 ) | ( x87 & ~n8693 ) | ( n8508 & ~n8693 ) ;
  assign n8832 = x87 & n8508 ;
  assign n8833 = ( ~n8513 & n8831 ) | ( ~n8513 & n8832 ) | ( n8831 & n8832 ) ;
  assign n8834 = ( n8513 & n8831 ) | ( n8513 & n8832 ) | ( n8831 & n8832 ) ;
  assign n8835 = ( n8513 & n8833 ) | ( n8513 & ~n8834 ) | ( n8833 & ~n8834 ) ;
  assign n8836 = ( x88 & n8830 ) | ( x88 & ~n8835 ) | ( n8830 & ~n8835 ) ;
  assign n8837 = ( x88 & n8514 ) | ( x88 & ~n8693 ) | ( n8514 & ~n8693 ) ;
  assign n8838 = x88 & n8514 ;
  assign n8839 = ( n8519 & n8837 ) | ( n8519 & n8838 ) | ( n8837 & n8838 ) ;
  assign n8840 = ( ~n8519 & n8837 ) | ( ~n8519 & n8838 ) | ( n8837 & n8838 ) ;
  assign n8841 = ( n8519 & ~n8839 ) | ( n8519 & n8840 ) | ( ~n8839 & n8840 ) ;
  assign n8842 = ( x89 & n8836 ) | ( x89 & ~n8841 ) | ( n8836 & ~n8841 ) ;
  assign n8843 = ( x89 & n8520 ) | ( x89 & ~n8693 ) | ( n8520 & ~n8693 ) ;
  assign n8844 = x89 & n8520 ;
  assign n8845 = ( ~n8525 & n8843 ) | ( ~n8525 & n8844 ) | ( n8843 & n8844 ) ;
  assign n8846 = ( n8525 & n8843 ) | ( n8525 & n8844 ) | ( n8843 & n8844 ) ;
  assign n8847 = ( n8525 & n8845 ) | ( n8525 & ~n8846 ) | ( n8845 & ~n8846 ) ;
  assign n8848 = ( x90 & n8842 ) | ( x90 & ~n8847 ) | ( n8842 & ~n8847 ) ;
  assign n8849 = ( x90 & n8526 ) | ( x90 & ~n8693 ) | ( n8526 & ~n8693 ) ;
  assign n8850 = x90 & n8526 ;
  assign n8851 = ( n8531 & n8849 ) | ( n8531 & n8850 ) | ( n8849 & n8850 ) ;
  assign n8852 = ( ~n8531 & n8849 ) | ( ~n8531 & n8850 ) | ( n8849 & n8850 ) ;
  assign n8853 = ( n8531 & ~n8851 ) | ( n8531 & n8852 ) | ( ~n8851 & n8852 ) ;
  assign n8854 = ( x91 & n8848 ) | ( x91 & ~n8853 ) | ( n8848 & ~n8853 ) ;
  assign n8855 = ( x91 & n8532 ) | ( x91 & ~n8693 ) | ( n8532 & ~n8693 ) ;
  assign n8856 = x91 & n8532 ;
  assign n8857 = ( ~n8537 & n8855 ) | ( ~n8537 & n8856 ) | ( n8855 & n8856 ) ;
  assign n8858 = ( n8537 & n8855 ) | ( n8537 & n8856 ) | ( n8855 & n8856 ) ;
  assign n8859 = ( n8537 & n8857 ) | ( n8537 & ~n8858 ) | ( n8857 & ~n8858 ) ;
  assign n8860 = ( x92 & n8854 ) | ( x92 & ~n8859 ) | ( n8854 & ~n8859 ) ;
  assign n8861 = ( x92 & n8538 ) | ( x92 & ~n8693 ) | ( n8538 & ~n8693 ) ;
  assign n8862 = x92 & n8538 ;
  assign n8863 = ( n8543 & n8861 ) | ( n8543 & n8862 ) | ( n8861 & n8862 ) ;
  assign n8864 = ( ~n8543 & n8861 ) | ( ~n8543 & n8862 ) | ( n8861 & n8862 ) ;
  assign n8865 = ( n8543 & ~n8863 ) | ( n8543 & n8864 ) | ( ~n8863 & n8864 ) ;
  assign n8866 = ( x93 & n8860 ) | ( x93 & ~n8865 ) | ( n8860 & ~n8865 ) ;
  assign n8867 = ( x93 & n8544 ) | ( x93 & ~n8693 ) | ( n8544 & ~n8693 ) ;
  assign n8868 = x93 & n8544 ;
  assign n8869 = ( ~n8549 & n8867 ) | ( ~n8549 & n8868 ) | ( n8867 & n8868 ) ;
  assign n8870 = ( n8549 & n8867 ) | ( n8549 & n8868 ) | ( n8867 & n8868 ) ;
  assign n8871 = ( n8549 & n8869 ) | ( n8549 & ~n8870 ) | ( n8869 & ~n8870 ) ;
  assign n8872 = ( x94 & n8866 ) | ( x94 & ~n8871 ) | ( n8866 & ~n8871 ) ;
  assign n8873 = ( x94 & n8550 ) | ( x94 & ~n8693 ) | ( n8550 & ~n8693 ) ;
  assign n8874 = x94 & n8550 ;
  assign n8875 = ( n8555 & n8873 ) | ( n8555 & n8874 ) | ( n8873 & n8874 ) ;
  assign n8876 = ( ~n8555 & n8873 ) | ( ~n8555 & n8874 ) | ( n8873 & n8874 ) ;
  assign n8877 = ( n8555 & ~n8875 ) | ( n8555 & n8876 ) | ( ~n8875 & n8876 ) ;
  assign n8878 = ( x95 & n8872 ) | ( x95 & ~n8877 ) | ( n8872 & ~n8877 ) ;
  assign n8879 = ( x95 & n8556 ) | ( x95 & ~n8693 ) | ( n8556 & ~n8693 ) ;
  assign n8880 = x95 & n8556 ;
  assign n8881 = ( ~n8561 & n8879 ) | ( ~n8561 & n8880 ) | ( n8879 & n8880 ) ;
  assign n8882 = ( n8561 & n8879 ) | ( n8561 & n8880 ) | ( n8879 & n8880 ) ;
  assign n8883 = ( n8561 & n8881 ) | ( n8561 & ~n8882 ) | ( n8881 & ~n8882 ) ;
  assign n8884 = ( x96 & n8878 ) | ( x96 & ~n8883 ) | ( n8878 & ~n8883 ) ;
  assign n8885 = ( x96 & n8562 ) | ( x96 & ~n8693 ) | ( n8562 & ~n8693 ) ;
  assign n8886 = x96 & n8562 ;
  assign n8887 = ( n8567 & n8885 ) | ( n8567 & n8886 ) | ( n8885 & n8886 ) ;
  assign n8888 = ( ~n8567 & n8885 ) | ( ~n8567 & n8886 ) | ( n8885 & n8886 ) ;
  assign n8889 = ( n8567 & ~n8887 ) | ( n8567 & n8888 ) | ( ~n8887 & n8888 ) ;
  assign n8890 = ( x97 & n8884 ) | ( x97 & ~n8889 ) | ( n8884 & ~n8889 ) ;
  assign n8891 = ( x97 & n8568 ) | ( x97 & ~n8693 ) | ( n8568 & ~n8693 ) ;
  assign n8892 = x97 & n8568 ;
  assign n8893 = ( ~n8573 & n8891 ) | ( ~n8573 & n8892 ) | ( n8891 & n8892 ) ;
  assign n8894 = ( n8573 & n8891 ) | ( n8573 & n8892 ) | ( n8891 & n8892 ) ;
  assign n8895 = ( n8573 & n8893 ) | ( n8573 & ~n8894 ) | ( n8893 & ~n8894 ) ;
  assign n8896 = ( x98 & n8890 ) | ( x98 & ~n8895 ) | ( n8890 & ~n8895 ) ;
  assign n8897 = ( x98 & n8574 ) | ( x98 & ~n8693 ) | ( n8574 & ~n8693 ) ;
  assign n8898 = x98 & n8574 ;
  assign n8899 = ( n8579 & n8897 ) | ( n8579 & n8898 ) | ( n8897 & n8898 ) ;
  assign n8900 = ( ~n8579 & n8897 ) | ( ~n8579 & n8898 ) | ( n8897 & n8898 ) ;
  assign n8901 = ( n8579 & ~n8899 ) | ( n8579 & n8900 ) | ( ~n8899 & n8900 ) ;
  assign n8902 = ( x99 & n8896 ) | ( x99 & ~n8901 ) | ( n8896 & ~n8901 ) ;
  assign n8903 = ( x99 & n8580 ) | ( x99 & ~n8693 ) | ( n8580 & ~n8693 ) ;
  assign n8904 = x99 & n8580 ;
  assign n8905 = ( ~n8585 & n8903 ) | ( ~n8585 & n8904 ) | ( n8903 & n8904 ) ;
  assign n8906 = ( n8585 & n8903 ) | ( n8585 & n8904 ) | ( n8903 & n8904 ) ;
  assign n8907 = ( n8585 & n8905 ) | ( n8585 & ~n8906 ) | ( n8905 & ~n8906 ) ;
  assign n8908 = ( x100 & n8902 ) | ( x100 & ~n8907 ) | ( n8902 & ~n8907 ) ;
  assign n8909 = ( x100 & n8586 ) | ( x100 & ~n8693 ) | ( n8586 & ~n8693 ) ;
  assign n8910 = x100 & n8586 ;
  assign n8911 = ( n8591 & n8909 ) | ( n8591 & n8910 ) | ( n8909 & n8910 ) ;
  assign n8912 = ( ~n8591 & n8909 ) | ( ~n8591 & n8910 ) | ( n8909 & n8910 ) ;
  assign n8913 = ( n8591 & ~n8911 ) | ( n8591 & n8912 ) | ( ~n8911 & n8912 ) ;
  assign n8914 = ( x101 & n8908 ) | ( x101 & ~n8913 ) | ( n8908 & ~n8913 ) ;
  assign n8915 = ( x101 & n8592 ) | ( x101 & ~n8693 ) | ( n8592 & ~n8693 ) ;
  assign n8916 = x101 & n8592 ;
  assign n8917 = ( ~n8597 & n8915 ) | ( ~n8597 & n8916 ) | ( n8915 & n8916 ) ;
  assign n8918 = ( n8597 & n8915 ) | ( n8597 & n8916 ) | ( n8915 & n8916 ) ;
  assign n8919 = ( n8597 & n8917 ) | ( n8597 & ~n8918 ) | ( n8917 & ~n8918 ) ;
  assign n8920 = ( x102 & n8914 ) | ( x102 & ~n8919 ) | ( n8914 & ~n8919 ) ;
  assign n8921 = ( x102 & n8598 ) | ( x102 & ~n8693 ) | ( n8598 & ~n8693 ) ;
  assign n8922 = x102 & n8598 ;
  assign n8923 = ( n8603 & n8921 ) | ( n8603 & n8922 ) | ( n8921 & n8922 ) ;
  assign n8924 = ( ~n8603 & n8921 ) | ( ~n8603 & n8922 ) | ( n8921 & n8922 ) ;
  assign n8925 = ( n8603 & ~n8923 ) | ( n8603 & n8924 ) | ( ~n8923 & n8924 ) ;
  assign n8926 = ( x103 & n8920 ) | ( x103 & ~n8925 ) | ( n8920 & ~n8925 ) ;
  assign n8927 = ( x103 & n8604 ) | ( x103 & ~n8693 ) | ( n8604 & ~n8693 ) ;
  assign n8928 = x103 & n8604 ;
  assign n8929 = ( ~n8609 & n8927 ) | ( ~n8609 & n8928 ) | ( n8927 & n8928 ) ;
  assign n8930 = ( n8609 & n8927 ) | ( n8609 & n8928 ) | ( n8927 & n8928 ) ;
  assign n8931 = ( n8609 & n8929 ) | ( n8609 & ~n8930 ) | ( n8929 & ~n8930 ) ;
  assign n8932 = ( x104 & n8926 ) | ( x104 & ~n8931 ) | ( n8926 & ~n8931 ) ;
  assign n8933 = ( x104 & n8610 ) | ( x104 & ~n8693 ) | ( n8610 & ~n8693 ) ;
  assign n8934 = x104 & n8610 ;
  assign n8935 = ( n8615 & n8933 ) | ( n8615 & n8934 ) | ( n8933 & n8934 ) ;
  assign n8936 = ( ~n8615 & n8933 ) | ( ~n8615 & n8934 ) | ( n8933 & n8934 ) ;
  assign n8937 = ( n8615 & ~n8935 ) | ( n8615 & n8936 ) | ( ~n8935 & n8936 ) ;
  assign n8938 = ( x105 & n8932 ) | ( x105 & ~n8937 ) | ( n8932 & ~n8937 ) ;
  assign n8939 = ( x105 & n8616 ) | ( x105 & ~n8693 ) | ( n8616 & ~n8693 ) ;
  assign n8940 = x105 & n8616 ;
  assign n8941 = ( ~n8621 & n8939 ) | ( ~n8621 & n8940 ) | ( n8939 & n8940 ) ;
  assign n8942 = ( n8621 & n8939 ) | ( n8621 & n8940 ) | ( n8939 & n8940 ) ;
  assign n8943 = ( n8621 & n8941 ) | ( n8621 & ~n8942 ) | ( n8941 & ~n8942 ) ;
  assign n8944 = ( x106 & n8938 ) | ( x106 & ~n8943 ) | ( n8938 & ~n8943 ) ;
  assign n8945 = ( x106 & n8622 ) | ( x106 & ~n8693 ) | ( n8622 & ~n8693 ) ;
  assign n8946 = x106 & n8622 ;
  assign n8947 = ( n8627 & n8945 ) | ( n8627 & n8946 ) | ( n8945 & n8946 ) ;
  assign n8948 = ( ~n8627 & n8945 ) | ( ~n8627 & n8946 ) | ( n8945 & n8946 ) ;
  assign n8949 = ( n8627 & ~n8947 ) | ( n8627 & n8948 ) | ( ~n8947 & n8948 ) ;
  assign n8950 = ( x107 & n8944 ) | ( x107 & ~n8949 ) | ( n8944 & ~n8949 ) ;
  assign n8951 = ( x107 & n8628 ) | ( x107 & ~n8693 ) | ( n8628 & ~n8693 ) ;
  assign n8952 = x107 & n8628 ;
  assign n8953 = ( ~n8633 & n8951 ) | ( ~n8633 & n8952 ) | ( n8951 & n8952 ) ;
  assign n8954 = ( n8633 & n8951 ) | ( n8633 & n8952 ) | ( n8951 & n8952 ) ;
  assign n8955 = ( n8633 & n8953 ) | ( n8633 & ~n8954 ) | ( n8953 & ~n8954 ) ;
  assign n8956 = ( x108 & n8950 ) | ( x108 & ~n8955 ) | ( n8950 & ~n8955 ) ;
  assign n8957 = ( x108 & n8634 ) | ( x108 & ~n8693 ) | ( n8634 & ~n8693 ) ;
  assign n8958 = x108 & n8634 ;
  assign n8959 = ( n8639 & n8957 ) | ( n8639 & n8958 ) | ( n8957 & n8958 ) ;
  assign n8960 = ( ~n8639 & n8957 ) | ( ~n8639 & n8958 ) | ( n8957 & n8958 ) ;
  assign n8961 = ( n8639 & ~n8959 ) | ( n8639 & n8960 ) | ( ~n8959 & n8960 ) ;
  assign n8962 = ( x109 & n8956 ) | ( x109 & ~n8961 ) | ( n8956 & ~n8961 ) ;
  assign n8963 = ( x109 & n8640 ) | ( x109 & ~n8693 ) | ( n8640 & ~n8693 ) ;
  assign n8964 = x109 & n8640 ;
  assign n8965 = ( ~n8645 & n8963 ) | ( ~n8645 & n8964 ) | ( n8963 & n8964 ) ;
  assign n8966 = ( n8645 & n8963 ) | ( n8645 & n8964 ) | ( n8963 & n8964 ) ;
  assign n8967 = ( n8645 & n8965 ) | ( n8645 & ~n8966 ) | ( n8965 & ~n8966 ) ;
  assign n8968 = ( x110 & n8962 ) | ( x110 & ~n8967 ) | ( n8962 & ~n8967 ) ;
  assign n8969 = ( x110 & n8646 ) | ( x110 & ~n8693 ) | ( n8646 & ~n8693 ) ;
  assign n8970 = x110 & n8646 ;
  assign n8971 = ( n8651 & n8969 ) | ( n8651 & n8970 ) | ( n8969 & n8970 ) ;
  assign n8972 = ( ~n8651 & n8969 ) | ( ~n8651 & n8970 ) | ( n8969 & n8970 ) ;
  assign n8973 = ( n8651 & ~n8971 ) | ( n8651 & n8972 ) | ( ~n8971 & n8972 ) ;
  assign n8974 = ( x111 & n8968 ) | ( x111 & ~n8973 ) | ( n8968 & ~n8973 ) ;
  assign n8975 = ( x111 & n8652 ) | ( x111 & ~n8693 ) | ( n8652 & ~n8693 ) ;
  assign n8976 = x111 & n8652 ;
  assign n8977 = ( ~n8657 & n8975 ) | ( ~n8657 & n8976 ) | ( n8975 & n8976 ) ;
  assign n8978 = ( n8657 & n8975 ) | ( n8657 & n8976 ) | ( n8975 & n8976 ) ;
  assign n8979 = ( n8657 & n8977 ) | ( n8657 & ~n8978 ) | ( n8977 & ~n8978 ) ;
  assign n8980 = ( x112 & n8974 ) | ( x112 & ~n8979 ) | ( n8974 & ~n8979 ) ;
  assign n8981 = ( x112 & n8658 ) | ( x112 & ~n8693 ) | ( n8658 & ~n8693 ) ;
  assign n8982 = x112 & n8658 ;
  assign n8983 = ( n8663 & n8981 ) | ( n8663 & n8982 ) | ( n8981 & n8982 ) ;
  assign n8984 = ( ~n8663 & n8981 ) | ( ~n8663 & n8982 ) | ( n8981 & n8982 ) ;
  assign n8985 = ( n8663 & ~n8983 ) | ( n8663 & n8984 ) | ( ~n8983 & n8984 ) ;
  assign n8986 = ( x113 & n8980 ) | ( x113 & ~n8985 ) | ( n8980 & ~n8985 ) ;
  assign n8987 = ( x113 & n8664 ) | ( x113 & ~n8693 ) | ( n8664 & ~n8693 ) ;
  assign n8988 = x113 & n8664 ;
  assign n8989 = ( ~n8669 & n8987 ) | ( ~n8669 & n8988 ) | ( n8987 & n8988 ) ;
  assign n8990 = ( n8669 & n8987 ) | ( n8669 & n8988 ) | ( n8987 & n8988 ) ;
  assign n8991 = ( n8669 & n8989 ) | ( n8669 & ~n8990 ) | ( n8989 & ~n8990 ) ;
  assign n8992 = ( x114 & n8986 ) | ( x114 & ~n8991 ) | ( n8986 & ~n8991 ) ;
  assign n8993 = ( x114 & n8670 ) | ( x114 & ~n8693 ) | ( n8670 & ~n8693 ) ;
  assign n8994 = x114 & n8670 ;
  assign n8995 = ( n8675 & n8993 ) | ( n8675 & n8994 ) | ( n8993 & n8994 ) ;
  assign n8996 = ( ~n8675 & n8993 ) | ( ~n8675 & n8994 ) | ( n8993 & n8994 ) ;
  assign n8997 = ( n8675 & ~n8995 ) | ( n8675 & n8996 ) | ( ~n8995 & n8996 ) ;
  assign n8998 = ( x115 & n8992 ) | ( x115 & ~n8997 ) | ( n8992 & ~n8997 ) ;
  assign n8999 = ( x115 & n8676 ) | ( x115 & ~n8693 ) | ( n8676 & ~n8693 ) ;
  assign n9000 = x115 & n8676 ;
  assign n9001 = ( ~n8681 & n8999 ) | ( ~n8681 & n9000 ) | ( n8999 & n9000 ) ;
  assign n9002 = ( n8681 & n8999 ) | ( n8681 & n9000 ) | ( n8999 & n9000 ) ;
  assign n9003 = ( n8681 & n9001 ) | ( n8681 & ~n9002 ) | ( n9001 & ~n9002 ) ;
  assign n9004 = ( x116 & n8998 ) | ( x116 & ~n9003 ) | ( n8998 & ~n9003 ) ;
  assign n9005 = ( x116 & n8682 ) | ( x116 & ~n8693 ) | ( n8682 & ~n8693 ) ;
  assign n9006 = x116 & n8682 ;
  assign n9007 = ( ~n8687 & n9005 ) | ( ~n8687 & n9006 ) | ( n9005 & n9006 ) ;
  assign n9008 = ( n8687 & n9005 ) | ( n8687 & n9006 ) | ( n9005 & n9006 ) ;
  assign n9009 = ( n8687 & n9007 ) | ( n8687 & ~n9008 ) | ( n9007 & ~n9008 ) ;
  assign n9010 = ( x117 & n9004 ) | ( x117 & ~n9009 ) | ( n9004 & ~n9009 ) ;
  assign n9011 = x118 | n9010 ;
  assign n9012 = ( x118 & n139 ) | ( x118 & n9010 ) | ( n139 & n9010 ) ;
  assign n9013 = ( n8691 & ~n9011 ) | ( n8691 & n9012 ) | ( ~n9011 & n9012 ) ;
  assign n9014 = ( x118 & ~n8691 ) | ( x118 & n9010 ) | ( ~n8691 & n9010 ) ;
  assign n9015 = n139 | n9014 ;
  assign n9016 = ( x9 & ~x64 ) | ( x9 & n9015 ) | ( ~x64 & n9015 ) ;
  assign n9017 = ~x9 & n9015 ;
  assign n9018 = ( n8697 & n9016 ) | ( n8697 & ~n9017 ) | ( n9016 & ~n9017 ) ;
  assign n9019 = ~x8 & x64 ;
  assign n9020 = ( x65 & ~n9018 ) | ( x65 & n9019 ) | ( ~n9018 & n9019 ) ;
  assign n9021 = ( x65 & n8697 ) | ( x65 & ~n9015 ) | ( n8697 & ~n9015 ) ;
  assign n9022 = x65 & n8697 ;
  assign n9023 = ( n8696 & n9021 ) | ( n8696 & n9022 ) | ( n9021 & n9022 ) ;
  assign n9024 = ( ~n8696 & n9021 ) | ( ~n8696 & n9022 ) | ( n9021 & n9022 ) ;
  assign n9025 = ( n8696 & ~n9023 ) | ( n8696 & n9024 ) | ( ~n9023 & n9024 ) ;
  assign n9026 = ( x66 & n9020 ) | ( x66 & ~n9025 ) | ( n9020 & ~n9025 ) ;
  assign n9027 = ( x66 & n8698 ) | ( x66 & ~n9015 ) | ( n8698 & ~n9015 ) ;
  assign n9028 = x66 & n8698 ;
  assign n9029 = ( n8703 & n9027 ) | ( n8703 & n9028 ) | ( n9027 & n9028 ) ;
  assign n9030 = ( ~n8703 & n9027 ) | ( ~n8703 & n9028 ) | ( n9027 & n9028 ) ;
  assign n9031 = ( n8703 & ~n9029 ) | ( n8703 & n9030 ) | ( ~n9029 & n9030 ) ;
  assign n9032 = ( x67 & n9026 ) | ( x67 & ~n9031 ) | ( n9026 & ~n9031 ) ;
  assign n9033 = ( x67 & n8704 ) | ( x67 & ~n9015 ) | ( n8704 & ~n9015 ) ;
  assign n9034 = x67 & n8704 ;
  assign n9035 = ( ~n8709 & n9033 ) | ( ~n8709 & n9034 ) | ( n9033 & n9034 ) ;
  assign n9036 = ( n8709 & n9033 ) | ( n8709 & n9034 ) | ( n9033 & n9034 ) ;
  assign n9037 = ( n8709 & n9035 ) | ( n8709 & ~n9036 ) | ( n9035 & ~n9036 ) ;
  assign n9038 = ( x68 & n9032 ) | ( x68 & ~n9037 ) | ( n9032 & ~n9037 ) ;
  assign n9039 = ( x68 & n8710 ) | ( x68 & ~n9015 ) | ( n8710 & ~n9015 ) ;
  assign n9040 = x68 & n8710 ;
  assign n9041 = ( n8715 & n9039 ) | ( n8715 & n9040 ) | ( n9039 & n9040 ) ;
  assign n9042 = ( ~n8715 & n9039 ) | ( ~n8715 & n9040 ) | ( n9039 & n9040 ) ;
  assign n9043 = ( n8715 & ~n9041 ) | ( n8715 & n9042 ) | ( ~n9041 & n9042 ) ;
  assign n9044 = ( x69 & n9038 ) | ( x69 & ~n9043 ) | ( n9038 & ~n9043 ) ;
  assign n9045 = ( x69 & n8716 ) | ( x69 & ~n9015 ) | ( n8716 & ~n9015 ) ;
  assign n9046 = x69 & n8716 ;
  assign n9047 = ( ~n8721 & n9045 ) | ( ~n8721 & n9046 ) | ( n9045 & n9046 ) ;
  assign n9048 = ( n8721 & n9045 ) | ( n8721 & n9046 ) | ( n9045 & n9046 ) ;
  assign n9049 = ( n8721 & n9047 ) | ( n8721 & ~n9048 ) | ( n9047 & ~n9048 ) ;
  assign n9050 = ( x70 & n9044 ) | ( x70 & ~n9049 ) | ( n9044 & ~n9049 ) ;
  assign n9051 = ( x70 & n8722 ) | ( x70 & ~n9015 ) | ( n8722 & ~n9015 ) ;
  assign n9052 = x70 & n8722 ;
  assign n9053 = ( n8727 & n9051 ) | ( n8727 & n9052 ) | ( n9051 & n9052 ) ;
  assign n9054 = ( ~n8727 & n9051 ) | ( ~n8727 & n9052 ) | ( n9051 & n9052 ) ;
  assign n9055 = ( n8727 & ~n9053 ) | ( n8727 & n9054 ) | ( ~n9053 & n9054 ) ;
  assign n9056 = ( x71 & n9050 ) | ( x71 & ~n9055 ) | ( n9050 & ~n9055 ) ;
  assign n9057 = ( x71 & n8728 ) | ( x71 & ~n9015 ) | ( n8728 & ~n9015 ) ;
  assign n9058 = x71 & n8728 ;
  assign n9059 = ( ~n8733 & n9057 ) | ( ~n8733 & n9058 ) | ( n9057 & n9058 ) ;
  assign n9060 = ( n8733 & n9057 ) | ( n8733 & n9058 ) | ( n9057 & n9058 ) ;
  assign n9061 = ( n8733 & n9059 ) | ( n8733 & ~n9060 ) | ( n9059 & ~n9060 ) ;
  assign n9062 = ( x72 & n9056 ) | ( x72 & ~n9061 ) | ( n9056 & ~n9061 ) ;
  assign n9063 = ( x72 & n8734 ) | ( x72 & ~n9015 ) | ( n8734 & ~n9015 ) ;
  assign n9064 = x72 & n8734 ;
  assign n9065 = ( n8739 & n9063 ) | ( n8739 & n9064 ) | ( n9063 & n9064 ) ;
  assign n9066 = ( ~n8739 & n9063 ) | ( ~n8739 & n9064 ) | ( n9063 & n9064 ) ;
  assign n9067 = ( n8739 & ~n9065 ) | ( n8739 & n9066 ) | ( ~n9065 & n9066 ) ;
  assign n9068 = ( x73 & n9062 ) | ( x73 & ~n9067 ) | ( n9062 & ~n9067 ) ;
  assign n9069 = ( x73 & n8740 ) | ( x73 & ~n9015 ) | ( n8740 & ~n9015 ) ;
  assign n9070 = x73 & n8740 ;
  assign n9071 = ( ~n8745 & n9069 ) | ( ~n8745 & n9070 ) | ( n9069 & n9070 ) ;
  assign n9072 = ( n8745 & n9069 ) | ( n8745 & n9070 ) | ( n9069 & n9070 ) ;
  assign n9073 = ( n8745 & n9071 ) | ( n8745 & ~n9072 ) | ( n9071 & ~n9072 ) ;
  assign n9074 = ( x74 & n9068 ) | ( x74 & ~n9073 ) | ( n9068 & ~n9073 ) ;
  assign n9075 = ( x74 & n8746 ) | ( x74 & ~n9015 ) | ( n8746 & ~n9015 ) ;
  assign n9076 = x74 & n8746 ;
  assign n9077 = ( n8751 & n9075 ) | ( n8751 & n9076 ) | ( n9075 & n9076 ) ;
  assign n9078 = ( ~n8751 & n9075 ) | ( ~n8751 & n9076 ) | ( n9075 & n9076 ) ;
  assign n9079 = ( n8751 & ~n9077 ) | ( n8751 & n9078 ) | ( ~n9077 & n9078 ) ;
  assign n9080 = ( x75 & n9074 ) | ( x75 & ~n9079 ) | ( n9074 & ~n9079 ) ;
  assign n9081 = ( x75 & n8752 ) | ( x75 & ~n9015 ) | ( n8752 & ~n9015 ) ;
  assign n9082 = x75 & n8752 ;
  assign n9083 = ( ~n8757 & n9081 ) | ( ~n8757 & n9082 ) | ( n9081 & n9082 ) ;
  assign n9084 = ( n8757 & n9081 ) | ( n8757 & n9082 ) | ( n9081 & n9082 ) ;
  assign n9085 = ( n8757 & n9083 ) | ( n8757 & ~n9084 ) | ( n9083 & ~n9084 ) ;
  assign n9086 = ( x76 & n9080 ) | ( x76 & ~n9085 ) | ( n9080 & ~n9085 ) ;
  assign n9087 = ( x76 & n8758 ) | ( x76 & ~n9015 ) | ( n8758 & ~n9015 ) ;
  assign n9088 = x76 & n8758 ;
  assign n9089 = ( n8763 & n9087 ) | ( n8763 & n9088 ) | ( n9087 & n9088 ) ;
  assign n9090 = ( ~n8763 & n9087 ) | ( ~n8763 & n9088 ) | ( n9087 & n9088 ) ;
  assign n9091 = ( n8763 & ~n9089 ) | ( n8763 & n9090 ) | ( ~n9089 & n9090 ) ;
  assign n9092 = ( x77 & n9086 ) | ( x77 & ~n9091 ) | ( n9086 & ~n9091 ) ;
  assign n9093 = ( x77 & n8764 ) | ( x77 & ~n9015 ) | ( n8764 & ~n9015 ) ;
  assign n9094 = x77 & n8764 ;
  assign n9095 = ( ~n8769 & n9093 ) | ( ~n8769 & n9094 ) | ( n9093 & n9094 ) ;
  assign n9096 = ( n8769 & n9093 ) | ( n8769 & n9094 ) | ( n9093 & n9094 ) ;
  assign n9097 = ( n8769 & n9095 ) | ( n8769 & ~n9096 ) | ( n9095 & ~n9096 ) ;
  assign n9098 = ( x78 & n9092 ) | ( x78 & ~n9097 ) | ( n9092 & ~n9097 ) ;
  assign n9099 = ( x78 & n8770 ) | ( x78 & ~n9015 ) | ( n8770 & ~n9015 ) ;
  assign n9100 = x78 & n8770 ;
  assign n9101 = ( n8775 & n9099 ) | ( n8775 & n9100 ) | ( n9099 & n9100 ) ;
  assign n9102 = ( ~n8775 & n9099 ) | ( ~n8775 & n9100 ) | ( n9099 & n9100 ) ;
  assign n9103 = ( n8775 & ~n9101 ) | ( n8775 & n9102 ) | ( ~n9101 & n9102 ) ;
  assign n9104 = ( x79 & n9098 ) | ( x79 & ~n9103 ) | ( n9098 & ~n9103 ) ;
  assign n9105 = ( x79 & n8776 ) | ( x79 & ~n9015 ) | ( n8776 & ~n9015 ) ;
  assign n9106 = x79 & n8776 ;
  assign n9107 = ( ~n8781 & n9105 ) | ( ~n8781 & n9106 ) | ( n9105 & n9106 ) ;
  assign n9108 = ( n8781 & n9105 ) | ( n8781 & n9106 ) | ( n9105 & n9106 ) ;
  assign n9109 = ( n8781 & n9107 ) | ( n8781 & ~n9108 ) | ( n9107 & ~n9108 ) ;
  assign n9110 = ( x80 & n9104 ) | ( x80 & ~n9109 ) | ( n9104 & ~n9109 ) ;
  assign n9111 = ( x80 & n8782 ) | ( x80 & ~n9015 ) | ( n8782 & ~n9015 ) ;
  assign n9112 = x80 & n8782 ;
  assign n9113 = ( n8787 & n9111 ) | ( n8787 & n9112 ) | ( n9111 & n9112 ) ;
  assign n9114 = ( ~n8787 & n9111 ) | ( ~n8787 & n9112 ) | ( n9111 & n9112 ) ;
  assign n9115 = ( n8787 & ~n9113 ) | ( n8787 & n9114 ) | ( ~n9113 & n9114 ) ;
  assign n9116 = ( x81 & n9110 ) | ( x81 & ~n9115 ) | ( n9110 & ~n9115 ) ;
  assign n9117 = ( x81 & n8788 ) | ( x81 & ~n9015 ) | ( n8788 & ~n9015 ) ;
  assign n9118 = x81 & n8788 ;
  assign n9119 = ( ~n8793 & n9117 ) | ( ~n8793 & n9118 ) | ( n9117 & n9118 ) ;
  assign n9120 = ( n8793 & n9117 ) | ( n8793 & n9118 ) | ( n9117 & n9118 ) ;
  assign n9121 = ( n8793 & n9119 ) | ( n8793 & ~n9120 ) | ( n9119 & ~n9120 ) ;
  assign n9122 = ( x82 & n9116 ) | ( x82 & ~n9121 ) | ( n9116 & ~n9121 ) ;
  assign n9123 = ( x82 & n8794 ) | ( x82 & ~n9015 ) | ( n8794 & ~n9015 ) ;
  assign n9124 = x82 & n8794 ;
  assign n9125 = ( n8799 & n9123 ) | ( n8799 & n9124 ) | ( n9123 & n9124 ) ;
  assign n9126 = ( ~n8799 & n9123 ) | ( ~n8799 & n9124 ) | ( n9123 & n9124 ) ;
  assign n9127 = ( n8799 & ~n9125 ) | ( n8799 & n9126 ) | ( ~n9125 & n9126 ) ;
  assign n9128 = ( x83 & n9122 ) | ( x83 & ~n9127 ) | ( n9122 & ~n9127 ) ;
  assign n9129 = ( x83 & n8800 ) | ( x83 & ~n9015 ) | ( n8800 & ~n9015 ) ;
  assign n9130 = x83 & n8800 ;
  assign n9131 = ( ~n8805 & n9129 ) | ( ~n8805 & n9130 ) | ( n9129 & n9130 ) ;
  assign n9132 = ( n8805 & n9129 ) | ( n8805 & n9130 ) | ( n9129 & n9130 ) ;
  assign n9133 = ( n8805 & n9131 ) | ( n8805 & ~n9132 ) | ( n9131 & ~n9132 ) ;
  assign n9134 = ( x84 & n9128 ) | ( x84 & ~n9133 ) | ( n9128 & ~n9133 ) ;
  assign n9135 = ( x84 & n8806 ) | ( x84 & ~n9015 ) | ( n8806 & ~n9015 ) ;
  assign n9136 = x84 & n8806 ;
  assign n9137 = ( n8811 & n9135 ) | ( n8811 & n9136 ) | ( n9135 & n9136 ) ;
  assign n9138 = ( ~n8811 & n9135 ) | ( ~n8811 & n9136 ) | ( n9135 & n9136 ) ;
  assign n9139 = ( n8811 & ~n9137 ) | ( n8811 & n9138 ) | ( ~n9137 & n9138 ) ;
  assign n9140 = ( x85 & n9134 ) | ( x85 & ~n9139 ) | ( n9134 & ~n9139 ) ;
  assign n9141 = ( x85 & n8812 ) | ( x85 & ~n9015 ) | ( n8812 & ~n9015 ) ;
  assign n9142 = x85 & n8812 ;
  assign n9143 = ( ~n8817 & n9141 ) | ( ~n8817 & n9142 ) | ( n9141 & n9142 ) ;
  assign n9144 = ( n8817 & n9141 ) | ( n8817 & n9142 ) | ( n9141 & n9142 ) ;
  assign n9145 = ( n8817 & n9143 ) | ( n8817 & ~n9144 ) | ( n9143 & ~n9144 ) ;
  assign n9146 = ( x86 & n9140 ) | ( x86 & ~n9145 ) | ( n9140 & ~n9145 ) ;
  assign n9147 = ( x86 & n8818 ) | ( x86 & ~n9015 ) | ( n8818 & ~n9015 ) ;
  assign n9148 = x86 & n8818 ;
  assign n9149 = ( n8823 & n9147 ) | ( n8823 & n9148 ) | ( n9147 & n9148 ) ;
  assign n9150 = ( ~n8823 & n9147 ) | ( ~n8823 & n9148 ) | ( n9147 & n9148 ) ;
  assign n9151 = ( n8823 & ~n9149 ) | ( n8823 & n9150 ) | ( ~n9149 & n9150 ) ;
  assign n9152 = ( x87 & n9146 ) | ( x87 & ~n9151 ) | ( n9146 & ~n9151 ) ;
  assign n9153 = ( x87 & n8824 ) | ( x87 & ~n9015 ) | ( n8824 & ~n9015 ) ;
  assign n9154 = x87 & n8824 ;
  assign n9155 = ( ~n8829 & n9153 ) | ( ~n8829 & n9154 ) | ( n9153 & n9154 ) ;
  assign n9156 = ( n8829 & n9153 ) | ( n8829 & n9154 ) | ( n9153 & n9154 ) ;
  assign n9157 = ( n8829 & n9155 ) | ( n8829 & ~n9156 ) | ( n9155 & ~n9156 ) ;
  assign n9158 = ( x88 & n9152 ) | ( x88 & ~n9157 ) | ( n9152 & ~n9157 ) ;
  assign n9159 = ( x88 & n8830 ) | ( x88 & ~n9015 ) | ( n8830 & ~n9015 ) ;
  assign n9160 = x88 & n8830 ;
  assign n9161 = ( n8835 & n9159 ) | ( n8835 & n9160 ) | ( n9159 & n9160 ) ;
  assign n9162 = ( ~n8835 & n9159 ) | ( ~n8835 & n9160 ) | ( n9159 & n9160 ) ;
  assign n9163 = ( n8835 & ~n9161 ) | ( n8835 & n9162 ) | ( ~n9161 & n9162 ) ;
  assign n9164 = ( x89 & n9158 ) | ( x89 & ~n9163 ) | ( n9158 & ~n9163 ) ;
  assign n9165 = ( x89 & n8836 ) | ( x89 & ~n9015 ) | ( n8836 & ~n9015 ) ;
  assign n9166 = x89 & n8836 ;
  assign n9167 = ( ~n8841 & n9165 ) | ( ~n8841 & n9166 ) | ( n9165 & n9166 ) ;
  assign n9168 = ( n8841 & n9165 ) | ( n8841 & n9166 ) | ( n9165 & n9166 ) ;
  assign n9169 = ( n8841 & n9167 ) | ( n8841 & ~n9168 ) | ( n9167 & ~n9168 ) ;
  assign n9170 = ( x90 & n9164 ) | ( x90 & ~n9169 ) | ( n9164 & ~n9169 ) ;
  assign n9171 = ( x90 & n8842 ) | ( x90 & ~n9015 ) | ( n8842 & ~n9015 ) ;
  assign n9172 = x90 & n8842 ;
  assign n9173 = ( n8847 & n9171 ) | ( n8847 & n9172 ) | ( n9171 & n9172 ) ;
  assign n9174 = ( ~n8847 & n9171 ) | ( ~n8847 & n9172 ) | ( n9171 & n9172 ) ;
  assign n9175 = ( n8847 & ~n9173 ) | ( n8847 & n9174 ) | ( ~n9173 & n9174 ) ;
  assign n9176 = ( x91 & n9170 ) | ( x91 & ~n9175 ) | ( n9170 & ~n9175 ) ;
  assign n9177 = ( x91 & n8848 ) | ( x91 & ~n9015 ) | ( n8848 & ~n9015 ) ;
  assign n9178 = x91 & n8848 ;
  assign n9179 = ( ~n8853 & n9177 ) | ( ~n8853 & n9178 ) | ( n9177 & n9178 ) ;
  assign n9180 = ( n8853 & n9177 ) | ( n8853 & n9178 ) | ( n9177 & n9178 ) ;
  assign n9181 = ( n8853 & n9179 ) | ( n8853 & ~n9180 ) | ( n9179 & ~n9180 ) ;
  assign n9182 = ( x92 & n9176 ) | ( x92 & ~n9181 ) | ( n9176 & ~n9181 ) ;
  assign n9183 = ( x92 & n8854 ) | ( x92 & ~n9015 ) | ( n8854 & ~n9015 ) ;
  assign n9184 = x92 & n8854 ;
  assign n9185 = ( n8859 & n9183 ) | ( n8859 & n9184 ) | ( n9183 & n9184 ) ;
  assign n9186 = ( ~n8859 & n9183 ) | ( ~n8859 & n9184 ) | ( n9183 & n9184 ) ;
  assign n9187 = ( n8859 & ~n9185 ) | ( n8859 & n9186 ) | ( ~n9185 & n9186 ) ;
  assign n9188 = ( x93 & n9182 ) | ( x93 & ~n9187 ) | ( n9182 & ~n9187 ) ;
  assign n9189 = ( x93 & n8860 ) | ( x93 & ~n9015 ) | ( n8860 & ~n9015 ) ;
  assign n9190 = x93 & n8860 ;
  assign n9191 = ( ~n8865 & n9189 ) | ( ~n8865 & n9190 ) | ( n9189 & n9190 ) ;
  assign n9192 = ( n8865 & n9189 ) | ( n8865 & n9190 ) | ( n9189 & n9190 ) ;
  assign n9193 = ( n8865 & n9191 ) | ( n8865 & ~n9192 ) | ( n9191 & ~n9192 ) ;
  assign n9194 = ( x94 & n9188 ) | ( x94 & ~n9193 ) | ( n9188 & ~n9193 ) ;
  assign n9195 = ( x94 & n8866 ) | ( x94 & ~n9015 ) | ( n8866 & ~n9015 ) ;
  assign n9196 = x94 & n8866 ;
  assign n9197 = ( n8871 & n9195 ) | ( n8871 & n9196 ) | ( n9195 & n9196 ) ;
  assign n9198 = ( ~n8871 & n9195 ) | ( ~n8871 & n9196 ) | ( n9195 & n9196 ) ;
  assign n9199 = ( n8871 & ~n9197 ) | ( n8871 & n9198 ) | ( ~n9197 & n9198 ) ;
  assign n9200 = ( x95 & n9194 ) | ( x95 & ~n9199 ) | ( n9194 & ~n9199 ) ;
  assign n9201 = ( x95 & n8872 ) | ( x95 & ~n9015 ) | ( n8872 & ~n9015 ) ;
  assign n9202 = x95 & n8872 ;
  assign n9203 = ( ~n8877 & n9201 ) | ( ~n8877 & n9202 ) | ( n9201 & n9202 ) ;
  assign n9204 = ( n8877 & n9201 ) | ( n8877 & n9202 ) | ( n9201 & n9202 ) ;
  assign n9205 = ( n8877 & n9203 ) | ( n8877 & ~n9204 ) | ( n9203 & ~n9204 ) ;
  assign n9206 = ( x96 & n9200 ) | ( x96 & ~n9205 ) | ( n9200 & ~n9205 ) ;
  assign n9207 = ( x96 & n8878 ) | ( x96 & ~n9015 ) | ( n8878 & ~n9015 ) ;
  assign n9208 = x96 & n8878 ;
  assign n9209 = ( n8883 & n9207 ) | ( n8883 & n9208 ) | ( n9207 & n9208 ) ;
  assign n9210 = ( ~n8883 & n9207 ) | ( ~n8883 & n9208 ) | ( n9207 & n9208 ) ;
  assign n9211 = ( n8883 & ~n9209 ) | ( n8883 & n9210 ) | ( ~n9209 & n9210 ) ;
  assign n9212 = ( x97 & n9206 ) | ( x97 & ~n9211 ) | ( n9206 & ~n9211 ) ;
  assign n9213 = ( x97 & n8884 ) | ( x97 & ~n9015 ) | ( n8884 & ~n9015 ) ;
  assign n9214 = x97 & n8884 ;
  assign n9215 = ( ~n8889 & n9213 ) | ( ~n8889 & n9214 ) | ( n9213 & n9214 ) ;
  assign n9216 = ( n8889 & n9213 ) | ( n8889 & n9214 ) | ( n9213 & n9214 ) ;
  assign n9217 = ( n8889 & n9215 ) | ( n8889 & ~n9216 ) | ( n9215 & ~n9216 ) ;
  assign n9218 = ( x98 & n9212 ) | ( x98 & ~n9217 ) | ( n9212 & ~n9217 ) ;
  assign n9219 = ( x98 & n8890 ) | ( x98 & ~n9015 ) | ( n8890 & ~n9015 ) ;
  assign n9220 = x98 & n8890 ;
  assign n9221 = ( n8895 & n9219 ) | ( n8895 & n9220 ) | ( n9219 & n9220 ) ;
  assign n9222 = ( ~n8895 & n9219 ) | ( ~n8895 & n9220 ) | ( n9219 & n9220 ) ;
  assign n9223 = ( n8895 & ~n9221 ) | ( n8895 & n9222 ) | ( ~n9221 & n9222 ) ;
  assign n9224 = ( x99 & n9218 ) | ( x99 & ~n9223 ) | ( n9218 & ~n9223 ) ;
  assign n9225 = ( x99 & n8896 ) | ( x99 & ~n9015 ) | ( n8896 & ~n9015 ) ;
  assign n9226 = x99 & n8896 ;
  assign n9227 = ( ~n8901 & n9225 ) | ( ~n8901 & n9226 ) | ( n9225 & n9226 ) ;
  assign n9228 = ( n8901 & n9225 ) | ( n8901 & n9226 ) | ( n9225 & n9226 ) ;
  assign n9229 = ( n8901 & n9227 ) | ( n8901 & ~n9228 ) | ( n9227 & ~n9228 ) ;
  assign n9230 = ( x100 & n9224 ) | ( x100 & ~n9229 ) | ( n9224 & ~n9229 ) ;
  assign n9231 = ( x100 & n8902 ) | ( x100 & ~n9015 ) | ( n8902 & ~n9015 ) ;
  assign n9232 = x100 & n8902 ;
  assign n9233 = ( n8907 & n9231 ) | ( n8907 & n9232 ) | ( n9231 & n9232 ) ;
  assign n9234 = ( ~n8907 & n9231 ) | ( ~n8907 & n9232 ) | ( n9231 & n9232 ) ;
  assign n9235 = ( n8907 & ~n9233 ) | ( n8907 & n9234 ) | ( ~n9233 & n9234 ) ;
  assign n9236 = ( x101 & n9230 ) | ( x101 & ~n9235 ) | ( n9230 & ~n9235 ) ;
  assign n9237 = ( x101 & n8908 ) | ( x101 & ~n9015 ) | ( n8908 & ~n9015 ) ;
  assign n9238 = x101 & n8908 ;
  assign n9239 = ( ~n8913 & n9237 ) | ( ~n8913 & n9238 ) | ( n9237 & n9238 ) ;
  assign n9240 = ( n8913 & n9237 ) | ( n8913 & n9238 ) | ( n9237 & n9238 ) ;
  assign n9241 = ( n8913 & n9239 ) | ( n8913 & ~n9240 ) | ( n9239 & ~n9240 ) ;
  assign n9242 = ( x102 & n9236 ) | ( x102 & ~n9241 ) | ( n9236 & ~n9241 ) ;
  assign n9243 = ( x102 & n8914 ) | ( x102 & ~n9015 ) | ( n8914 & ~n9015 ) ;
  assign n9244 = x102 & n8914 ;
  assign n9245 = ( n8919 & n9243 ) | ( n8919 & n9244 ) | ( n9243 & n9244 ) ;
  assign n9246 = ( ~n8919 & n9243 ) | ( ~n8919 & n9244 ) | ( n9243 & n9244 ) ;
  assign n9247 = ( n8919 & ~n9245 ) | ( n8919 & n9246 ) | ( ~n9245 & n9246 ) ;
  assign n9248 = ( x103 & n9242 ) | ( x103 & ~n9247 ) | ( n9242 & ~n9247 ) ;
  assign n9249 = ( x103 & n8920 ) | ( x103 & ~n9015 ) | ( n8920 & ~n9015 ) ;
  assign n9250 = x103 & n8920 ;
  assign n9251 = ( ~n8925 & n9249 ) | ( ~n8925 & n9250 ) | ( n9249 & n9250 ) ;
  assign n9252 = ( n8925 & n9249 ) | ( n8925 & n9250 ) | ( n9249 & n9250 ) ;
  assign n9253 = ( n8925 & n9251 ) | ( n8925 & ~n9252 ) | ( n9251 & ~n9252 ) ;
  assign n9254 = ( x104 & n9248 ) | ( x104 & ~n9253 ) | ( n9248 & ~n9253 ) ;
  assign n9255 = ( x104 & n8926 ) | ( x104 & ~n9015 ) | ( n8926 & ~n9015 ) ;
  assign n9256 = x104 & n8926 ;
  assign n9257 = ( n8931 & n9255 ) | ( n8931 & n9256 ) | ( n9255 & n9256 ) ;
  assign n9258 = ( ~n8931 & n9255 ) | ( ~n8931 & n9256 ) | ( n9255 & n9256 ) ;
  assign n9259 = ( n8931 & ~n9257 ) | ( n8931 & n9258 ) | ( ~n9257 & n9258 ) ;
  assign n9260 = ( x105 & n9254 ) | ( x105 & ~n9259 ) | ( n9254 & ~n9259 ) ;
  assign n9261 = ( x105 & n8932 ) | ( x105 & ~n9015 ) | ( n8932 & ~n9015 ) ;
  assign n9262 = x105 & n8932 ;
  assign n9263 = ( ~n8937 & n9261 ) | ( ~n8937 & n9262 ) | ( n9261 & n9262 ) ;
  assign n9264 = ( n8937 & n9261 ) | ( n8937 & n9262 ) | ( n9261 & n9262 ) ;
  assign n9265 = ( n8937 & n9263 ) | ( n8937 & ~n9264 ) | ( n9263 & ~n9264 ) ;
  assign n9266 = ( x106 & n9260 ) | ( x106 & ~n9265 ) | ( n9260 & ~n9265 ) ;
  assign n9267 = ( x106 & n8938 ) | ( x106 & ~n9015 ) | ( n8938 & ~n9015 ) ;
  assign n9268 = x106 & n8938 ;
  assign n9269 = ( n8943 & n9267 ) | ( n8943 & n9268 ) | ( n9267 & n9268 ) ;
  assign n9270 = ( ~n8943 & n9267 ) | ( ~n8943 & n9268 ) | ( n9267 & n9268 ) ;
  assign n9271 = ( n8943 & ~n9269 ) | ( n8943 & n9270 ) | ( ~n9269 & n9270 ) ;
  assign n9272 = ( x107 & n9266 ) | ( x107 & ~n9271 ) | ( n9266 & ~n9271 ) ;
  assign n9273 = ( x107 & n8944 ) | ( x107 & ~n9015 ) | ( n8944 & ~n9015 ) ;
  assign n9274 = x107 & n8944 ;
  assign n9275 = ( ~n8949 & n9273 ) | ( ~n8949 & n9274 ) | ( n9273 & n9274 ) ;
  assign n9276 = ( n8949 & n9273 ) | ( n8949 & n9274 ) | ( n9273 & n9274 ) ;
  assign n9277 = ( n8949 & n9275 ) | ( n8949 & ~n9276 ) | ( n9275 & ~n9276 ) ;
  assign n9278 = ( x108 & n9272 ) | ( x108 & ~n9277 ) | ( n9272 & ~n9277 ) ;
  assign n9279 = ( x108 & n8950 ) | ( x108 & ~n9015 ) | ( n8950 & ~n9015 ) ;
  assign n9280 = x108 & n8950 ;
  assign n9281 = ( n8955 & n9279 ) | ( n8955 & n9280 ) | ( n9279 & n9280 ) ;
  assign n9282 = ( ~n8955 & n9279 ) | ( ~n8955 & n9280 ) | ( n9279 & n9280 ) ;
  assign n9283 = ( n8955 & ~n9281 ) | ( n8955 & n9282 ) | ( ~n9281 & n9282 ) ;
  assign n9284 = ( x109 & n9278 ) | ( x109 & ~n9283 ) | ( n9278 & ~n9283 ) ;
  assign n9285 = ( x109 & n8956 ) | ( x109 & ~n9015 ) | ( n8956 & ~n9015 ) ;
  assign n9286 = x109 & n8956 ;
  assign n9287 = ( ~n8961 & n9285 ) | ( ~n8961 & n9286 ) | ( n9285 & n9286 ) ;
  assign n9288 = ( n8961 & n9285 ) | ( n8961 & n9286 ) | ( n9285 & n9286 ) ;
  assign n9289 = ( n8961 & n9287 ) | ( n8961 & ~n9288 ) | ( n9287 & ~n9288 ) ;
  assign n9290 = ( x110 & n9284 ) | ( x110 & ~n9289 ) | ( n9284 & ~n9289 ) ;
  assign n9291 = ( x110 & n8962 ) | ( x110 & ~n9015 ) | ( n8962 & ~n9015 ) ;
  assign n9292 = x110 & n8962 ;
  assign n9293 = ( n8967 & n9291 ) | ( n8967 & n9292 ) | ( n9291 & n9292 ) ;
  assign n9294 = ( ~n8967 & n9291 ) | ( ~n8967 & n9292 ) | ( n9291 & n9292 ) ;
  assign n9295 = ( n8967 & ~n9293 ) | ( n8967 & n9294 ) | ( ~n9293 & n9294 ) ;
  assign n9296 = ( x111 & n9290 ) | ( x111 & ~n9295 ) | ( n9290 & ~n9295 ) ;
  assign n9297 = ( x111 & n8968 ) | ( x111 & ~n9015 ) | ( n8968 & ~n9015 ) ;
  assign n9298 = x111 & n8968 ;
  assign n9299 = ( ~n8973 & n9297 ) | ( ~n8973 & n9298 ) | ( n9297 & n9298 ) ;
  assign n9300 = ( n8973 & n9297 ) | ( n8973 & n9298 ) | ( n9297 & n9298 ) ;
  assign n9301 = ( n8973 & n9299 ) | ( n8973 & ~n9300 ) | ( n9299 & ~n9300 ) ;
  assign n9302 = ( x112 & n9296 ) | ( x112 & ~n9301 ) | ( n9296 & ~n9301 ) ;
  assign n9303 = ( x112 & n8974 ) | ( x112 & ~n9015 ) | ( n8974 & ~n9015 ) ;
  assign n9304 = x112 & n8974 ;
  assign n9305 = ( n8979 & n9303 ) | ( n8979 & n9304 ) | ( n9303 & n9304 ) ;
  assign n9306 = ( ~n8979 & n9303 ) | ( ~n8979 & n9304 ) | ( n9303 & n9304 ) ;
  assign n9307 = ( n8979 & ~n9305 ) | ( n8979 & n9306 ) | ( ~n9305 & n9306 ) ;
  assign n9308 = ( x113 & n9302 ) | ( x113 & ~n9307 ) | ( n9302 & ~n9307 ) ;
  assign n9309 = ( x113 & n8980 ) | ( x113 & ~n9015 ) | ( n8980 & ~n9015 ) ;
  assign n9310 = x113 & n8980 ;
  assign n9311 = ( ~n8985 & n9309 ) | ( ~n8985 & n9310 ) | ( n9309 & n9310 ) ;
  assign n9312 = ( n8985 & n9309 ) | ( n8985 & n9310 ) | ( n9309 & n9310 ) ;
  assign n9313 = ( n8985 & n9311 ) | ( n8985 & ~n9312 ) | ( n9311 & ~n9312 ) ;
  assign n9314 = ( x114 & n9308 ) | ( x114 & ~n9313 ) | ( n9308 & ~n9313 ) ;
  assign n9315 = ( x114 & n8986 ) | ( x114 & ~n9015 ) | ( n8986 & ~n9015 ) ;
  assign n9316 = x114 & n8986 ;
  assign n9317 = ( n8991 & n9315 ) | ( n8991 & n9316 ) | ( n9315 & n9316 ) ;
  assign n9318 = ( ~n8991 & n9315 ) | ( ~n8991 & n9316 ) | ( n9315 & n9316 ) ;
  assign n9319 = ( n8991 & ~n9317 ) | ( n8991 & n9318 ) | ( ~n9317 & n9318 ) ;
  assign n9320 = ( x115 & n9314 ) | ( x115 & ~n9319 ) | ( n9314 & ~n9319 ) ;
  assign n9321 = ( x115 & n8992 ) | ( x115 & ~n9015 ) | ( n8992 & ~n9015 ) ;
  assign n9322 = x115 & n8992 ;
  assign n9323 = ( ~n8997 & n9321 ) | ( ~n8997 & n9322 ) | ( n9321 & n9322 ) ;
  assign n9324 = ( n8997 & n9321 ) | ( n8997 & n9322 ) | ( n9321 & n9322 ) ;
  assign n9325 = ( n8997 & n9323 ) | ( n8997 & ~n9324 ) | ( n9323 & ~n9324 ) ;
  assign n9326 = ( x116 & n9320 ) | ( x116 & ~n9325 ) | ( n9320 & ~n9325 ) ;
  assign n9327 = ( x116 & n8998 ) | ( x116 & ~n9015 ) | ( n8998 & ~n9015 ) ;
  assign n9328 = x116 & n8998 ;
  assign n9329 = ( n9003 & n9327 ) | ( n9003 & n9328 ) | ( n9327 & n9328 ) ;
  assign n9330 = ( ~n9003 & n9327 ) | ( ~n9003 & n9328 ) | ( n9327 & n9328 ) ;
  assign n9331 = ( n9003 & ~n9329 ) | ( n9003 & n9330 ) | ( ~n9329 & n9330 ) ;
  assign n9332 = ( x117 & n9326 ) | ( x117 & ~n9331 ) | ( n9326 & ~n9331 ) ;
  assign n9333 = ( x117 & n9004 ) | ( x117 & ~n9015 ) | ( n9004 & ~n9015 ) ;
  assign n9334 = x117 & n9004 ;
  assign n9335 = ( n9009 & n9333 ) | ( n9009 & n9334 ) | ( n9333 & n9334 ) ;
  assign n9336 = ( ~n9009 & n9333 ) | ( ~n9009 & n9334 ) | ( n9333 & n9334 ) ;
  assign n9337 = ( n9009 & ~n9335 ) | ( n9009 & n9336 ) | ( ~n9335 & n9336 ) ;
  assign n9338 = ( x118 & n9332 ) | ( x118 & ~n9337 ) | ( n9332 & ~n9337 ) ;
  assign n9339 = x119 | n9338 ;
  assign n9340 = ( x119 & n138 ) | ( x119 & n9338 ) | ( n138 & n9338 ) ;
  assign n9341 = ( n9013 & ~n9339 ) | ( n9013 & n9340 ) | ( ~n9339 & n9340 ) ;
  assign n9342 = ( x119 & ~n9013 ) | ( x119 & n9338 ) | ( ~n9013 & n9338 ) ;
  assign n9343 = n138 | n9342 ;
  assign n9344 = ( x8 & ~x64 ) | ( x8 & n9343 ) | ( ~x64 & n9343 ) ;
  assign n9345 = ~x8 & n9343 ;
  assign n9346 = ( n9019 & n9344 ) | ( n9019 & ~n9345 ) | ( n9344 & ~n9345 ) ;
  assign n9347 = ~x7 & x64 ;
  assign n9348 = ( x65 & ~n9346 ) | ( x65 & n9347 ) | ( ~n9346 & n9347 ) ;
  assign n9349 = ( x65 & n9019 ) | ( x65 & ~n9343 ) | ( n9019 & ~n9343 ) ;
  assign n9350 = x65 & n9019 ;
  assign n9351 = ( n9018 & n9349 ) | ( n9018 & n9350 ) | ( n9349 & n9350 ) ;
  assign n9352 = ( ~n9018 & n9349 ) | ( ~n9018 & n9350 ) | ( n9349 & n9350 ) ;
  assign n9353 = ( n9018 & ~n9351 ) | ( n9018 & n9352 ) | ( ~n9351 & n9352 ) ;
  assign n9354 = ( x66 & n9348 ) | ( x66 & ~n9353 ) | ( n9348 & ~n9353 ) ;
  assign n9355 = ( x66 & n9020 ) | ( x66 & ~n9343 ) | ( n9020 & ~n9343 ) ;
  assign n9356 = x66 & n9020 ;
  assign n9357 = ( n9025 & n9355 ) | ( n9025 & n9356 ) | ( n9355 & n9356 ) ;
  assign n9358 = ( ~n9025 & n9355 ) | ( ~n9025 & n9356 ) | ( n9355 & n9356 ) ;
  assign n9359 = ( n9025 & ~n9357 ) | ( n9025 & n9358 ) | ( ~n9357 & n9358 ) ;
  assign n9360 = ( x67 & n9354 ) | ( x67 & ~n9359 ) | ( n9354 & ~n9359 ) ;
  assign n9361 = ( x67 & n9026 ) | ( x67 & ~n9343 ) | ( n9026 & ~n9343 ) ;
  assign n9362 = x67 & n9026 ;
  assign n9363 = ( ~n9031 & n9361 ) | ( ~n9031 & n9362 ) | ( n9361 & n9362 ) ;
  assign n9364 = ( n9031 & n9361 ) | ( n9031 & n9362 ) | ( n9361 & n9362 ) ;
  assign n9365 = ( n9031 & n9363 ) | ( n9031 & ~n9364 ) | ( n9363 & ~n9364 ) ;
  assign n9366 = ( x68 & n9360 ) | ( x68 & ~n9365 ) | ( n9360 & ~n9365 ) ;
  assign n9367 = ( x68 & n9032 ) | ( x68 & ~n9343 ) | ( n9032 & ~n9343 ) ;
  assign n9368 = x68 & n9032 ;
  assign n9369 = ( n9037 & n9367 ) | ( n9037 & n9368 ) | ( n9367 & n9368 ) ;
  assign n9370 = ( ~n9037 & n9367 ) | ( ~n9037 & n9368 ) | ( n9367 & n9368 ) ;
  assign n9371 = ( n9037 & ~n9369 ) | ( n9037 & n9370 ) | ( ~n9369 & n9370 ) ;
  assign n9372 = ( x69 & n9366 ) | ( x69 & ~n9371 ) | ( n9366 & ~n9371 ) ;
  assign n9373 = ( x69 & n9038 ) | ( x69 & ~n9343 ) | ( n9038 & ~n9343 ) ;
  assign n9374 = x69 & n9038 ;
  assign n9375 = ( ~n9043 & n9373 ) | ( ~n9043 & n9374 ) | ( n9373 & n9374 ) ;
  assign n9376 = ( n9043 & n9373 ) | ( n9043 & n9374 ) | ( n9373 & n9374 ) ;
  assign n9377 = ( n9043 & n9375 ) | ( n9043 & ~n9376 ) | ( n9375 & ~n9376 ) ;
  assign n9378 = ( x70 & n9372 ) | ( x70 & ~n9377 ) | ( n9372 & ~n9377 ) ;
  assign n9379 = ( x70 & n9044 ) | ( x70 & ~n9343 ) | ( n9044 & ~n9343 ) ;
  assign n9380 = x70 & n9044 ;
  assign n9381 = ( n9049 & n9379 ) | ( n9049 & n9380 ) | ( n9379 & n9380 ) ;
  assign n9382 = ( ~n9049 & n9379 ) | ( ~n9049 & n9380 ) | ( n9379 & n9380 ) ;
  assign n9383 = ( n9049 & ~n9381 ) | ( n9049 & n9382 ) | ( ~n9381 & n9382 ) ;
  assign n9384 = ( x71 & n9378 ) | ( x71 & ~n9383 ) | ( n9378 & ~n9383 ) ;
  assign n9385 = ( x71 & n9050 ) | ( x71 & ~n9343 ) | ( n9050 & ~n9343 ) ;
  assign n9386 = x71 & n9050 ;
  assign n9387 = ( ~n9055 & n9385 ) | ( ~n9055 & n9386 ) | ( n9385 & n9386 ) ;
  assign n9388 = ( n9055 & n9385 ) | ( n9055 & n9386 ) | ( n9385 & n9386 ) ;
  assign n9389 = ( n9055 & n9387 ) | ( n9055 & ~n9388 ) | ( n9387 & ~n9388 ) ;
  assign n9390 = ( x72 & n9384 ) | ( x72 & ~n9389 ) | ( n9384 & ~n9389 ) ;
  assign n9391 = ( x72 & n9056 ) | ( x72 & ~n9343 ) | ( n9056 & ~n9343 ) ;
  assign n9392 = x72 & n9056 ;
  assign n9393 = ( n9061 & n9391 ) | ( n9061 & n9392 ) | ( n9391 & n9392 ) ;
  assign n9394 = ( ~n9061 & n9391 ) | ( ~n9061 & n9392 ) | ( n9391 & n9392 ) ;
  assign n9395 = ( n9061 & ~n9393 ) | ( n9061 & n9394 ) | ( ~n9393 & n9394 ) ;
  assign n9396 = ( x73 & n9390 ) | ( x73 & ~n9395 ) | ( n9390 & ~n9395 ) ;
  assign n9397 = ( x73 & n9062 ) | ( x73 & ~n9343 ) | ( n9062 & ~n9343 ) ;
  assign n9398 = x73 & n9062 ;
  assign n9399 = ( ~n9067 & n9397 ) | ( ~n9067 & n9398 ) | ( n9397 & n9398 ) ;
  assign n9400 = ( n9067 & n9397 ) | ( n9067 & n9398 ) | ( n9397 & n9398 ) ;
  assign n9401 = ( n9067 & n9399 ) | ( n9067 & ~n9400 ) | ( n9399 & ~n9400 ) ;
  assign n9402 = ( x74 & n9396 ) | ( x74 & ~n9401 ) | ( n9396 & ~n9401 ) ;
  assign n9403 = ( x74 & n9068 ) | ( x74 & ~n9343 ) | ( n9068 & ~n9343 ) ;
  assign n9404 = x74 & n9068 ;
  assign n9405 = ( n9073 & n9403 ) | ( n9073 & n9404 ) | ( n9403 & n9404 ) ;
  assign n9406 = ( ~n9073 & n9403 ) | ( ~n9073 & n9404 ) | ( n9403 & n9404 ) ;
  assign n9407 = ( n9073 & ~n9405 ) | ( n9073 & n9406 ) | ( ~n9405 & n9406 ) ;
  assign n9408 = ( x75 & n9402 ) | ( x75 & ~n9407 ) | ( n9402 & ~n9407 ) ;
  assign n9409 = ( x75 & n9074 ) | ( x75 & ~n9343 ) | ( n9074 & ~n9343 ) ;
  assign n9410 = x75 & n9074 ;
  assign n9411 = ( ~n9079 & n9409 ) | ( ~n9079 & n9410 ) | ( n9409 & n9410 ) ;
  assign n9412 = ( n9079 & n9409 ) | ( n9079 & n9410 ) | ( n9409 & n9410 ) ;
  assign n9413 = ( n9079 & n9411 ) | ( n9079 & ~n9412 ) | ( n9411 & ~n9412 ) ;
  assign n9414 = ( x76 & n9408 ) | ( x76 & ~n9413 ) | ( n9408 & ~n9413 ) ;
  assign n9415 = ( x76 & n9080 ) | ( x76 & ~n9343 ) | ( n9080 & ~n9343 ) ;
  assign n9416 = x76 & n9080 ;
  assign n9417 = ( n9085 & n9415 ) | ( n9085 & n9416 ) | ( n9415 & n9416 ) ;
  assign n9418 = ( ~n9085 & n9415 ) | ( ~n9085 & n9416 ) | ( n9415 & n9416 ) ;
  assign n9419 = ( n9085 & ~n9417 ) | ( n9085 & n9418 ) | ( ~n9417 & n9418 ) ;
  assign n9420 = ( x77 & n9414 ) | ( x77 & ~n9419 ) | ( n9414 & ~n9419 ) ;
  assign n9421 = ( x77 & n9086 ) | ( x77 & ~n9343 ) | ( n9086 & ~n9343 ) ;
  assign n9422 = x77 & n9086 ;
  assign n9423 = ( ~n9091 & n9421 ) | ( ~n9091 & n9422 ) | ( n9421 & n9422 ) ;
  assign n9424 = ( n9091 & n9421 ) | ( n9091 & n9422 ) | ( n9421 & n9422 ) ;
  assign n9425 = ( n9091 & n9423 ) | ( n9091 & ~n9424 ) | ( n9423 & ~n9424 ) ;
  assign n9426 = ( x78 & n9420 ) | ( x78 & ~n9425 ) | ( n9420 & ~n9425 ) ;
  assign n9427 = ( x78 & n9092 ) | ( x78 & ~n9343 ) | ( n9092 & ~n9343 ) ;
  assign n9428 = x78 & n9092 ;
  assign n9429 = ( n9097 & n9427 ) | ( n9097 & n9428 ) | ( n9427 & n9428 ) ;
  assign n9430 = ( ~n9097 & n9427 ) | ( ~n9097 & n9428 ) | ( n9427 & n9428 ) ;
  assign n9431 = ( n9097 & ~n9429 ) | ( n9097 & n9430 ) | ( ~n9429 & n9430 ) ;
  assign n9432 = ( x79 & n9426 ) | ( x79 & ~n9431 ) | ( n9426 & ~n9431 ) ;
  assign n9433 = ( x79 & n9098 ) | ( x79 & ~n9343 ) | ( n9098 & ~n9343 ) ;
  assign n9434 = x79 & n9098 ;
  assign n9435 = ( ~n9103 & n9433 ) | ( ~n9103 & n9434 ) | ( n9433 & n9434 ) ;
  assign n9436 = ( n9103 & n9433 ) | ( n9103 & n9434 ) | ( n9433 & n9434 ) ;
  assign n9437 = ( n9103 & n9435 ) | ( n9103 & ~n9436 ) | ( n9435 & ~n9436 ) ;
  assign n9438 = ( x80 & n9432 ) | ( x80 & ~n9437 ) | ( n9432 & ~n9437 ) ;
  assign n9439 = ( x80 & n9104 ) | ( x80 & ~n9343 ) | ( n9104 & ~n9343 ) ;
  assign n9440 = x80 & n9104 ;
  assign n9441 = ( n9109 & n9439 ) | ( n9109 & n9440 ) | ( n9439 & n9440 ) ;
  assign n9442 = ( ~n9109 & n9439 ) | ( ~n9109 & n9440 ) | ( n9439 & n9440 ) ;
  assign n9443 = ( n9109 & ~n9441 ) | ( n9109 & n9442 ) | ( ~n9441 & n9442 ) ;
  assign n9444 = ( x81 & n9438 ) | ( x81 & ~n9443 ) | ( n9438 & ~n9443 ) ;
  assign n9445 = ( x81 & n9110 ) | ( x81 & ~n9343 ) | ( n9110 & ~n9343 ) ;
  assign n9446 = x81 & n9110 ;
  assign n9447 = ( ~n9115 & n9445 ) | ( ~n9115 & n9446 ) | ( n9445 & n9446 ) ;
  assign n9448 = ( n9115 & n9445 ) | ( n9115 & n9446 ) | ( n9445 & n9446 ) ;
  assign n9449 = ( n9115 & n9447 ) | ( n9115 & ~n9448 ) | ( n9447 & ~n9448 ) ;
  assign n9450 = ( x82 & n9444 ) | ( x82 & ~n9449 ) | ( n9444 & ~n9449 ) ;
  assign n9451 = ( x82 & n9116 ) | ( x82 & ~n9343 ) | ( n9116 & ~n9343 ) ;
  assign n9452 = x82 & n9116 ;
  assign n9453 = ( n9121 & n9451 ) | ( n9121 & n9452 ) | ( n9451 & n9452 ) ;
  assign n9454 = ( ~n9121 & n9451 ) | ( ~n9121 & n9452 ) | ( n9451 & n9452 ) ;
  assign n9455 = ( n9121 & ~n9453 ) | ( n9121 & n9454 ) | ( ~n9453 & n9454 ) ;
  assign n9456 = ( x83 & n9450 ) | ( x83 & ~n9455 ) | ( n9450 & ~n9455 ) ;
  assign n9457 = ( x83 & n9122 ) | ( x83 & ~n9343 ) | ( n9122 & ~n9343 ) ;
  assign n9458 = x83 & n9122 ;
  assign n9459 = ( ~n9127 & n9457 ) | ( ~n9127 & n9458 ) | ( n9457 & n9458 ) ;
  assign n9460 = ( n9127 & n9457 ) | ( n9127 & n9458 ) | ( n9457 & n9458 ) ;
  assign n9461 = ( n9127 & n9459 ) | ( n9127 & ~n9460 ) | ( n9459 & ~n9460 ) ;
  assign n9462 = ( x84 & n9456 ) | ( x84 & ~n9461 ) | ( n9456 & ~n9461 ) ;
  assign n9463 = ( x84 & n9128 ) | ( x84 & ~n9343 ) | ( n9128 & ~n9343 ) ;
  assign n9464 = x84 & n9128 ;
  assign n9465 = ( n9133 & n9463 ) | ( n9133 & n9464 ) | ( n9463 & n9464 ) ;
  assign n9466 = ( ~n9133 & n9463 ) | ( ~n9133 & n9464 ) | ( n9463 & n9464 ) ;
  assign n9467 = ( n9133 & ~n9465 ) | ( n9133 & n9466 ) | ( ~n9465 & n9466 ) ;
  assign n9468 = ( x85 & n9462 ) | ( x85 & ~n9467 ) | ( n9462 & ~n9467 ) ;
  assign n9469 = ( x85 & n9134 ) | ( x85 & ~n9343 ) | ( n9134 & ~n9343 ) ;
  assign n9470 = x85 & n9134 ;
  assign n9471 = ( ~n9139 & n9469 ) | ( ~n9139 & n9470 ) | ( n9469 & n9470 ) ;
  assign n9472 = ( n9139 & n9469 ) | ( n9139 & n9470 ) | ( n9469 & n9470 ) ;
  assign n9473 = ( n9139 & n9471 ) | ( n9139 & ~n9472 ) | ( n9471 & ~n9472 ) ;
  assign n9474 = ( x86 & n9468 ) | ( x86 & ~n9473 ) | ( n9468 & ~n9473 ) ;
  assign n9475 = ( x86 & n9140 ) | ( x86 & ~n9343 ) | ( n9140 & ~n9343 ) ;
  assign n9476 = x86 & n9140 ;
  assign n9477 = ( n9145 & n9475 ) | ( n9145 & n9476 ) | ( n9475 & n9476 ) ;
  assign n9478 = ( ~n9145 & n9475 ) | ( ~n9145 & n9476 ) | ( n9475 & n9476 ) ;
  assign n9479 = ( n9145 & ~n9477 ) | ( n9145 & n9478 ) | ( ~n9477 & n9478 ) ;
  assign n9480 = ( x87 & n9474 ) | ( x87 & ~n9479 ) | ( n9474 & ~n9479 ) ;
  assign n9481 = ( x87 & n9146 ) | ( x87 & ~n9343 ) | ( n9146 & ~n9343 ) ;
  assign n9482 = x87 & n9146 ;
  assign n9483 = ( ~n9151 & n9481 ) | ( ~n9151 & n9482 ) | ( n9481 & n9482 ) ;
  assign n9484 = ( n9151 & n9481 ) | ( n9151 & n9482 ) | ( n9481 & n9482 ) ;
  assign n9485 = ( n9151 & n9483 ) | ( n9151 & ~n9484 ) | ( n9483 & ~n9484 ) ;
  assign n9486 = ( x88 & n9480 ) | ( x88 & ~n9485 ) | ( n9480 & ~n9485 ) ;
  assign n9487 = ( x88 & n9152 ) | ( x88 & ~n9343 ) | ( n9152 & ~n9343 ) ;
  assign n9488 = x88 & n9152 ;
  assign n9489 = ( n9157 & n9487 ) | ( n9157 & n9488 ) | ( n9487 & n9488 ) ;
  assign n9490 = ( ~n9157 & n9487 ) | ( ~n9157 & n9488 ) | ( n9487 & n9488 ) ;
  assign n9491 = ( n9157 & ~n9489 ) | ( n9157 & n9490 ) | ( ~n9489 & n9490 ) ;
  assign n9492 = ( x89 & n9486 ) | ( x89 & ~n9491 ) | ( n9486 & ~n9491 ) ;
  assign n9493 = ( x89 & n9158 ) | ( x89 & ~n9343 ) | ( n9158 & ~n9343 ) ;
  assign n9494 = x89 & n9158 ;
  assign n9495 = ( ~n9163 & n9493 ) | ( ~n9163 & n9494 ) | ( n9493 & n9494 ) ;
  assign n9496 = ( n9163 & n9493 ) | ( n9163 & n9494 ) | ( n9493 & n9494 ) ;
  assign n9497 = ( n9163 & n9495 ) | ( n9163 & ~n9496 ) | ( n9495 & ~n9496 ) ;
  assign n9498 = ( x90 & n9492 ) | ( x90 & ~n9497 ) | ( n9492 & ~n9497 ) ;
  assign n9499 = ( x90 & n9164 ) | ( x90 & ~n9343 ) | ( n9164 & ~n9343 ) ;
  assign n9500 = x90 & n9164 ;
  assign n9501 = ( n9169 & n9499 ) | ( n9169 & n9500 ) | ( n9499 & n9500 ) ;
  assign n9502 = ( ~n9169 & n9499 ) | ( ~n9169 & n9500 ) | ( n9499 & n9500 ) ;
  assign n9503 = ( n9169 & ~n9501 ) | ( n9169 & n9502 ) | ( ~n9501 & n9502 ) ;
  assign n9504 = ( x91 & n9498 ) | ( x91 & ~n9503 ) | ( n9498 & ~n9503 ) ;
  assign n9505 = ( x91 & n9170 ) | ( x91 & ~n9343 ) | ( n9170 & ~n9343 ) ;
  assign n9506 = x91 & n9170 ;
  assign n9507 = ( ~n9175 & n9505 ) | ( ~n9175 & n9506 ) | ( n9505 & n9506 ) ;
  assign n9508 = ( n9175 & n9505 ) | ( n9175 & n9506 ) | ( n9505 & n9506 ) ;
  assign n9509 = ( n9175 & n9507 ) | ( n9175 & ~n9508 ) | ( n9507 & ~n9508 ) ;
  assign n9510 = ( x92 & n9504 ) | ( x92 & ~n9509 ) | ( n9504 & ~n9509 ) ;
  assign n9511 = ( x92 & n9176 ) | ( x92 & ~n9343 ) | ( n9176 & ~n9343 ) ;
  assign n9512 = x92 & n9176 ;
  assign n9513 = ( n9181 & n9511 ) | ( n9181 & n9512 ) | ( n9511 & n9512 ) ;
  assign n9514 = ( ~n9181 & n9511 ) | ( ~n9181 & n9512 ) | ( n9511 & n9512 ) ;
  assign n9515 = ( n9181 & ~n9513 ) | ( n9181 & n9514 ) | ( ~n9513 & n9514 ) ;
  assign n9516 = ( x93 & n9510 ) | ( x93 & ~n9515 ) | ( n9510 & ~n9515 ) ;
  assign n9517 = ( x93 & n9182 ) | ( x93 & ~n9343 ) | ( n9182 & ~n9343 ) ;
  assign n9518 = x93 & n9182 ;
  assign n9519 = ( ~n9187 & n9517 ) | ( ~n9187 & n9518 ) | ( n9517 & n9518 ) ;
  assign n9520 = ( n9187 & n9517 ) | ( n9187 & n9518 ) | ( n9517 & n9518 ) ;
  assign n9521 = ( n9187 & n9519 ) | ( n9187 & ~n9520 ) | ( n9519 & ~n9520 ) ;
  assign n9522 = ( x94 & n9516 ) | ( x94 & ~n9521 ) | ( n9516 & ~n9521 ) ;
  assign n9523 = ( x94 & n9188 ) | ( x94 & ~n9343 ) | ( n9188 & ~n9343 ) ;
  assign n9524 = x94 & n9188 ;
  assign n9525 = ( n9193 & n9523 ) | ( n9193 & n9524 ) | ( n9523 & n9524 ) ;
  assign n9526 = ( ~n9193 & n9523 ) | ( ~n9193 & n9524 ) | ( n9523 & n9524 ) ;
  assign n9527 = ( n9193 & ~n9525 ) | ( n9193 & n9526 ) | ( ~n9525 & n9526 ) ;
  assign n9528 = ( x95 & n9522 ) | ( x95 & ~n9527 ) | ( n9522 & ~n9527 ) ;
  assign n9529 = ( x95 & n9194 ) | ( x95 & ~n9343 ) | ( n9194 & ~n9343 ) ;
  assign n9530 = x95 & n9194 ;
  assign n9531 = ( ~n9199 & n9529 ) | ( ~n9199 & n9530 ) | ( n9529 & n9530 ) ;
  assign n9532 = ( n9199 & n9529 ) | ( n9199 & n9530 ) | ( n9529 & n9530 ) ;
  assign n9533 = ( n9199 & n9531 ) | ( n9199 & ~n9532 ) | ( n9531 & ~n9532 ) ;
  assign n9534 = ( x96 & n9528 ) | ( x96 & ~n9533 ) | ( n9528 & ~n9533 ) ;
  assign n9535 = ( x96 & n9200 ) | ( x96 & ~n9343 ) | ( n9200 & ~n9343 ) ;
  assign n9536 = x96 & n9200 ;
  assign n9537 = ( n9205 & n9535 ) | ( n9205 & n9536 ) | ( n9535 & n9536 ) ;
  assign n9538 = ( ~n9205 & n9535 ) | ( ~n9205 & n9536 ) | ( n9535 & n9536 ) ;
  assign n9539 = ( n9205 & ~n9537 ) | ( n9205 & n9538 ) | ( ~n9537 & n9538 ) ;
  assign n9540 = ( x97 & n9534 ) | ( x97 & ~n9539 ) | ( n9534 & ~n9539 ) ;
  assign n9541 = ( x97 & n9206 ) | ( x97 & ~n9343 ) | ( n9206 & ~n9343 ) ;
  assign n9542 = x97 & n9206 ;
  assign n9543 = ( ~n9211 & n9541 ) | ( ~n9211 & n9542 ) | ( n9541 & n9542 ) ;
  assign n9544 = ( n9211 & n9541 ) | ( n9211 & n9542 ) | ( n9541 & n9542 ) ;
  assign n9545 = ( n9211 & n9543 ) | ( n9211 & ~n9544 ) | ( n9543 & ~n9544 ) ;
  assign n9546 = ( x98 & n9540 ) | ( x98 & ~n9545 ) | ( n9540 & ~n9545 ) ;
  assign n9547 = ( x98 & n9212 ) | ( x98 & ~n9343 ) | ( n9212 & ~n9343 ) ;
  assign n9548 = x98 & n9212 ;
  assign n9549 = ( n9217 & n9547 ) | ( n9217 & n9548 ) | ( n9547 & n9548 ) ;
  assign n9550 = ( ~n9217 & n9547 ) | ( ~n9217 & n9548 ) | ( n9547 & n9548 ) ;
  assign n9551 = ( n9217 & ~n9549 ) | ( n9217 & n9550 ) | ( ~n9549 & n9550 ) ;
  assign n9552 = ( x99 & n9546 ) | ( x99 & ~n9551 ) | ( n9546 & ~n9551 ) ;
  assign n9553 = ( x99 & n9218 ) | ( x99 & ~n9343 ) | ( n9218 & ~n9343 ) ;
  assign n9554 = x99 & n9218 ;
  assign n9555 = ( ~n9223 & n9553 ) | ( ~n9223 & n9554 ) | ( n9553 & n9554 ) ;
  assign n9556 = ( n9223 & n9553 ) | ( n9223 & n9554 ) | ( n9553 & n9554 ) ;
  assign n9557 = ( n9223 & n9555 ) | ( n9223 & ~n9556 ) | ( n9555 & ~n9556 ) ;
  assign n9558 = ( x100 & n9552 ) | ( x100 & ~n9557 ) | ( n9552 & ~n9557 ) ;
  assign n9559 = ( x100 & n9224 ) | ( x100 & ~n9343 ) | ( n9224 & ~n9343 ) ;
  assign n9560 = x100 & n9224 ;
  assign n9561 = ( n9229 & n9559 ) | ( n9229 & n9560 ) | ( n9559 & n9560 ) ;
  assign n9562 = ( ~n9229 & n9559 ) | ( ~n9229 & n9560 ) | ( n9559 & n9560 ) ;
  assign n9563 = ( n9229 & ~n9561 ) | ( n9229 & n9562 ) | ( ~n9561 & n9562 ) ;
  assign n9564 = ( x101 & n9558 ) | ( x101 & ~n9563 ) | ( n9558 & ~n9563 ) ;
  assign n9565 = ( x101 & n9230 ) | ( x101 & ~n9343 ) | ( n9230 & ~n9343 ) ;
  assign n9566 = x101 & n9230 ;
  assign n9567 = ( ~n9235 & n9565 ) | ( ~n9235 & n9566 ) | ( n9565 & n9566 ) ;
  assign n9568 = ( n9235 & n9565 ) | ( n9235 & n9566 ) | ( n9565 & n9566 ) ;
  assign n9569 = ( n9235 & n9567 ) | ( n9235 & ~n9568 ) | ( n9567 & ~n9568 ) ;
  assign n9570 = ( x102 & n9564 ) | ( x102 & ~n9569 ) | ( n9564 & ~n9569 ) ;
  assign n9571 = ( x102 & n9236 ) | ( x102 & ~n9343 ) | ( n9236 & ~n9343 ) ;
  assign n9572 = x102 & n9236 ;
  assign n9573 = ( n9241 & n9571 ) | ( n9241 & n9572 ) | ( n9571 & n9572 ) ;
  assign n9574 = ( ~n9241 & n9571 ) | ( ~n9241 & n9572 ) | ( n9571 & n9572 ) ;
  assign n9575 = ( n9241 & ~n9573 ) | ( n9241 & n9574 ) | ( ~n9573 & n9574 ) ;
  assign n9576 = ( x103 & n9570 ) | ( x103 & ~n9575 ) | ( n9570 & ~n9575 ) ;
  assign n9577 = ( x103 & n9242 ) | ( x103 & ~n9343 ) | ( n9242 & ~n9343 ) ;
  assign n9578 = x103 & n9242 ;
  assign n9579 = ( ~n9247 & n9577 ) | ( ~n9247 & n9578 ) | ( n9577 & n9578 ) ;
  assign n9580 = ( n9247 & n9577 ) | ( n9247 & n9578 ) | ( n9577 & n9578 ) ;
  assign n9581 = ( n9247 & n9579 ) | ( n9247 & ~n9580 ) | ( n9579 & ~n9580 ) ;
  assign n9582 = ( x104 & n9576 ) | ( x104 & ~n9581 ) | ( n9576 & ~n9581 ) ;
  assign n9583 = ( x104 & n9248 ) | ( x104 & ~n9343 ) | ( n9248 & ~n9343 ) ;
  assign n9584 = x104 & n9248 ;
  assign n9585 = ( n9253 & n9583 ) | ( n9253 & n9584 ) | ( n9583 & n9584 ) ;
  assign n9586 = ( ~n9253 & n9583 ) | ( ~n9253 & n9584 ) | ( n9583 & n9584 ) ;
  assign n9587 = ( n9253 & ~n9585 ) | ( n9253 & n9586 ) | ( ~n9585 & n9586 ) ;
  assign n9588 = ( x105 & n9582 ) | ( x105 & ~n9587 ) | ( n9582 & ~n9587 ) ;
  assign n9589 = ( x105 & n9254 ) | ( x105 & ~n9343 ) | ( n9254 & ~n9343 ) ;
  assign n9590 = x105 & n9254 ;
  assign n9591 = ( ~n9259 & n9589 ) | ( ~n9259 & n9590 ) | ( n9589 & n9590 ) ;
  assign n9592 = ( n9259 & n9589 ) | ( n9259 & n9590 ) | ( n9589 & n9590 ) ;
  assign n9593 = ( n9259 & n9591 ) | ( n9259 & ~n9592 ) | ( n9591 & ~n9592 ) ;
  assign n9594 = ( x106 & n9588 ) | ( x106 & ~n9593 ) | ( n9588 & ~n9593 ) ;
  assign n9595 = ( x106 & n9260 ) | ( x106 & ~n9343 ) | ( n9260 & ~n9343 ) ;
  assign n9596 = x106 & n9260 ;
  assign n9597 = ( n9265 & n9595 ) | ( n9265 & n9596 ) | ( n9595 & n9596 ) ;
  assign n9598 = ( ~n9265 & n9595 ) | ( ~n9265 & n9596 ) | ( n9595 & n9596 ) ;
  assign n9599 = ( n9265 & ~n9597 ) | ( n9265 & n9598 ) | ( ~n9597 & n9598 ) ;
  assign n9600 = ( x107 & n9594 ) | ( x107 & ~n9599 ) | ( n9594 & ~n9599 ) ;
  assign n9601 = ( x107 & n9266 ) | ( x107 & ~n9343 ) | ( n9266 & ~n9343 ) ;
  assign n9602 = x107 & n9266 ;
  assign n9603 = ( ~n9271 & n9601 ) | ( ~n9271 & n9602 ) | ( n9601 & n9602 ) ;
  assign n9604 = ( n9271 & n9601 ) | ( n9271 & n9602 ) | ( n9601 & n9602 ) ;
  assign n9605 = ( n9271 & n9603 ) | ( n9271 & ~n9604 ) | ( n9603 & ~n9604 ) ;
  assign n9606 = ( x108 & n9600 ) | ( x108 & ~n9605 ) | ( n9600 & ~n9605 ) ;
  assign n9607 = ( x108 & n9272 ) | ( x108 & ~n9343 ) | ( n9272 & ~n9343 ) ;
  assign n9608 = x108 & n9272 ;
  assign n9609 = ( n9277 & n9607 ) | ( n9277 & n9608 ) | ( n9607 & n9608 ) ;
  assign n9610 = ( ~n9277 & n9607 ) | ( ~n9277 & n9608 ) | ( n9607 & n9608 ) ;
  assign n9611 = ( n9277 & ~n9609 ) | ( n9277 & n9610 ) | ( ~n9609 & n9610 ) ;
  assign n9612 = ( x109 & n9606 ) | ( x109 & ~n9611 ) | ( n9606 & ~n9611 ) ;
  assign n9613 = ( x109 & n9278 ) | ( x109 & ~n9343 ) | ( n9278 & ~n9343 ) ;
  assign n9614 = x109 & n9278 ;
  assign n9615 = ( ~n9283 & n9613 ) | ( ~n9283 & n9614 ) | ( n9613 & n9614 ) ;
  assign n9616 = ( n9283 & n9613 ) | ( n9283 & n9614 ) | ( n9613 & n9614 ) ;
  assign n9617 = ( n9283 & n9615 ) | ( n9283 & ~n9616 ) | ( n9615 & ~n9616 ) ;
  assign n9618 = ( x110 & n9612 ) | ( x110 & ~n9617 ) | ( n9612 & ~n9617 ) ;
  assign n9619 = ( x110 & n9284 ) | ( x110 & ~n9343 ) | ( n9284 & ~n9343 ) ;
  assign n9620 = x110 & n9284 ;
  assign n9621 = ( n9289 & n9619 ) | ( n9289 & n9620 ) | ( n9619 & n9620 ) ;
  assign n9622 = ( ~n9289 & n9619 ) | ( ~n9289 & n9620 ) | ( n9619 & n9620 ) ;
  assign n9623 = ( n9289 & ~n9621 ) | ( n9289 & n9622 ) | ( ~n9621 & n9622 ) ;
  assign n9624 = ( x111 & n9618 ) | ( x111 & ~n9623 ) | ( n9618 & ~n9623 ) ;
  assign n9625 = ( x111 & n9290 ) | ( x111 & ~n9343 ) | ( n9290 & ~n9343 ) ;
  assign n9626 = x111 & n9290 ;
  assign n9627 = ( ~n9295 & n9625 ) | ( ~n9295 & n9626 ) | ( n9625 & n9626 ) ;
  assign n9628 = ( n9295 & n9625 ) | ( n9295 & n9626 ) | ( n9625 & n9626 ) ;
  assign n9629 = ( n9295 & n9627 ) | ( n9295 & ~n9628 ) | ( n9627 & ~n9628 ) ;
  assign n9630 = ( x112 & n9624 ) | ( x112 & ~n9629 ) | ( n9624 & ~n9629 ) ;
  assign n9631 = ( x112 & n9296 ) | ( x112 & ~n9343 ) | ( n9296 & ~n9343 ) ;
  assign n9632 = x112 & n9296 ;
  assign n9633 = ( n9301 & n9631 ) | ( n9301 & n9632 ) | ( n9631 & n9632 ) ;
  assign n9634 = ( ~n9301 & n9631 ) | ( ~n9301 & n9632 ) | ( n9631 & n9632 ) ;
  assign n9635 = ( n9301 & ~n9633 ) | ( n9301 & n9634 ) | ( ~n9633 & n9634 ) ;
  assign n9636 = ( x113 & n9630 ) | ( x113 & ~n9635 ) | ( n9630 & ~n9635 ) ;
  assign n9637 = ( x113 & n9302 ) | ( x113 & ~n9343 ) | ( n9302 & ~n9343 ) ;
  assign n9638 = x113 & n9302 ;
  assign n9639 = ( ~n9307 & n9637 ) | ( ~n9307 & n9638 ) | ( n9637 & n9638 ) ;
  assign n9640 = ( n9307 & n9637 ) | ( n9307 & n9638 ) | ( n9637 & n9638 ) ;
  assign n9641 = ( n9307 & n9639 ) | ( n9307 & ~n9640 ) | ( n9639 & ~n9640 ) ;
  assign n9642 = ( x114 & n9636 ) | ( x114 & ~n9641 ) | ( n9636 & ~n9641 ) ;
  assign n9643 = ( x114 & n9308 ) | ( x114 & ~n9343 ) | ( n9308 & ~n9343 ) ;
  assign n9644 = x114 & n9308 ;
  assign n9645 = ( n9313 & n9643 ) | ( n9313 & n9644 ) | ( n9643 & n9644 ) ;
  assign n9646 = ( ~n9313 & n9643 ) | ( ~n9313 & n9644 ) | ( n9643 & n9644 ) ;
  assign n9647 = ( n9313 & ~n9645 ) | ( n9313 & n9646 ) | ( ~n9645 & n9646 ) ;
  assign n9648 = ( x115 & n9642 ) | ( x115 & ~n9647 ) | ( n9642 & ~n9647 ) ;
  assign n9649 = ( x115 & n9314 ) | ( x115 & ~n9343 ) | ( n9314 & ~n9343 ) ;
  assign n9650 = x115 & n9314 ;
  assign n9651 = ( ~n9319 & n9649 ) | ( ~n9319 & n9650 ) | ( n9649 & n9650 ) ;
  assign n9652 = ( n9319 & n9649 ) | ( n9319 & n9650 ) | ( n9649 & n9650 ) ;
  assign n9653 = ( n9319 & n9651 ) | ( n9319 & ~n9652 ) | ( n9651 & ~n9652 ) ;
  assign n9654 = ( x116 & n9648 ) | ( x116 & ~n9653 ) | ( n9648 & ~n9653 ) ;
  assign n9655 = ( x116 & n9320 ) | ( x116 & ~n9343 ) | ( n9320 & ~n9343 ) ;
  assign n9656 = x116 & n9320 ;
  assign n9657 = ( n9325 & n9655 ) | ( n9325 & n9656 ) | ( n9655 & n9656 ) ;
  assign n9658 = ( ~n9325 & n9655 ) | ( ~n9325 & n9656 ) | ( n9655 & n9656 ) ;
  assign n9659 = ( n9325 & ~n9657 ) | ( n9325 & n9658 ) | ( ~n9657 & n9658 ) ;
  assign n9660 = ( x117 & n9654 ) | ( x117 & ~n9659 ) | ( n9654 & ~n9659 ) ;
  assign n9661 = ( x117 & n9326 ) | ( x117 & ~n9343 ) | ( n9326 & ~n9343 ) ;
  assign n9662 = x117 & n9326 ;
  assign n9663 = ( ~n9331 & n9661 ) | ( ~n9331 & n9662 ) | ( n9661 & n9662 ) ;
  assign n9664 = ( n9331 & n9661 ) | ( n9331 & n9662 ) | ( n9661 & n9662 ) ;
  assign n9665 = ( n9331 & n9663 ) | ( n9331 & ~n9664 ) | ( n9663 & ~n9664 ) ;
  assign n9666 = ( x118 & n9660 ) | ( x118 & ~n9665 ) | ( n9660 & ~n9665 ) ;
  assign n9667 = ( x118 & n9332 ) | ( x118 & ~n9343 ) | ( n9332 & ~n9343 ) ;
  assign n9668 = x118 & n9332 ;
  assign n9669 = ( ~n9337 & n9667 ) | ( ~n9337 & n9668 ) | ( n9667 & n9668 ) ;
  assign n9670 = ( n9337 & n9667 ) | ( n9337 & n9668 ) | ( n9667 & n9668 ) ;
  assign n9671 = ( n9337 & n9669 ) | ( n9337 & ~n9670 ) | ( n9669 & ~n9670 ) ;
  assign n9672 = ( x119 & n9666 ) | ( x119 & ~n9671 ) | ( n9666 & ~n9671 ) ;
  assign n9673 = x120 | n9672 ;
  assign n9674 = ( x120 & n137 ) | ( x120 & n9672 ) | ( n137 & n9672 ) ;
  assign n9675 = ( n9341 & ~n9673 ) | ( n9341 & n9674 ) | ( ~n9673 & n9674 ) ;
  assign n9676 = ( x120 & ~n9341 ) | ( x120 & n9672 ) | ( ~n9341 & n9672 ) ;
  assign n9677 = n137 | n9676 ;
  assign n9678 = ( x7 & ~x64 ) | ( x7 & n9677 ) | ( ~x64 & n9677 ) ;
  assign n9679 = ~x7 & n9677 ;
  assign n9680 = ( n9347 & n9678 ) | ( n9347 & ~n9679 ) | ( n9678 & ~n9679 ) ;
  assign n9681 = ~x6 & x64 ;
  assign n9682 = ( x65 & ~n9680 ) | ( x65 & n9681 ) | ( ~n9680 & n9681 ) ;
  assign n9683 = ( x65 & n9347 ) | ( x65 & ~n9677 ) | ( n9347 & ~n9677 ) ;
  assign n9684 = x65 & n9347 ;
  assign n9685 = ( n9346 & n9683 ) | ( n9346 & n9684 ) | ( n9683 & n9684 ) ;
  assign n9686 = ( ~n9346 & n9683 ) | ( ~n9346 & n9684 ) | ( n9683 & n9684 ) ;
  assign n9687 = ( n9346 & ~n9685 ) | ( n9346 & n9686 ) | ( ~n9685 & n9686 ) ;
  assign n9688 = ( x66 & n9682 ) | ( x66 & ~n9687 ) | ( n9682 & ~n9687 ) ;
  assign n9689 = ( x66 & n9348 ) | ( x66 & ~n9677 ) | ( n9348 & ~n9677 ) ;
  assign n9690 = x66 & n9348 ;
  assign n9691 = ( n9353 & n9689 ) | ( n9353 & n9690 ) | ( n9689 & n9690 ) ;
  assign n9692 = ( ~n9353 & n9689 ) | ( ~n9353 & n9690 ) | ( n9689 & n9690 ) ;
  assign n9693 = ( n9353 & ~n9691 ) | ( n9353 & n9692 ) | ( ~n9691 & n9692 ) ;
  assign n9694 = ( x67 & n9688 ) | ( x67 & ~n9693 ) | ( n9688 & ~n9693 ) ;
  assign n9695 = ( x67 & n9354 ) | ( x67 & ~n9677 ) | ( n9354 & ~n9677 ) ;
  assign n9696 = x67 & n9354 ;
  assign n9697 = ( ~n9359 & n9695 ) | ( ~n9359 & n9696 ) | ( n9695 & n9696 ) ;
  assign n9698 = ( n9359 & n9695 ) | ( n9359 & n9696 ) | ( n9695 & n9696 ) ;
  assign n9699 = ( n9359 & n9697 ) | ( n9359 & ~n9698 ) | ( n9697 & ~n9698 ) ;
  assign n9700 = ( x68 & n9694 ) | ( x68 & ~n9699 ) | ( n9694 & ~n9699 ) ;
  assign n9701 = ( x68 & n9360 ) | ( x68 & ~n9677 ) | ( n9360 & ~n9677 ) ;
  assign n9702 = x68 & n9360 ;
  assign n9703 = ( n9365 & n9701 ) | ( n9365 & n9702 ) | ( n9701 & n9702 ) ;
  assign n9704 = ( ~n9365 & n9701 ) | ( ~n9365 & n9702 ) | ( n9701 & n9702 ) ;
  assign n9705 = ( n9365 & ~n9703 ) | ( n9365 & n9704 ) | ( ~n9703 & n9704 ) ;
  assign n9706 = ( x69 & n9700 ) | ( x69 & ~n9705 ) | ( n9700 & ~n9705 ) ;
  assign n9707 = ( x69 & n9366 ) | ( x69 & ~n9677 ) | ( n9366 & ~n9677 ) ;
  assign n9708 = x69 & n9366 ;
  assign n9709 = ( ~n9371 & n9707 ) | ( ~n9371 & n9708 ) | ( n9707 & n9708 ) ;
  assign n9710 = ( n9371 & n9707 ) | ( n9371 & n9708 ) | ( n9707 & n9708 ) ;
  assign n9711 = ( n9371 & n9709 ) | ( n9371 & ~n9710 ) | ( n9709 & ~n9710 ) ;
  assign n9712 = ( x70 & n9706 ) | ( x70 & ~n9711 ) | ( n9706 & ~n9711 ) ;
  assign n9713 = ( x70 & n9372 ) | ( x70 & ~n9677 ) | ( n9372 & ~n9677 ) ;
  assign n9714 = x70 & n9372 ;
  assign n9715 = ( n9377 & n9713 ) | ( n9377 & n9714 ) | ( n9713 & n9714 ) ;
  assign n9716 = ( ~n9377 & n9713 ) | ( ~n9377 & n9714 ) | ( n9713 & n9714 ) ;
  assign n9717 = ( n9377 & ~n9715 ) | ( n9377 & n9716 ) | ( ~n9715 & n9716 ) ;
  assign n9718 = ( x71 & n9712 ) | ( x71 & ~n9717 ) | ( n9712 & ~n9717 ) ;
  assign n9719 = ( x71 & n9378 ) | ( x71 & ~n9677 ) | ( n9378 & ~n9677 ) ;
  assign n9720 = x71 & n9378 ;
  assign n9721 = ( ~n9383 & n9719 ) | ( ~n9383 & n9720 ) | ( n9719 & n9720 ) ;
  assign n9722 = ( n9383 & n9719 ) | ( n9383 & n9720 ) | ( n9719 & n9720 ) ;
  assign n9723 = ( n9383 & n9721 ) | ( n9383 & ~n9722 ) | ( n9721 & ~n9722 ) ;
  assign n9724 = ( x72 & n9718 ) | ( x72 & ~n9723 ) | ( n9718 & ~n9723 ) ;
  assign n9725 = ( x72 & n9384 ) | ( x72 & ~n9677 ) | ( n9384 & ~n9677 ) ;
  assign n9726 = x72 & n9384 ;
  assign n9727 = ( n9389 & n9725 ) | ( n9389 & n9726 ) | ( n9725 & n9726 ) ;
  assign n9728 = ( ~n9389 & n9725 ) | ( ~n9389 & n9726 ) | ( n9725 & n9726 ) ;
  assign n9729 = ( n9389 & ~n9727 ) | ( n9389 & n9728 ) | ( ~n9727 & n9728 ) ;
  assign n9730 = ( x73 & n9724 ) | ( x73 & ~n9729 ) | ( n9724 & ~n9729 ) ;
  assign n9731 = ( x73 & n9390 ) | ( x73 & ~n9677 ) | ( n9390 & ~n9677 ) ;
  assign n9732 = x73 & n9390 ;
  assign n9733 = ( ~n9395 & n9731 ) | ( ~n9395 & n9732 ) | ( n9731 & n9732 ) ;
  assign n9734 = ( n9395 & n9731 ) | ( n9395 & n9732 ) | ( n9731 & n9732 ) ;
  assign n9735 = ( n9395 & n9733 ) | ( n9395 & ~n9734 ) | ( n9733 & ~n9734 ) ;
  assign n9736 = ( x74 & n9730 ) | ( x74 & ~n9735 ) | ( n9730 & ~n9735 ) ;
  assign n9737 = ( x74 & n9396 ) | ( x74 & ~n9677 ) | ( n9396 & ~n9677 ) ;
  assign n9738 = x74 & n9396 ;
  assign n9739 = ( n9401 & n9737 ) | ( n9401 & n9738 ) | ( n9737 & n9738 ) ;
  assign n9740 = ( ~n9401 & n9737 ) | ( ~n9401 & n9738 ) | ( n9737 & n9738 ) ;
  assign n9741 = ( n9401 & ~n9739 ) | ( n9401 & n9740 ) | ( ~n9739 & n9740 ) ;
  assign n9742 = ( x75 & n9736 ) | ( x75 & ~n9741 ) | ( n9736 & ~n9741 ) ;
  assign n9743 = ( x75 & n9402 ) | ( x75 & ~n9677 ) | ( n9402 & ~n9677 ) ;
  assign n9744 = x75 & n9402 ;
  assign n9745 = ( ~n9407 & n9743 ) | ( ~n9407 & n9744 ) | ( n9743 & n9744 ) ;
  assign n9746 = ( n9407 & n9743 ) | ( n9407 & n9744 ) | ( n9743 & n9744 ) ;
  assign n9747 = ( n9407 & n9745 ) | ( n9407 & ~n9746 ) | ( n9745 & ~n9746 ) ;
  assign n9748 = ( x76 & n9742 ) | ( x76 & ~n9747 ) | ( n9742 & ~n9747 ) ;
  assign n9749 = ( x76 & n9408 ) | ( x76 & ~n9677 ) | ( n9408 & ~n9677 ) ;
  assign n9750 = x76 & n9408 ;
  assign n9751 = ( n9413 & n9749 ) | ( n9413 & n9750 ) | ( n9749 & n9750 ) ;
  assign n9752 = ( ~n9413 & n9749 ) | ( ~n9413 & n9750 ) | ( n9749 & n9750 ) ;
  assign n9753 = ( n9413 & ~n9751 ) | ( n9413 & n9752 ) | ( ~n9751 & n9752 ) ;
  assign n9754 = ( x77 & n9748 ) | ( x77 & ~n9753 ) | ( n9748 & ~n9753 ) ;
  assign n9755 = ( x77 & n9414 ) | ( x77 & ~n9677 ) | ( n9414 & ~n9677 ) ;
  assign n9756 = x77 & n9414 ;
  assign n9757 = ( ~n9419 & n9755 ) | ( ~n9419 & n9756 ) | ( n9755 & n9756 ) ;
  assign n9758 = ( n9419 & n9755 ) | ( n9419 & n9756 ) | ( n9755 & n9756 ) ;
  assign n9759 = ( n9419 & n9757 ) | ( n9419 & ~n9758 ) | ( n9757 & ~n9758 ) ;
  assign n9760 = ( x78 & n9754 ) | ( x78 & ~n9759 ) | ( n9754 & ~n9759 ) ;
  assign n9761 = ( x78 & n9420 ) | ( x78 & ~n9677 ) | ( n9420 & ~n9677 ) ;
  assign n9762 = x78 & n9420 ;
  assign n9763 = ( n9425 & n9761 ) | ( n9425 & n9762 ) | ( n9761 & n9762 ) ;
  assign n9764 = ( ~n9425 & n9761 ) | ( ~n9425 & n9762 ) | ( n9761 & n9762 ) ;
  assign n9765 = ( n9425 & ~n9763 ) | ( n9425 & n9764 ) | ( ~n9763 & n9764 ) ;
  assign n9766 = ( x79 & n9760 ) | ( x79 & ~n9765 ) | ( n9760 & ~n9765 ) ;
  assign n9767 = ( x79 & n9426 ) | ( x79 & ~n9677 ) | ( n9426 & ~n9677 ) ;
  assign n9768 = x79 & n9426 ;
  assign n9769 = ( ~n9431 & n9767 ) | ( ~n9431 & n9768 ) | ( n9767 & n9768 ) ;
  assign n9770 = ( n9431 & n9767 ) | ( n9431 & n9768 ) | ( n9767 & n9768 ) ;
  assign n9771 = ( n9431 & n9769 ) | ( n9431 & ~n9770 ) | ( n9769 & ~n9770 ) ;
  assign n9772 = ( x80 & n9766 ) | ( x80 & ~n9771 ) | ( n9766 & ~n9771 ) ;
  assign n9773 = ( x80 & n9432 ) | ( x80 & ~n9677 ) | ( n9432 & ~n9677 ) ;
  assign n9774 = x80 & n9432 ;
  assign n9775 = ( n9437 & n9773 ) | ( n9437 & n9774 ) | ( n9773 & n9774 ) ;
  assign n9776 = ( ~n9437 & n9773 ) | ( ~n9437 & n9774 ) | ( n9773 & n9774 ) ;
  assign n9777 = ( n9437 & ~n9775 ) | ( n9437 & n9776 ) | ( ~n9775 & n9776 ) ;
  assign n9778 = ( x81 & n9772 ) | ( x81 & ~n9777 ) | ( n9772 & ~n9777 ) ;
  assign n9779 = ( x81 & n9438 ) | ( x81 & ~n9677 ) | ( n9438 & ~n9677 ) ;
  assign n9780 = x81 & n9438 ;
  assign n9781 = ( ~n9443 & n9779 ) | ( ~n9443 & n9780 ) | ( n9779 & n9780 ) ;
  assign n9782 = ( n9443 & n9779 ) | ( n9443 & n9780 ) | ( n9779 & n9780 ) ;
  assign n9783 = ( n9443 & n9781 ) | ( n9443 & ~n9782 ) | ( n9781 & ~n9782 ) ;
  assign n9784 = ( x82 & n9778 ) | ( x82 & ~n9783 ) | ( n9778 & ~n9783 ) ;
  assign n9785 = ( x82 & n9444 ) | ( x82 & ~n9677 ) | ( n9444 & ~n9677 ) ;
  assign n9786 = x82 & n9444 ;
  assign n9787 = ( n9449 & n9785 ) | ( n9449 & n9786 ) | ( n9785 & n9786 ) ;
  assign n9788 = ( ~n9449 & n9785 ) | ( ~n9449 & n9786 ) | ( n9785 & n9786 ) ;
  assign n9789 = ( n9449 & ~n9787 ) | ( n9449 & n9788 ) | ( ~n9787 & n9788 ) ;
  assign n9790 = ( x83 & n9784 ) | ( x83 & ~n9789 ) | ( n9784 & ~n9789 ) ;
  assign n9791 = ( x83 & n9450 ) | ( x83 & ~n9677 ) | ( n9450 & ~n9677 ) ;
  assign n9792 = x83 & n9450 ;
  assign n9793 = ( ~n9455 & n9791 ) | ( ~n9455 & n9792 ) | ( n9791 & n9792 ) ;
  assign n9794 = ( n9455 & n9791 ) | ( n9455 & n9792 ) | ( n9791 & n9792 ) ;
  assign n9795 = ( n9455 & n9793 ) | ( n9455 & ~n9794 ) | ( n9793 & ~n9794 ) ;
  assign n9796 = ( x84 & n9790 ) | ( x84 & ~n9795 ) | ( n9790 & ~n9795 ) ;
  assign n9797 = ( x84 & n9456 ) | ( x84 & ~n9677 ) | ( n9456 & ~n9677 ) ;
  assign n9798 = x84 & n9456 ;
  assign n9799 = ( n9461 & n9797 ) | ( n9461 & n9798 ) | ( n9797 & n9798 ) ;
  assign n9800 = ( ~n9461 & n9797 ) | ( ~n9461 & n9798 ) | ( n9797 & n9798 ) ;
  assign n9801 = ( n9461 & ~n9799 ) | ( n9461 & n9800 ) | ( ~n9799 & n9800 ) ;
  assign n9802 = ( x85 & n9796 ) | ( x85 & ~n9801 ) | ( n9796 & ~n9801 ) ;
  assign n9803 = ( x85 & n9462 ) | ( x85 & ~n9677 ) | ( n9462 & ~n9677 ) ;
  assign n9804 = x85 & n9462 ;
  assign n9805 = ( ~n9467 & n9803 ) | ( ~n9467 & n9804 ) | ( n9803 & n9804 ) ;
  assign n9806 = ( n9467 & n9803 ) | ( n9467 & n9804 ) | ( n9803 & n9804 ) ;
  assign n9807 = ( n9467 & n9805 ) | ( n9467 & ~n9806 ) | ( n9805 & ~n9806 ) ;
  assign n9808 = ( x86 & n9802 ) | ( x86 & ~n9807 ) | ( n9802 & ~n9807 ) ;
  assign n9809 = ( x86 & n9468 ) | ( x86 & ~n9677 ) | ( n9468 & ~n9677 ) ;
  assign n9810 = x86 & n9468 ;
  assign n9811 = ( n9473 & n9809 ) | ( n9473 & n9810 ) | ( n9809 & n9810 ) ;
  assign n9812 = ( ~n9473 & n9809 ) | ( ~n9473 & n9810 ) | ( n9809 & n9810 ) ;
  assign n9813 = ( n9473 & ~n9811 ) | ( n9473 & n9812 ) | ( ~n9811 & n9812 ) ;
  assign n9814 = ( x87 & n9808 ) | ( x87 & ~n9813 ) | ( n9808 & ~n9813 ) ;
  assign n9815 = ( x87 & n9474 ) | ( x87 & ~n9677 ) | ( n9474 & ~n9677 ) ;
  assign n9816 = x87 & n9474 ;
  assign n9817 = ( ~n9479 & n9815 ) | ( ~n9479 & n9816 ) | ( n9815 & n9816 ) ;
  assign n9818 = ( n9479 & n9815 ) | ( n9479 & n9816 ) | ( n9815 & n9816 ) ;
  assign n9819 = ( n9479 & n9817 ) | ( n9479 & ~n9818 ) | ( n9817 & ~n9818 ) ;
  assign n9820 = ( x88 & n9814 ) | ( x88 & ~n9819 ) | ( n9814 & ~n9819 ) ;
  assign n9821 = ( x88 & n9480 ) | ( x88 & ~n9677 ) | ( n9480 & ~n9677 ) ;
  assign n9822 = x88 & n9480 ;
  assign n9823 = ( n9485 & n9821 ) | ( n9485 & n9822 ) | ( n9821 & n9822 ) ;
  assign n9824 = ( ~n9485 & n9821 ) | ( ~n9485 & n9822 ) | ( n9821 & n9822 ) ;
  assign n9825 = ( n9485 & ~n9823 ) | ( n9485 & n9824 ) | ( ~n9823 & n9824 ) ;
  assign n9826 = ( x89 & n9820 ) | ( x89 & ~n9825 ) | ( n9820 & ~n9825 ) ;
  assign n9827 = ( x89 & n9486 ) | ( x89 & ~n9677 ) | ( n9486 & ~n9677 ) ;
  assign n9828 = x89 & n9486 ;
  assign n9829 = ( ~n9491 & n9827 ) | ( ~n9491 & n9828 ) | ( n9827 & n9828 ) ;
  assign n9830 = ( n9491 & n9827 ) | ( n9491 & n9828 ) | ( n9827 & n9828 ) ;
  assign n9831 = ( n9491 & n9829 ) | ( n9491 & ~n9830 ) | ( n9829 & ~n9830 ) ;
  assign n9832 = ( x90 & n9826 ) | ( x90 & ~n9831 ) | ( n9826 & ~n9831 ) ;
  assign n9833 = ( x90 & n9492 ) | ( x90 & ~n9677 ) | ( n9492 & ~n9677 ) ;
  assign n9834 = x90 & n9492 ;
  assign n9835 = ( n9497 & n9833 ) | ( n9497 & n9834 ) | ( n9833 & n9834 ) ;
  assign n9836 = ( ~n9497 & n9833 ) | ( ~n9497 & n9834 ) | ( n9833 & n9834 ) ;
  assign n9837 = ( n9497 & ~n9835 ) | ( n9497 & n9836 ) | ( ~n9835 & n9836 ) ;
  assign n9838 = ( x91 & n9832 ) | ( x91 & ~n9837 ) | ( n9832 & ~n9837 ) ;
  assign n9839 = ( x91 & n9498 ) | ( x91 & ~n9677 ) | ( n9498 & ~n9677 ) ;
  assign n9840 = x91 & n9498 ;
  assign n9841 = ( ~n9503 & n9839 ) | ( ~n9503 & n9840 ) | ( n9839 & n9840 ) ;
  assign n9842 = ( n9503 & n9839 ) | ( n9503 & n9840 ) | ( n9839 & n9840 ) ;
  assign n9843 = ( n9503 & n9841 ) | ( n9503 & ~n9842 ) | ( n9841 & ~n9842 ) ;
  assign n9844 = ( x92 & n9838 ) | ( x92 & ~n9843 ) | ( n9838 & ~n9843 ) ;
  assign n9845 = ( x92 & n9504 ) | ( x92 & ~n9677 ) | ( n9504 & ~n9677 ) ;
  assign n9846 = x92 & n9504 ;
  assign n9847 = ( n9509 & n9845 ) | ( n9509 & n9846 ) | ( n9845 & n9846 ) ;
  assign n9848 = ( ~n9509 & n9845 ) | ( ~n9509 & n9846 ) | ( n9845 & n9846 ) ;
  assign n9849 = ( n9509 & ~n9847 ) | ( n9509 & n9848 ) | ( ~n9847 & n9848 ) ;
  assign n9850 = ( x93 & n9844 ) | ( x93 & ~n9849 ) | ( n9844 & ~n9849 ) ;
  assign n9851 = ( x93 & n9510 ) | ( x93 & ~n9677 ) | ( n9510 & ~n9677 ) ;
  assign n9852 = x93 & n9510 ;
  assign n9853 = ( ~n9515 & n9851 ) | ( ~n9515 & n9852 ) | ( n9851 & n9852 ) ;
  assign n9854 = ( n9515 & n9851 ) | ( n9515 & n9852 ) | ( n9851 & n9852 ) ;
  assign n9855 = ( n9515 & n9853 ) | ( n9515 & ~n9854 ) | ( n9853 & ~n9854 ) ;
  assign n9856 = ( x94 & n9850 ) | ( x94 & ~n9855 ) | ( n9850 & ~n9855 ) ;
  assign n9857 = ( x94 & n9516 ) | ( x94 & ~n9677 ) | ( n9516 & ~n9677 ) ;
  assign n9858 = x94 & n9516 ;
  assign n9859 = ( n9521 & n9857 ) | ( n9521 & n9858 ) | ( n9857 & n9858 ) ;
  assign n9860 = ( ~n9521 & n9857 ) | ( ~n9521 & n9858 ) | ( n9857 & n9858 ) ;
  assign n9861 = ( n9521 & ~n9859 ) | ( n9521 & n9860 ) | ( ~n9859 & n9860 ) ;
  assign n9862 = ( x95 & n9856 ) | ( x95 & ~n9861 ) | ( n9856 & ~n9861 ) ;
  assign n9863 = ( x95 & n9522 ) | ( x95 & ~n9677 ) | ( n9522 & ~n9677 ) ;
  assign n9864 = x95 & n9522 ;
  assign n9865 = ( ~n9527 & n9863 ) | ( ~n9527 & n9864 ) | ( n9863 & n9864 ) ;
  assign n9866 = ( n9527 & n9863 ) | ( n9527 & n9864 ) | ( n9863 & n9864 ) ;
  assign n9867 = ( n9527 & n9865 ) | ( n9527 & ~n9866 ) | ( n9865 & ~n9866 ) ;
  assign n9868 = ( x96 & n9862 ) | ( x96 & ~n9867 ) | ( n9862 & ~n9867 ) ;
  assign n9869 = ( x96 & n9528 ) | ( x96 & ~n9677 ) | ( n9528 & ~n9677 ) ;
  assign n9870 = x96 & n9528 ;
  assign n9871 = ( n9533 & n9869 ) | ( n9533 & n9870 ) | ( n9869 & n9870 ) ;
  assign n9872 = ( ~n9533 & n9869 ) | ( ~n9533 & n9870 ) | ( n9869 & n9870 ) ;
  assign n9873 = ( n9533 & ~n9871 ) | ( n9533 & n9872 ) | ( ~n9871 & n9872 ) ;
  assign n9874 = ( x97 & n9868 ) | ( x97 & ~n9873 ) | ( n9868 & ~n9873 ) ;
  assign n9875 = ( x97 & n9534 ) | ( x97 & ~n9677 ) | ( n9534 & ~n9677 ) ;
  assign n9876 = x97 & n9534 ;
  assign n9877 = ( ~n9539 & n9875 ) | ( ~n9539 & n9876 ) | ( n9875 & n9876 ) ;
  assign n9878 = ( n9539 & n9875 ) | ( n9539 & n9876 ) | ( n9875 & n9876 ) ;
  assign n9879 = ( n9539 & n9877 ) | ( n9539 & ~n9878 ) | ( n9877 & ~n9878 ) ;
  assign n9880 = ( x98 & n9874 ) | ( x98 & ~n9879 ) | ( n9874 & ~n9879 ) ;
  assign n9881 = ( x98 & n9540 ) | ( x98 & ~n9677 ) | ( n9540 & ~n9677 ) ;
  assign n9882 = x98 & n9540 ;
  assign n9883 = ( n9545 & n9881 ) | ( n9545 & n9882 ) | ( n9881 & n9882 ) ;
  assign n9884 = ( ~n9545 & n9881 ) | ( ~n9545 & n9882 ) | ( n9881 & n9882 ) ;
  assign n9885 = ( n9545 & ~n9883 ) | ( n9545 & n9884 ) | ( ~n9883 & n9884 ) ;
  assign n9886 = ( x99 & n9880 ) | ( x99 & ~n9885 ) | ( n9880 & ~n9885 ) ;
  assign n9887 = ( x99 & n9546 ) | ( x99 & ~n9677 ) | ( n9546 & ~n9677 ) ;
  assign n9888 = x99 & n9546 ;
  assign n9889 = ( ~n9551 & n9887 ) | ( ~n9551 & n9888 ) | ( n9887 & n9888 ) ;
  assign n9890 = ( n9551 & n9887 ) | ( n9551 & n9888 ) | ( n9887 & n9888 ) ;
  assign n9891 = ( n9551 & n9889 ) | ( n9551 & ~n9890 ) | ( n9889 & ~n9890 ) ;
  assign n9892 = ( x100 & n9886 ) | ( x100 & ~n9891 ) | ( n9886 & ~n9891 ) ;
  assign n9893 = ( x100 & n9552 ) | ( x100 & ~n9677 ) | ( n9552 & ~n9677 ) ;
  assign n9894 = x100 & n9552 ;
  assign n9895 = ( n9557 & n9893 ) | ( n9557 & n9894 ) | ( n9893 & n9894 ) ;
  assign n9896 = ( ~n9557 & n9893 ) | ( ~n9557 & n9894 ) | ( n9893 & n9894 ) ;
  assign n9897 = ( n9557 & ~n9895 ) | ( n9557 & n9896 ) | ( ~n9895 & n9896 ) ;
  assign n9898 = ( x101 & n9892 ) | ( x101 & ~n9897 ) | ( n9892 & ~n9897 ) ;
  assign n9899 = ( x101 & n9558 ) | ( x101 & ~n9677 ) | ( n9558 & ~n9677 ) ;
  assign n9900 = x101 & n9558 ;
  assign n9901 = ( ~n9563 & n9899 ) | ( ~n9563 & n9900 ) | ( n9899 & n9900 ) ;
  assign n9902 = ( n9563 & n9899 ) | ( n9563 & n9900 ) | ( n9899 & n9900 ) ;
  assign n9903 = ( n9563 & n9901 ) | ( n9563 & ~n9902 ) | ( n9901 & ~n9902 ) ;
  assign n9904 = ( x102 & n9898 ) | ( x102 & ~n9903 ) | ( n9898 & ~n9903 ) ;
  assign n9905 = ( x102 & n9564 ) | ( x102 & ~n9677 ) | ( n9564 & ~n9677 ) ;
  assign n9906 = x102 & n9564 ;
  assign n9907 = ( n9569 & n9905 ) | ( n9569 & n9906 ) | ( n9905 & n9906 ) ;
  assign n9908 = ( ~n9569 & n9905 ) | ( ~n9569 & n9906 ) | ( n9905 & n9906 ) ;
  assign n9909 = ( n9569 & ~n9907 ) | ( n9569 & n9908 ) | ( ~n9907 & n9908 ) ;
  assign n9910 = ( x103 & n9904 ) | ( x103 & ~n9909 ) | ( n9904 & ~n9909 ) ;
  assign n9911 = ( x103 & n9570 ) | ( x103 & ~n9677 ) | ( n9570 & ~n9677 ) ;
  assign n9912 = x103 & n9570 ;
  assign n9913 = ( ~n9575 & n9911 ) | ( ~n9575 & n9912 ) | ( n9911 & n9912 ) ;
  assign n9914 = ( n9575 & n9911 ) | ( n9575 & n9912 ) | ( n9911 & n9912 ) ;
  assign n9915 = ( n9575 & n9913 ) | ( n9575 & ~n9914 ) | ( n9913 & ~n9914 ) ;
  assign n9916 = ( x104 & n9910 ) | ( x104 & ~n9915 ) | ( n9910 & ~n9915 ) ;
  assign n9917 = ( x104 & n9576 ) | ( x104 & ~n9677 ) | ( n9576 & ~n9677 ) ;
  assign n9918 = x104 & n9576 ;
  assign n9919 = ( n9581 & n9917 ) | ( n9581 & n9918 ) | ( n9917 & n9918 ) ;
  assign n9920 = ( ~n9581 & n9917 ) | ( ~n9581 & n9918 ) | ( n9917 & n9918 ) ;
  assign n9921 = ( n9581 & ~n9919 ) | ( n9581 & n9920 ) | ( ~n9919 & n9920 ) ;
  assign n9922 = ( x105 & n9916 ) | ( x105 & ~n9921 ) | ( n9916 & ~n9921 ) ;
  assign n9923 = ( x105 & n9582 ) | ( x105 & ~n9677 ) | ( n9582 & ~n9677 ) ;
  assign n9924 = x105 & n9582 ;
  assign n9925 = ( ~n9587 & n9923 ) | ( ~n9587 & n9924 ) | ( n9923 & n9924 ) ;
  assign n9926 = ( n9587 & n9923 ) | ( n9587 & n9924 ) | ( n9923 & n9924 ) ;
  assign n9927 = ( n9587 & n9925 ) | ( n9587 & ~n9926 ) | ( n9925 & ~n9926 ) ;
  assign n9928 = ( x106 & n9922 ) | ( x106 & ~n9927 ) | ( n9922 & ~n9927 ) ;
  assign n9929 = ( x106 & n9588 ) | ( x106 & ~n9677 ) | ( n9588 & ~n9677 ) ;
  assign n9930 = x106 & n9588 ;
  assign n9931 = ( n9593 & n9929 ) | ( n9593 & n9930 ) | ( n9929 & n9930 ) ;
  assign n9932 = ( ~n9593 & n9929 ) | ( ~n9593 & n9930 ) | ( n9929 & n9930 ) ;
  assign n9933 = ( n9593 & ~n9931 ) | ( n9593 & n9932 ) | ( ~n9931 & n9932 ) ;
  assign n9934 = ( x107 & n9928 ) | ( x107 & ~n9933 ) | ( n9928 & ~n9933 ) ;
  assign n9935 = ( x107 & n9594 ) | ( x107 & ~n9677 ) | ( n9594 & ~n9677 ) ;
  assign n9936 = x107 & n9594 ;
  assign n9937 = ( ~n9599 & n9935 ) | ( ~n9599 & n9936 ) | ( n9935 & n9936 ) ;
  assign n9938 = ( n9599 & n9935 ) | ( n9599 & n9936 ) | ( n9935 & n9936 ) ;
  assign n9939 = ( n9599 & n9937 ) | ( n9599 & ~n9938 ) | ( n9937 & ~n9938 ) ;
  assign n9940 = ( x108 & n9934 ) | ( x108 & ~n9939 ) | ( n9934 & ~n9939 ) ;
  assign n9941 = ( x108 & n9600 ) | ( x108 & ~n9677 ) | ( n9600 & ~n9677 ) ;
  assign n9942 = x108 & n9600 ;
  assign n9943 = ( n9605 & n9941 ) | ( n9605 & n9942 ) | ( n9941 & n9942 ) ;
  assign n9944 = ( ~n9605 & n9941 ) | ( ~n9605 & n9942 ) | ( n9941 & n9942 ) ;
  assign n9945 = ( n9605 & ~n9943 ) | ( n9605 & n9944 ) | ( ~n9943 & n9944 ) ;
  assign n9946 = ( x109 & n9940 ) | ( x109 & ~n9945 ) | ( n9940 & ~n9945 ) ;
  assign n9947 = ( x109 & n9606 ) | ( x109 & ~n9677 ) | ( n9606 & ~n9677 ) ;
  assign n9948 = x109 & n9606 ;
  assign n9949 = ( ~n9611 & n9947 ) | ( ~n9611 & n9948 ) | ( n9947 & n9948 ) ;
  assign n9950 = ( n9611 & n9947 ) | ( n9611 & n9948 ) | ( n9947 & n9948 ) ;
  assign n9951 = ( n9611 & n9949 ) | ( n9611 & ~n9950 ) | ( n9949 & ~n9950 ) ;
  assign n9952 = ( x110 & n9946 ) | ( x110 & ~n9951 ) | ( n9946 & ~n9951 ) ;
  assign n9953 = ( x110 & n9612 ) | ( x110 & ~n9677 ) | ( n9612 & ~n9677 ) ;
  assign n9954 = x110 & n9612 ;
  assign n9955 = ( n9617 & n9953 ) | ( n9617 & n9954 ) | ( n9953 & n9954 ) ;
  assign n9956 = ( ~n9617 & n9953 ) | ( ~n9617 & n9954 ) | ( n9953 & n9954 ) ;
  assign n9957 = ( n9617 & ~n9955 ) | ( n9617 & n9956 ) | ( ~n9955 & n9956 ) ;
  assign n9958 = ( x111 & n9952 ) | ( x111 & ~n9957 ) | ( n9952 & ~n9957 ) ;
  assign n9959 = ( x111 & n9618 ) | ( x111 & ~n9677 ) | ( n9618 & ~n9677 ) ;
  assign n9960 = x111 & n9618 ;
  assign n9961 = ( ~n9623 & n9959 ) | ( ~n9623 & n9960 ) | ( n9959 & n9960 ) ;
  assign n9962 = ( n9623 & n9959 ) | ( n9623 & n9960 ) | ( n9959 & n9960 ) ;
  assign n9963 = ( n9623 & n9961 ) | ( n9623 & ~n9962 ) | ( n9961 & ~n9962 ) ;
  assign n9964 = ( x112 & n9958 ) | ( x112 & ~n9963 ) | ( n9958 & ~n9963 ) ;
  assign n9965 = ( x112 & n9624 ) | ( x112 & ~n9677 ) | ( n9624 & ~n9677 ) ;
  assign n9966 = x112 & n9624 ;
  assign n9967 = ( n9629 & n9965 ) | ( n9629 & n9966 ) | ( n9965 & n9966 ) ;
  assign n9968 = ( ~n9629 & n9965 ) | ( ~n9629 & n9966 ) | ( n9965 & n9966 ) ;
  assign n9969 = ( n9629 & ~n9967 ) | ( n9629 & n9968 ) | ( ~n9967 & n9968 ) ;
  assign n9970 = ( x113 & n9964 ) | ( x113 & ~n9969 ) | ( n9964 & ~n9969 ) ;
  assign n9971 = ( x113 & n9630 ) | ( x113 & ~n9677 ) | ( n9630 & ~n9677 ) ;
  assign n9972 = x113 & n9630 ;
  assign n9973 = ( ~n9635 & n9971 ) | ( ~n9635 & n9972 ) | ( n9971 & n9972 ) ;
  assign n9974 = ( n9635 & n9971 ) | ( n9635 & n9972 ) | ( n9971 & n9972 ) ;
  assign n9975 = ( n9635 & n9973 ) | ( n9635 & ~n9974 ) | ( n9973 & ~n9974 ) ;
  assign n9976 = ( x114 & n9970 ) | ( x114 & ~n9975 ) | ( n9970 & ~n9975 ) ;
  assign n9977 = ( x114 & n9636 ) | ( x114 & ~n9677 ) | ( n9636 & ~n9677 ) ;
  assign n9978 = x114 & n9636 ;
  assign n9979 = ( n9641 & n9977 ) | ( n9641 & n9978 ) | ( n9977 & n9978 ) ;
  assign n9980 = ( ~n9641 & n9977 ) | ( ~n9641 & n9978 ) | ( n9977 & n9978 ) ;
  assign n9981 = ( n9641 & ~n9979 ) | ( n9641 & n9980 ) | ( ~n9979 & n9980 ) ;
  assign n9982 = ( x115 & n9976 ) | ( x115 & ~n9981 ) | ( n9976 & ~n9981 ) ;
  assign n9983 = ( x115 & n9642 ) | ( x115 & ~n9677 ) | ( n9642 & ~n9677 ) ;
  assign n9984 = x115 & n9642 ;
  assign n9985 = ( ~n9647 & n9983 ) | ( ~n9647 & n9984 ) | ( n9983 & n9984 ) ;
  assign n9986 = ( n9647 & n9983 ) | ( n9647 & n9984 ) | ( n9983 & n9984 ) ;
  assign n9987 = ( n9647 & n9985 ) | ( n9647 & ~n9986 ) | ( n9985 & ~n9986 ) ;
  assign n9988 = ( x116 & n9982 ) | ( x116 & ~n9987 ) | ( n9982 & ~n9987 ) ;
  assign n9989 = ( x116 & n9648 ) | ( x116 & ~n9677 ) | ( n9648 & ~n9677 ) ;
  assign n9990 = x116 & n9648 ;
  assign n9991 = ( n9653 & n9989 ) | ( n9653 & n9990 ) | ( n9989 & n9990 ) ;
  assign n9992 = ( ~n9653 & n9989 ) | ( ~n9653 & n9990 ) | ( n9989 & n9990 ) ;
  assign n9993 = ( n9653 & ~n9991 ) | ( n9653 & n9992 ) | ( ~n9991 & n9992 ) ;
  assign n9994 = ( x117 & n9988 ) | ( x117 & ~n9993 ) | ( n9988 & ~n9993 ) ;
  assign n9995 = ( x117 & n9654 ) | ( x117 & ~n9677 ) | ( n9654 & ~n9677 ) ;
  assign n9996 = x117 & n9654 ;
  assign n9997 = ( ~n9659 & n9995 ) | ( ~n9659 & n9996 ) | ( n9995 & n9996 ) ;
  assign n9998 = ( n9659 & n9995 ) | ( n9659 & n9996 ) | ( n9995 & n9996 ) ;
  assign n9999 = ( n9659 & n9997 ) | ( n9659 & ~n9998 ) | ( n9997 & ~n9998 ) ;
  assign n10000 = ( x118 & n9994 ) | ( x118 & ~n9999 ) | ( n9994 & ~n9999 ) ;
  assign n10001 = ( x118 & n9660 ) | ( x118 & ~n9677 ) | ( n9660 & ~n9677 ) ;
  assign n10002 = x118 & n9660 ;
  assign n10003 = ( n9665 & n10001 ) | ( n9665 & n10002 ) | ( n10001 & n10002 ) ;
  assign n10004 = ( ~n9665 & n10001 ) | ( ~n9665 & n10002 ) | ( n10001 & n10002 ) ;
  assign n10005 = ( n9665 & ~n10003 ) | ( n9665 & n10004 ) | ( ~n10003 & n10004 ) ;
  assign n10006 = ( x119 & n10000 ) | ( x119 & ~n10005 ) | ( n10000 & ~n10005 ) ;
  assign n10007 = ( x119 & n9666 ) | ( x119 & ~n9677 ) | ( n9666 & ~n9677 ) ;
  assign n10008 = x119 & n9666 ;
  assign n10009 = ( n9671 & n10007 ) | ( n9671 & n10008 ) | ( n10007 & n10008 ) ;
  assign n10010 = ( ~n9671 & n10007 ) | ( ~n9671 & n10008 ) | ( n10007 & n10008 ) ;
  assign n10011 = ( n9671 & ~n10009 ) | ( n9671 & n10010 ) | ( ~n10009 & n10010 ) ;
  assign n10012 = ( x120 & n10006 ) | ( x120 & ~n10011 ) | ( n10006 & ~n10011 ) ;
  assign n10013 = x121 | n10012 ;
  assign n10014 = ( x121 & n136 ) | ( x121 & n10012 ) | ( n136 & n10012 ) ;
  assign n10015 = ( n9675 & ~n10013 ) | ( n9675 & n10014 ) | ( ~n10013 & n10014 ) ;
  assign n10016 = ( x121 & ~n9675 ) | ( x121 & n10012 ) | ( ~n9675 & n10012 ) ;
  assign n10017 = n136 | n10016 ;
  assign n10018 = ( x6 & ~x64 ) | ( x6 & n10017 ) | ( ~x64 & n10017 ) ;
  assign n10019 = ~x6 & n10017 ;
  assign n10020 = ( n9681 & n10018 ) | ( n9681 & ~n10019 ) | ( n10018 & ~n10019 ) ;
  assign n10021 = ~x5 & x64 ;
  assign n10022 = ( x65 & ~n10020 ) | ( x65 & n10021 ) | ( ~n10020 & n10021 ) ;
  assign n10023 = ( x65 & n9681 ) | ( x65 & ~n10017 ) | ( n9681 & ~n10017 ) ;
  assign n10024 = x65 & n9681 ;
  assign n10025 = ( n9680 & n10023 ) | ( n9680 & n10024 ) | ( n10023 & n10024 ) ;
  assign n10026 = ( ~n9680 & n10023 ) | ( ~n9680 & n10024 ) | ( n10023 & n10024 ) ;
  assign n10027 = ( n9680 & ~n10025 ) | ( n9680 & n10026 ) | ( ~n10025 & n10026 ) ;
  assign n10028 = ( x66 & n10022 ) | ( x66 & ~n10027 ) | ( n10022 & ~n10027 ) ;
  assign n10029 = ( x66 & n9682 ) | ( x66 & ~n10017 ) | ( n9682 & ~n10017 ) ;
  assign n10030 = x66 & n9682 ;
  assign n10031 = ( n9687 & n10029 ) | ( n9687 & n10030 ) | ( n10029 & n10030 ) ;
  assign n10032 = ( ~n9687 & n10029 ) | ( ~n9687 & n10030 ) | ( n10029 & n10030 ) ;
  assign n10033 = ( n9687 & ~n10031 ) | ( n9687 & n10032 ) | ( ~n10031 & n10032 ) ;
  assign n10034 = ( x67 & n10028 ) | ( x67 & ~n10033 ) | ( n10028 & ~n10033 ) ;
  assign n10035 = ( x67 & n9688 ) | ( x67 & ~n10017 ) | ( n9688 & ~n10017 ) ;
  assign n10036 = x67 & n9688 ;
  assign n10037 = ( ~n9693 & n10035 ) | ( ~n9693 & n10036 ) | ( n10035 & n10036 ) ;
  assign n10038 = ( n9693 & n10035 ) | ( n9693 & n10036 ) | ( n10035 & n10036 ) ;
  assign n10039 = ( n9693 & n10037 ) | ( n9693 & ~n10038 ) | ( n10037 & ~n10038 ) ;
  assign n10040 = ( x68 & n10034 ) | ( x68 & ~n10039 ) | ( n10034 & ~n10039 ) ;
  assign n10041 = ( x68 & n9694 ) | ( x68 & ~n10017 ) | ( n9694 & ~n10017 ) ;
  assign n10042 = x68 & n9694 ;
  assign n10043 = ( n9699 & n10041 ) | ( n9699 & n10042 ) | ( n10041 & n10042 ) ;
  assign n10044 = ( ~n9699 & n10041 ) | ( ~n9699 & n10042 ) | ( n10041 & n10042 ) ;
  assign n10045 = ( n9699 & ~n10043 ) | ( n9699 & n10044 ) | ( ~n10043 & n10044 ) ;
  assign n10046 = ( x69 & n10040 ) | ( x69 & ~n10045 ) | ( n10040 & ~n10045 ) ;
  assign n10047 = ( x69 & n9700 ) | ( x69 & ~n10017 ) | ( n9700 & ~n10017 ) ;
  assign n10048 = x69 & n9700 ;
  assign n10049 = ( ~n9705 & n10047 ) | ( ~n9705 & n10048 ) | ( n10047 & n10048 ) ;
  assign n10050 = ( n9705 & n10047 ) | ( n9705 & n10048 ) | ( n10047 & n10048 ) ;
  assign n10051 = ( n9705 & n10049 ) | ( n9705 & ~n10050 ) | ( n10049 & ~n10050 ) ;
  assign n10052 = ( x70 & n10046 ) | ( x70 & ~n10051 ) | ( n10046 & ~n10051 ) ;
  assign n10053 = ( x70 & n9706 ) | ( x70 & ~n10017 ) | ( n9706 & ~n10017 ) ;
  assign n10054 = x70 & n9706 ;
  assign n10055 = ( n9711 & n10053 ) | ( n9711 & n10054 ) | ( n10053 & n10054 ) ;
  assign n10056 = ( ~n9711 & n10053 ) | ( ~n9711 & n10054 ) | ( n10053 & n10054 ) ;
  assign n10057 = ( n9711 & ~n10055 ) | ( n9711 & n10056 ) | ( ~n10055 & n10056 ) ;
  assign n10058 = ( x71 & n10052 ) | ( x71 & ~n10057 ) | ( n10052 & ~n10057 ) ;
  assign n10059 = ( x71 & n9712 ) | ( x71 & ~n10017 ) | ( n9712 & ~n10017 ) ;
  assign n10060 = x71 & n9712 ;
  assign n10061 = ( ~n9717 & n10059 ) | ( ~n9717 & n10060 ) | ( n10059 & n10060 ) ;
  assign n10062 = ( n9717 & n10059 ) | ( n9717 & n10060 ) | ( n10059 & n10060 ) ;
  assign n10063 = ( n9717 & n10061 ) | ( n9717 & ~n10062 ) | ( n10061 & ~n10062 ) ;
  assign n10064 = ( x72 & n10058 ) | ( x72 & ~n10063 ) | ( n10058 & ~n10063 ) ;
  assign n10065 = ( x72 & n9718 ) | ( x72 & ~n10017 ) | ( n9718 & ~n10017 ) ;
  assign n10066 = x72 & n9718 ;
  assign n10067 = ( n9723 & n10065 ) | ( n9723 & n10066 ) | ( n10065 & n10066 ) ;
  assign n10068 = ( ~n9723 & n10065 ) | ( ~n9723 & n10066 ) | ( n10065 & n10066 ) ;
  assign n10069 = ( n9723 & ~n10067 ) | ( n9723 & n10068 ) | ( ~n10067 & n10068 ) ;
  assign n10070 = ( x73 & n10064 ) | ( x73 & ~n10069 ) | ( n10064 & ~n10069 ) ;
  assign n10071 = ( x73 & n9724 ) | ( x73 & ~n10017 ) | ( n9724 & ~n10017 ) ;
  assign n10072 = x73 & n9724 ;
  assign n10073 = ( ~n9729 & n10071 ) | ( ~n9729 & n10072 ) | ( n10071 & n10072 ) ;
  assign n10074 = ( n9729 & n10071 ) | ( n9729 & n10072 ) | ( n10071 & n10072 ) ;
  assign n10075 = ( n9729 & n10073 ) | ( n9729 & ~n10074 ) | ( n10073 & ~n10074 ) ;
  assign n10076 = ( x74 & n10070 ) | ( x74 & ~n10075 ) | ( n10070 & ~n10075 ) ;
  assign n10077 = ( x74 & n9730 ) | ( x74 & ~n10017 ) | ( n9730 & ~n10017 ) ;
  assign n10078 = x74 & n9730 ;
  assign n10079 = ( n9735 & n10077 ) | ( n9735 & n10078 ) | ( n10077 & n10078 ) ;
  assign n10080 = ( ~n9735 & n10077 ) | ( ~n9735 & n10078 ) | ( n10077 & n10078 ) ;
  assign n10081 = ( n9735 & ~n10079 ) | ( n9735 & n10080 ) | ( ~n10079 & n10080 ) ;
  assign n10082 = ( x75 & n10076 ) | ( x75 & ~n10081 ) | ( n10076 & ~n10081 ) ;
  assign n10083 = ( x75 & n9736 ) | ( x75 & ~n10017 ) | ( n9736 & ~n10017 ) ;
  assign n10084 = x75 & n9736 ;
  assign n10085 = ( ~n9741 & n10083 ) | ( ~n9741 & n10084 ) | ( n10083 & n10084 ) ;
  assign n10086 = ( n9741 & n10083 ) | ( n9741 & n10084 ) | ( n10083 & n10084 ) ;
  assign n10087 = ( n9741 & n10085 ) | ( n9741 & ~n10086 ) | ( n10085 & ~n10086 ) ;
  assign n10088 = ( x76 & n10082 ) | ( x76 & ~n10087 ) | ( n10082 & ~n10087 ) ;
  assign n10089 = ( x76 & n9742 ) | ( x76 & ~n10017 ) | ( n9742 & ~n10017 ) ;
  assign n10090 = x76 & n9742 ;
  assign n10091 = ( n9747 & n10089 ) | ( n9747 & n10090 ) | ( n10089 & n10090 ) ;
  assign n10092 = ( ~n9747 & n10089 ) | ( ~n9747 & n10090 ) | ( n10089 & n10090 ) ;
  assign n10093 = ( n9747 & ~n10091 ) | ( n9747 & n10092 ) | ( ~n10091 & n10092 ) ;
  assign n10094 = ( x77 & n10088 ) | ( x77 & ~n10093 ) | ( n10088 & ~n10093 ) ;
  assign n10095 = ( x77 & n9748 ) | ( x77 & ~n10017 ) | ( n9748 & ~n10017 ) ;
  assign n10096 = x77 & n9748 ;
  assign n10097 = ( ~n9753 & n10095 ) | ( ~n9753 & n10096 ) | ( n10095 & n10096 ) ;
  assign n10098 = ( n9753 & n10095 ) | ( n9753 & n10096 ) | ( n10095 & n10096 ) ;
  assign n10099 = ( n9753 & n10097 ) | ( n9753 & ~n10098 ) | ( n10097 & ~n10098 ) ;
  assign n10100 = ( x78 & n10094 ) | ( x78 & ~n10099 ) | ( n10094 & ~n10099 ) ;
  assign n10101 = ( x78 & n9754 ) | ( x78 & ~n10017 ) | ( n9754 & ~n10017 ) ;
  assign n10102 = x78 & n9754 ;
  assign n10103 = ( n9759 & n10101 ) | ( n9759 & n10102 ) | ( n10101 & n10102 ) ;
  assign n10104 = ( ~n9759 & n10101 ) | ( ~n9759 & n10102 ) | ( n10101 & n10102 ) ;
  assign n10105 = ( n9759 & ~n10103 ) | ( n9759 & n10104 ) | ( ~n10103 & n10104 ) ;
  assign n10106 = ( x79 & n10100 ) | ( x79 & ~n10105 ) | ( n10100 & ~n10105 ) ;
  assign n10107 = ( x79 & n9760 ) | ( x79 & ~n10017 ) | ( n9760 & ~n10017 ) ;
  assign n10108 = x79 & n9760 ;
  assign n10109 = ( ~n9765 & n10107 ) | ( ~n9765 & n10108 ) | ( n10107 & n10108 ) ;
  assign n10110 = ( n9765 & n10107 ) | ( n9765 & n10108 ) | ( n10107 & n10108 ) ;
  assign n10111 = ( n9765 & n10109 ) | ( n9765 & ~n10110 ) | ( n10109 & ~n10110 ) ;
  assign n10112 = ( x80 & n10106 ) | ( x80 & ~n10111 ) | ( n10106 & ~n10111 ) ;
  assign n10113 = ( x80 & n9766 ) | ( x80 & ~n10017 ) | ( n9766 & ~n10017 ) ;
  assign n10114 = x80 & n9766 ;
  assign n10115 = ( n9771 & n10113 ) | ( n9771 & n10114 ) | ( n10113 & n10114 ) ;
  assign n10116 = ( ~n9771 & n10113 ) | ( ~n9771 & n10114 ) | ( n10113 & n10114 ) ;
  assign n10117 = ( n9771 & ~n10115 ) | ( n9771 & n10116 ) | ( ~n10115 & n10116 ) ;
  assign n10118 = ( x81 & n10112 ) | ( x81 & ~n10117 ) | ( n10112 & ~n10117 ) ;
  assign n10119 = ( x81 & n9772 ) | ( x81 & ~n10017 ) | ( n9772 & ~n10017 ) ;
  assign n10120 = x81 & n9772 ;
  assign n10121 = ( ~n9777 & n10119 ) | ( ~n9777 & n10120 ) | ( n10119 & n10120 ) ;
  assign n10122 = ( n9777 & n10119 ) | ( n9777 & n10120 ) | ( n10119 & n10120 ) ;
  assign n10123 = ( n9777 & n10121 ) | ( n9777 & ~n10122 ) | ( n10121 & ~n10122 ) ;
  assign n10124 = ( x82 & n10118 ) | ( x82 & ~n10123 ) | ( n10118 & ~n10123 ) ;
  assign n10125 = ( x82 & n9778 ) | ( x82 & ~n10017 ) | ( n9778 & ~n10017 ) ;
  assign n10126 = x82 & n9778 ;
  assign n10127 = ( n9783 & n10125 ) | ( n9783 & n10126 ) | ( n10125 & n10126 ) ;
  assign n10128 = ( ~n9783 & n10125 ) | ( ~n9783 & n10126 ) | ( n10125 & n10126 ) ;
  assign n10129 = ( n9783 & ~n10127 ) | ( n9783 & n10128 ) | ( ~n10127 & n10128 ) ;
  assign n10130 = ( x83 & n10124 ) | ( x83 & ~n10129 ) | ( n10124 & ~n10129 ) ;
  assign n10131 = ( x83 & n9784 ) | ( x83 & ~n10017 ) | ( n9784 & ~n10017 ) ;
  assign n10132 = x83 & n9784 ;
  assign n10133 = ( ~n9789 & n10131 ) | ( ~n9789 & n10132 ) | ( n10131 & n10132 ) ;
  assign n10134 = ( n9789 & n10131 ) | ( n9789 & n10132 ) | ( n10131 & n10132 ) ;
  assign n10135 = ( n9789 & n10133 ) | ( n9789 & ~n10134 ) | ( n10133 & ~n10134 ) ;
  assign n10136 = ( x84 & n10130 ) | ( x84 & ~n10135 ) | ( n10130 & ~n10135 ) ;
  assign n10137 = ( x84 & n9790 ) | ( x84 & ~n10017 ) | ( n9790 & ~n10017 ) ;
  assign n10138 = x84 & n9790 ;
  assign n10139 = ( n9795 & n10137 ) | ( n9795 & n10138 ) | ( n10137 & n10138 ) ;
  assign n10140 = ( ~n9795 & n10137 ) | ( ~n9795 & n10138 ) | ( n10137 & n10138 ) ;
  assign n10141 = ( n9795 & ~n10139 ) | ( n9795 & n10140 ) | ( ~n10139 & n10140 ) ;
  assign n10142 = ( x85 & n10136 ) | ( x85 & ~n10141 ) | ( n10136 & ~n10141 ) ;
  assign n10143 = ( x85 & n9796 ) | ( x85 & ~n10017 ) | ( n9796 & ~n10017 ) ;
  assign n10144 = x85 & n9796 ;
  assign n10145 = ( ~n9801 & n10143 ) | ( ~n9801 & n10144 ) | ( n10143 & n10144 ) ;
  assign n10146 = ( n9801 & n10143 ) | ( n9801 & n10144 ) | ( n10143 & n10144 ) ;
  assign n10147 = ( n9801 & n10145 ) | ( n9801 & ~n10146 ) | ( n10145 & ~n10146 ) ;
  assign n10148 = ( x86 & n10142 ) | ( x86 & ~n10147 ) | ( n10142 & ~n10147 ) ;
  assign n10149 = ( x86 & n9802 ) | ( x86 & ~n10017 ) | ( n9802 & ~n10017 ) ;
  assign n10150 = x86 & n9802 ;
  assign n10151 = ( n9807 & n10149 ) | ( n9807 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10152 = ( ~n9807 & n10149 ) | ( ~n9807 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10153 = ( n9807 & ~n10151 ) | ( n9807 & n10152 ) | ( ~n10151 & n10152 ) ;
  assign n10154 = ( x87 & n10148 ) | ( x87 & ~n10153 ) | ( n10148 & ~n10153 ) ;
  assign n10155 = ( x87 & n9808 ) | ( x87 & ~n10017 ) | ( n9808 & ~n10017 ) ;
  assign n10156 = x87 & n9808 ;
  assign n10157 = ( ~n9813 & n10155 ) | ( ~n9813 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10158 = ( n9813 & n10155 ) | ( n9813 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10159 = ( n9813 & n10157 ) | ( n9813 & ~n10158 ) | ( n10157 & ~n10158 ) ;
  assign n10160 = ( x88 & n10154 ) | ( x88 & ~n10159 ) | ( n10154 & ~n10159 ) ;
  assign n10161 = ( x88 & n9814 ) | ( x88 & ~n10017 ) | ( n9814 & ~n10017 ) ;
  assign n10162 = x88 & n9814 ;
  assign n10163 = ( n9819 & n10161 ) | ( n9819 & n10162 ) | ( n10161 & n10162 ) ;
  assign n10164 = ( ~n9819 & n10161 ) | ( ~n9819 & n10162 ) | ( n10161 & n10162 ) ;
  assign n10165 = ( n9819 & ~n10163 ) | ( n9819 & n10164 ) | ( ~n10163 & n10164 ) ;
  assign n10166 = ( x89 & n10160 ) | ( x89 & ~n10165 ) | ( n10160 & ~n10165 ) ;
  assign n10167 = ( x89 & n9820 ) | ( x89 & ~n10017 ) | ( n9820 & ~n10017 ) ;
  assign n10168 = x89 & n9820 ;
  assign n10169 = ( ~n9825 & n10167 ) | ( ~n9825 & n10168 ) | ( n10167 & n10168 ) ;
  assign n10170 = ( n9825 & n10167 ) | ( n9825 & n10168 ) | ( n10167 & n10168 ) ;
  assign n10171 = ( n9825 & n10169 ) | ( n9825 & ~n10170 ) | ( n10169 & ~n10170 ) ;
  assign n10172 = ( x90 & n10166 ) | ( x90 & ~n10171 ) | ( n10166 & ~n10171 ) ;
  assign n10173 = ( x90 & n9826 ) | ( x90 & ~n10017 ) | ( n9826 & ~n10017 ) ;
  assign n10174 = x90 & n9826 ;
  assign n10175 = ( n9831 & n10173 ) | ( n9831 & n10174 ) | ( n10173 & n10174 ) ;
  assign n10176 = ( ~n9831 & n10173 ) | ( ~n9831 & n10174 ) | ( n10173 & n10174 ) ;
  assign n10177 = ( n9831 & ~n10175 ) | ( n9831 & n10176 ) | ( ~n10175 & n10176 ) ;
  assign n10178 = ( x91 & n10172 ) | ( x91 & ~n10177 ) | ( n10172 & ~n10177 ) ;
  assign n10179 = ( x91 & n9832 ) | ( x91 & ~n10017 ) | ( n9832 & ~n10017 ) ;
  assign n10180 = x91 & n9832 ;
  assign n10181 = ( ~n9837 & n10179 ) | ( ~n9837 & n10180 ) | ( n10179 & n10180 ) ;
  assign n10182 = ( n9837 & n10179 ) | ( n9837 & n10180 ) | ( n10179 & n10180 ) ;
  assign n10183 = ( n9837 & n10181 ) | ( n9837 & ~n10182 ) | ( n10181 & ~n10182 ) ;
  assign n10184 = ( x92 & n10178 ) | ( x92 & ~n10183 ) | ( n10178 & ~n10183 ) ;
  assign n10185 = ( x92 & n9838 ) | ( x92 & ~n10017 ) | ( n9838 & ~n10017 ) ;
  assign n10186 = x92 & n9838 ;
  assign n10187 = ( n9843 & n10185 ) | ( n9843 & n10186 ) | ( n10185 & n10186 ) ;
  assign n10188 = ( ~n9843 & n10185 ) | ( ~n9843 & n10186 ) | ( n10185 & n10186 ) ;
  assign n10189 = ( n9843 & ~n10187 ) | ( n9843 & n10188 ) | ( ~n10187 & n10188 ) ;
  assign n10190 = ( x93 & n10184 ) | ( x93 & ~n10189 ) | ( n10184 & ~n10189 ) ;
  assign n10191 = ( x93 & n9844 ) | ( x93 & ~n10017 ) | ( n9844 & ~n10017 ) ;
  assign n10192 = x93 & n9844 ;
  assign n10193 = ( ~n9849 & n10191 ) | ( ~n9849 & n10192 ) | ( n10191 & n10192 ) ;
  assign n10194 = ( n9849 & n10191 ) | ( n9849 & n10192 ) | ( n10191 & n10192 ) ;
  assign n10195 = ( n9849 & n10193 ) | ( n9849 & ~n10194 ) | ( n10193 & ~n10194 ) ;
  assign n10196 = ( x94 & n10190 ) | ( x94 & ~n10195 ) | ( n10190 & ~n10195 ) ;
  assign n10197 = ( x94 & n9850 ) | ( x94 & ~n10017 ) | ( n9850 & ~n10017 ) ;
  assign n10198 = x94 & n9850 ;
  assign n10199 = ( n9855 & n10197 ) | ( n9855 & n10198 ) | ( n10197 & n10198 ) ;
  assign n10200 = ( ~n9855 & n10197 ) | ( ~n9855 & n10198 ) | ( n10197 & n10198 ) ;
  assign n10201 = ( n9855 & ~n10199 ) | ( n9855 & n10200 ) | ( ~n10199 & n10200 ) ;
  assign n10202 = ( x95 & n10196 ) | ( x95 & ~n10201 ) | ( n10196 & ~n10201 ) ;
  assign n10203 = ( x95 & n9856 ) | ( x95 & ~n10017 ) | ( n9856 & ~n10017 ) ;
  assign n10204 = x95 & n9856 ;
  assign n10205 = ( ~n9861 & n10203 ) | ( ~n9861 & n10204 ) | ( n10203 & n10204 ) ;
  assign n10206 = ( n9861 & n10203 ) | ( n9861 & n10204 ) | ( n10203 & n10204 ) ;
  assign n10207 = ( n9861 & n10205 ) | ( n9861 & ~n10206 ) | ( n10205 & ~n10206 ) ;
  assign n10208 = ( x96 & n10202 ) | ( x96 & ~n10207 ) | ( n10202 & ~n10207 ) ;
  assign n10209 = ( x96 & n9862 ) | ( x96 & ~n10017 ) | ( n9862 & ~n10017 ) ;
  assign n10210 = x96 & n9862 ;
  assign n10211 = ( n9867 & n10209 ) | ( n9867 & n10210 ) | ( n10209 & n10210 ) ;
  assign n10212 = ( ~n9867 & n10209 ) | ( ~n9867 & n10210 ) | ( n10209 & n10210 ) ;
  assign n10213 = ( n9867 & ~n10211 ) | ( n9867 & n10212 ) | ( ~n10211 & n10212 ) ;
  assign n10214 = ( x97 & n10208 ) | ( x97 & ~n10213 ) | ( n10208 & ~n10213 ) ;
  assign n10215 = ( x97 & n9868 ) | ( x97 & ~n10017 ) | ( n9868 & ~n10017 ) ;
  assign n10216 = x97 & n9868 ;
  assign n10217 = ( ~n9873 & n10215 ) | ( ~n9873 & n10216 ) | ( n10215 & n10216 ) ;
  assign n10218 = ( n9873 & n10215 ) | ( n9873 & n10216 ) | ( n10215 & n10216 ) ;
  assign n10219 = ( n9873 & n10217 ) | ( n9873 & ~n10218 ) | ( n10217 & ~n10218 ) ;
  assign n10220 = ( x98 & n10214 ) | ( x98 & ~n10219 ) | ( n10214 & ~n10219 ) ;
  assign n10221 = ( x98 & n9874 ) | ( x98 & ~n10017 ) | ( n9874 & ~n10017 ) ;
  assign n10222 = x98 & n9874 ;
  assign n10223 = ( n9879 & n10221 ) | ( n9879 & n10222 ) | ( n10221 & n10222 ) ;
  assign n10224 = ( ~n9879 & n10221 ) | ( ~n9879 & n10222 ) | ( n10221 & n10222 ) ;
  assign n10225 = ( n9879 & ~n10223 ) | ( n9879 & n10224 ) | ( ~n10223 & n10224 ) ;
  assign n10226 = ( x99 & n10220 ) | ( x99 & ~n10225 ) | ( n10220 & ~n10225 ) ;
  assign n10227 = ( x99 & n9880 ) | ( x99 & ~n10017 ) | ( n9880 & ~n10017 ) ;
  assign n10228 = x99 & n9880 ;
  assign n10229 = ( ~n9885 & n10227 ) | ( ~n9885 & n10228 ) | ( n10227 & n10228 ) ;
  assign n10230 = ( n9885 & n10227 ) | ( n9885 & n10228 ) | ( n10227 & n10228 ) ;
  assign n10231 = ( n9885 & n10229 ) | ( n9885 & ~n10230 ) | ( n10229 & ~n10230 ) ;
  assign n10232 = ( x100 & n10226 ) | ( x100 & ~n10231 ) | ( n10226 & ~n10231 ) ;
  assign n10233 = ( x100 & n9886 ) | ( x100 & ~n10017 ) | ( n9886 & ~n10017 ) ;
  assign n10234 = x100 & n9886 ;
  assign n10235 = ( n9891 & n10233 ) | ( n9891 & n10234 ) | ( n10233 & n10234 ) ;
  assign n10236 = ( ~n9891 & n10233 ) | ( ~n9891 & n10234 ) | ( n10233 & n10234 ) ;
  assign n10237 = ( n9891 & ~n10235 ) | ( n9891 & n10236 ) | ( ~n10235 & n10236 ) ;
  assign n10238 = ( x101 & n10232 ) | ( x101 & ~n10237 ) | ( n10232 & ~n10237 ) ;
  assign n10239 = ( x101 & n9892 ) | ( x101 & ~n10017 ) | ( n9892 & ~n10017 ) ;
  assign n10240 = x101 & n9892 ;
  assign n10241 = ( ~n9897 & n10239 ) | ( ~n9897 & n10240 ) | ( n10239 & n10240 ) ;
  assign n10242 = ( n9897 & n10239 ) | ( n9897 & n10240 ) | ( n10239 & n10240 ) ;
  assign n10243 = ( n9897 & n10241 ) | ( n9897 & ~n10242 ) | ( n10241 & ~n10242 ) ;
  assign n10244 = ( x102 & n10238 ) | ( x102 & ~n10243 ) | ( n10238 & ~n10243 ) ;
  assign n10245 = ( x102 & n9898 ) | ( x102 & ~n10017 ) | ( n9898 & ~n10017 ) ;
  assign n10246 = x102 & n9898 ;
  assign n10247 = ( n9903 & n10245 ) | ( n9903 & n10246 ) | ( n10245 & n10246 ) ;
  assign n10248 = ( ~n9903 & n10245 ) | ( ~n9903 & n10246 ) | ( n10245 & n10246 ) ;
  assign n10249 = ( n9903 & ~n10247 ) | ( n9903 & n10248 ) | ( ~n10247 & n10248 ) ;
  assign n10250 = ( x103 & n10244 ) | ( x103 & ~n10249 ) | ( n10244 & ~n10249 ) ;
  assign n10251 = ( x103 & n9904 ) | ( x103 & ~n10017 ) | ( n9904 & ~n10017 ) ;
  assign n10252 = x103 & n9904 ;
  assign n10253 = ( ~n9909 & n10251 ) | ( ~n9909 & n10252 ) | ( n10251 & n10252 ) ;
  assign n10254 = ( n9909 & n10251 ) | ( n9909 & n10252 ) | ( n10251 & n10252 ) ;
  assign n10255 = ( n9909 & n10253 ) | ( n9909 & ~n10254 ) | ( n10253 & ~n10254 ) ;
  assign n10256 = ( x104 & n10250 ) | ( x104 & ~n10255 ) | ( n10250 & ~n10255 ) ;
  assign n10257 = ( x104 & n9910 ) | ( x104 & ~n10017 ) | ( n9910 & ~n10017 ) ;
  assign n10258 = x104 & n9910 ;
  assign n10259 = ( n9915 & n10257 ) | ( n9915 & n10258 ) | ( n10257 & n10258 ) ;
  assign n10260 = ( ~n9915 & n10257 ) | ( ~n9915 & n10258 ) | ( n10257 & n10258 ) ;
  assign n10261 = ( n9915 & ~n10259 ) | ( n9915 & n10260 ) | ( ~n10259 & n10260 ) ;
  assign n10262 = ( x105 & n10256 ) | ( x105 & ~n10261 ) | ( n10256 & ~n10261 ) ;
  assign n10263 = ( x105 & n9916 ) | ( x105 & ~n10017 ) | ( n9916 & ~n10017 ) ;
  assign n10264 = x105 & n9916 ;
  assign n10265 = ( ~n9921 & n10263 ) | ( ~n9921 & n10264 ) | ( n10263 & n10264 ) ;
  assign n10266 = ( n9921 & n10263 ) | ( n9921 & n10264 ) | ( n10263 & n10264 ) ;
  assign n10267 = ( n9921 & n10265 ) | ( n9921 & ~n10266 ) | ( n10265 & ~n10266 ) ;
  assign n10268 = ( x106 & n10262 ) | ( x106 & ~n10267 ) | ( n10262 & ~n10267 ) ;
  assign n10269 = ( x106 & n9922 ) | ( x106 & ~n10017 ) | ( n9922 & ~n10017 ) ;
  assign n10270 = x106 & n9922 ;
  assign n10271 = ( n9927 & n10269 ) | ( n9927 & n10270 ) | ( n10269 & n10270 ) ;
  assign n10272 = ( ~n9927 & n10269 ) | ( ~n9927 & n10270 ) | ( n10269 & n10270 ) ;
  assign n10273 = ( n9927 & ~n10271 ) | ( n9927 & n10272 ) | ( ~n10271 & n10272 ) ;
  assign n10274 = ( x107 & n10268 ) | ( x107 & ~n10273 ) | ( n10268 & ~n10273 ) ;
  assign n10275 = ( x107 & n9928 ) | ( x107 & ~n10017 ) | ( n9928 & ~n10017 ) ;
  assign n10276 = x107 & n9928 ;
  assign n10277 = ( ~n9933 & n10275 ) | ( ~n9933 & n10276 ) | ( n10275 & n10276 ) ;
  assign n10278 = ( n9933 & n10275 ) | ( n9933 & n10276 ) | ( n10275 & n10276 ) ;
  assign n10279 = ( n9933 & n10277 ) | ( n9933 & ~n10278 ) | ( n10277 & ~n10278 ) ;
  assign n10280 = ( x108 & n10274 ) | ( x108 & ~n10279 ) | ( n10274 & ~n10279 ) ;
  assign n10281 = ( x108 & n9934 ) | ( x108 & ~n10017 ) | ( n9934 & ~n10017 ) ;
  assign n10282 = x108 & n9934 ;
  assign n10283 = ( n9939 & n10281 ) | ( n9939 & n10282 ) | ( n10281 & n10282 ) ;
  assign n10284 = ( ~n9939 & n10281 ) | ( ~n9939 & n10282 ) | ( n10281 & n10282 ) ;
  assign n10285 = ( n9939 & ~n10283 ) | ( n9939 & n10284 ) | ( ~n10283 & n10284 ) ;
  assign n10286 = ( x109 & n10280 ) | ( x109 & ~n10285 ) | ( n10280 & ~n10285 ) ;
  assign n10287 = ( x109 & n9940 ) | ( x109 & ~n10017 ) | ( n9940 & ~n10017 ) ;
  assign n10288 = x109 & n9940 ;
  assign n10289 = ( ~n9945 & n10287 ) | ( ~n9945 & n10288 ) | ( n10287 & n10288 ) ;
  assign n10290 = ( n9945 & n10287 ) | ( n9945 & n10288 ) | ( n10287 & n10288 ) ;
  assign n10291 = ( n9945 & n10289 ) | ( n9945 & ~n10290 ) | ( n10289 & ~n10290 ) ;
  assign n10292 = ( x110 & n10286 ) | ( x110 & ~n10291 ) | ( n10286 & ~n10291 ) ;
  assign n10293 = ( x110 & n9946 ) | ( x110 & ~n10017 ) | ( n9946 & ~n10017 ) ;
  assign n10294 = x110 & n9946 ;
  assign n10295 = ( n9951 & n10293 ) | ( n9951 & n10294 ) | ( n10293 & n10294 ) ;
  assign n10296 = ( ~n9951 & n10293 ) | ( ~n9951 & n10294 ) | ( n10293 & n10294 ) ;
  assign n10297 = ( n9951 & ~n10295 ) | ( n9951 & n10296 ) | ( ~n10295 & n10296 ) ;
  assign n10298 = ( x111 & n10292 ) | ( x111 & ~n10297 ) | ( n10292 & ~n10297 ) ;
  assign n10299 = ( x111 & n9952 ) | ( x111 & ~n10017 ) | ( n9952 & ~n10017 ) ;
  assign n10300 = x111 & n9952 ;
  assign n10301 = ( ~n9957 & n10299 ) | ( ~n9957 & n10300 ) | ( n10299 & n10300 ) ;
  assign n10302 = ( n9957 & n10299 ) | ( n9957 & n10300 ) | ( n10299 & n10300 ) ;
  assign n10303 = ( n9957 & n10301 ) | ( n9957 & ~n10302 ) | ( n10301 & ~n10302 ) ;
  assign n10304 = ( x112 & n10298 ) | ( x112 & ~n10303 ) | ( n10298 & ~n10303 ) ;
  assign n10305 = ( x112 & n9958 ) | ( x112 & ~n10017 ) | ( n9958 & ~n10017 ) ;
  assign n10306 = x112 & n9958 ;
  assign n10307 = ( n9963 & n10305 ) | ( n9963 & n10306 ) | ( n10305 & n10306 ) ;
  assign n10308 = ( ~n9963 & n10305 ) | ( ~n9963 & n10306 ) | ( n10305 & n10306 ) ;
  assign n10309 = ( n9963 & ~n10307 ) | ( n9963 & n10308 ) | ( ~n10307 & n10308 ) ;
  assign n10310 = ( x113 & n10304 ) | ( x113 & ~n10309 ) | ( n10304 & ~n10309 ) ;
  assign n10311 = ( x113 & n9964 ) | ( x113 & ~n10017 ) | ( n9964 & ~n10017 ) ;
  assign n10312 = x113 & n9964 ;
  assign n10313 = ( ~n9969 & n10311 ) | ( ~n9969 & n10312 ) | ( n10311 & n10312 ) ;
  assign n10314 = ( n9969 & n10311 ) | ( n9969 & n10312 ) | ( n10311 & n10312 ) ;
  assign n10315 = ( n9969 & n10313 ) | ( n9969 & ~n10314 ) | ( n10313 & ~n10314 ) ;
  assign n10316 = ( x114 & n10310 ) | ( x114 & ~n10315 ) | ( n10310 & ~n10315 ) ;
  assign n10317 = ( x114 & n9970 ) | ( x114 & ~n10017 ) | ( n9970 & ~n10017 ) ;
  assign n10318 = x114 & n9970 ;
  assign n10319 = ( n9975 & n10317 ) | ( n9975 & n10318 ) | ( n10317 & n10318 ) ;
  assign n10320 = ( ~n9975 & n10317 ) | ( ~n9975 & n10318 ) | ( n10317 & n10318 ) ;
  assign n10321 = ( n9975 & ~n10319 ) | ( n9975 & n10320 ) | ( ~n10319 & n10320 ) ;
  assign n10322 = ( x115 & n10316 ) | ( x115 & ~n10321 ) | ( n10316 & ~n10321 ) ;
  assign n10323 = ( x115 & n9976 ) | ( x115 & ~n10017 ) | ( n9976 & ~n10017 ) ;
  assign n10324 = x115 & n9976 ;
  assign n10325 = ( ~n9981 & n10323 ) | ( ~n9981 & n10324 ) | ( n10323 & n10324 ) ;
  assign n10326 = ( n9981 & n10323 ) | ( n9981 & n10324 ) | ( n10323 & n10324 ) ;
  assign n10327 = ( n9981 & n10325 ) | ( n9981 & ~n10326 ) | ( n10325 & ~n10326 ) ;
  assign n10328 = ( x116 & n10322 ) | ( x116 & ~n10327 ) | ( n10322 & ~n10327 ) ;
  assign n10329 = ( x116 & n9982 ) | ( x116 & ~n10017 ) | ( n9982 & ~n10017 ) ;
  assign n10330 = x116 & n9982 ;
  assign n10331 = ( n9987 & n10329 ) | ( n9987 & n10330 ) | ( n10329 & n10330 ) ;
  assign n10332 = ( ~n9987 & n10329 ) | ( ~n9987 & n10330 ) | ( n10329 & n10330 ) ;
  assign n10333 = ( n9987 & ~n10331 ) | ( n9987 & n10332 ) | ( ~n10331 & n10332 ) ;
  assign n10334 = ( x117 & n10328 ) | ( x117 & ~n10333 ) | ( n10328 & ~n10333 ) ;
  assign n10335 = ( x117 & n9988 ) | ( x117 & ~n10017 ) | ( n9988 & ~n10017 ) ;
  assign n10336 = x117 & n9988 ;
  assign n10337 = ( ~n9993 & n10335 ) | ( ~n9993 & n10336 ) | ( n10335 & n10336 ) ;
  assign n10338 = ( n9993 & n10335 ) | ( n9993 & n10336 ) | ( n10335 & n10336 ) ;
  assign n10339 = ( n9993 & n10337 ) | ( n9993 & ~n10338 ) | ( n10337 & ~n10338 ) ;
  assign n10340 = ( x118 & n10334 ) | ( x118 & ~n10339 ) | ( n10334 & ~n10339 ) ;
  assign n10341 = ( x118 & n9994 ) | ( x118 & ~n10017 ) | ( n9994 & ~n10017 ) ;
  assign n10342 = x118 & n9994 ;
  assign n10343 = ( n9999 & n10341 ) | ( n9999 & n10342 ) | ( n10341 & n10342 ) ;
  assign n10344 = ( ~n9999 & n10341 ) | ( ~n9999 & n10342 ) | ( n10341 & n10342 ) ;
  assign n10345 = ( n9999 & ~n10343 ) | ( n9999 & n10344 ) | ( ~n10343 & n10344 ) ;
  assign n10346 = ( x119 & n10340 ) | ( x119 & ~n10345 ) | ( n10340 & ~n10345 ) ;
  assign n10347 = ( x119 & n10000 ) | ( x119 & ~n10017 ) | ( n10000 & ~n10017 ) ;
  assign n10348 = x119 & n10000 ;
  assign n10349 = ( ~n10005 & n10347 ) | ( ~n10005 & n10348 ) | ( n10347 & n10348 ) ;
  assign n10350 = ( n10005 & n10347 ) | ( n10005 & n10348 ) | ( n10347 & n10348 ) ;
  assign n10351 = ( n10005 & n10349 ) | ( n10005 & ~n10350 ) | ( n10349 & ~n10350 ) ;
  assign n10352 = ( x120 & n10346 ) | ( x120 & ~n10351 ) | ( n10346 & ~n10351 ) ;
  assign n10353 = ( x120 & n10006 ) | ( x120 & ~n10017 ) | ( n10006 & ~n10017 ) ;
  assign n10354 = x120 & n10006 ;
  assign n10355 = ( ~n10011 & n10353 ) | ( ~n10011 & n10354 ) | ( n10353 & n10354 ) ;
  assign n10356 = ( n10011 & n10353 ) | ( n10011 & n10354 ) | ( n10353 & n10354 ) ;
  assign n10357 = ( n10011 & n10355 ) | ( n10011 & ~n10356 ) | ( n10355 & ~n10356 ) ;
  assign n10358 = ( x121 & n10352 ) | ( x121 & ~n10357 ) | ( n10352 & ~n10357 ) ;
  assign n10359 = x122 | n10358 ;
  assign n10360 = ( x122 & n135 ) | ( x122 & n10358 ) | ( n135 & n10358 ) ;
  assign n10361 = ( n10015 & ~n10359 ) | ( n10015 & n10360 ) | ( ~n10359 & n10360 ) ;
  assign n10362 = ( x122 & ~n10015 ) | ( x122 & n10358 ) | ( ~n10015 & n10358 ) ;
  assign n10363 = n135 | n10362 ;
  assign n10364 = ( x5 & ~x64 ) | ( x5 & n10363 ) | ( ~x64 & n10363 ) ;
  assign n10365 = ~x5 & n10363 ;
  assign n10366 = ( n10021 & n10364 ) | ( n10021 & ~n10365 ) | ( n10364 & ~n10365 ) ;
  assign n10367 = ~x4 & x64 ;
  assign n10368 = ( x65 & ~n10366 ) | ( x65 & n10367 ) | ( ~n10366 & n10367 ) ;
  assign n10369 = ( x65 & n10021 ) | ( x65 & ~n10363 ) | ( n10021 & ~n10363 ) ;
  assign n10370 = x65 & n10021 ;
  assign n10371 = ( n10020 & n10369 ) | ( n10020 & n10370 ) | ( n10369 & n10370 ) ;
  assign n10372 = ( ~n10020 & n10369 ) | ( ~n10020 & n10370 ) | ( n10369 & n10370 ) ;
  assign n10373 = ( n10020 & ~n10371 ) | ( n10020 & n10372 ) | ( ~n10371 & n10372 ) ;
  assign n10374 = ( x66 & n10368 ) | ( x66 & ~n10373 ) | ( n10368 & ~n10373 ) ;
  assign n10375 = ( x66 & n10022 ) | ( x66 & ~n10363 ) | ( n10022 & ~n10363 ) ;
  assign n10376 = x66 & n10022 ;
  assign n10377 = ( n10027 & n10375 ) | ( n10027 & n10376 ) | ( n10375 & n10376 ) ;
  assign n10378 = ( ~n10027 & n10375 ) | ( ~n10027 & n10376 ) | ( n10375 & n10376 ) ;
  assign n10379 = ( n10027 & ~n10377 ) | ( n10027 & n10378 ) | ( ~n10377 & n10378 ) ;
  assign n10380 = ( x67 & n10374 ) | ( x67 & ~n10379 ) | ( n10374 & ~n10379 ) ;
  assign n10381 = ( x67 & n10028 ) | ( x67 & ~n10363 ) | ( n10028 & ~n10363 ) ;
  assign n10382 = x67 & n10028 ;
  assign n10383 = ( ~n10033 & n10381 ) | ( ~n10033 & n10382 ) | ( n10381 & n10382 ) ;
  assign n10384 = ( n10033 & n10381 ) | ( n10033 & n10382 ) | ( n10381 & n10382 ) ;
  assign n10385 = ( n10033 & n10383 ) | ( n10033 & ~n10384 ) | ( n10383 & ~n10384 ) ;
  assign n10386 = ( x68 & n10380 ) | ( x68 & ~n10385 ) | ( n10380 & ~n10385 ) ;
  assign n10387 = ( x68 & n10034 ) | ( x68 & ~n10363 ) | ( n10034 & ~n10363 ) ;
  assign n10388 = x68 & n10034 ;
  assign n10389 = ( n10039 & n10387 ) | ( n10039 & n10388 ) | ( n10387 & n10388 ) ;
  assign n10390 = ( ~n10039 & n10387 ) | ( ~n10039 & n10388 ) | ( n10387 & n10388 ) ;
  assign n10391 = ( n10039 & ~n10389 ) | ( n10039 & n10390 ) | ( ~n10389 & n10390 ) ;
  assign n10392 = ( x69 & n10386 ) | ( x69 & ~n10391 ) | ( n10386 & ~n10391 ) ;
  assign n10393 = ( x69 & n10040 ) | ( x69 & ~n10363 ) | ( n10040 & ~n10363 ) ;
  assign n10394 = x69 & n10040 ;
  assign n10395 = ( ~n10045 & n10393 ) | ( ~n10045 & n10394 ) | ( n10393 & n10394 ) ;
  assign n10396 = ( n10045 & n10393 ) | ( n10045 & n10394 ) | ( n10393 & n10394 ) ;
  assign n10397 = ( n10045 & n10395 ) | ( n10045 & ~n10396 ) | ( n10395 & ~n10396 ) ;
  assign n10398 = ( x70 & n10392 ) | ( x70 & ~n10397 ) | ( n10392 & ~n10397 ) ;
  assign n10399 = ( x70 & n10046 ) | ( x70 & ~n10363 ) | ( n10046 & ~n10363 ) ;
  assign n10400 = x70 & n10046 ;
  assign n10401 = ( n10051 & n10399 ) | ( n10051 & n10400 ) | ( n10399 & n10400 ) ;
  assign n10402 = ( ~n10051 & n10399 ) | ( ~n10051 & n10400 ) | ( n10399 & n10400 ) ;
  assign n10403 = ( n10051 & ~n10401 ) | ( n10051 & n10402 ) | ( ~n10401 & n10402 ) ;
  assign n10404 = ( x71 & n10398 ) | ( x71 & ~n10403 ) | ( n10398 & ~n10403 ) ;
  assign n10405 = ( x71 & n10052 ) | ( x71 & ~n10363 ) | ( n10052 & ~n10363 ) ;
  assign n10406 = x71 & n10052 ;
  assign n10407 = ( ~n10057 & n10405 ) | ( ~n10057 & n10406 ) | ( n10405 & n10406 ) ;
  assign n10408 = ( n10057 & n10405 ) | ( n10057 & n10406 ) | ( n10405 & n10406 ) ;
  assign n10409 = ( n10057 & n10407 ) | ( n10057 & ~n10408 ) | ( n10407 & ~n10408 ) ;
  assign n10410 = ( x72 & n10404 ) | ( x72 & ~n10409 ) | ( n10404 & ~n10409 ) ;
  assign n10411 = ( x72 & n10058 ) | ( x72 & ~n10363 ) | ( n10058 & ~n10363 ) ;
  assign n10412 = x72 & n10058 ;
  assign n10413 = ( n10063 & n10411 ) | ( n10063 & n10412 ) | ( n10411 & n10412 ) ;
  assign n10414 = ( ~n10063 & n10411 ) | ( ~n10063 & n10412 ) | ( n10411 & n10412 ) ;
  assign n10415 = ( n10063 & ~n10413 ) | ( n10063 & n10414 ) | ( ~n10413 & n10414 ) ;
  assign n10416 = ( x73 & n10410 ) | ( x73 & ~n10415 ) | ( n10410 & ~n10415 ) ;
  assign n10417 = ( x73 & n10064 ) | ( x73 & ~n10363 ) | ( n10064 & ~n10363 ) ;
  assign n10418 = x73 & n10064 ;
  assign n10419 = ( ~n10069 & n10417 ) | ( ~n10069 & n10418 ) | ( n10417 & n10418 ) ;
  assign n10420 = ( n10069 & n10417 ) | ( n10069 & n10418 ) | ( n10417 & n10418 ) ;
  assign n10421 = ( n10069 & n10419 ) | ( n10069 & ~n10420 ) | ( n10419 & ~n10420 ) ;
  assign n10422 = ( x74 & n10416 ) | ( x74 & ~n10421 ) | ( n10416 & ~n10421 ) ;
  assign n10423 = ( x74 & n10070 ) | ( x74 & ~n10363 ) | ( n10070 & ~n10363 ) ;
  assign n10424 = x74 & n10070 ;
  assign n10425 = ( n10075 & n10423 ) | ( n10075 & n10424 ) | ( n10423 & n10424 ) ;
  assign n10426 = ( ~n10075 & n10423 ) | ( ~n10075 & n10424 ) | ( n10423 & n10424 ) ;
  assign n10427 = ( n10075 & ~n10425 ) | ( n10075 & n10426 ) | ( ~n10425 & n10426 ) ;
  assign n10428 = ( x75 & n10422 ) | ( x75 & ~n10427 ) | ( n10422 & ~n10427 ) ;
  assign n10429 = ( x75 & n10076 ) | ( x75 & ~n10363 ) | ( n10076 & ~n10363 ) ;
  assign n10430 = x75 & n10076 ;
  assign n10431 = ( ~n10081 & n10429 ) | ( ~n10081 & n10430 ) | ( n10429 & n10430 ) ;
  assign n10432 = ( n10081 & n10429 ) | ( n10081 & n10430 ) | ( n10429 & n10430 ) ;
  assign n10433 = ( n10081 & n10431 ) | ( n10081 & ~n10432 ) | ( n10431 & ~n10432 ) ;
  assign n10434 = ( x76 & n10428 ) | ( x76 & ~n10433 ) | ( n10428 & ~n10433 ) ;
  assign n10435 = ( x76 & n10082 ) | ( x76 & ~n10363 ) | ( n10082 & ~n10363 ) ;
  assign n10436 = x76 & n10082 ;
  assign n10437 = ( n10087 & n10435 ) | ( n10087 & n10436 ) | ( n10435 & n10436 ) ;
  assign n10438 = ( ~n10087 & n10435 ) | ( ~n10087 & n10436 ) | ( n10435 & n10436 ) ;
  assign n10439 = ( n10087 & ~n10437 ) | ( n10087 & n10438 ) | ( ~n10437 & n10438 ) ;
  assign n10440 = ( x77 & n10434 ) | ( x77 & ~n10439 ) | ( n10434 & ~n10439 ) ;
  assign n10441 = ( x77 & n10088 ) | ( x77 & ~n10363 ) | ( n10088 & ~n10363 ) ;
  assign n10442 = x77 & n10088 ;
  assign n10443 = ( ~n10093 & n10441 ) | ( ~n10093 & n10442 ) | ( n10441 & n10442 ) ;
  assign n10444 = ( n10093 & n10441 ) | ( n10093 & n10442 ) | ( n10441 & n10442 ) ;
  assign n10445 = ( n10093 & n10443 ) | ( n10093 & ~n10444 ) | ( n10443 & ~n10444 ) ;
  assign n10446 = ( x78 & n10440 ) | ( x78 & ~n10445 ) | ( n10440 & ~n10445 ) ;
  assign n10447 = ( x78 & n10094 ) | ( x78 & ~n10363 ) | ( n10094 & ~n10363 ) ;
  assign n10448 = x78 & n10094 ;
  assign n10449 = ( n10099 & n10447 ) | ( n10099 & n10448 ) | ( n10447 & n10448 ) ;
  assign n10450 = ( ~n10099 & n10447 ) | ( ~n10099 & n10448 ) | ( n10447 & n10448 ) ;
  assign n10451 = ( n10099 & ~n10449 ) | ( n10099 & n10450 ) | ( ~n10449 & n10450 ) ;
  assign n10452 = ( x79 & n10446 ) | ( x79 & ~n10451 ) | ( n10446 & ~n10451 ) ;
  assign n10453 = ( x79 & n10100 ) | ( x79 & ~n10363 ) | ( n10100 & ~n10363 ) ;
  assign n10454 = x79 & n10100 ;
  assign n10455 = ( ~n10105 & n10453 ) | ( ~n10105 & n10454 ) | ( n10453 & n10454 ) ;
  assign n10456 = ( n10105 & n10453 ) | ( n10105 & n10454 ) | ( n10453 & n10454 ) ;
  assign n10457 = ( n10105 & n10455 ) | ( n10105 & ~n10456 ) | ( n10455 & ~n10456 ) ;
  assign n10458 = ( x80 & n10452 ) | ( x80 & ~n10457 ) | ( n10452 & ~n10457 ) ;
  assign n10459 = ( x80 & n10106 ) | ( x80 & ~n10363 ) | ( n10106 & ~n10363 ) ;
  assign n10460 = x80 & n10106 ;
  assign n10461 = ( n10111 & n10459 ) | ( n10111 & n10460 ) | ( n10459 & n10460 ) ;
  assign n10462 = ( ~n10111 & n10459 ) | ( ~n10111 & n10460 ) | ( n10459 & n10460 ) ;
  assign n10463 = ( n10111 & ~n10461 ) | ( n10111 & n10462 ) | ( ~n10461 & n10462 ) ;
  assign n10464 = ( x81 & n10458 ) | ( x81 & ~n10463 ) | ( n10458 & ~n10463 ) ;
  assign n10465 = ( x81 & n10112 ) | ( x81 & ~n10363 ) | ( n10112 & ~n10363 ) ;
  assign n10466 = x81 & n10112 ;
  assign n10467 = ( ~n10117 & n10465 ) | ( ~n10117 & n10466 ) | ( n10465 & n10466 ) ;
  assign n10468 = ( n10117 & n10465 ) | ( n10117 & n10466 ) | ( n10465 & n10466 ) ;
  assign n10469 = ( n10117 & n10467 ) | ( n10117 & ~n10468 ) | ( n10467 & ~n10468 ) ;
  assign n10470 = ( x82 & n10464 ) | ( x82 & ~n10469 ) | ( n10464 & ~n10469 ) ;
  assign n10471 = ( x82 & n10118 ) | ( x82 & ~n10363 ) | ( n10118 & ~n10363 ) ;
  assign n10472 = x82 & n10118 ;
  assign n10473 = ( n10123 & n10471 ) | ( n10123 & n10472 ) | ( n10471 & n10472 ) ;
  assign n10474 = ( ~n10123 & n10471 ) | ( ~n10123 & n10472 ) | ( n10471 & n10472 ) ;
  assign n10475 = ( n10123 & ~n10473 ) | ( n10123 & n10474 ) | ( ~n10473 & n10474 ) ;
  assign n10476 = ( x83 & n10470 ) | ( x83 & ~n10475 ) | ( n10470 & ~n10475 ) ;
  assign n10477 = ( x83 & n10124 ) | ( x83 & ~n10363 ) | ( n10124 & ~n10363 ) ;
  assign n10478 = x83 & n10124 ;
  assign n10479 = ( ~n10129 & n10477 ) | ( ~n10129 & n10478 ) | ( n10477 & n10478 ) ;
  assign n10480 = ( n10129 & n10477 ) | ( n10129 & n10478 ) | ( n10477 & n10478 ) ;
  assign n10481 = ( n10129 & n10479 ) | ( n10129 & ~n10480 ) | ( n10479 & ~n10480 ) ;
  assign n10482 = ( x84 & n10476 ) | ( x84 & ~n10481 ) | ( n10476 & ~n10481 ) ;
  assign n10483 = ( x84 & n10130 ) | ( x84 & ~n10363 ) | ( n10130 & ~n10363 ) ;
  assign n10484 = x84 & n10130 ;
  assign n10485 = ( n10135 & n10483 ) | ( n10135 & n10484 ) | ( n10483 & n10484 ) ;
  assign n10486 = ( ~n10135 & n10483 ) | ( ~n10135 & n10484 ) | ( n10483 & n10484 ) ;
  assign n10487 = ( n10135 & ~n10485 ) | ( n10135 & n10486 ) | ( ~n10485 & n10486 ) ;
  assign n10488 = ( x85 & n10482 ) | ( x85 & ~n10487 ) | ( n10482 & ~n10487 ) ;
  assign n10489 = ( x85 & n10136 ) | ( x85 & ~n10363 ) | ( n10136 & ~n10363 ) ;
  assign n10490 = x85 & n10136 ;
  assign n10491 = ( ~n10141 & n10489 ) | ( ~n10141 & n10490 ) | ( n10489 & n10490 ) ;
  assign n10492 = ( n10141 & n10489 ) | ( n10141 & n10490 ) | ( n10489 & n10490 ) ;
  assign n10493 = ( n10141 & n10491 ) | ( n10141 & ~n10492 ) | ( n10491 & ~n10492 ) ;
  assign n10494 = ( x86 & n10488 ) | ( x86 & ~n10493 ) | ( n10488 & ~n10493 ) ;
  assign n10495 = ( x86 & n10142 ) | ( x86 & ~n10363 ) | ( n10142 & ~n10363 ) ;
  assign n10496 = x86 & n10142 ;
  assign n10497 = ( n10147 & n10495 ) | ( n10147 & n10496 ) | ( n10495 & n10496 ) ;
  assign n10498 = ( ~n10147 & n10495 ) | ( ~n10147 & n10496 ) | ( n10495 & n10496 ) ;
  assign n10499 = ( n10147 & ~n10497 ) | ( n10147 & n10498 ) | ( ~n10497 & n10498 ) ;
  assign n10500 = ( x87 & n10494 ) | ( x87 & ~n10499 ) | ( n10494 & ~n10499 ) ;
  assign n10501 = ( x87 & n10148 ) | ( x87 & ~n10363 ) | ( n10148 & ~n10363 ) ;
  assign n10502 = x87 & n10148 ;
  assign n10503 = ( ~n10153 & n10501 ) | ( ~n10153 & n10502 ) | ( n10501 & n10502 ) ;
  assign n10504 = ( n10153 & n10501 ) | ( n10153 & n10502 ) | ( n10501 & n10502 ) ;
  assign n10505 = ( n10153 & n10503 ) | ( n10153 & ~n10504 ) | ( n10503 & ~n10504 ) ;
  assign n10506 = ( x88 & n10500 ) | ( x88 & ~n10505 ) | ( n10500 & ~n10505 ) ;
  assign n10507 = ( x88 & n10154 ) | ( x88 & ~n10363 ) | ( n10154 & ~n10363 ) ;
  assign n10508 = x88 & n10154 ;
  assign n10509 = ( n10159 & n10507 ) | ( n10159 & n10508 ) | ( n10507 & n10508 ) ;
  assign n10510 = ( ~n10159 & n10507 ) | ( ~n10159 & n10508 ) | ( n10507 & n10508 ) ;
  assign n10511 = ( n10159 & ~n10509 ) | ( n10159 & n10510 ) | ( ~n10509 & n10510 ) ;
  assign n10512 = ( x89 & n10506 ) | ( x89 & ~n10511 ) | ( n10506 & ~n10511 ) ;
  assign n10513 = ( x89 & n10160 ) | ( x89 & ~n10363 ) | ( n10160 & ~n10363 ) ;
  assign n10514 = x89 & n10160 ;
  assign n10515 = ( ~n10165 & n10513 ) | ( ~n10165 & n10514 ) | ( n10513 & n10514 ) ;
  assign n10516 = ( n10165 & n10513 ) | ( n10165 & n10514 ) | ( n10513 & n10514 ) ;
  assign n10517 = ( n10165 & n10515 ) | ( n10165 & ~n10516 ) | ( n10515 & ~n10516 ) ;
  assign n10518 = ( x90 & n10512 ) | ( x90 & ~n10517 ) | ( n10512 & ~n10517 ) ;
  assign n10519 = ( x90 & n10166 ) | ( x90 & ~n10363 ) | ( n10166 & ~n10363 ) ;
  assign n10520 = x90 & n10166 ;
  assign n10521 = ( n10171 & n10519 ) | ( n10171 & n10520 ) | ( n10519 & n10520 ) ;
  assign n10522 = ( ~n10171 & n10519 ) | ( ~n10171 & n10520 ) | ( n10519 & n10520 ) ;
  assign n10523 = ( n10171 & ~n10521 ) | ( n10171 & n10522 ) | ( ~n10521 & n10522 ) ;
  assign n10524 = ( x91 & n10518 ) | ( x91 & ~n10523 ) | ( n10518 & ~n10523 ) ;
  assign n10525 = ( x91 & n10172 ) | ( x91 & ~n10363 ) | ( n10172 & ~n10363 ) ;
  assign n10526 = x91 & n10172 ;
  assign n10527 = ( ~n10177 & n10525 ) | ( ~n10177 & n10526 ) | ( n10525 & n10526 ) ;
  assign n10528 = ( n10177 & n10525 ) | ( n10177 & n10526 ) | ( n10525 & n10526 ) ;
  assign n10529 = ( n10177 & n10527 ) | ( n10177 & ~n10528 ) | ( n10527 & ~n10528 ) ;
  assign n10530 = ( x92 & n10524 ) | ( x92 & ~n10529 ) | ( n10524 & ~n10529 ) ;
  assign n10531 = ( x92 & n10178 ) | ( x92 & ~n10363 ) | ( n10178 & ~n10363 ) ;
  assign n10532 = x92 & n10178 ;
  assign n10533 = ( n10183 & n10531 ) | ( n10183 & n10532 ) | ( n10531 & n10532 ) ;
  assign n10534 = ( ~n10183 & n10531 ) | ( ~n10183 & n10532 ) | ( n10531 & n10532 ) ;
  assign n10535 = ( n10183 & ~n10533 ) | ( n10183 & n10534 ) | ( ~n10533 & n10534 ) ;
  assign n10536 = ( x93 & n10530 ) | ( x93 & ~n10535 ) | ( n10530 & ~n10535 ) ;
  assign n10537 = ( x93 & n10184 ) | ( x93 & ~n10363 ) | ( n10184 & ~n10363 ) ;
  assign n10538 = x93 & n10184 ;
  assign n10539 = ( ~n10189 & n10537 ) | ( ~n10189 & n10538 ) | ( n10537 & n10538 ) ;
  assign n10540 = ( n10189 & n10537 ) | ( n10189 & n10538 ) | ( n10537 & n10538 ) ;
  assign n10541 = ( n10189 & n10539 ) | ( n10189 & ~n10540 ) | ( n10539 & ~n10540 ) ;
  assign n10542 = ( x94 & n10536 ) | ( x94 & ~n10541 ) | ( n10536 & ~n10541 ) ;
  assign n10543 = ( x94 & n10190 ) | ( x94 & ~n10363 ) | ( n10190 & ~n10363 ) ;
  assign n10544 = x94 & n10190 ;
  assign n10545 = ( n10195 & n10543 ) | ( n10195 & n10544 ) | ( n10543 & n10544 ) ;
  assign n10546 = ( ~n10195 & n10543 ) | ( ~n10195 & n10544 ) | ( n10543 & n10544 ) ;
  assign n10547 = ( n10195 & ~n10545 ) | ( n10195 & n10546 ) | ( ~n10545 & n10546 ) ;
  assign n10548 = ( x95 & n10542 ) | ( x95 & ~n10547 ) | ( n10542 & ~n10547 ) ;
  assign n10549 = ( x95 & n10196 ) | ( x95 & ~n10363 ) | ( n10196 & ~n10363 ) ;
  assign n10550 = x95 & n10196 ;
  assign n10551 = ( ~n10201 & n10549 ) | ( ~n10201 & n10550 ) | ( n10549 & n10550 ) ;
  assign n10552 = ( n10201 & n10549 ) | ( n10201 & n10550 ) | ( n10549 & n10550 ) ;
  assign n10553 = ( n10201 & n10551 ) | ( n10201 & ~n10552 ) | ( n10551 & ~n10552 ) ;
  assign n10554 = ( x96 & n10548 ) | ( x96 & ~n10553 ) | ( n10548 & ~n10553 ) ;
  assign n10555 = ( x96 & n10202 ) | ( x96 & ~n10363 ) | ( n10202 & ~n10363 ) ;
  assign n10556 = x96 & n10202 ;
  assign n10557 = ( n10207 & n10555 ) | ( n10207 & n10556 ) | ( n10555 & n10556 ) ;
  assign n10558 = ( ~n10207 & n10555 ) | ( ~n10207 & n10556 ) | ( n10555 & n10556 ) ;
  assign n10559 = ( n10207 & ~n10557 ) | ( n10207 & n10558 ) | ( ~n10557 & n10558 ) ;
  assign n10560 = ( x97 & n10554 ) | ( x97 & ~n10559 ) | ( n10554 & ~n10559 ) ;
  assign n10561 = ( x97 & n10208 ) | ( x97 & ~n10363 ) | ( n10208 & ~n10363 ) ;
  assign n10562 = x97 & n10208 ;
  assign n10563 = ( ~n10213 & n10561 ) | ( ~n10213 & n10562 ) | ( n10561 & n10562 ) ;
  assign n10564 = ( n10213 & n10561 ) | ( n10213 & n10562 ) | ( n10561 & n10562 ) ;
  assign n10565 = ( n10213 & n10563 ) | ( n10213 & ~n10564 ) | ( n10563 & ~n10564 ) ;
  assign n10566 = ( x98 & n10560 ) | ( x98 & ~n10565 ) | ( n10560 & ~n10565 ) ;
  assign n10567 = ( x98 & n10214 ) | ( x98 & ~n10363 ) | ( n10214 & ~n10363 ) ;
  assign n10568 = x98 & n10214 ;
  assign n10569 = ( n10219 & n10567 ) | ( n10219 & n10568 ) | ( n10567 & n10568 ) ;
  assign n10570 = ( ~n10219 & n10567 ) | ( ~n10219 & n10568 ) | ( n10567 & n10568 ) ;
  assign n10571 = ( n10219 & ~n10569 ) | ( n10219 & n10570 ) | ( ~n10569 & n10570 ) ;
  assign n10572 = ( x99 & n10566 ) | ( x99 & ~n10571 ) | ( n10566 & ~n10571 ) ;
  assign n10573 = ( x99 & n10220 ) | ( x99 & ~n10363 ) | ( n10220 & ~n10363 ) ;
  assign n10574 = x99 & n10220 ;
  assign n10575 = ( ~n10225 & n10573 ) | ( ~n10225 & n10574 ) | ( n10573 & n10574 ) ;
  assign n10576 = ( n10225 & n10573 ) | ( n10225 & n10574 ) | ( n10573 & n10574 ) ;
  assign n10577 = ( n10225 & n10575 ) | ( n10225 & ~n10576 ) | ( n10575 & ~n10576 ) ;
  assign n10578 = ( x100 & n10572 ) | ( x100 & ~n10577 ) | ( n10572 & ~n10577 ) ;
  assign n10579 = ( x100 & n10226 ) | ( x100 & ~n10363 ) | ( n10226 & ~n10363 ) ;
  assign n10580 = x100 & n10226 ;
  assign n10581 = ( n10231 & n10579 ) | ( n10231 & n10580 ) | ( n10579 & n10580 ) ;
  assign n10582 = ( ~n10231 & n10579 ) | ( ~n10231 & n10580 ) | ( n10579 & n10580 ) ;
  assign n10583 = ( n10231 & ~n10581 ) | ( n10231 & n10582 ) | ( ~n10581 & n10582 ) ;
  assign n10584 = ( x101 & n10578 ) | ( x101 & ~n10583 ) | ( n10578 & ~n10583 ) ;
  assign n10585 = ( x101 & n10232 ) | ( x101 & ~n10363 ) | ( n10232 & ~n10363 ) ;
  assign n10586 = x101 & n10232 ;
  assign n10587 = ( ~n10237 & n10585 ) | ( ~n10237 & n10586 ) | ( n10585 & n10586 ) ;
  assign n10588 = ( n10237 & n10585 ) | ( n10237 & n10586 ) | ( n10585 & n10586 ) ;
  assign n10589 = ( n10237 & n10587 ) | ( n10237 & ~n10588 ) | ( n10587 & ~n10588 ) ;
  assign n10590 = ( x102 & n10584 ) | ( x102 & ~n10589 ) | ( n10584 & ~n10589 ) ;
  assign n10591 = ( x102 & n10238 ) | ( x102 & ~n10363 ) | ( n10238 & ~n10363 ) ;
  assign n10592 = x102 & n10238 ;
  assign n10593 = ( n10243 & n10591 ) | ( n10243 & n10592 ) | ( n10591 & n10592 ) ;
  assign n10594 = ( ~n10243 & n10591 ) | ( ~n10243 & n10592 ) | ( n10591 & n10592 ) ;
  assign n10595 = ( n10243 & ~n10593 ) | ( n10243 & n10594 ) | ( ~n10593 & n10594 ) ;
  assign n10596 = ( x103 & n10590 ) | ( x103 & ~n10595 ) | ( n10590 & ~n10595 ) ;
  assign n10597 = ( x103 & n10244 ) | ( x103 & ~n10363 ) | ( n10244 & ~n10363 ) ;
  assign n10598 = x103 & n10244 ;
  assign n10599 = ( ~n10249 & n10597 ) | ( ~n10249 & n10598 ) | ( n10597 & n10598 ) ;
  assign n10600 = ( n10249 & n10597 ) | ( n10249 & n10598 ) | ( n10597 & n10598 ) ;
  assign n10601 = ( n10249 & n10599 ) | ( n10249 & ~n10600 ) | ( n10599 & ~n10600 ) ;
  assign n10602 = ( x104 & n10596 ) | ( x104 & ~n10601 ) | ( n10596 & ~n10601 ) ;
  assign n10603 = ( x104 & n10250 ) | ( x104 & ~n10363 ) | ( n10250 & ~n10363 ) ;
  assign n10604 = x104 & n10250 ;
  assign n10605 = ( n10255 & n10603 ) | ( n10255 & n10604 ) | ( n10603 & n10604 ) ;
  assign n10606 = ( ~n10255 & n10603 ) | ( ~n10255 & n10604 ) | ( n10603 & n10604 ) ;
  assign n10607 = ( n10255 & ~n10605 ) | ( n10255 & n10606 ) | ( ~n10605 & n10606 ) ;
  assign n10608 = ( x105 & n10602 ) | ( x105 & ~n10607 ) | ( n10602 & ~n10607 ) ;
  assign n10609 = ( x105 & n10256 ) | ( x105 & ~n10363 ) | ( n10256 & ~n10363 ) ;
  assign n10610 = x105 & n10256 ;
  assign n10611 = ( ~n10261 & n10609 ) | ( ~n10261 & n10610 ) | ( n10609 & n10610 ) ;
  assign n10612 = ( n10261 & n10609 ) | ( n10261 & n10610 ) | ( n10609 & n10610 ) ;
  assign n10613 = ( n10261 & n10611 ) | ( n10261 & ~n10612 ) | ( n10611 & ~n10612 ) ;
  assign n10614 = ( x106 & n10608 ) | ( x106 & ~n10613 ) | ( n10608 & ~n10613 ) ;
  assign n10615 = ( x106 & n10262 ) | ( x106 & ~n10363 ) | ( n10262 & ~n10363 ) ;
  assign n10616 = x106 & n10262 ;
  assign n10617 = ( n10267 & n10615 ) | ( n10267 & n10616 ) | ( n10615 & n10616 ) ;
  assign n10618 = ( ~n10267 & n10615 ) | ( ~n10267 & n10616 ) | ( n10615 & n10616 ) ;
  assign n10619 = ( n10267 & ~n10617 ) | ( n10267 & n10618 ) | ( ~n10617 & n10618 ) ;
  assign n10620 = ( x107 & n10614 ) | ( x107 & ~n10619 ) | ( n10614 & ~n10619 ) ;
  assign n10621 = ( x107 & n10268 ) | ( x107 & ~n10363 ) | ( n10268 & ~n10363 ) ;
  assign n10622 = x107 & n10268 ;
  assign n10623 = ( ~n10273 & n10621 ) | ( ~n10273 & n10622 ) | ( n10621 & n10622 ) ;
  assign n10624 = ( n10273 & n10621 ) | ( n10273 & n10622 ) | ( n10621 & n10622 ) ;
  assign n10625 = ( n10273 & n10623 ) | ( n10273 & ~n10624 ) | ( n10623 & ~n10624 ) ;
  assign n10626 = ( x108 & n10620 ) | ( x108 & ~n10625 ) | ( n10620 & ~n10625 ) ;
  assign n10627 = ( x108 & n10274 ) | ( x108 & ~n10363 ) | ( n10274 & ~n10363 ) ;
  assign n10628 = x108 & n10274 ;
  assign n10629 = ( n10279 & n10627 ) | ( n10279 & n10628 ) | ( n10627 & n10628 ) ;
  assign n10630 = ( ~n10279 & n10627 ) | ( ~n10279 & n10628 ) | ( n10627 & n10628 ) ;
  assign n10631 = ( n10279 & ~n10629 ) | ( n10279 & n10630 ) | ( ~n10629 & n10630 ) ;
  assign n10632 = ( x109 & n10626 ) | ( x109 & ~n10631 ) | ( n10626 & ~n10631 ) ;
  assign n10633 = ( x109 & n10280 ) | ( x109 & ~n10363 ) | ( n10280 & ~n10363 ) ;
  assign n10634 = x109 & n10280 ;
  assign n10635 = ( ~n10285 & n10633 ) | ( ~n10285 & n10634 ) | ( n10633 & n10634 ) ;
  assign n10636 = ( n10285 & n10633 ) | ( n10285 & n10634 ) | ( n10633 & n10634 ) ;
  assign n10637 = ( n10285 & n10635 ) | ( n10285 & ~n10636 ) | ( n10635 & ~n10636 ) ;
  assign n10638 = ( x110 & n10632 ) | ( x110 & ~n10637 ) | ( n10632 & ~n10637 ) ;
  assign n10639 = ( x110 & n10286 ) | ( x110 & ~n10363 ) | ( n10286 & ~n10363 ) ;
  assign n10640 = x110 & n10286 ;
  assign n10641 = ( n10291 & n10639 ) | ( n10291 & n10640 ) | ( n10639 & n10640 ) ;
  assign n10642 = ( ~n10291 & n10639 ) | ( ~n10291 & n10640 ) | ( n10639 & n10640 ) ;
  assign n10643 = ( n10291 & ~n10641 ) | ( n10291 & n10642 ) | ( ~n10641 & n10642 ) ;
  assign n10644 = ( x111 & n10638 ) | ( x111 & ~n10643 ) | ( n10638 & ~n10643 ) ;
  assign n10645 = ( x111 & n10292 ) | ( x111 & ~n10363 ) | ( n10292 & ~n10363 ) ;
  assign n10646 = x111 & n10292 ;
  assign n10647 = ( ~n10297 & n10645 ) | ( ~n10297 & n10646 ) | ( n10645 & n10646 ) ;
  assign n10648 = ( n10297 & n10645 ) | ( n10297 & n10646 ) | ( n10645 & n10646 ) ;
  assign n10649 = ( n10297 & n10647 ) | ( n10297 & ~n10648 ) | ( n10647 & ~n10648 ) ;
  assign n10650 = ( x112 & n10644 ) | ( x112 & ~n10649 ) | ( n10644 & ~n10649 ) ;
  assign n10651 = ( x112 & n10298 ) | ( x112 & ~n10363 ) | ( n10298 & ~n10363 ) ;
  assign n10652 = x112 & n10298 ;
  assign n10653 = ( n10303 & n10651 ) | ( n10303 & n10652 ) | ( n10651 & n10652 ) ;
  assign n10654 = ( ~n10303 & n10651 ) | ( ~n10303 & n10652 ) | ( n10651 & n10652 ) ;
  assign n10655 = ( n10303 & ~n10653 ) | ( n10303 & n10654 ) | ( ~n10653 & n10654 ) ;
  assign n10656 = ( x113 & n10650 ) | ( x113 & ~n10655 ) | ( n10650 & ~n10655 ) ;
  assign n10657 = ( x113 & n10304 ) | ( x113 & ~n10363 ) | ( n10304 & ~n10363 ) ;
  assign n10658 = x113 & n10304 ;
  assign n10659 = ( ~n10309 & n10657 ) | ( ~n10309 & n10658 ) | ( n10657 & n10658 ) ;
  assign n10660 = ( n10309 & n10657 ) | ( n10309 & n10658 ) | ( n10657 & n10658 ) ;
  assign n10661 = ( n10309 & n10659 ) | ( n10309 & ~n10660 ) | ( n10659 & ~n10660 ) ;
  assign n10662 = ( x114 & n10656 ) | ( x114 & ~n10661 ) | ( n10656 & ~n10661 ) ;
  assign n10663 = ( x114 & n10310 ) | ( x114 & ~n10363 ) | ( n10310 & ~n10363 ) ;
  assign n10664 = x114 & n10310 ;
  assign n10665 = ( n10315 & n10663 ) | ( n10315 & n10664 ) | ( n10663 & n10664 ) ;
  assign n10666 = ( ~n10315 & n10663 ) | ( ~n10315 & n10664 ) | ( n10663 & n10664 ) ;
  assign n10667 = ( n10315 & ~n10665 ) | ( n10315 & n10666 ) | ( ~n10665 & n10666 ) ;
  assign n10668 = ( x115 & n10662 ) | ( x115 & ~n10667 ) | ( n10662 & ~n10667 ) ;
  assign n10669 = ( x115 & n10316 ) | ( x115 & ~n10363 ) | ( n10316 & ~n10363 ) ;
  assign n10670 = x115 & n10316 ;
  assign n10671 = ( ~n10321 & n10669 ) | ( ~n10321 & n10670 ) | ( n10669 & n10670 ) ;
  assign n10672 = ( n10321 & n10669 ) | ( n10321 & n10670 ) | ( n10669 & n10670 ) ;
  assign n10673 = ( n10321 & n10671 ) | ( n10321 & ~n10672 ) | ( n10671 & ~n10672 ) ;
  assign n10674 = ( x116 & n10668 ) | ( x116 & ~n10673 ) | ( n10668 & ~n10673 ) ;
  assign n10675 = ( x116 & n10322 ) | ( x116 & ~n10363 ) | ( n10322 & ~n10363 ) ;
  assign n10676 = x116 & n10322 ;
  assign n10677 = ( n10327 & n10675 ) | ( n10327 & n10676 ) | ( n10675 & n10676 ) ;
  assign n10678 = ( ~n10327 & n10675 ) | ( ~n10327 & n10676 ) | ( n10675 & n10676 ) ;
  assign n10679 = ( n10327 & ~n10677 ) | ( n10327 & n10678 ) | ( ~n10677 & n10678 ) ;
  assign n10680 = ( x117 & n10674 ) | ( x117 & ~n10679 ) | ( n10674 & ~n10679 ) ;
  assign n10681 = ( x117 & n10328 ) | ( x117 & ~n10363 ) | ( n10328 & ~n10363 ) ;
  assign n10682 = x117 & n10328 ;
  assign n10683 = ( ~n10333 & n10681 ) | ( ~n10333 & n10682 ) | ( n10681 & n10682 ) ;
  assign n10684 = ( n10333 & n10681 ) | ( n10333 & n10682 ) | ( n10681 & n10682 ) ;
  assign n10685 = ( n10333 & n10683 ) | ( n10333 & ~n10684 ) | ( n10683 & ~n10684 ) ;
  assign n10686 = ( x118 & n10680 ) | ( x118 & ~n10685 ) | ( n10680 & ~n10685 ) ;
  assign n10687 = ( x118 & n10334 ) | ( x118 & ~n10363 ) | ( n10334 & ~n10363 ) ;
  assign n10688 = x118 & n10334 ;
  assign n10689 = ( n10339 & n10687 ) | ( n10339 & n10688 ) | ( n10687 & n10688 ) ;
  assign n10690 = ( ~n10339 & n10687 ) | ( ~n10339 & n10688 ) | ( n10687 & n10688 ) ;
  assign n10691 = ( n10339 & ~n10689 ) | ( n10339 & n10690 ) | ( ~n10689 & n10690 ) ;
  assign n10692 = ( x119 & n10686 ) | ( x119 & ~n10691 ) | ( n10686 & ~n10691 ) ;
  assign n10693 = ( x119 & n10340 ) | ( x119 & ~n10363 ) | ( n10340 & ~n10363 ) ;
  assign n10694 = x119 & n10340 ;
  assign n10695 = ( ~n10345 & n10693 ) | ( ~n10345 & n10694 ) | ( n10693 & n10694 ) ;
  assign n10696 = ( n10345 & n10693 ) | ( n10345 & n10694 ) | ( n10693 & n10694 ) ;
  assign n10697 = ( n10345 & n10695 ) | ( n10345 & ~n10696 ) | ( n10695 & ~n10696 ) ;
  assign n10698 = ( x120 & n10692 ) | ( x120 & ~n10697 ) | ( n10692 & ~n10697 ) ;
  assign n10699 = ( x120 & n10346 ) | ( x120 & ~n10363 ) | ( n10346 & ~n10363 ) ;
  assign n10700 = x120 & n10346 ;
  assign n10701 = ( n10351 & n10699 ) | ( n10351 & n10700 ) | ( n10699 & n10700 ) ;
  assign n10702 = ( ~n10351 & n10699 ) | ( ~n10351 & n10700 ) | ( n10699 & n10700 ) ;
  assign n10703 = ( n10351 & ~n10701 ) | ( n10351 & n10702 ) | ( ~n10701 & n10702 ) ;
  assign n10704 = ( x121 & n10698 ) | ( x121 & ~n10703 ) | ( n10698 & ~n10703 ) ;
  assign n10705 = ( x121 & n10352 ) | ( x121 & ~n10363 ) | ( n10352 & ~n10363 ) ;
  assign n10706 = x121 & n10352 ;
  assign n10707 = ( n10357 & n10705 ) | ( n10357 & n10706 ) | ( n10705 & n10706 ) ;
  assign n10708 = ( ~n10357 & n10705 ) | ( ~n10357 & n10706 ) | ( n10705 & n10706 ) ;
  assign n10709 = ( n10357 & ~n10707 ) | ( n10357 & n10708 ) | ( ~n10707 & n10708 ) ;
  assign n10710 = ( x122 & n10704 ) | ( x122 & ~n10709 ) | ( n10704 & ~n10709 ) ;
  assign n10711 = x123 | n10710 ;
  assign n10712 = ( x123 & n134 ) | ( x123 & n10710 ) | ( n134 & n10710 ) ;
  assign n10713 = ( n10361 & ~n10711 ) | ( n10361 & n10712 ) | ( ~n10711 & n10712 ) ;
  assign n10714 = ( x123 & ~n10361 ) | ( x123 & n10710 ) | ( ~n10361 & n10710 ) ;
  assign n10715 = n134 | n10714 ;
  assign n10716 = ( x4 & ~x64 ) | ( x4 & n10715 ) | ( ~x64 & n10715 ) ;
  assign n10717 = ~x4 & n10715 ;
  assign n10718 = ( n10367 & n10716 ) | ( n10367 & ~n10717 ) | ( n10716 & ~n10717 ) ;
  assign n10719 = ~x3 & x64 ;
  assign n10720 = ( x65 & ~n10718 ) | ( x65 & n10719 ) | ( ~n10718 & n10719 ) ;
  assign n10721 = ( x65 & n10367 ) | ( x65 & ~n10715 ) | ( n10367 & ~n10715 ) ;
  assign n10722 = x65 & n10367 ;
  assign n10723 = ( n10366 & n10721 ) | ( n10366 & n10722 ) | ( n10721 & n10722 ) ;
  assign n10724 = ( ~n10366 & n10721 ) | ( ~n10366 & n10722 ) | ( n10721 & n10722 ) ;
  assign n10725 = ( n10366 & ~n10723 ) | ( n10366 & n10724 ) | ( ~n10723 & n10724 ) ;
  assign n10726 = ( x66 & n10720 ) | ( x66 & ~n10725 ) | ( n10720 & ~n10725 ) ;
  assign n10727 = ( x66 & n10368 ) | ( x66 & ~n10715 ) | ( n10368 & ~n10715 ) ;
  assign n10728 = x66 & n10368 ;
  assign n10729 = ( n10373 & n10727 ) | ( n10373 & n10728 ) | ( n10727 & n10728 ) ;
  assign n10730 = ( ~n10373 & n10727 ) | ( ~n10373 & n10728 ) | ( n10727 & n10728 ) ;
  assign n10731 = ( n10373 & ~n10729 ) | ( n10373 & n10730 ) | ( ~n10729 & n10730 ) ;
  assign n10732 = ( x67 & n10726 ) | ( x67 & ~n10731 ) | ( n10726 & ~n10731 ) ;
  assign n10733 = ( x67 & n10374 ) | ( x67 & ~n10715 ) | ( n10374 & ~n10715 ) ;
  assign n10734 = x67 & n10374 ;
  assign n10735 = ( ~n10379 & n10733 ) | ( ~n10379 & n10734 ) | ( n10733 & n10734 ) ;
  assign n10736 = ( n10379 & n10733 ) | ( n10379 & n10734 ) | ( n10733 & n10734 ) ;
  assign n10737 = ( n10379 & n10735 ) | ( n10379 & ~n10736 ) | ( n10735 & ~n10736 ) ;
  assign n10738 = ( x68 & n10732 ) | ( x68 & ~n10737 ) | ( n10732 & ~n10737 ) ;
  assign n10739 = ( x68 & n10380 ) | ( x68 & ~n10715 ) | ( n10380 & ~n10715 ) ;
  assign n10740 = x68 & n10380 ;
  assign n10741 = ( n10385 & n10739 ) | ( n10385 & n10740 ) | ( n10739 & n10740 ) ;
  assign n10742 = ( ~n10385 & n10739 ) | ( ~n10385 & n10740 ) | ( n10739 & n10740 ) ;
  assign n10743 = ( n10385 & ~n10741 ) | ( n10385 & n10742 ) | ( ~n10741 & n10742 ) ;
  assign n10744 = ( x69 & n10738 ) | ( x69 & ~n10743 ) | ( n10738 & ~n10743 ) ;
  assign n10745 = ( x69 & n10386 ) | ( x69 & ~n10715 ) | ( n10386 & ~n10715 ) ;
  assign n10746 = x69 & n10386 ;
  assign n10747 = ( ~n10391 & n10745 ) | ( ~n10391 & n10746 ) | ( n10745 & n10746 ) ;
  assign n10748 = ( n10391 & n10745 ) | ( n10391 & n10746 ) | ( n10745 & n10746 ) ;
  assign n10749 = ( n10391 & n10747 ) | ( n10391 & ~n10748 ) | ( n10747 & ~n10748 ) ;
  assign n10750 = ( x70 & n10744 ) | ( x70 & ~n10749 ) | ( n10744 & ~n10749 ) ;
  assign n10751 = ( x70 & n10392 ) | ( x70 & ~n10715 ) | ( n10392 & ~n10715 ) ;
  assign n10752 = x70 & n10392 ;
  assign n10753 = ( n10397 & n10751 ) | ( n10397 & n10752 ) | ( n10751 & n10752 ) ;
  assign n10754 = ( ~n10397 & n10751 ) | ( ~n10397 & n10752 ) | ( n10751 & n10752 ) ;
  assign n10755 = ( n10397 & ~n10753 ) | ( n10397 & n10754 ) | ( ~n10753 & n10754 ) ;
  assign n10756 = ( x71 & n10750 ) | ( x71 & ~n10755 ) | ( n10750 & ~n10755 ) ;
  assign n10757 = ( x71 & n10398 ) | ( x71 & ~n10715 ) | ( n10398 & ~n10715 ) ;
  assign n10758 = x71 & n10398 ;
  assign n10759 = ( ~n10403 & n10757 ) | ( ~n10403 & n10758 ) | ( n10757 & n10758 ) ;
  assign n10760 = ( n10403 & n10757 ) | ( n10403 & n10758 ) | ( n10757 & n10758 ) ;
  assign n10761 = ( n10403 & n10759 ) | ( n10403 & ~n10760 ) | ( n10759 & ~n10760 ) ;
  assign n10762 = ( x72 & n10756 ) | ( x72 & ~n10761 ) | ( n10756 & ~n10761 ) ;
  assign n10763 = ( x72 & n10404 ) | ( x72 & ~n10715 ) | ( n10404 & ~n10715 ) ;
  assign n10764 = x72 & n10404 ;
  assign n10765 = ( n10409 & n10763 ) | ( n10409 & n10764 ) | ( n10763 & n10764 ) ;
  assign n10766 = ( ~n10409 & n10763 ) | ( ~n10409 & n10764 ) | ( n10763 & n10764 ) ;
  assign n10767 = ( n10409 & ~n10765 ) | ( n10409 & n10766 ) | ( ~n10765 & n10766 ) ;
  assign n10768 = ( x73 & n10762 ) | ( x73 & ~n10767 ) | ( n10762 & ~n10767 ) ;
  assign n10769 = ( x73 & n10410 ) | ( x73 & ~n10715 ) | ( n10410 & ~n10715 ) ;
  assign n10770 = x73 & n10410 ;
  assign n10771 = ( ~n10415 & n10769 ) | ( ~n10415 & n10770 ) | ( n10769 & n10770 ) ;
  assign n10772 = ( n10415 & n10769 ) | ( n10415 & n10770 ) | ( n10769 & n10770 ) ;
  assign n10773 = ( n10415 & n10771 ) | ( n10415 & ~n10772 ) | ( n10771 & ~n10772 ) ;
  assign n10774 = ( x74 & n10768 ) | ( x74 & ~n10773 ) | ( n10768 & ~n10773 ) ;
  assign n10775 = ( x74 & n10416 ) | ( x74 & ~n10715 ) | ( n10416 & ~n10715 ) ;
  assign n10776 = x74 & n10416 ;
  assign n10777 = ( n10421 & n10775 ) | ( n10421 & n10776 ) | ( n10775 & n10776 ) ;
  assign n10778 = ( ~n10421 & n10775 ) | ( ~n10421 & n10776 ) | ( n10775 & n10776 ) ;
  assign n10779 = ( n10421 & ~n10777 ) | ( n10421 & n10778 ) | ( ~n10777 & n10778 ) ;
  assign n10780 = ( x75 & n10774 ) | ( x75 & ~n10779 ) | ( n10774 & ~n10779 ) ;
  assign n10781 = ( x75 & n10422 ) | ( x75 & ~n10715 ) | ( n10422 & ~n10715 ) ;
  assign n10782 = x75 & n10422 ;
  assign n10783 = ( ~n10427 & n10781 ) | ( ~n10427 & n10782 ) | ( n10781 & n10782 ) ;
  assign n10784 = ( n10427 & n10781 ) | ( n10427 & n10782 ) | ( n10781 & n10782 ) ;
  assign n10785 = ( n10427 & n10783 ) | ( n10427 & ~n10784 ) | ( n10783 & ~n10784 ) ;
  assign n10786 = ( x76 & n10780 ) | ( x76 & ~n10785 ) | ( n10780 & ~n10785 ) ;
  assign n10787 = ( x76 & n10428 ) | ( x76 & ~n10715 ) | ( n10428 & ~n10715 ) ;
  assign n10788 = x76 & n10428 ;
  assign n10789 = ( n10433 & n10787 ) | ( n10433 & n10788 ) | ( n10787 & n10788 ) ;
  assign n10790 = ( ~n10433 & n10787 ) | ( ~n10433 & n10788 ) | ( n10787 & n10788 ) ;
  assign n10791 = ( n10433 & ~n10789 ) | ( n10433 & n10790 ) | ( ~n10789 & n10790 ) ;
  assign n10792 = ( x77 & n10786 ) | ( x77 & ~n10791 ) | ( n10786 & ~n10791 ) ;
  assign n10793 = ( x77 & n10434 ) | ( x77 & ~n10715 ) | ( n10434 & ~n10715 ) ;
  assign n10794 = x77 & n10434 ;
  assign n10795 = ( ~n10439 & n10793 ) | ( ~n10439 & n10794 ) | ( n10793 & n10794 ) ;
  assign n10796 = ( n10439 & n10793 ) | ( n10439 & n10794 ) | ( n10793 & n10794 ) ;
  assign n10797 = ( n10439 & n10795 ) | ( n10439 & ~n10796 ) | ( n10795 & ~n10796 ) ;
  assign n10798 = ( x78 & n10792 ) | ( x78 & ~n10797 ) | ( n10792 & ~n10797 ) ;
  assign n10799 = ( x78 & n10440 ) | ( x78 & ~n10715 ) | ( n10440 & ~n10715 ) ;
  assign n10800 = x78 & n10440 ;
  assign n10801 = ( n10445 & n10799 ) | ( n10445 & n10800 ) | ( n10799 & n10800 ) ;
  assign n10802 = ( ~n10445 & n10799 ) | ( ~n10445 & n10800 ) | ( n10799 & n10800 ) ;
  assign n10803 = ( n10445 & ~n10801 ) | ( n10445 & n10802 ) | ( ~n10801 & n10802 ) ;
  assign n10804 = ( x79 & n10798 ) | ( x79 & ~n10803 ) | ( n10798 & ~n10803 ) ;
  assign n10805 = ( x79 & n10446 ) | ( x79 & ~n10715 ) | ( n10446 & ~n10715 ) ;
  assign n10806 = x79 & n10446 ;
  assign n10807 = ( ~n10451 & n10805 ) | ( ~n10451 & n10806 ) | ( n10805 & n10806 ) ;
  assign n10808 = ( n10451 & n10805 ) | ( n10451 & n10806 ) | ( n10805 & n10806 ) ;
  assign n10809 = ( n10451 & n10807 ) | ( n10451 & ~n10808 ) | ( n10807 & ~n10808 ) ;
  assign n10810 = ( x80 & n10804 ) | ( x80 & ~n10809 ) | ( n10804 & ~n10809 ) ;
  assign n10811 = ( x80 & n10452 ) | ( x80 & ~n10715 ) | ( n10452 & ~n10715 ) ;
  assign n10812 = x80 & n10452 ;
  assign n10813 = ( n10457 & n10811 ) | ( n10457 & n10812 ) | ( n10811 & n10812 ) ;
  assign n10814 = ( ~n10457 & n10811 ) | ( ~n10457 & n10812 ) | ( n10811 & n10812 ) ;
  assign n10815 = ( n10457 & ~n10813 ) | ( n10457 & n10814 ) | ( ~n10813 & n10814 ) ;
  assign n10816 = ( x81 & n10810 ) | ( x81 & ~n10815 ) | ( n10810 & ~n10815 ) ;
  assign n10817 = ( x81 & n10458 ) | ( x81 & ~n10715 ) | ( n10458 & ~n10715 ) ;
  assign n10818 = x81 & n10458 ;
  assign n10819 = ( ~n10463 & n10817 ) | ( ~n10463 & n10818 ) | ( n10817 & n10818 ) ;
  assign n10820 = ( n10463 & n10817 ) | ( n10463 & n10818 ) | ( n10817 & n10818 ) ;
  assign n10821 = ( n10463 & n10819 ) | ( n10463 & ~n10820 ) | ( n10819 & ~n10820 ) ;
  assign n10822 = ( x82 & n10816 ) | ( x82 & ~n10821 ) | ( n10816 & ~n10821 ) ;
  assign n10823 = ( x82 & n10464 ) | ( x82 & ~n10715 ) | ( n10464 & ~n10715 ) ;
  assign n10824 = x82 & n10464 ;
  assign n10825 = ( n10469 & n10823 ) | ( n10469 & n10824 ) | ( n10823 & n10824 ) ;
  assign n10826 = ( ~n10469 & n10823 ) | ( ~n10469 & n10824 ) | ( n10823 & n10824 ) ;
  assign n10827 = ( n10469 & ~n10825 ) | ( n10469 & n10826 ) | ( ~n10825 & n10826 ) ;
  assign n10828 = ( x83 & n10822 ) | ( x83 & ~n10827 ) | ( n10822 & ~n10827 ) ;
  assign n10829 = ( x83 & n10470 ) | ( x83 & ~n10715 ) | ( n10470 & ~n10715 ) ;
  assign n10830 = x83 & n10470 ;
  assign n10831 = ( ~n10475 & n10829 ) | ( ~n10475 & n10830 ) | ( n10829 & n10830 ) ;
  assign n10832 = ( n10475 & n10829 ) | ( n10475 & n10830 ) | ( n10829 & n10830 ) ;
  assign n10833 = ( n10475 & n10831 ) | ( n10475 & ~n10832 ) | ( n10831 & ~n10832 ) ;
  assign n10834 = ( x84 & n10828 ) | ( x84 & ~n10833 ) | ( n10828 & ~n10833 ) ;
  assign n10835 = ( x84 & n10476 ) | ( x84 & ~n10715 ) | ( n10476 & ~n10715 ) ;
  assign n10836 = x84 & n10476 ;
  assign n10837 = ( n10481 & n10835 ) | ( n10481 & n10836 ) | ( n10835 & n10836 ) ;
  assign n10838 = ( ~n10481 & n10835 ) | ( ~n10481 & n10836 ) | ( n10835 & n10836 ) ;
  assign n10839 = ( n10481 & ~n10837 ) | ( n10481 & n10838 ) | ( ~n10837 & n10838 ) ;
  assign n10840 = ( x85 & n10834 ) | ( x85 & ~n10839 ) | ( n10834 & ~n10839 ) ;
  assign n10841 = ( x85 & n10482 ) | ( x85 & ~n10715 ) | ( n10482 & ~n10715 ) ;
  assign n10842 = x85 & n10482 ;
  assign n10843 = ( ~n10487 & n10841 ) | ( ~n10487 & n10842 ) | ( n10841 & n10842 ) ;
  assign n10844 = ( n10487 & n10841 ) | ( n10487 & n10842 ) | ( n10841 & n10842 ) ;
  assign n10845 = ( n10487 & n10843 ) | ( n10487 & ~n10844 ) | ( n10843 & ~n10844 ) ;
  assign n10846 = ( x86 & n10840 ) | ( x86 & ~n10845 ) | ( n10840 & ~n10845 ) ;
  assign n10847 = ( x86 & n10488 ) | ( x86 & ~n10715 ) | ( n10488 & ~n10715 ) ;
  assign n10848 = x86 & n10488 ;
  assign n10849 = ( n10493 & n10847 ) | ( n10493 & n10848 ) | ( n10847 & n10848 ) ;
  assign n10850 = ( ~n10493 & n10847 ) | ( ~n10493 & n10848 ) | ( n10847 & n10848 ) ;
  assign n10851 = ( n10493 & ~n10849 ) | ( n10493 & n10850 ) | ( ~n10849 & n10850 ) ;
  assign n10852 = ( x87 & n10846 ) | ( x87 & ~n10851 ) | ( n10846 & ~n10851 ) ;
  assign n10853 = ( x87 & n10494 ) | ( x87 & ~n10715 ) | ( n10494 & ~n10715 ) ;
  assign n10854 = x87 & n10494 ;
  assign n10855 = ( ~n10499 & n10853 ) | ( ~n10499 & n10854 ) | ( n10853 & n10854 ) ;
  assign n10856 = ( n10499 & n10853 ) | ( n10499 & n10854 ) | ( n10853 & n10854 ) ;
  assign n10857 = ( n10499 & n10855 ) | ( n10499 & ~n10856 ) | ( n10855 & ~n10856 ) ;
  assign n10858 = ( x88 & n10852 ) | ( x88 & ~n10857 ) | ( n10852 & ~n10857 ) ;
  assign n10859 = ( x88 & n10500 ) | ( x88 & ~n10715 ) | ( n10500 & ~n10715 ) ;
  assign n10860 = x88 & n10500 ;
  assign n10861 = ( n10505 & n10859 ) | ( n10505 & n10860 ) | ( n10859 & n10860 ) ;
  assign n10862 = ( ~n10505 & n10859 ) | ( ~n10505 & n10860 ) | ( n10859 & n10860 ) ;
  assign n10863 = ( n10505 & ~n10861 ) | ( n10505 & n10862 ) | ( ~n10861 & n10862 ) ;
  assign n10864 = ( x89 & n10858 ) | ( x89 & ~n10863 ) | ( n10858 & ~n10863 ) ;
  assign n10865 = ( x89 & n10506 ) | ( x89 & ~n10715 ) | ( n10506 & ~n10715 ) ;
  assign n10866 = x89 & n10506 ;
  assign n10867 = ( ~n10511 & n10865 ) | ( ~n10511 & n10866 ) | ( n10865 & n10866 ) ;
  assign n10868 = ( n10511 & n10865 ) | ( n10511 & n10866 ) | ( n10865 & n10866 ) ;
  assign n10869 = ( n10511 & n10867 ) | ( n10511 & ~n10868 ) | ( n10867 & ~n10868 ) ;
  assign n10870 = ( x90 & n10864 ) | ( x90 & ~n10869 ) | ( n10864 & ~n10869 ) ;
  assign n10871 = ( x90 & n10512 ) | ( x90 & ~n10715 ) | ( n10512 & ~n10715 ) ;
  assign n10872 = x90 & n10512 ;
  assign n10873 = ( n10517 & n10871 ) | ( n10517 & n10872 ) | ( n10871 & n10872 ) ;
  assign n10874 = ( ~n10517 & n10871 ) | ( ~n10517 & n10872 ) | ( n10871 & n10872 ) ;
  assign n10875 = ( n10517 & ~n10873 ) | ( n10517 & n10874 ) | ( ~n10873 & n10874 ) ;
  assign n10876 = ( x91 & n10870 ) | ( x91 & ~n10875 ) | ( n10870 & ~n10875 ) ;
  assign n10877 = ( x91 & n10518 ) | ( x91 & ~n10715 ) | ( n10518 & ~n10715 ) ;
  assign n10878 = x91 & n10518 ;
  assign n10879 = ( ~n10523 & n10877 ) | ( ~n10523 & n10878 ) | ( n10877 & n10878 ) ;
  assign n10880 = ( n10523 & n10877 ) | ( n10523 & n10878 ) | ( n10877 & n10878 ) ;
  assign n10881 = ( n10523 & n10879 ) | ( n10523 & ~n10880 ) | ( n10879 & ~n10880 ) ;
  assign n10882 = ( x92 & n10876 ) | ( x92 & ~n10881 ) | ( n10876 & ~n10881 ) ;
  assign n10883 = ( x92 & n10524 ) | ( x92 & ~n10715 ) | ( n10524 & ~n10715 ) ;
  assign n10884 = x92 & n10524 ;
  assign n10885 = ( n10529 & n10883 ) | ( n10529 & n10884 ) | ( n10883 & n10884 ) ;
  assign n10886 = ( ~n10529 & n10883 ) | ( ~n10529 & n10884 ) | ( n10883 & n10884 ) ;
  assign n10887 = ( n10529 & ~n10885 ) | ( n10529 & n10886 ) | ( ~n10885 & n10886 ) ;
  assign n10888 = ( x93 & n10882 ) | ( x93 & ~n10887 ) | ( n10882 & ~n10887 ) ;
  assign n10889 = ( x93 & n10530 ) | ( x93 & ~n10715 ) | ( n10530 & ~n10715 ) ;
  assign n10890 = x93 & n10530 ;
  assign n10891 = ( ~n10535 & n10889 ) | ( ~n10535 & n10890 ) | ( n10889 & n10890 ) ;
  assign n10892 = ( n10535 & n10889 ) | ( n10535 & n10890 ) | ( n10889 & n10890 ) ;
  assign n10893 = ( n10535 & n10891 ) | ( n10535 & ~n10892 ) | ( n10891 & ~n10892 ) ;
  assign n10894 = ( x94 & n10888 ) | ( x94 & ~n10893 ) | ( n10888 & ~n10893 ) ;
  assign n10895 = ( x94 & n10536 ) | ( x94 & ~n10715 ) | ( n10536 & ~n10715 ) ;
  assign n10896 = x94 & n10536 ;
  assign n10897 = ( n10541 & n10895 ) | ( n10541 & n10896 ) | ( n10895 & n10896 ) ;
  assign n10898 = ( ~n10541 & n10895 ) | ( ~n10541 & n10896 ) | ( n10895 & n10896 ) ;
  assign n10899 = ( n10541 & ~n10897 ) | ( n10541 & n10898 ) | ( ~n10897 & n10898 ) ;
  assign n10900 = ( x95 & n10894 ) | ( x95 & ~n10899 ) | ( n10894 & ~n10899 ) ;
  assign n10901 = ( x95 & n10542 ) | ( x95 & ~n10715 ) | ( n10542 & ~n10715 ) ;
  assign n10902 = x95 & n10542 ;
  assign n10903 = ( ~n10547 & n10901 ) | ( ~n10547 & n10902 ) | ( n10901 & n10902 ) ;
  assign n10904 = ( n10547 & n10901 ) | ( n10547 & n10902 ) | ( n10901 & n10902 ) ;
  assign n10905 = ( n10547 & n10903 ) | ( n10547 & ~n10904 ) | ( n10903 & ~n10904 ) ;
  assign n10906 = ( x96 & n10900 ) | ( x96 & ~n10905 ) | ( n10900 & ~n10905 ) ;
  assign n10907 = ( x96 & n10548 ) | ( x96 & ~n10715 ) | ( n10548 & ~n10715 ) ;
  assign n10908 = x96 & n10548 ;
  assign n10909 = ( n10553 & n10907 ) | ( n10553 & n10908 ) | ( n10907 & n10908 ) ;
  assign n10910 = ( ~n10553 & n10907 ) | ( ~n10553 & n10908 ) | ( n10907 & n10908 ) ;
  assign n10911 = ( n10553 & ~n10909 ) | ( n10553 & n10910 ) | ( ~n10909 & n10910 ) ;
  assign n10912 = ( x97 & n10906 ) | ( x97 & ~n10911 ) | ( n10906 & ~n10911 ) ;
  assign n10913 = ( x97 & n10554 ) | ( x97 & ~n10715 ) | ( n10554 & ~n10715 ) ;
  assign n10914 = x97 & n10554 ;
  assign n10915 = ( ~n10559 & n10913 ) | ( ~n10559 & n10914 ) | ( n10913 & n10914 ) ;
  assign n10916 = ( n10559 & n10913 ) | ( n10559 & n10914 ) | ( n10913 & n10914 ) ;
  assign n10917 = ( n10559 & n10915 ) | ( n10559 & ~n10916 ) | ( n10915 & ~n10916 ) ;
  assign n10918 = ( x98 & n10912 ) | ( x98 & ~n10917 ) | ( n10912 & ~n10917 ) ;
  assign n10919 = ( x98 & n10560 ) | ( x98 & ~n10715 ) | ( n10560 & ~n10715 ) ;
  assign n10920 = x98 & n10560 ;
  assign n10921 = ( n10565 & n10919 ) | ( n10565 & n10920 ) | ( n10919 & n10920 ) ;
  assign n10922 = ( ~n10565 & n10919 ) | ( ~n10565 & n10920 ) | ( n10919 & n10920 ) ;
  assign n10923 = ( n10565 & ~n10921 ) | ( n10565 & n10922 ) | ( ~n10921 & n10922 ) ;
  assign n10924 = ( x99 & n10918 ) | ( x99 & ~n10923 ) | ( n10918 & ~n10923 ) ;
  assign n10925 = ( x99 & n10566 ) | ( x99 & ~n10715 ) | ( n10566 & ~n10715 ) ;
  assign n10926 = x99 & n10566 ;
  assign n10927 = ( ~n10571 & n10925 ) | ( ~n10571 & n10926 ) | ( n10925 & n10926 ) ;
  assign n10928 = ( n10571 & n10925 ) | ( n10571 & n10926 ) | ( n10925 & n10926 ) ;
  assign n10929 = ( n10571 & n10927 ) | ( n10571 & ~n10928 ) | ( n10927 & ~n10928 ) ;
  assign n10930 = ( x100 & n10924 ) | ( x100 & ~n10929 ) | ( n10924 & ~n10929 ) ;
  assign n10931 = ( x100 & n10572 ) | ( x100 & ~n10715 ) | ( n10572 & ~n10715 ) ;
  assign n10932 = x100 & n10572 ;
  assign n10933 = ( n10577 & n10931 ) | ( n10577 & n10932 ) | ( n10931 & n10932 ) ;
  assign n10934 = ( ~n10577 & n10931 ) | ( ~n10577 & n10932 ) | ( n10931 & n10932 ) ;
  assign n10935 = ( n10577 & ~n10933 ) | ( n10577 & n10934 ) | ( ~n10933 & n10934 ) ;
  assign n10936 = ( x101 & n10930 ) | ( x101 & ~n10935 ) | ( n10930 & ~n10935 ) ;
  assign n10937 = ( x101 & n10578 ) | ( x101 & ~n10715 ) | ( n10578 & ~n10715 ) ;
  assign n10938 = x101 & n10578 ;
  assign n10939 = ( ~n10583 & n10937 ) | ( ~n10583 & n10938 ) | ( n10937 & n10938 ) ;
  assign n10940 = ( n10583 & n10937 ) | ( n10583 & n10938 ) | ( n10937 & n10938 ) ;
  assign n10941 = ( n10583 & n10939 ) | ( n10583 & ~n10940 ) | ( n10939 & ~n10940 ) ;
  assign n10942 = ( x102 & n10936 ) | ( x102 & ~n10941 ) | ( n10936 & ~n10941 ) ;
  assign n10943 = ( x102 & n10584 ) | ( x102 & ~n10715 ) | ( n10584 & ~n10715 ) ;
  assign n10944 = x102 & n10584 ;
  assign n10945 = ( n10589 & n10943 ) | ( n10589 & n10944 ) | ( n10943 & n10944 ) ;
  assign n10946 = ( ~n10589 & n10943 ) | ( ~n10589 & n10944 ) | ( n10943 & n10944 ) ;
  assign n10947 = ( n10589 & ~n10945 ) | ( n10589 & n10946 ) | ( ~n10945 & n10946 ) ;
  assign n10948 = ( x103 & n10942 ) | ( x103 & ~n10947 ) | ( n10942 & ~n10947 ) ;
  assign n10949 = ( x103 & n10590 ) | ( x103 & ~n10715 ) | ( n10590 & ~n10715 ) ;
  assign n10950 = x103 & n10590 ;
  assign n10951 = ( ~n10595 & n10949 ) | ( ~n10595 & n10950 ) | ( n10949 & n10950 ) ;
  assign n10952 = ( n10595 & n10949 ) | ( n10595 & n10950 ) | ( n10949 & n10950 ) ;
  assign n10953 = ( n10595 & n10951 ) | ( n10595 & ~n10952 ) | ( n10951 & ~n10952 ) ;
  assign n10954 = ( x104 & n10948 ) | ( x104 & ~n10953 ) | ( n10948 & ~n10953 ) ;
  assign n10955 = ( x104 & n10596 ) | ( x104 & ~n10715 ) | ( n10596 & ~n10715 ) ;
  assign n10956 = x104 & n10596 ;
  assign n10957 = ( n10601 & n10955 ) | ( n10601 & n10956 ) | ( n10955 & n10956 ) ;
  assign n10958 = ( ~n10601 & n10955 ) | ( ~n10601 & n10956 ) | ( n10955 & n10956 ) ;
  assign n10959 = ( n10601 & ~n10957 ) | ( n10601 & n10958 ) | ( ~n10957 & n10958 ) ;
  assign n10960 = ( x105 & n10954 ) | ( x105 & ~n10959 ) | ( n10954 & ~n10959 ) ;
  assign n10961 = ( x105 & n10602 ) | ( x105 & ~n10715 ) | ( n10602 & ~n10715 ) ;
  assign n10962 = x105 & n10602 ;
  assign n10963 = ( ~n10607 & n10961 ) | ( ~n10607 & n10962 ) | ( n10961 & n10962 ) ;
  assign n10964 = ( n10607 & n10961 ) | ( n10607 & n10962 ) | ( n10961 & n10962 ) ;
  assign n10965 = ( n10607 & n10963 ) | ( n10607 & ~n10964 ) | ( n10963 & ~n10964 ) ;
  assign n10966 = ( x106 & n10960 ) | ( x106 & ~n10965 ) | ( n10960 & ~n10965 ) ;
  assign n10967 = ( x106 & n10608 ) | ( x106 & ~n10715 ) | ( n10608 & ~n10715 ) ;
  assign n10968 = x106 & n10608 ;
  assign n10969 = ( n10613 & n10967 ) | ( n10613 & n10968 ) | ( n10967 & n10968 ) ;
  assign n10970 = ( ~n10613 & n10967 ) | ( ~n10613 & n10968 ) | ( n10967 & n10968 ) ;
  assign n10971 = ( n10613 & ~n10969 ) | ( n10613 & n10970 ) | ( ~n10969 & n10970 ) ;
  assign n10972 = ( x107 & n10966 ) | ( x107 & ~n10971 ) | ( n10966 & ~n10971 ) ;
  assign n10973 = ( x107 & n10614 ) | ( x107 & ~n10715 ) | ( n10614 & ~n10715 ) ;
  assign n10974 = x107 & n10614 ;
  assign n10975 = ( ~n10619 & n10973 ) | ( ~n10619 & n10974 ) | ( n10973 & n10974 ) ;
  assign n10976 = ( n10619 & n10973 ) | ( n10619 & n10974 ) | ( n10973 & n10974 ) ;
  assign n10977 = ( n10619 & n10975 ) | ( n10619 & ~n10976 ) | ( n10975 & ~n10976 ) ;
  assign n10978 = ( x108 & n10972 ) | ( x108 & ~n10977 ) | ( n10972 & ~n10977 ) ;
  assign n10979 = ( x108 & n10620 ) | ( x108 & ~n10715 ) | ( n10620 & ~n10715 ) ;
  assign n10980 = x108 & n10620 ;
  assign n10981 = ( n10625 & n10979 ) | ( n10625 & n10980 ) | ( n10979 & n10980 ) ;
  assign n10982 = ( ~n10625 & n10979 ) | ( ~n10625 & n10980 ) | ( n10979 & n10980 ) ;
  assign n10983 = ( n10625 & ~n10981 ) | ( n10625 & n10982 ) | ( ~n10981 & n10982 ) ;
  assign n10984 = ( x109 & n10978 ) | ( x109 & ~n10983 ) | ( n10978 & ~n10983 ) ;
  assign n10985 = ( x109 & n10626 ) | ( x109 & ~n10715 ) | ( n10626 & ~n10715 ) ;
  assign n10986 = x109 & n10626 ;
  assign n10987 = ( ~n10631 & n10985 ) | ( ~n10631 & n10986 ) | ( n10985 & n10986 ) ;
  assign n10988 = ( n10631 & n10985 ) | ( n10631 & n10986 ) | ( n10985 & n10986 ) ;
  assign n10989 = ( n10631 & n10987 ) | ( n10631 & ~n10988 ) | ( n10987 & ~n10988 ) ;
  assign n10990 = ( x110 & n10984 ) | ( x110 & ~n10989 ) | ( n10984 & ~n10989 ) ;
  assign n10991 = ( x110 & n10632 ) | ( x110 & ~n10715 ) | ( n10632 & ~n10715 ) ;
  assign n10992 = x110 & n10632 ;
  assign n10993 = ( n10637 & n10991 ) | ( n10637 & n10992 ) | ( n10991 & n10992 ) ;
  assign n10994 = ( ~n10637 & n10991 ) | ( ~n10637 & n10992 ) | ( n10991 & n10992 ) ;
  assign n10995 = ( n10637 & ~n10993 ) | ( n10637 & n10994 ) | ( ~n10993 & n10994 ) ;
  assign n10996 = ( x111 & n10990 ) | ( x111 & ~n10995 ) | ( n10990 & ~n10995 ) ;
  assign n10997 = ( x111 & n10638 ) | ( x111 & ~n10715 ) | ( n10638 & ~n10715 ) ;
  assign n10998 = x111 & n10638 ;
  assign n10999 = ( ~n10643 & n10997 ) | ( ~n10643 & n10998 ) | ( n10997 & n10998 ) ;
  assign n11000 = ( n10643 & n10997 ) | ( n10643 & n10998 ) | ( n10997 & n10998 ) ;
  assign n11001 = ( n10643 & n10999 ) | ( n10643 & ~n11000 ) | ( n10999 & ~n11000 ) ;
  assign n11002 = ( x112 & n10996 ) | ( x112 & ~n11001 ) | ( n10996 & ~n11001 ) ;
  assign n11003 = ( x112 & n10644 ) | ( x112 & ~n10715 ) | ( n10644 & ~n10715 ) ;
  assign n11004 = x112 & n10644 ;
  assign n11005 = ( n10649 & n11003 ) | ( n10649 & n11004 ) | ( n11003 & n11004 ) ;
  assign n11006 = ( ~n10649 & n11003 ) | ( ~n10649 & n11004 ) | ( n11003 & n11004 ) ;
  assign n11007 = ( n10649 & ~n11005 ) | ( n10649 & n11006 ) | ( ~n11005 & n11006 ) ;
  assign n11008 = ( x113 & n11002 ) | ( x113 & ~n11007 ) | ( n11002 & ~n11007 ) ;
  assign n11009 = ( x113 & n10650 ) | ( x113 & ~n10715 ) | ( n10650 & ~n10715 ) ;
  assign n11010 = x113 & n10650 ;
  assign n11011 = ( ~n10655 & n11009 ) | ( ~n10655 & n11010 ) | ( n11009 & n11010 ) ;
  assign n11012 = ( n10655 & n11009 ) | ( n10655 & n11010 ) | ( n11009 & n11010 ) ;
  assign n11013 = ( n10655 & n11011 ) | ( n10655 & ~n11012 ) | ( n11011 & ~n11012 ) ;
  assign n11014 = ( x114 & n11008 ) | ( x114 & ~n11013 ) | ( n11008 & ~n11013 ) ;
  assign n11015 = ( x114 & n10656 ) | ( x114 & ~n10715 ) | ( n10656 & ~n10715 ) ;
  assign n11016 = x114 & n10656 ;
  assign n11017 = ( n10661 & n11015 ) | ( n10661 & n11016 ) | ( n11015 & n11016 ) ;
  assign n11018 = ( ~n10661 & n11015 ) | ( ~n10661 & n11016 ) | ( n11015 & n11016 ) ;
  assign n11019 = ( n10661 & ~n11017 ) | ( n10661 & n11018 ) | ( ~n11017 & n11018 ) ;
  assign n11020 = ( x115 & n11014 ) | ( x115 & ~n11019 ) | ( n11014 & ~n11019 ) ;
  assign n11021 = ( x115 & n10662 ) | ( x115 & ~n10715 ) | ( n10662 & ~n10715 ) ;
  assign n11022 = x115 & n10662 ;
  assign n11023 = ( ~n10667 & n11021 ) | ( ~n10667 & n11022 ) | ( n11021 & n11022 ) ;
  assign n11024 = ( n10667 & n11021 ) | ( n10667 & n11022 ) | ( n11021 & n11022 ) ;
  assign n11025 = ( n10667 & n11023 ) | ( n10667 & ~n11024 ) | ( n11023 & ~n11024 ) ;
  assign n11026 = ( x116 & n11020 ) | ( x116 & ~n11025 ) | ( n11020 & ~n11025 ) ;
  assign n11027 = ( x116 & n10668 ) | ( x116 & ~n10715 ) | ( n10668 & ~n10715 ) ;
  assign n11028 = x116 & n10668 ;
  assign n11029 = ( n10673 & n11027 ) | ( n10673 & n11028 ) | ( n11027 & n11028 ) ;
  assign n11030 = ( ~n10673 & n11027 ) | ( ~n10673 & n11028 ) | ( n11027 & n11028 ) ;
  assign n11031 = ( n10673 & ~n11029 ) | ( n10673 & n11030 ) | ( ~n11029 & n11030 ) ;
  assign n11032 = ( x117 & n11026 ) | ( x117 & ~n11031 ) | ( n11026 & ~n11031 ) ;
  assign n11033 = ( x117 & n10674 ) | ( x117 & ~n10715 ) | ( n10674 & ~n10715 ) ;
  assign n11034 = x117 & n10674 ;
  assign n11035 = ( ~n10679 & n11033 ) | ( ~n10679 & n11034 ) | ( n11033 & n11034 ) ;
  assign n11036 = ( n10679 & n11033 ) | ( n10679 & n11034 ) | ( n11033 & n11034 ) ;
  assign n11037 = ( n10679 & n11035 ) | ( n10679 & ~n11036 ) | ( n11035 & ~n11036 ) ;
  assign n11038 = ( x118 & n11032 ) | ( x118 & ~n11037 ) | ( n11032 & ~n11037 ) ;
  assign n11039 = ( x118 & n10680 ) | ( x118 & ~n10715 ) | ( n10680 & ~n10715 ) ;
  assign n11040 = x118 & n10680 ;
  assign n11041 = ( n10685 & n11039 ) | ( n10685 & n11040 ) | ( n11039 & n11040 ) ;
  assign n11042 = ( ~n10685 & n11039 ) | ( ~n10685 & n11040 ) | ( n11039 & n11040 ) ;
  assign n11043 = ( n10685 & ~n11041 ) | ( n10685 & n11042 ) | ( ~n11041 & n11042 ) ;
  assign n11044 = ( x119 & n11038 ) | ( x119 & ~n11043 ) | ( n11038 & ~n11043 ) ;
  assign n11045 = ( x119 & n10686 ) | ( x119 & ~n10715 ) | ( n10686 & ~n10715 ) ;
  assign n11046 = x119 & n10686 ;
  assign n11047 = ( ~n10691 & n11045 ) | ( ~n10691 & n11046 ) | ( n11045 & n11046 ) ;
  assign n11048 = ( n10691 & n11045 ) | ( n10691 & n11046 ) | ( n11045 & n11046 ) ;
  assign n11049 = ( n10691 & n11047 ) | ( n10691 & ~n11048 ) | ( n11047 & ~n11048 ) ;
  assign n11050 = ( x120 & n11044 ) | ( x120 & ~n11049 ) | ( n11044 & ~n11049 ) ;
  assign n11051 = ( x120 & n10692 ) | ( x120 & ~n10715 ) | ( n10692 & ~n10715 ) ;
  assign n11052 = x120 & n10692 ;
  assign n11053 = ( n10697 & n11051 ) | ( n10697 & n11052 ) | ( n11051 & n11052 ) ;
  assign n11054 = ( ~n10697 & n11051 ) | ( ~n10697 & n11052 ) | ( n11051 & n11052 ) ;
  assign n11055 = ( n10697 & ~n11053 ) | ( n10697 & n11054 ) | ( ~n11053 & n11054 ) ;
  assign n11056 = ( x121 & n11050 ) | ( x121 & ~n11055 ) | ( n11050 & ~n11055 ) ;
  assign n11057 = ( x121 & n10698 ) | ( x121 & ~n10715 ) | ( n10698 & ~n10715 ) ;
  assign n11058 = x121 & n10698 ;
  assign n11059 = ( ~n10703 & n11057 ) | ( ~n10703 & n11058 ) | ( n11057 & n11058 ) ;
  assign n11060 = ( n10703 & n11057 ) | ( n10703 & n11058 ) | ( n11057 & n11058 ) ;
  assign n11061 = ( n10703 & n11059 ) | ( n10703 & ~n11060 ) | ( n11059 & ~n11060 ) ;
  assign n11062 = ( x122 & n11056 ) | ( x122 & ~n11061 ) | ( n11056 & ~n11061 ) ;
  assign n11063 = ( x122 & n10704 ) | ( x122 & ~n10715 ) | ( n10704 & ~n10715 ) ;
  assign n11064 = x122 & n10704 ;
  assign n11065 = ( ~n10709 & n11063 ) | ( ~n10709 & n11064 ) | ( n11063 & n11064 ) ;
  assign n11066 = ( n10709 & n11063 ) | ( n10709 & n11064 ) | ( n11063 & n11064 ) ;
  assign n11067 = ( n10709 & n11065 ) | ( n10709 & ~n11066 ) | ( n11065 & ~n11066 ) ;
  assign n11068 = ( x123 & n11062 ) | ( x123 & ~n11067 ) | ( n11062 & ~n11067 ) ;
  assign n11069 = x124 | n11068 ;
  assign n11070 = ( x124 & n133 ) | ( x124 & n11068 ) | ( n133 & n11068 ) ;
  assign n11071 = ( n10713 & ~n11069 ) | ( n10713 & n11070 ) | ( ~n11069 & n11070 ) ;
  assign n11072 = ( x124 & ~n10713 ) | ( x124 & n11068 ) | ( ~n10713 & n11068 ) ;
  assign n11073 = n133 | n11072 ;
  assign n11074 = ( x3 & ~x64 ) | ( x3 & n11073 ) | ( ~x64 & n11073 ) ;
  assign n11075 = ~x3 & n11073 ;
  assign n11076 = ( n10719 & n11074 ) | ( n10719 & ~n11075 ) | ( n11074 & ~n11075 ) ;
  assign n11077 = ~x2 & x64 ;
  assign n11078 = ( x65 & ~n11076 ) | ( x65 & n11077 ) | ( ~n11076 & n11077 ) ;
  assign n11079 = ( x65 & n10719 ) | ( x65 & ~n11073 ) | ( n10719 & ~n11073 ) ;
  assign n11080 = x65 & n10719 ;
  assign n11081 = ( n10718 & n11079 ) | ( n10718 & n11080 ) | ( n11079 & n11080 ) ;
  assign n11082 = ( ~n10718 & n11079 ) | ( ~n10718 & n11080 ) | ( n11079 & n11080 ) ;
  assign n11083 = ( n10718 & ~n11081 ) | ( n10718 & n11082 ) | ( ~n11081 & n11082 ) ;
  assign n11084 = ( x66 & n11078 ) | ( x66 & ~n11083 ) | ( n11078 & ~n11083 ) ;
  assign n11085 = ( x66 & n10720 ) | ( x66 & ~n11073 ) | ( n10720 & ~n11073 ) ;
  assign n11086 = x66 & n10720 ;
  assign n11087 = ( n10725 & n11085 ) | ( n10725 & n11086 ) | ( n11085 & n11086 ) ;
  assign n11088 = ( ~n10725 & n11085 ) | ( ~n10725 & n11086 ) | ( n11085 & n11086 ) ;
  assign n11089 = ( n10725 & ~n11087 ) | ( n10725 & n11088 ) | ( ~n11087 & n11088 ) ;
  assign n11090 = ( x67 & n11084 ) | ( x67 & ~n11089 ) | ( n11084 & ~n11089 ) ;
  assign n11091 = ( x67 & n10726 ) | ( x67 & ~n11073 ) | ( n10726 & ~n11073 ) ;
  assign n11092 = x67 & n10726 ;
  assign n11093 = ( ~n10731 & n11091 ) | ( ~n10731 & n11092 ) | ( n11091 & n11092 ) ;
  assign n11094 = ( n10731 & n11091 ) | ( n10731 & n11092 ) | ( n11091 & n11092 ) ;
  assign n11095 = ( n10731 & n11093 ) | ( n10731 & ~n11094 ) | ( n11093 & ~n11094 ) ;
  assign n11096 = ( x68 & n11090 ) | ( x68 & ~n11095 ) | ( n11090 & ~n11095 ) ;
  assign n11097 = ( x68 & n10732 ) | ( x68 & ~n11073 ) | ( n10732 & ~n11073 ) ;
  assign n11098 = x68 & n10732 ;
  assign n11099 = ( n10737 & n11097 ) | ( n10737 & n11098 ) | ( n11097 & n11098 ) ;
  assign n11100 = ( ~n10737 & n11097 ) | ( ~n10737 & n11098 ) | ( n11097 & n11098 ) ;
  assign n11101 = ( n10737 & ~n11099 ) | ( n10737 & n11100 ) | ( ~n11099 & n11100 ) ;
  assign n11102 = ( x69 & n11096 ) | ( x69 & ~n11101 ) | ( n11096 & ~n11101 ) ;
  assign n11103 = ( x69 & n10738 ) | ( x69 & ~n11073 ) | ( n10738 & ~n11073 ) ;
  assign n11104 = x69 & n10738 ;
  assign n11105 = ( ~n10743 & n11103 ) | ( ~n10743 & n11104 ) | ( n11103 & n11104 ) ;
  assign n11106 = ( n10743 & n11103 ) | ( n10743 & n11104 ) | ( n11103 & n11104 ) ;
  assign n11107 = ( n10743 & n11105 ) | ( n10743 & ~n11106 ) | ( n11105 & ~n11106 ) ;
  assign n11108 = ( x70 & n11102 ) | ( x70 & ~n11107 ) | ( n11102 & ~n11107 ) ;
  assign n11109 = ( x70 & n10744 ) | ( x70 & ~n11073 ) | ( n10744 & ~n11073 ) ;
  assign n11110 = x70 & n10744 ;
  assign n11111 = ( n10749 & n11109 ) | ( n10749 & n11110 ) | ( n11109 & n11110 ) ;
  assign n11112 = ( ~n10749 & n11109 ) | ( ~n10749 & n11110 ) | ( n11109 & n11110 ) ;
  assign n11113 = ( n10749 & ~n11111 ) | ( n10749 & n11112 ) | ( ~n11111 & n11112 ) ;
  assign n11114 = ( x71 & n11108 ) | ( x71 & ~n11113 ) | ( n11108 & ~n11113 ) ;
  assign n11115 = ( x71 & n10750 ) | ( x71 & ~n11073 ) | ( n10750 & ~n11073 ) ;
  assign n11116 = x71 & n10750 ;
  assign n11117 = ( ~n10755 & n11115 ) | ( ~n10755 & n11116 ) | ( n11115 & n11116 ) ;
  assign n11118 = ( n10755 & n11115 ) | ( n10755 & n11116 ) | ( n11115 & n11116 ) ;
  assign n11119 = ( n10755 & n11117 ) | ( n10755 & ~n11118 ) | ( n11117 & ~n11118 ) ;
  assign n11120 = ( x72 & n11114 ) | ( x72 & ~n11119 ) | ( n11114 & ~n11119 ) ;
  assign n11121 = ( x72 & n10756 ) | ( x72 & ~n11073 ) | ( n10756 & ~n11073 ) ;
  assign n11122 = x72 & n10756 ;
  assign n11123 = ( n10761 & n11121 ) | ( n10761 & n11122 ) | ( n11121 & n11122 ) ;
  assign n11124 = ( ~n10761 & n11121 ) | ( ~n10761 & n11122 ) | ( n11121 & n11122 ) ;
  assign n11125 = ( n10761 & ~n11123 ) | ( n10761 & n11124 ) | ( ~n11123 & n11124 ) ;
  assign n11126 = ( x73 & n11120 ) | ( x73 & ~n11125 ) | ( n11120 & ~n11125 ) ;
  assign n11127 = ( x73 & n10762 ) | ( x73 & ~n11073 ) | ( n10762 & ~n11073 ) ;
  assign n11128 = x73 & n10762 ;
  assign n11129 = ( ~n10767 & n11127 ) | ( ~n10767 & n11128 ) | ( n11127 & n11128 ) ;
  assign n11130 = ( n10767 & n11127 ) | ( n10767 & n11128 ) | ( n11127 & n11128 ) ;
  assign n11131 = ( n10767 & n11129 ) | ( n10767 & ~n11130 ) | ( n11129 & ~n11130 ) ;
  assign n11132 = ( x74 & n11126 ) | ( x74 & ~n11131 ) | ( n11126 & ~n11131 ) ;
  assign n11133 = ( x74 & n10768 ) | ( x74 & ~n11073 ) | ( n10768 & ~n11073 ) ;
  assign n11134 = x74 & n10768 ;
  assign n11135 = ( n10773 & n11133 ) | ( n10773 & n11134 ) | ( n11133 & n11134 ) ;
  assign n11136 = ( ~n10773 & n11133 ) | ( ~n10773 & n11134 ) | ( n11133 & n11134 ) ;
  assign n11137 = ( n10773 & ~n11135 ) | ( n10773 & n11136 ) | ( ~n11135 & n11136 ) ;
  assign n11138 = ( x75 & n11132 ) | ( x75 & ~n11137 ) | ( n11132 & ~n11137 ) ;
  assign n11139 = ( x75 & n10774 ) | ( x75 & ~n11073 ) | ( n10774 & ~n11073 ) ;
  assign n11140 = x75 & n10774 ;
  assign n11141 = ( ~n10779 & n11139 ) | ( ~n10779 & n11140 ) | ( n11139 & n11140 ) ;
  assign n11142 = ( n10779 & n11139 ) | ( n10779 & n11140 ) | ( n11139 & n11140 ) ;
  assign n11143 = ( n10779 & n11141 ) | ( n10779 & ~n11142 ) | ( n11141 & ~n11142 ) ;
  assign n11144 = ( x76 & n11138 ) | ( x76 & ~n11143 ) | ( n11138 & ~n11143 ) ;
  assign n11145 = ( x76 & n10780 ) | ( x76 & ~n11073 ) | ( n10780 & ~n11073 ) ;
  assign n11146 = x76 & n10780 ;
  assign n11147 = ( n10785 & n11145 ) | ( n10785 & n11146 ) | ( n11145 & n11146 ) ;
  assign n11148 = ( ~n10785 & n11145 ) | ( ~n10785 & n11146 ) | ( n11145 & n11146 ) ;
  assign n11149 = ( n10785 & ~n11147 ) | ( n10785 & n11148 ) | ( ~n11147 & n11148 ) ;
  assign n11150 = ( x77 & n11144 ) | ( x77 & ~n11149 ) | ( n11144 & ~n11149 ) ;
  assign n11151 = ( x77 & n10786 ) | ( x77 & ~n11073 ) | ( n10786 & ~n11073 ) ;
  assign n11152 = x77 & n10786 ;
  assign n11153 = ( ~n10791 & n11151 ) | ( ~n10791 & n11152 ) | ( n11151 & n11152 ) ;
  assign n11154 = ( n10791 & n11151 ) | ( n10791 & n11152 ) | ( n11151 & n11152 ) ;
  assign n11155 = ( n10791 & n11153 ) | ( n10791 & ~n11154 ) | ( n11153 & ~n11154 ) ;
  assign n11156 = ( x78 & n11150 ) | ( x78 & ~n11155 ) | ( n11150 & ~n11155 ) ;
  assign n11157 = ( x78 & n10792 ) | ( x78 & ~n11073 ) | ( n10792 & ~n11073 ) ;
  assign n11158 = x78 & n10792 ;
  assign n11159 = ( n10797 & n11157 ) | ( n10797 & n11158 ) | ( n11157 & n11158 ) ;
  assign n11160 = ( ~n10797 & n11157 ) | ( ~n10797 & n11158 ) | ( n11157 & n11158 ) ;
  assign n11161 = ( n10797 & ~n11159 ) | ( n10797 & n11160 ) | ( ~n11159 & n11160 ) ;
  assign n11162 = ( x79 & n11156 ) | ( x79 & ~n11161 ) | ( n11156 & ~n11161 ) ;
  assign n11163 = ( x79 & n10798 ) | ( x79 & ~n11073 ) | ( n10798 & ~n11073 ) ;
  assign n11164 = x79 & n10798 ;
  assign n11165 = ( ~n10803 & n11163 ) | ( ~n10803 & n11164 ) | ( n11163 & n11164 ) ;
  assign n11166 = ( n10803 & n11163 ) | ( n10803 & n11164 ) | ( n11163 & n11164 ) ;
  assign n11167 = ( n10803 & n11165 ) | ( n10803 & ~n11166 ) | ( n11165 & ~n11166 ) ;
  assign n11168 = ( x80 & n11162 ) | ( x80 & ~n11167 ) | ( n11162 & ~n11167 ) ;
  assign n11169 = ( x80 & n10804 ) | ( x80 & ~n11073 ) | ( n10804 & ~n11073 ) ;
  assign n11170 = x80 & n10804 ;
  assign n11171 = ( n10809 & n11169 ) | ( n10809 & n11170 ) | ( n11169 & n11170 ) ;
  assign n11172 = ( ~n10809 & n11169 ) | ( ~n10809 & n11170 ) | ( n11169 & n11170 ) ;
  assign n11173 = ( n10809 & ~n11171 ) | ( n10809 & n11172 ) | ( ~n11171 & n11172 ) ;
  assign n11174 = ( x81 & n11168 ) | ( x81 & ~n11173 ) | ( n11168 & ~n11173 ) ;
  assign n11175 = ( x81 & n10810 ) | ( x81 & ~n11073 ) | ( n10810 & ~n11073 ) ;
  assign n11176 = x81 & n10810 ;
  assign n11177 = ( ~n10815 & n11175 ) | ( ~n10815 & n11176 ) | ( n11175 & n11176 ) ;
  assign n11178 = ( n10815 & n11175 ) | ( n10815 & n11176 ) | ( n11175 & n11176 ) ;
  assign n11179 = ( n10815 & n11177 ) | ( n10815 & ~n11178 ) | ( n11177 & ~n11178 ) ;
  assign n11180 = ( x82 & n11174 ) | ( x82 & ~n11179 ) | ( n11174 & ~n11179 ) ;
  assign n11181 = ( x82 & n10816 ) | ( x82 & ~n11073 ) | ( n10816 & ~n11073 ) ;
  assign n11182 = x82 & n10816 ;
  assign n11183 = ( n10821 & n11181 ) | ( n10821 & n11182 ) | ( n11181 & n11182 ) ;
  assign n11184 = ( ~n10821 & n11181 ) | ( ~n10821 & n11182 ) | ( n11181 & n11182 ) ;
  assign n11185 = ( n10821 & ~n11183 ) | ( n10821 & n11184 ) | ( ~n11183 & n11184 ) ;
  assign n11186 = ( x83 & n11180 ) | ( x83 & ~n11185 ) | ( n11180 & ~n11185 ) ;
  assign n11187 = ( x83 & n10822 ) | ( x83 & ~n11073 ) | ( n10822 & ~n11073 ) ;
  assign n11188 = x83 & n10822 ;
  assign n11189 = ( ~n10827 & n11187 ) | ( ~n10827 & n11188 ) | ( n11187 & n11188 ) ;
  assign n11190 = ( n10827 & n11187 ) | ( n10827 & n11188 ) | ( n11187 & n11188 ) ;
  assign n11191 = ( n10827 & n11189 ) | ( n10827 & ~n11190 ) | ( n11189 & ~n11190 ) ;
  assign n11192 = ( x84 & n11186 ) | ( x84 & ~n11191 ) | ( n11186 & ~n11191 ) ;
  assign n11193 = ( x84 & n10828 ) | ( x84 & ~n11073 ) | ( n10828 & ~n11073 ) ;
  assign n11194 = x84 & n10828 ;
  assign n11195 = ( n10833 & n11193 ) | ( n10833 & n11194 ) | ( n11193 & n11194 ) ;
  assign n11196 = ( ~n10833 & n11193 ) | ( ~n10833 & n11194 ) | ( n11193 & n11194 ) ;
  assign n11197 = ( n10833 & ~n11195 ) | ( n10833 & n11196 ) | ( ~n11195 & n11196 ) ;
  assign n11198 = ( x85 & n11192 ) | ( x85 & ~n11197 ) | ( n11192 & ~n11197 ) ;
  assign n11199 = ( x85 & n10834 ) | ( x85 & ~n11073 ) | ( n10834 & ~n11073 ) ;
  assign n11200 = x85 & n10834 ;
  assign n11201 = ( ~n10839 & n11199 ) | ( ~n10839 & n11200 ) | ( n11199 & n11200 ) ;
  assign n11202 = ( n10839 & n11199 ) | ( n10839 & n11200 ) | ( n11199 & n11200 ) ;
  assign n11203 = ( n10839 & n11201 ) | ( n10839 & ~n11202 ) | ( n11201 & ~n11202 ) ;
  assign n11204 = ( x86 & n11198 ) | ( x86 & ~n11203 ) | ( n11198 & ~n11203 ) ;
  assign n11205 = ( x86 & n10840 ) | ( x86 & ~n11073 ) | ( n10840 & ~n11073 ) ;
  assign n11206 = x86 & n10840 ;
  assign n11207 = ( n10845 & n11205 ) | ( n10845 & n11206 ) | ( n11205 & n11206 ) ;
  assign n11208 = ( ~n10845 & n11205 ) | ( ~n10845 & n11206 ) | ( n11205 & n11206 ) ;
  assign n11209 = ( n10845 & ~n11207 ) | ( n10845 & n11208 ) | ( ~n11207 & n11208 ) ;
  assign n11210 = ( x87 & n11204 ) | ( x87 & ~n11209 ) | ( n11204 & ~n11209 ) ;
  assign n11211 = ( x87 & n10846 ) | ( x87 & ~n11073 ) | ( n10846 & ~n11073 ) ;
  assign n11212 = x87 & n10846 ;
  assign n11213 = ( ~n10851 & n11211 ) | ( ~n10851 & n11212 ) | ( n11211 & n11212 ) ;
  assign n11214 = ( n10851 & n11211 ) | ( n10851 & n11212 ) | ( n11211 & n11212 ) ;
  assign n11215 = ( n10851 & n11213 ) | ( n10851 & ~n11214 ) | ( n11213 & ~n11214 ) ;
  assign n11216 = ( x88 & n11210 ) | ( x88 & ~n11215 ) | ( n11210 & ~n11215 ) ;
  assign n11217 = ( x88 & n10852 ) | ( x88 & ~n11073 ) | ( n10852 & ~n11073 ) ;
  assign n11218 = x88 & n10852 ;
  assign n11219 = ( n10857 & n11217 ) | ( n10857 & n11218 ) | ( n11217 & n11218 ) ;
  assign n11220 = ( ~n10857 & n11217 ) | ( ~n10857 & n11218 ) | ( n11217 & n11218 ) ;
  assign n11221 = ( n10857 & ~n11219 ) | ( n10857 & n11220 ) | ( ~n11219 & n11220 ) ;
  assign n11222 = ( x89 & n11216 ) | ( x89 & ~n11221 ) | ( n11216 & ~n11221 ) ;
  assign n11223 = ( x89 & n10858 ) | ( x89 & ~n11073 ) | ( n10858 & ~n11073 ) ;
  assign n11224 = x89 & n10858 ;
  assign n11225 = ( ~n10863 & n11223 ) | ( ~n10863 & n11224 ) | ( n11223 & n11224 ) ;
  assign n11226 = ( n10863 & n11223 ) | ( n10863 & n11224 ) | ( n11223 & n11224 ) ;
  assign n11227 = ( n10863 & n11225 ) | ( n10863 & ~n11226 ) | ( n11225 & ~n11226 ) ;
  assign n11228 = ( x90 & n11222 ) | ( x90 & ~n11227 ) | ( n11222 & ~n11227 ) ;
  assign n11229 = ( x90 & n10864 ) | ( x90 & ~n11073 ) | ( n10864 & ~n11073 ) ;
  assign n11230 = x90 & n10864 ;
  assign n11231 = ( n10869 & n11229 ) | ( n10869 & n11230 ) | ( n11229 & n11230 ) ;
  assign n11232 = ( ~n10869 & n11229 ) | ( ~n10869 & n11230 ) | ( n11229 & n11230 ) ;
  assign n11233 = ( n10869 & ~n11231 ) | ( n10869 & n11232 ) | ( ~n11231 & n11232 ) ;
  assign n11234 = ( x91 & n11228 ) | ( x91 & ~n11233 ) | ( n11228 & ~n11233 ) ;
  assign n11235 = ( x91 & n10870 ) | ( x91 & ~n11073 ) | ( n10870 & ~n11073 ) ;
  assign n11236 = x91 & n10870 ;
  assign n11237 = ( ~n10875 & n11235 ) | ( ~n10875 & n11236 ) | ( n11235 & n11236 ) ;
  assign n11238 = ( n10875 & n11235 ) | ( n10875 & n11236 ) | ( n11235 & n11236 ) ;
  assign n11239 = ( n10875 & n11237 ) | ( n10875 & ~n11238 ) | ( n11237 & ~n11238 ) ;
  assign n11240 = ( x92 & n11234 ) | ( x92 & ~n11239 ) | ( n11234 & ~n11239 ) ;
  assign n11241 = ( x92 & n10876 ) | ( x92 & ~n11073 ) | ( n10876 & ~n11073 ) ;
  assign n11242 = x92 & n10876 ;
  assign n11243 = ( n10881 & n11241 ) | ( n10881 & n11242 ) | ( n11241 & n11242 ) ;
  assign n11244 = ( ~n10881 & n11241 ) | ( ~n10881 & n11242 ) | ( n11241 & n11242 ) ;
  assign n11245 = ( n10881 & ~n11243 ) | ( n10881 & n11244 ) | ( ~n11243 & n11244 ) ;
  assign n11246 = ( x93 & n11240 ) | ( x93 & ~n11245 ) | ( n11240 & ~n11245 ) ;
  assign n11247 = ( x93 & n10882 ) | ( x93 & ~n11073 ) | ( n10882 & ~n11073 ) ;
  assign n11248 = x93 & n10882 ;
  assign n11249 = ( ~n10887 & n11247 ) | ( ~n10887 & n11248 ) | ( n11247 & n11248 ) ;
  assign n11250 = ( n10887 & n11247 ) | ( n10887 & n11248 ) | ( n11247 & n11248 ) ;
  assign n11251 = ( n10887 & n11249 ) | ( n10887 & ~n11250 ) | ( n11249 & ~n11250 ) ;
  assign n11252 = ( x94 & n11246 ) | ( x94 & ~n11251 ) | ( n11246 & ~n11251 ) ;
  assign n11253 = ( x94 & n10888 ) | ( x94 & ~n11073 ) | ( n10888 & ~n11073 ) ;
  assign n11254 = x94 & n10888 ;
  assign n11255 = ( n10893 & n11253 ) | ( n10893 & n11254 ) | ( n11253 & n11254 ) ;
  assign n11256 = ( ~n10893 & n11253 ) | ( ~n10893 & n11254 ) | ( n11253 & n11254 ) ;
  assign n11257 = ( n10893 & ~n11255 ) | ( n10893 & n11256 ) | ( ~n11255 & n11256 ) ;
  assign n11258 = ( x95 & n11252 ) | ( x95 & ~n11257 ) | ( n11252 & ~n11257 ) ;
  assign n11259 = ( x95 & n10894 ) | ( x95 & ~n11073 ) | ( n10894 & ~n11073 ) ;
  assign n11260 = x95 & n10894 ;
  assign n11261 = ( ~n10899 & n11259 ) | ( ~n10899 & n11260 ) | ( n11259 & n11260 ) ;
  assign n11262 = ( n10899 & n11259 ) | ( n10899 & n11260 ) | ( n11259 & n11260 ) ;
  assign n11263 = ( n10899 & n11261 ) | ( n10899 & ~n11262 ) | ( n11261 & ~n11262 ) ;
  assign n11264 = ( x96 & n11258 ) | ( x96 & ~n11263 ) | ( n11258 & ~n11263 ) ;
  assign n11265 = ( x96 & n10900 ) | ( x96 & ~n11073 ) | ( n10900 & ~n11073 ) ;
  assign n11266 = x96 & n10900 ;
  assign n11267 = ( n10905 & n11265 ) | ( n10905 & n11266 ) | ( n11265 & n11266 ) ;
  assign n11268 = ( ~n10905 & n11265 ) | ( ~n10905 & n11266 ) | ( n11265 & n11266 ) ;
  assign n11269 = ( n10905 & ~n11267 ) | ( n10905 & n11268 ) | ( ~n11267 & n11268 ) ;
  assign n11270 = ( x97 & n11264 ) | ( x97 & ~n11269 ) | ( n11264 & ~n11269 ) ;
  assign n11271 = ( x97 & n10906 ) | ( x97 & ~n11073 ) | ( n10906 & ~n11073 ) ;
  assign n11272 = x97 & n10906 ;
  assign n11273 = ( ~n10911 & n11271 ) | ( ~n10911 & n11272 ) | ( n11271 & n11272 ) ;
  assign n11274 = ( n10911 & n11271 ) | ( n10911 & n11272 ) | ( n11271 & n11272 ) ;
  assign n11275 = ( n10911 & n11273 ) | ( n10911 & ~n11274 ) | ( n11273 & ~n11274 ) ;
  assign n11276 = ( x98 & n11270 ) | ( x98 & ~n11275 ) | ( n11270 & ~n11275 ) ;
  assign n11277 = ( x98 & n10912 ) | ( x98 & ~n11073 ) | ( n10912 & ~n11073 ) ;
  assign n11278 = x98 & n10912 ;
  assign n11279 = ( n10917 & n11277 ) | ( n10917 & n11278 ) | ( n11277 & n11278 ) ;
  assign n11280 = ( ~n10917 & n11277 ) | ( ~n10917 & n11278 ) | ( n11277 & n11278 ) ;
  assign n11281 = ( n10917 & ~n11279 ) | ( n10917 & n11280 ) | ( ~n11279 & n11280 ) ;
  assign n11282 = ( x99 & n11276 ) | ( x99 & ~n11281 ) | ( n11276 & ~n11281 ) ;
  assign n11283 = ( x99 & n10918 ) | ( x99 & ~n11073 ) | ( n10918 & ~n11073 ) ;
  assign n11284 = x99 & n10918 ;
  assign n11285 = ( ~n10923 & n11283 ) | ( ~n10923 & n11284 ) | ( n11283 & n11284 ) ;
  assign n11286 = ( n10923 & n11283 ) | ( n10923 & n11284 ) | ( n11283 & n11284 ) ;
  assign n11287 = ( n10923 & n11285 ) | ( n10923 & ~n11286 ) | ( n11285 & ~n11286 ) ;
  assign n11288 = ( x100 & n11282 ) | ( x100 & ~n11287 ) | ( n11282 & ~n11287 ) ;
  assign n11289 = ( x100 & n10924 ) | ( x100 & ~n11073 ) | ( n10924 & ~n11073 ) ;
  assign n11290 = x100 & n10924 ;
  assign n11291 = ( n10929 & n11289 ) | ( n10929 & n11290 ) | ( n11289 & n11290 ) ;
  assign n11292 = ( ~n10929 & n11289 ) | ( ~n10929 & n11290 ) | ( n11289 & n11290 ) ;
  assign n11293 = ( n10929 & ~n11291 ) | ( n10929 & n11292 ) | ( ~n11291 & n11292 ) ;
  assign n11294 = ( x101 & n11288 ) | ( x101 & ~n11293 ) | ( n11288 & ~n11293 ) ;
  assign n11295 = ( x101 & n10930 ) | ( x101 & ~n11073 ) | ( n10930 & ~n11073 ) ;
  assign n11296 = x101 & n10930 ;
  assign n11297 = ( ~n10935 & n11295 ) | ( ~n10935 & n11296 ) | ( n11295 & n11296 ) ;
  assign n11298 = ( n10935 & n11295 ) | ( n10935 & n11296 ) | ( n11295 & n11296 ) ;
  assign n11299 = ( n10935 & n11297 ) | ( n10935 & ~n11298 ) | ( n11297 & ~n11298 ) ;
  assign n11300 = ( x102 & n11294 ) | ( x102 & ~n11299 ) | ( n11294 & ~n11299 ) ;
  assign n11301 = ( x102 & n10936 ) | ( x102 & ~n11073 ) | ( n10936 & ~n11073 ) ;
  assign n11302 = x102 & n10936 ;
  assign n11303 = ( n10941 & n11301 ) | ( n10941 & n11302 ) | ( n11301 & n11302 ) ;
  assign n11304 = ( ~n10941 & n11301 ) | ( ~n10941 & n11302 ) | ( n11301 & n11302 ) ;
  assign n11305 = ( n10941 & ~n11303 ) | ( n10941 & n11304 ) | ( ~n11303 & n11304 ) ;
  assign n11306 = ( x103 & n11300 ) | ( x103 & ~n11305 ) | ( n11300 & ~n11305 ) ;
  assign n11307 = ( x103 & n10942 ) | ( x103 & ~n11073 ) | ( n10942 & ~n11073 ) ;
  assign n11308 = x103 & n10942 ;
  assign n11309 = ( ~n10947 & n11307 ) | ( ~n10947 & n11308 ) | ( n11307 & n11308 ) ;
  assign n11310 = ( n10947 & n11307 ) | ( n10947 & n11308 ) | ( n11307 & n11308 ) ;
  assign n11311 = ( n10947 & n11309 ) | ( n10947 & ~n11310 ) | ( n11309 & ~n11310 ) ;
  assign n11312 = ( x104 & n11306 ) | ( x104 & ~n11311 ) | ( n11306 & ~n11311 ) ;
  assign n11313 = ( x104 & n10948 ) | ( x104 & ~n11073 ) | ( n10948 & ~n11073 ) ;
  assign n11314 = x104 & n10948 ;
  assign n11315 = ( n10953 & n11313 ) | ( n10953 & n11314 ) | ( n11313 & n11314 ) ;
  assign n11316 = ( ~n10953 & n11313 ) | ( ~n10953 & n11314 ) | ( n11313 & n11314 ) ;
  assign n11317 = ( n10953 & ~n11315 ) | ( n10953 & n11316 ) | ( ~n11315 & n11316 ) ;
  assign n11318 = ( x105 & n11312 ) | ( x105 & ~n11317 ) | ( n11312 & ~n11317 ) ;
  assign n11319 = ( x105 & n10954 ) | ( x105 & ~n11073 ) | ( n10954 & ~n11073 ) ;
  assign n11320 = x105 & n10954 ;
  assign n11321 = ( ~n10959 & n11319 ) | ( ~n10959 & n11320 ) | ( n11319 & n11320 ) ;
  assign n11322 = ( n10959 & n11319 ) | ( n10959 & n11320 ) | ( n11319 & n11320 ) ;
  assign n11323 = ( n10959 & n11321 ) | ( n10959 & ~n11322 ) | ( n11321 & ~n11322 ) ;
  assign n11324 = ( x106 & n11318 ) | ( x106 & ~n11323 ) | ( n11318 & ~n11323 ) ;
  assign n11325 = ( x106 & n10960 ) | ( x106 & ~n11073 ) | ( n10960 & ~n11073 ) ;
  assign n11326 = x106 & n10960 ;
  assign n11327 = ( n10965 & n11325 ) | ( n10965 & n11326 ) | ( n11325 & n11326 ) ;
  assign n11328 = ( ~n10965 & n11325 ) | ( ~n10965 & n11326 ) | ( n11325 & n11326 ) ;
  assign n11329 = ( n10965 & ~n11327 ) | ( n10965 & n11328 ) | ( ~n11327 & n11328 ) ;
  assign n11330 = ( x107 & n11324 ) | ( x107 & ~n11329 ) | ( n11324 & ~n11329 ) ;
  assign n11331 = ( x107 & n10966 ) | ( x107 & ~n11073 ) | ( n10966 & ~n11073 ) ;
  assign n11332 = x107 & n10966 ;
  assign n11333 = ( ~n10971 & n11331 ) | ( ~n10971 & n11332 ) | ( n11331 & n11332 ) ;
  assign n11334 = ( n10971 & n11331 ) | ( n10971 & n11332 ) | ( n11331 & n11332 ) ;
  assign n11335 = ( n10971 & n11333 ) | ( n10971 & ~n11334 ) | ( n11333 & ~n11334 ) ;
  assign n11336 = ( x108 & n11330 ) | ( x108 & ~n11335 ) | ( n11330 & ~n11335 ) ;
  assign n11337 = ( x108 & n10972 ) | ( x108 & ~n11073 ) | ( n10972 & ~n11073 ) ;
  assign n11338 = x108 & n10972 ;
  assign n11339 = ( n10977 & n11337 ) | ( n10977 & n11338 ) | ( n11337 & n11338 ) ;
  assign n11340 = ( ~n10977 & n11337 ) | ( ~n10977 & n11338 ) | ( n11337 & n11338 ) ;
  assign n11341 = ( n10977 & ~n11339 ) | ( n10977 & n11340 ) | ( ~n11339 & n11340 ) ;
  assign n11342 = ( x109 & n11336 ) | ( x109 & ~n11341 ) | ( n11336 & ~n11341 ) ;
  assign n11343 = ( x109 & n10978 ) | ( x109 & ~n11073 ) | ( n10978 & ~n11073 ) ;
  assign n11344 = x109 & n10978 ;
  assign n11345 = ( ~n10983 & n11343 ) | ( ~n10983 & n11344 ) | ( n11343 & n11344 ) ;
  assign n11346 = ( n10983 & n11343 ) | ( n10983 & n11344 ) | ( n11343 & n11344 ) ;
  assign n11347 = ( n10983 & n11345 ) | ( n10983 & ~n11346 ) | ( n11345 & ~n11346 ) ;
  assign n11348 = ( x110 & n11342 ) | ( x110 & ~n11347 ) | ( n11342 & ~n11347 ) ;
  assign n11349 = ( x110 & n10984 ) | ( x110 & ~n11073 ) | ( n10984 & ~n11073 ) ;
  assign n11350 = x110 & n10984 ;
  assign n11351 = ( n10989 & n11349 ) | ( n10989 & n11350 ) | ( n11349 & n11350 ) ;
  assign n11352 = ( ~n10989 & n11349 ) | ( ~n10989 & n11350 ) | ( n11349 & n11350 ) ;
  assign n11353 = ( n10989 & ~n11351 ) | ( n10989 & n11352 ) | ( ~n11351 & n11352 ) ;
  assign n11354 = ( x111 & n11348 ) | ( x111 & ~n11353 ) | ( n11348 & ~n11353 ) ;
  assign n11355 = ( x111 & n10990 ) | ( x111 & ~n11073 ) | ( n10990 & ~n11073 ) ;
  assign n11356 = x111 & n10990 ;
  assign n11357 = ( ~n10995 & n11355 ) | ( ~n10995 & n11356 ) | ( n11355 & n11356 ) ;
  assign n11358 = ( n10995 & n11355 ) | ( n10995 & n11356 ) | ( n11355 & n11356 ) ;
  assign n11359 = ( n10995 & n11357 ) | ( n10995 & ~n11358 ) | ( n11357 & ~n11358 ) ;
  assign n11360 = ( x112 & n11354 ) | ( x112 & ~n11359 ) | ( n11354 & ~n11359 ) ;
  assign n11361 = ( x112 & n10996 ) | ( x112 & ~n11073 ) | ( n10996 & ~n11073 ) ;
  assign n11362 = x112 & n10996 ;
  assign n11363 = ( n11001 & n11361 ) | ( n11001 & n11362 ) | ( n11361 & n11362 ) ;
  assign n11364 = ( ~n11001 & n11361 ) | ( ~n11001 & n11362 ) | ( n11361 & n11362 ) ;
  assign n11365 = ( n11001 & ~n11363 ) | ( n11001 & n11364 ) | ( ~n11363 & n11364 ) ;
  assign n11366 = ( x113 & n11360 ) | ( x113 & ~n11365 ) | ( n11360 & ~n11365 ) ;
  assign n11367 = ( x113 & n11002 ) | ( x113 & ~n11073 ) | ( n11002 & ~n11073 ) ;
  assign n11368 = x113 & n11002 ;
  assign n11369 = ( ~n11007 & n11367 ) | ( ~n11007 & n11368 ) | ( n11367 & n11368 ) ;
  assign n11370 = ( n11007 & n11367 ) | ( n11007 & n11368 ) | ( n11367 & n11368 ) ;
  assign n11371 = ( n11007 & n11369 ) | ( n11007 & ~n11370 ) | ( n11369 & ~n11370 ) ;
  assign n11372 = ( x114 & n11366 ) | ( x114 & ~n11371 ) | ( n11366 & ~n11371 ) ;
  assign n11373 = ( x114 & n11008 ) | ( x114 & ~n11073 ) | ( n11008 & ~n11073 ) ;
  assign n11374 = x114 & n11008 ;
  assign n11375 = ( n11013 & n11373 ) | ( n11013 & n11374 ) | ( n11373 & n11374 ) ;
  assign n11376 = ( ~n11013 & n11373 ) | ( ~n11013 & n11374 ) | ( n11373 & n11374 ) ;
  assign n11377 = ( n11013 & ~n11375 ) | ( n11013 & n11376 ) | ( ~n11375 & n11376 ) ;
  assign n11378 = ( x115 & n11372 ) | ( x115 & ~n11377 ) | ( n11372 & ~n11377 ) ;
  assign n11379 = ( x115 & n11014 ) | ( x115 & ~n11073 ) | ( n11014 & ~n11073 ) ;
  assign n11380 = x115 & n11014 ;
  assign n11381 = ( ~n11019 & n11379 ) | ( ~n11019 & n11380 ) | ( n11379 & n11380 ) ;
  assign n11382 = ( n11019 & n11379 ) | ( n11019 & n11380 ) | ( n11379 & n11380 ) ;
  assign n11383 = ( n11019 & n11381 ) | ( n11019 & ~n11382 ) | ( n11381 & ~n11382 ) ;
  assign n11384 = ( x116 & n11378 ) | ( x116 & ~n11383 ) | ( n11378 & ~n11383 ) ;
  assign n11385 = ( x116 & n11020 ) | ( x116 & ~n11073 ) | ( n11020 & ~n11073 ) ;
  assign n11386 = x116 & n11020 ;
  assign n11387 = ( n11025 & n11385 ) | ( n11025 & n11386 ) | ( n11385 & n11386 ) ;
  assign n11388 = ( ~n11025 & n11385 ) | ( ~n11025 & n11386 ) | ( n11385 & n11386 ) ;
  assign n11389 = ( n11025 & ~n11387 ) | ( n11025 & n11388 ) | ( ~n11387 & n11388 ) ;
  assign n11390 = ( x117 & n11384 ) | ( x117 & ~n11389 ) | ( n11384 & ~n11389 ) ;
  assign n11391 = ( x117 & n11026 ) | ( x117 & ~n11073 ) | ( n11026 & ~n11073 ) ;
  assign n11392 = x117 & n11026 ;
  assign n11393 = ( ~n11031 & n11391 ) | ( ~n11031 & n11392 ) | ( n11391 & n11392 ) ;
  assign n11394 = ( n11031 & n11391 ) | ( n11031 & n11392 ) | ( n11391 & n11392 ) ;
  assign n11395 = ( n11031 & n11393 ) | ( n11031 & ~n11394 ) | ( n11393 & ~n11394 ) ;
  assign n11396 = ( x118 & n11390 ) | ( x118 & ~n11395 ) | ( n11390 & ~n11395 ) ;
  assign n11397 = ( x118 & n11032 ) | ( x118 & ~n11073 ) | ( n11032 & ~n11073 ) ;
  assign n11398 = x118 & n11032 ;
  assign n11399 = ( n11037 & n11397 ) | ( n11037 & n11398 ) | ( n11397 & n11398 ) ;
  assign n11400 = ( ~n11037 & n11397 ) | ( ~n11037 & n11398 ) | ( n11397 & n11398 ) ;
  assign n11401 = ( n11037 & ~n11399 ) | ( n11037 & n11400 ) | ( ~n11399 & n11400 ) ;
  assign n11402 = ( x119 & n11396 ) | ( x119 & ~n11401 ) | ( n11396 & ~n11401 ) ;
  assign n11403 = ( x119 & n11038 ) | ( x119 & ~n11073 ) | ( n11038 & ~n11073 ) ;
  assign n11404 = x119 & n11038 ;
  assign n11405 = ( ~n11043 & n11403 ) | ( ~n11043 & n11404 ) | ( n11403 & n11404 ) ;
  assign n11406 = ( n11043 & n11403 ) | ( n11043 & n11404 ) | ( n11403 & n11404 ) ;
  assign n11407 = ( n11043 & n11405 ) | ( n11043 & ~n11406 ) | ( n11405 & ~n11406 ) ;
  assign n11408 = ( x120 & n11402 ) | ( x120 & ~n11407 ) | ( n11402 & ~n11407 ) ;
  assign n11409 = ( x120 & n11044 ) | ( x120 & ~n11073 ) | ( n11044 & ~n11073 ) ;
  assign n11410 = x120 & n11044 ;
  assign n11411 = ( n11049 & n11409 ) | ( n11049 & n11410 ) | ( n11409 & n11410 ) ;
  assign n11412 = ( ~n11049 & n11409 ) | ( ~n11049 & n11410 ) | ( n11409 & n11410 ) ;
  assign n11413 = ( n11049 & ~n11411 ) | ( n11049 & n11412 ) | ( ~n11411 & n11412 ) ;
  assign n11414 = ( x121 & n11408 ) | ( x121 & ~n11413 ) | ( n11408 & ~n11413 ) ;
  assign n11415 = ( x121 & n11050 ) | ( x121 & ~n11073 ) | ( n11050 & ~n11073 ) ;
  assign n11416 = x121 & n11050 ;
  assign n11417 = ( ~n11055 & n11415 ) | ( ~n11055 & n11416 ) | ( n11415 & n11416 ) ;
  assign n11418 = ( n11055 & n11415 ) | ( n11055 & n11416 ) | ( n11415 & n11416 ) ;
  assign n11419 = ( n11055 & n11417 ) | ( n11055 & ~n11418 ) | ( n11417 & ~n11418 ) ;
  assign n11420 = ( x122 & n11414 ) | ( x122 & ~n11419 ) | ( n11414 & ~n11419 ) ;
  assign n11421 = ( x122 & n11056 ) | ( x122 & ~n11073 ) | ( n11056 & ~n11073 ) ;
  assign n11422 = x122 & n11056 ;
  assign n11423 = ( n11061 & n11421 ) | ( n11061 & n11422 ) | ( n11421 & n11422 ) ;
  assign n11424 = ( ~n11061 & n11421 ) | ( ~n11061 & n11422 ) | ( n11421 & n11422 ) ;
  assign n11425 = ( n11061 & ~n11423 ) | ( n11061 & n11424 ) | ( ~n11423 & n11424 ) ;
  assign n11426 = ( x123 & n11420 ) | ( x123 & ~n11425 ) | ( n11420 & ~n11425 ) ;
  assign n11427 = ( x123 & n11062 ) | ( x123 & ~n11073 ) | ( n11062 & ~n11073 ) ;
  assign n11428 = x123 & n11062 ;
  assign n11429 = ( n11067 & n11427 ) | ( n11067 & n11428 ) | ( n11427 & n11428 ) ;
  assign n11430 = ( ~n11067 & n11427 ) | ( ~n11067 & n11428 ) | ( n11427 & n11428 ) ;
  assign n11431 = ( n11067 & ~n11429 ) | ( n11067 & n11430 ) | ( ~n11429 & n11430 ) ;
  assign n11432 = ( x124 & n11426 ) | ( x124 & ~n11431 ) | ( n11426 & ~n11431 ) ;
  assign n11433 = x125 | n11432 ;
  assign n11434 = ( x125 & n132 ) | ( x125 & n11432 ) | ( n132 & n11432 ) ;
  assign n11435 = ( n11071 & ~n11433 ) | ( n11071 & n11434 ) | ( ~n11433 & n11434 ) ;
  assign n11436 = ( x125 & ~n11071 ) | ( x125 & n11432 ) | ( ~n11071 & n11432 ) ;
  assign n11437 = n132 | n11436 ;
  assign n11438 = ( x2 & ~x64 ) | ( x2 & n11437 ) | ( ~x64 & n11437 ) ;
  assign n11439 = ~x2 & n11437 ;
  assign n11440 = ( n11077 & n11438 ) | ( n11077 & ~n11439 ) | ( n11438 & ~n11439 ) ;
  assign n11441 = ( x65 & n129 ) | ( x65 & ~n11440 ) | ( n129 & ~n11440 ) ;
  assign n11442 = ( x65 & n11077 ) | ( x65 & ~n11437 ) | ( n11077 & ~n11437 ) ;
  assign n11443 = x65 & n11077 ;
  assign n11444 = ( n11076 & n11442 ) | ( n11076 & n11443 ) | ( n11442 & n11443 ) ;
  assign n11445 = ( ~n11076 & n11442 ) | ( ~n11076 & n11443 ) | ( n11442 & n11443 ) ;
  assign n11446 = ( n11076 & ~n11444 ) | ( n11076 & n11445 ) | ( ~n11444 & n11445 ) ;
  assign n11447 = ( x66 & n11441 ) | ( x66 & ~n11446 ) | ( n11441 & ~n11446 ) ;
  assign n11448 = ( x66 & n11078 ) | ( x66 & ~n11437 ) | ( n11078 & ~n11437 ) ;
  assign n11449 = x66 & n11078 ;
  assign n11450 = ( n11083 & n11448 ) | ( n11083 & n11449 ) | ( n11448 & n11449 ) ;
  assign n11451 = ( ~n11083 & n11448 ) | ( ~n11083 & n11449 ) | ( n11448 & n11449 ) ;
  assign n11452 = ( n11083 & ~n11450 ) | ( n11083 & n11451 ) | ( ~n11450 & n11451 ) ;
  assign n11453 = ( x67 & n11447 ) | ( x67 & ~n11452 ) | ( n11447 & ~n11452 ) ;
  assign n11454 = ( x67 & n11084 ) | ( x67 & ~n11437 ) | ( n11084 & ~n11437 ) ;
  assign n11455 = x67 & n11084 ;
  assign n11456 = ( ~n11089 & n11454 ) | ( ~n11089 & n11455 ) | ( n11454 & n11455 ) ;
  assign n11457 = ( n11089 & n11454 ) | ( n11089 & n11455 ) | ( n11454 & n11455 ) ;
  assign n11458 = ( n11089 & n11456 ) | ( n11089 & ~n11457 ) | ( n11456 & ~n11457 ) ;
  assign n11459 = ( x68 & n11453 ) | ( x68 & ~n11458 ) | ( n11453 & ~n11458 ) ;
  assign n11460 = ( x68 & n11090 ) | ( x68 & ~n11437 ) | ( n11090 & ~n11437 ) ;
  assign n11461 = x68 & n11090 ;
  assign n11462 = ( n11095 & n11460 ) | ( n11095 & n11461 ) | ( n11460 & n11461 ) ;
  assign n11463 = ( ~n11095 & n11460 ) | ( ~n11095 & n11461 ) | ( n11460 & n11461 ) ;
  assign n11464 = ( n11095 & ~n11462 ) | ( n11095 & n11463 ) | ( ~n11462 & n11463 ) ;
  assign n11465 = ( x69 & n11459 ) | ( x69 & ~n11464 ) | ( n11459 & ~n11464 ) ;
  assign n11466 = ( x69 & n11096 ) | ( x69 & ~n11437 ) | ( n11096 & ~n11437 ) ;
  assign n11467 = x69 & n11096 ;
  assign n11468 = ( ~n11101 & n11466 ) | ( ~n11101 & n11467 ) | ( n11466 & n11467 ) ;
  assign n11469 = ( n11101 & n11466 ) | ( n11101 & n11467 ) | ( n11466 & n11467 ) ;
  assign n11470 = ( n11101 & n11468 ) | ( n11101 & ~n11469 ) | ( n11468 & ~n11469 ) ;
  assign n11471 = ( x70 & n11465 ) | ( x70 & ~n11470 ) | ( n11465 & ~n11470 ) ;
  assign n11472 = ( x70 & n11102 ) | ( x70 & ~n11437 ) | ( n11102 & ~n11437 ) ;
  assign n11473 = x70 & n11102 ;
  assign n11474 = ( n11107 & n11472 ) | ( n11107 & n11473 ) | ( n11472 & n11473 ) ;
  assign n11475 = ( ~n11107 & n11472 ) | ( ~n11107 & n11473 ) | ( n11472 & n11473 ) ;
  assign n11476 = ( n11107 & ~n11474 ) | ( n11107 & n11475 ) | ( ~n11474 & n11475 ) ;
  assign n11477 = ( x71 & n11471 ) | ( x71 & ~n11476 ) | ( n11471 & ~n11476 ) ;
  assign n11478 = ( x71 & n11108 ) | ( x71 & ~n11437 ) | ( n11108 & ~n11437 ) ;
  assign n11479 = x71 & n11108 ;
  assign n11480 = ( ~n11113 & n11478 ) | ( ~n11113 & n11479 ) | ( n11478 & n11479 ) ;
  assign n11481 = ( n11113 & n11478 ) | ( n11113 & n11479 ) | ( n11478 & n11479 ) ;
  assign n11482 = ( n11113 & n11480 ) | ( n11113 & ~n11481 ) | ( n11480 & ~n11481 ) ;
  assign n11483 = ( x72 & n11477 ) | ( x72 & ~n11482 ) | ( n11477 & ~n11482 ) ;
  assign n11484 = ( x72 & n11114 ) | ( x72 & ~n11437 ) | ( n11114 & ~n11437 ) ;
  assign n11485 = x72 & n11114 ;
  assign n11486 = ( n11119 & n11484 ) | ( n11119 & n11485 ) | ( n11484 & n11485 ) ;
  assign n11487 = ( ~n11119 & n11484 ) | ( ~n11119 & n11485 ) | ( n11484 & n11485 ) ;
  assign n11488 = ( n11119 & ~n11486 ) | ( n11119 & n11487 ) | ( ~n11486 & n11487 ) ;
  assign n11489 = ( x73 & n11483 ) | ( x73 & ~n11488 ) | ( n11483 & ~n11488 ) ;
  assign n11490 = ( x73 & n11120 ) | ( x73 & ~n11437 ) | ( n11120 & ~n11437 ) ;
  assign n11491 = x73 & n11120 ;
  assign n11492 = ( ~n11125 & n11490 ) | ( ~n11125 & n11491 ) | ( n11490 & n11491 ) ;
  assign n11493 = ( n11125 & n11490 ) | ( n11125 & n11491 ) | ( n11490 & n11491 ) ;
  assign n11494 = ( n11125 & n11492 ) | ( n11125 & ~n11493 ) | ( n11492 & ~n11493 ) ;
  assign n11495 = ( x74 & n11489 ) | ( x74 & ~n11494 ) | ( n11489 & ~n11494 ) ;
  assign n11496 = ( x74 & n11126 ) | ( x74 & ~n11437 ) | ( n11126 & ~n11437 ) ;
  assign n11497 = x74 & n11126 ;
  assign n11498 = ( n11131 & n11496 ) | ( n11131 & n11497 ) | ( n11496 & n11497 ) ;
  assign n11499 = ( ~n11131 & n11496 ) | ( ~n11131 & n11497 ) | ( n11496 & n11497 ) ;
  assign n11500 = ( n11131 & ~n11498 ) | ( n11131 & n11499 ) | ( ~n11498 & n11499 ) ;
  assign n11501 = ( x75 & n11495 ) | ( x75 & ~n11500 ) | ( n11495 & ~n11500 ) ;
  assign n11502 = ( x75 & n11132 ) | ( x75 & ~n11437 ) | ( n11132 & ~n11437 ) ;
  assign n11503 = x75 & n11132 ;
  assign n11504 = ( ~n11137 & n11502 ) | ( ~n11137 & n11503 ) | ( n11502 & n11503 ) ;
  assign n11505 = ( n11137 & n11502 ) | ( n11137 & n11503 ) | ( n11502 & n11503 ) ;
  assign n11506 = ( n11137 & n11504 ) | ( n11137 & ~n11505 ) | ( n11504 & ~n11505 ) ;
  assign n11507 = ( x76 & n11501 ) | ( x76 & ~n11506 ) | ( n11501 & ~n11506 ) ;
  assign n11508 = ( x76 & n11138 ) | ( x76 & ~n11437 ) | ( n11138 & ~n11437 ) ;
  assign n11509 = x76 & n11138 ;
  assign n11510 = ( n11143 & n11508 ) | ( n11143 & n11509 ) | ( n11508 & n11509 ) ;
  assign n11511 = ( ~n11143 & n11508 ) | ( ~n11143 & n11509 ) | ( n11508 & n11509 ) ;
  assign n11512 = ( n11143 & ~n11510 ) | ( n11143 & n11511 ) | ( ~n11510 & n11511 ) ;
  assign n11513 = ( x77 & n11507 ) | ( x77 & ~n11512 ) | ( n11507 & ~n11512 ) ;
  assign n11514 = ( x77 & n11144 ) | ( x77 & ~n11437 ) | ( n11144 & ~n11437 ) ;
  assign n11515 = x77 & n11144 ;
  assign n11516 = ( ~n11149 & n11514 ) | ( ~n11149 & n11515 ) | ( n11514 & n11515 ) ;
  assign n11517 = ( n11149 & n11514 ) | ( n11149 & n11515 ) | ( n11514 & n11515 ) ;
  assign n11518 = ( n11149 & n11516 ) | ( n11149 & ~n11517 ) | ( n11516 & ~n11517 ) ;
  assign n11519 = ( x78 & n11513 ) | ( x78 & ~n11518 ) | ( n11513 & ~n11518 ) ;
  assign n11520 = ( x78 & n11150 ) | ( x78 & ~n11437 ) | ( n11150 & ~n11437 ) ;
  assign n11521 = x78 & n11150 ;
  assign n11522 = ( n11155 & n11520 ) | ( n11155 & n11521 ) | ( n11520 & n11521 ) ;
  assign n11523 = ( ~n11155 & n11520 ) | ( ~n11155 & n11521 ) | ( n11520 & n11521 ) ;
  assign n11524 = ( n11155 & ~n11522 ) | ( n11155 & n11523 ) | ( ~n11522 & n11523 ) ;
  assign n11525 = ( x79 & n11519 ) | ( x79 & ~n11524 ) | ( n11519 & ~n11524 ) ;
  assign n11526 = ( x79 & n11156 ) | ( x79 & ~n11437 ) | ( n11156 & ~n11437 ) ;
  assign n11527 = x79 & n11156 ;
  assign n11528 = ( ~n11161 & n11526 ) | ( ~n11161 & n11527 ) | ( n11526 & n11527 ) ;
  assign n11529 = ( n11161 & n11526 ) | ( n11161 & n11527 ) | ( n11526 & n11527 ) ;
  assign n11530 = ( n11161 & n11528 ) | ( n11161 & ~n11529 ) | ( n11528 & ~n11529 ) ;
  assign n11531 = ( x80 & n11525 ) | ( x80 & ~n11530 ) | ( n11525 & ~n11530 ) ;
  assign n11532 = ( x80 & n11162 ) | ( x80 & ~n11437 ) | ( n11162 & ~n11437 ) ;
  assign n11533 = x80 & n11162 ;
  assign n11534 = ( n11167 & n11532 ) | ( n11167 & n11533 ) | ( n11532 & n11533 ) ;
  assign n11535 = ( ~n11167 & n11532 ) | ( ~n11167 & n11533 ) | ( n11532 & n11533 ) ;
  assign n11536 = ( n11167 & ~n11534 ) | ( n11167 & n11535 ) | ( ~n11534 & n11535 ) ;
  assign n11537 = ( x81 & n11531 ) | ( x81 & ~n11536 ) | ( n11531 & ~n11536 ) ;
  assign n11538 = ( x81 & n11168 ) | ( x81 & ~n11437 ) | ( n11168 & ~n11437 ) ;
  assign n11539 = x81 & n11168 ;
  assign n11540 = ( ~n11173 & n11538 ) | ( ~n11173 & n11539 ) | ( n11538 & n11539 ) ;
  assign n11541 = ( n11173 & n11538 ) | ( n11173 & n11539 ) | ( n11538 & n11539 ) ;
  assign n11542 = ( n11173 & n11540 ) | ( n11173 & ~n11541 ) | ( n11540 & ~n11541 ) ;
  assign n11543 = ( x82 & n11537 ) | ( x82 & ~n11542 ) | ( n11537 & ~n11542 ) ;
  assign n11544 = ( x82 & n11174 ) | ( x82 & ~n11437 ) | ( n11174 & ~n11437 ) ;
  assign n11545 = x82 & n11174 ;
  assign n11546 = ( n11179 & n11544 ) | ( n11179 & n11545 ) | ( n11544 & n11545 ) ;
  assign n11547 = ( ~n11179 & n11544 ) | ( ~n11179 & n11545 ) | ( n11544 & n11545 ) ;
  assign n11548 = ( n11179 & ~n11546 ) | ( n11179 & n11547 ) | ( ~n11546 & n11547 ) ;
  assign n11549 = ( x83 & n11543 ) | ( x83 & ~n11548 ) | ( n11543 & ~n11548 ) ;
  assign n11550 = ( x83 & n11180 ) | ( x83 & ~n11437 ) | ( n11180 & ~n11437 ) ;
  assign n11551 = x83 & n11180 ;
  assign n11552 = ( ~n11185 & n11550 ) | ( ~n11185 & n11551 ) | ( n11550 & n11551 ) ;
  assign n11553 = ( n11185 & n11550 ) | ( n11185 & n11551 ) | ( n11550 & n11551 ) ;
  assign n11554 = ( n11185 & n11552 ) | ( n11185 & ~n11553 ) | ( n11552 & ~n11553 ) ;
  assign n11555 = ( x84 & n11549 ) | ( x84 & ~n11554 ) | ( n11549 & ~n11554 ) ;
  assign n11556 = ( x84 & n11186 ) | ( x84 & ~n11437 ) | ( n11186 & ~n11437 ) ;
  assign n11557 = x84 & n11186 ;
  assign n11558 = ( n11191 & n11556 ) | ( n11191 & n11557 ) | ( n11556 & n11557 ) ;
  assign n11559 = ( ~n11191 & n11556 ) | ( ~n11191 & n11557 ) | ( n11556 & n11557 ) ;
  assign n11560 = ( n11191 & ~n11558 ) | ( n11191 & n11559 ) | ( ~n11558 & n11559 ) ;
  assign n11561 = ( x85 & n11555 ) | ( x85 & ~n11560 ) | ( n11555 & ~n11560 ) ;
  assign n11562 = ( x85 & n11192 ) | ( x85 & ~n11437 ) | ( n11192 & ~n11437 ) ;
  assign n11563 = x85 & n11192 ;
  assign n11564 = ( ~n11197 & n11562 ) | ( ~n11197 & n11563 ) | ( n11562 & n11563 ) ;
  assign n11565 = ( n11197 & n11562 ) | ( n11197 & n11563 ) | ( n11562 & n11563 ) ;
  assign n11566 = ( n11197 & n11564 ) | ( n11197 & ~n11565 ) | ( n11564 & ~n11565 ) ;
  assign n11567 = ( x86 & n11561 ) | ( x86 & ~n11566 ) | ( n11561 & ~n11566 ) ;
  assign n11568 = ( x86 & n11198 ) | ( x86 & ~n11437 ) | ( n11198 & ~n11437 ) ;
  assign n11569 = x86 & n11198 ;
  assign n11570 = ( n11203 & n11568 ) | ( n11203 & n11569 ) | ( n11568 & n11569 ) ;
  assign n11571 = ( ~n11203 & n11568 ) | ( ~n11203 & n11569 ) | ( n11568 & n11569 ) ;
  assign n11572 = ( n11203 & ~n11570 ) | ( n11203 & n11571 ) | ( ~n11570 & n11571 ) ;
  assign n11573 = ( x87 & n11567 ) | ( x87 & ~n11572 ) | ( n11567 & ~n11572 ) ;
  assign n11574 = ( x87 & n11204 ) | ( x87 & ~n11437 ) | ( n11204 & ~n11437 ) ;
  assign n11575 = x87 & n11204 ;
  assign n11576 = ( ~n11209 & n11574 ) | ( ~n11209 & n11575 ) | ( n11574 & n11575 ) ;
  assign n11577 = ( n11209 & n11574 ) | ( n11209 & n11575 ) | ( n11574 & n11575 ) ;
  assign n11578 = ( n11209 & n11576 ) | ( n11209 & ~n11577 ) | ( n11576 & ~n11577 ) ;
  assign n11579 = ( x88 & n11573 ) | ( x88 & ~n11578 ) | ( n11573 & ~n11578 ) ;
  assign n11580 = ( x88 & n11210 ) | ( x88 & ~n11437 ) | ( n11210 & ~n11437 ) ;
  assign n11581 = x88 & n11210 ;
  assign n11582 = ( n11215 & n11580 ) | ( n11215 & n11581 ) | ( n11580 & n11581 ) ;
  assign n11583 = ( ~n11215 & n11580 ) | ( ~n11215 & n11581 ) | ( n11580 & n11581 ) ;
  assign n11584 = ( n11215 & ~n11582 ) | ( n11215 & n11583 ) | ( ~n11582 & n11583 ) ;
  assign n11585 = ( x89 & n11579 ) | ( x89 & ~n11584 ) | ( n11579 & ~n11584 ) ;
  assign n11586 = ( x89 & n11216 ) | ( x89 & ~n11437 ) | ( n11216 & ~n11437 ) ;
  assign n11587 = x89 & n11216 ;
  assign n11588 = ( ~n11221 & n11586 ) | ( ~n11221 & n11587 ) | ( n11586 & n11587 ) ;
  assign n11589 = ( n11221 & n11586 ) | ( n11221 & n11587 ) | ( n11586 & n11587 ) ;
  assign n11590 = ( n11221 & n11588 ) | ( n11221 & ~n11589 ) | ( n11588 & ~n11589 ) ;
  assign n11591 = ( x90 & n11585 ) | ( x90 & ~n11590 ) | ( n11585 & ~n11590 ) ;
  assign n11592 = ( x90 & n11222 ) | ( x90 & ~n11437 ) | ( n11222 & ~n11437 ) ;
  assign n11593 = x90 & n11222 ;
  assign n11594 = ( n11227 & n11592 ) | ( n11227 & n11593 ) | ( n11592 & n11593 ) ;
  assign n11595 = ( ~n11227 & n11592 ) | ( ~n11227 & n11593 ) | ( n11592 & n11593 ) ;
  assign n11596 = ( n11227 & ~n11594 ) | ( n11227 & n11595 ) | ( ~n11594 & n11595 ) ;
  assign n11597 = ( x91 & n11591 ) | ( x91 & ~n11596 ) | ( n11591 & ~n11596 ) ;
  assign n11598 = ( x91 & n11228 ) | ( x91 & ~n11437 ) | ( n11228 & ~n11437 ) ;
  assign n11599 = x91 & n11228 ;
  assign n11600 = ( ~n11233 & n11598 ) | ( ~n11233 & n11599 ) | ( n11598 & n11599 ) ;
  assign n11601 = ( n11233 & n11598 ) | ( n11233 & n11599 ) | ( n11598 & n11599 ) ;
  assign n11602 = ( n11233 & n11600 ) | ( n11233 & ~n11601 ) | ( n11600 & ~n11601 ) ;
  assign n11603 = ( x92 & n11597 ) | ( x92 & ~n11602 ) | ( n11597 & ~n11602 ) ;
  assign n11604 = ( x92 & n11234 ) | ( x92 & ~n11437 ) | ( n11234 & ~n11437 ) ;
  assign n11605 = x92 & n11234 ;
  assign n11606 = ( n11239 & n11604 ) | ( n11239 & n11605 ) | ( n11604 & n11605 ) ;
  assign n11607 = ( ~n11239 & n11604 ) | ( ~n11239 & n11605 ) | ( n11604 & n11605 ) ;
  assign n11608 = ( n11239 & ~n11606 ) | ( n11239 & n11607 ) | ( ~n11606 & n11607 ) ;
  assign n11609 = ( x93 & n11603 ) | ( x93 & ~n11608 ) | ( n11603 & ~n11608 ) ;
  assign n11610 = ( x93 & n11240 ) | ( x93 & ~n11437 ) | ( n11240 & ~n11437 ) ;
  assign n11611 = x93 & n11240 ;
  assign n11612 = ( ~n11245 & n11610 ) | ( ~n11245 & n11611 ) | ( n11610 & n11611 ) ;
  assign n11613 = ( n11245 & n11610 ) | ( n11245 & n11611 ) | ( n11610 & n11611 ) ;
  assign n11614 = ( n11245 & n11612 ) | ( n11245 & ~n11613 ) | ( n11612 & ~n11613 ) ;
  assign n11615 = ( x94 & n11609 ) | ( x94 & ~n11614 ) | ( n11609 & ~n11614 ) ;
  assign n11616 = ( x94 & n11246 ) | ( x94 & ~n11437 ) | ( n11246 & ~n11437 ) ;
  assign n11617 = x94 & n11246 ;
  assign n11618 = ( n11251 & n11616 ) | ( n11251 & n11617 ) | ( n11616 & n11617 ) ;
  assign n11619 = ( ~n11251 & n11616 ) | ( ~n11251 & n11617 ) | ( n11616 & n11617 ) ;
  assign n11620 = ( n11251 & ~n11618 ) | ( n11251 & n11619 ) | ( ~n11618 & n11619 ) ;
  assign n11621 = ( x95 & n11615 ) | ( x95 & ~n11620 ) | ( n11615 & ~n11620 ) ;
  assign n11622 = ( x95 & n11252 ) | ( x95 & ~n11437 ) | ( n11252 & ~n11437 ) ;
  assign n11623 = x95 & n11252 ;
  assign n11624 = ( ~n11257 & n11622 ) | ( ~n11257 & n11623 ) | ( n11622 & n11623 ) ;
  assign n11625 = ( n11257 & n11622 ) | ( n11257 & n11623 ) | ( n11622 & n11623 ) ;
  assign n11626 = ( n11257 & n11624 ) | ( n11257 & ~n11625 ) | ( n11624 & ~n11625 ) ;
  assign n11627 = ( x96 & n11621 ) | ( x96 & ~n11626 ) | ( n11621 & ~n11626 ) ;
  assign n11628 = ( x96 & n11258 ) | ( x96 & ~n11437 ) | ( n11258 & ~n11437 ) ;
  assign n11629 = x96 & n11258 ;
  assign n11630 = ( n11263 & n11628 ) | ( n11263 & n11629 ) | ( n11628 & n11629 ) ;
  assign n11631 = ( ~n11263 & n11628 ) | ( ~n11263 & n11629 ) | ( n11628 & n11629 ) ;
  assign n11632 = ( n11263 & ~n11630 ) | ( n11263 & n11631 ) | ( ~n11630 & n11631 ) ;
  assign n11633 = ( x97 & n11627 ) | ( x97 & ~n11632 ) | ( n11627 & ~n11632 ) ;
  assign n11634 = ( x97 & n11264 ) | ( x97 & ~n11437 ) | ( n11264 & ~n11437 ) ;
  assign n11635 = x97 & n11264 ;
  assign n11636 = ( ~n11269 & n11634 ) | ( ~n11269 & n11635 ) | ( n11634 & n11635 ) ;
  assign n11637 = ( n11269 & n11634 ) | ( n11269 & n11635 ) | ( n11634 & n11635 ) ;
  assign n11638 = ( n11269 & n11636 ) | ( n11269 & ~n11637 ) | ( n11636 & ~n11637 ) ;
  assign n11639 = ( x98 & n11633 ) | ( x98 & ~n11638 ) | ( n11633 & ~n11638 ) ;
  assign n11640 = ( x98 & n11270 ) | ( x98 & ~n11437 ) | ( n11270 & ~n11437 ) ;
  assign n11641 = x98 & n11270 ;
  assign n11642 = ( n11275 & n11640 ) | ( n11275 & n11641 ) | ( n11640 & n11641 ) ;
  assign n11643 = ( ~n11275 & n11640 ) | ( ~n11275 & n11641 ) | ( n11640 & n11641 ) ;
  assign n11644 = ( n11275 & ~n11642 ) | ( n11275 & n11643 ) | ( ~n11642 & n11643 ) ;
  assign n11645 = ( x99 & n11639 ) | ( x99 & ~n11644 ) | ( n11639 & ~n11644 ) ;
  assign n11646 = ( x99 & n11276 ) | ( x99 & ~n11437 ) | ( n11276 & ~n11437 ) ;
  assign n11647 = x99 & n11276 ;
  assign n11648 = ( ~n11281 & n11646 ) | ( ~n11281 & n11647 ) | ( n11646 & n11647 ) ;
  assign n11649 = ( n11281 & n11646 ) | ( n11281 & n11647 ) | ( n11646 & n11647 ) ;
  assign n11650 = ( n11281 & n11648 ) | ( n11281 & ~n11649 ) | ( n11648 & ~n11649 ) ;
  assign n11651 = ( x100 & n11645 ) | ( x100 & ~n11650 ) | ( n11645 & ~n11650 ) ;
  assign n11652 = ( x100 & n11282 ) | ( x100 & ~n11437 ) | ( n11282 & ~n11437 ) ;
  assign n11653 = x100 & n11282 ;
  assign n11654 = ( n11287 & n11652 ) | ( n11287 & n11653 ) | ( n11652 & n11653 ) ;
  assign n11655 = ( ~n11287 & n11652 ) | ( ~n11287 & n11653 ) | ( n11652 & n11653 ) ;
  assign n11656 = ( n11287 & ~n11654 ) | ( n11287 & n11655 ) | ( ~n11654 & n11655 ) ;
  assign n11657 = ( x101 & n11651 ) | ( x101 & ~n11656 ) | ( n11651 & ~n11656 ) ;
  assign n11658 = ( x101 & n11288 ) | ( x101 & ~n11437 ) | ( n11288 & ~n11437 ) ;
  assign n11659 = x101 & n11288 ;
  assign n11660 = ( ~n11293 & n11658 ) | ( ~n11293 & n11659 ) | ( n11658 & n11659 ) ;
  assign n11661 = ( n11293 & n11658 ) | ( n11293 & n11659 ) | ( n11658 & n11659 ) ;
  assign n11662 = ( n11293 & n11660 ) | ( n11293 & ~n11661 ) | ( n11660 & ~n11661 ) ;
  assign n11663 = ( x102 & n11657 ) | ( x102 & ~n11662 ) | ( n11657 & ~n11662 ) ;
  assign n11664 = ( x102 & n11294 ) | ( x102 & ~n11437 ) | ( n11294 & ~n11437 ) ;
  assign n11665 = x102 & n11294 ;
  assign n11666 = ( n11299 & n11664 ) | ( n11299 & n11665 ) | ( n11664 & n11665 ) ;
  assign n11667 = ( ~n11299 & n11664 ) | ( ~n11299 & n11665 ) | ( n11664 & n11665 ) ;
  assign n11668 = ( n11299 & ~n11666 ) | ( n11299 & n11667 ) | ( ~n11666 & n11667 ) ;
  assign n11669 = ( x103 & n11663 ) | ( x103 & ~n11668 ) | ( n11663 & ~n11668 ) ;
  assign n11670 = ( x103 & n11300 ) | ( x103 & ~n11437 ) | ( n11300 & ~n11437 ) ;
  assign n11671 = x103 & n11300 ;
  assign n11672 = ( ~n11305 & n11670 ) | ( ~n11305 & n11671 ) | ( n11670 & n11671 ) ;
  assign n11673 = ( n11305 & n11670 ) | ( n11305 & n11671 ) | ( n11670 & n11671 ) ;
  assign n11674 = ( n11305 & n11672 ) | ( n11305 & ~n11673 ) | ( n11672 & ~n11673 ) ;
  assign n11675 = ( x104 & n11669 ) | ( x104 & ~n11674 ) | ( n11669 & ~n11674 ) ;
  assign n11676 = ( x104 & n11306 ) | ( x104 & ~n11437 ) | ( n11306 & ~n11437 ) ;
  assign n11677 = x104 & n11306 ;
  assign n11678 = ( n11311 & n11676 ) | ( n11311 & n11677 ) | ( n11676 & n11677 ) ;
  assign n11679 = ( ~n11311 & n11676 ) | ( ~n11311 & n11677 ) | ( n11676 & n11677 ) ;
  assign n11680 = ( n11311 & ~n11678 ) | ( n11311 & n11679 ) | ( ~n11678 & n11679 ) ;
  assign n11681 = ( x105 & n11675 ) | ( x105 & ~n11680 ) | ( n11675 & ~n11680 ) ;
  assign n11682 = ( x105 & n11312 ) | ( x105 & ~n11437 ) | ( n11312 & ~n11437 ) ;
  assign n11683 = x105 & n11312 ;
  assign n11684 = ( ~n11317 & n11682 ) | ( ~n11317 & n11683 ) | ( n11682 & n11683 ) ;
  assign n11685 = ( n11317 & n11682 ) | ( n11317 & n11683 ) | ( n11682 & n11683 ) ;
  assign n11686 = ( n11317 & n11684 ) | ( n11317 & ~n11685 ) | ( n11684 & ~n11685 ) ;
  assign n11687 = ( x106 & n11681 ) | ( x106 & ~n11686 ) | ( n11681 & ~n11686 ) ;
  assign n11688 = ( x106 & n11318 ) | ( x106 & ~n11437 ) | ( n11318 & ~n11437 ) ;
  assign n11689 = x106 & n11318 ;
  assign n11690 = ( n11323 & n11688 ) | ( n11323 & n11689 ) | ( n11688 & n11689 ) ;
  assign n11691 = ( ~n11323 & n11688 ) | ( ~n11323 & n11689 ) | ( n11688 & n11689 ) ;
  assign n11692 = ( n11323 & ~n11690 ) | ( n11323 & n11691 ) | ( ~n11690 & n11691 ) ;
  assign n11693 = ( x107 & n11687 ) | ( x107 & ~n11692 ) | ( n11687 & ~n11692 ) ;
  assign n11694 = ( x107 & n11324 ) | ( x107 & ~n11437 ) | ( n11324 & ~n11437 ) ;
  assign n11695 = x107 & n11324 ;
  assign n11696 = ( ~n11329 & n11694 ) | ( ~n11329 & n11695 ) | ( n11694 & n11695 ) ;
  assign n11697 = ( n11329 & n11694 ) | ( n11329 & n11695 ) | ( n11694 & n11695 ) ;
  assign n11698 = ( n11329 & n11696 ) | ( n11329 & ~n11697 ) | ( n11696 & ~n11697 ) ;
  assign n11699 = ( x108 & n11693 ) | ( x108 & ~n11698 ) | ( n11693 & ~n11698 ) ;
  assign n11700 = ( x108 & n11330 ) | ( x108 & ~n11437 ) | ( n11330 & ~n11437 ) ;
  assign n11701 = x108 & n11330 ;
  assign n11702 = ( n11335 & n11700 ) | ( n11335 & n11701 ) | ( n11700 & n11701 ) ;
  assign n11703 = ( ~n11335 & n11700 ) | ( ~n11335 & n11701 ) | ( n11700 & n11701 ) ;
  assign n11704 = ( n11335 & ~n11702 ) | ( n11335 & n11703 ) | ( ~n11702 & n11703 ) ;
  assign n11705 = ( x109 & n11699 ) | ( x109 & ~n11704 ) | ( n11699 & ~n11704 ) ;
  assign n11706 = ( x109 & n11336 ) | ( x109 & ~n11437 ) | ( n11336 & ~n11437 ) ;
  assign n11707 = x109 & n11336 ;
  assign n11708 = ( ~n11341 & n11706 ) | ( ~n11341 & n11707 ) | ( n11706 & n11707 ) ;
  assign n11709 = ( n11341 & n11706 ) | ( n11341 & n11707 ) | ( n11706 & n11707 ) ;
  assign n11710 = ( n11341 & n11708 ) | ( n11341 & ~n11709 ) | ( n11708 & ~n11709 ) ;
  assign n11711 = ( x110 & n11705 ) | ( x110 & ~n11710 ) | ( n11705 & ~n11710 ) ;
  assign n11712 = ( x110 & n11342 ) | ( x110 & ~n11437 ) | ( n11342 & ~n11437 ) ;
  assign n11713 = x110 & n11342 ;
  assign n11714 = ( n11347 & n11712 ) | ( n11347 & n11713 ) | ( n11712 & n11713 ) ;
  assign n11715 = ( ~n11347 & n11712 ) | ( ~n11347 & n11713 ) | ( n11712 & n11713 ) ;
  assign n11716 = ( n11347 & ~n11714 ) | ( n11347 & n11715 ) | ( ~n11714 & n11715 ) ;
  assign n11717 = ( x111 & n11711 ) | ( x111 & ~n11716 ) | ( n11711 & ~n11716 ) ;
  assign n11718 = ( x111 & n11348 ) | ( x111 & ~n11437 ) | ( n11348 & ~n11437 ) ;
  assign n11719 = x111 & n11348 ;
  assign n11720 = ( ~n11353 & n11718 ) | ( ~n11353 & n11719 ) | ( n11718 & n11719 ) ;
  assign n11721 = ( n11353 & n11718 ) | ( n11353 & n11719 ) | ( n11718 & n11719 ) ;
  assign n11722 = ( n11353 & n11720 ) | ( n11353 & ~n11721 ) | ( n11720 & ~n11721 ) ;
  assign n11723 = ( x112 & n11717 ) | ( x112 & ~n11722 ) | ( n11717 & ~n11722 ) ;
  assign n11724 = ( x112 & n11354 ) | ( x112 & ~n11437 ) | ( n11354 & ~n11437 ) ;
  assign n11725 = x112 & n11354 ;
  assign n11726 = ( n11359 & n11724 ) | ( n11359 & n11725 ) | ( n11724 & n11725 ) ;
  assign n11727 = ( ~n11359 & n11724 ) | ( ~n11359 & n11725 ) | ( n11724 & n11725 ) ;
  assign n11728 = ( n11359 & ~n11726 ) | ( n11359 & n11727 ) | ( ~n11726 & n11727 ) ;
  assign n11729 = ( x113 & n11723 ) | ( x113 & ~n11728 ) | ( n11723 & ~n11728 ) ;
  assign n11730 = ( x113 & n11360 ) | ( x113 & ~n11437 ) | ( n11360 & ~n11437 ) ;
  assign n11731 = x113 & n11360 ;
  assign n11732 = ( ~n11365 & n11730 ) | ( ~n11365 & n11731 ) | ( n11730 & n11731 ) ;
  assign n11733 = ( n11365 & n11730 ) | ( n11365 & n11731 ) | ( n11730 & n11731 ) ;
  assign n11734 = ( n11365 & n11732 ) | ( n11365 & ~n11733 ) | ( n11732 & ~n11733 ) ;
  assign n11735 = ( x114 & n11729 ) | ( x114 & ~n11734 ) | ( n11729 & ~n11734 ) ;
  assign n11736 = ( x114 & n11366 ) | ( x114 & ~n11437 ) | ( n11366 & ~n11437 ) ;
  assign n11737 = x114 & n11366 ;
  assign n11738 = ( n11371 & n11736 ) | ( n11371 & n11737 ) | ( n11736 & n11737 ) ;
  assign n11739 = ( ~n11371 & n11736 ) | ( ~n11371 & n11737 ) | ( n11736 & n11737 ) ;
  assign n11740 = ( n11371 & ~n11738 ) | ( n11371 & n11739 ) | ( ~n11738 & n11739 ) ;
  assign n11741 = ( x115 & n11735 ) | ( x115 & ~n11740 ) | ( n11735 & ~n11740 ) ;
  assign n11742 = ( x115 & n11372 ) | ( x115 & ~n11437 ) | ( n11372 & ~n11437 ) ;
  assign n11743 = x115 & n11372 ;
  assign n11744 = ( ~n11377 & n11742 ) | ( ~n11377 & n11743 ) | ( n11742 & n11743 ) ;
  assign n11745 = ( n11377 & n11742 ) | ( n11377 & n11743 ) | ( n11742 & n11743 ) ;
  assign n11746 = ( n11377 & n11744 ) | ( n11377 & ~n11745 ) | ( n11744 & ~n11745 ) ;
  assign n11747 = ( x116 & n11741 ) | ( x116 & ~n11746 ) | ( n11741 & ~n11746 ) ;
  assign n11748 = ( x116 & n11378 ) | ( x116 & ~n11437 ) | ( n11378 & ~n11437 ) ;
  assign n11749 = x116 & n11378 ;
  assign n11750 = ( n11383 & n11748 ) | ( n11383 & n11749 ) | ( n11748 & n11749 ) ;
  assign n11751 = ( ~n11383 & n11748 ) | ( ~n11383 & n11749 ) | ( n11748 & n11749 ) ;
  assign n11752 = ( n11383 & ~n11750 ) | ( n11383 & n11751 ) | ( ~n11750 & n11751 ) ;
  assign n11753 = ( x117 & n11747 ) | ( x117 & ~n11752 ) | ( n11747 & ~n11752 ) ;
  assign n11754 = ( x117 & n11384 ) | ( x117 & ~n11437 ) | ( n11384 & ~n11437 ) ;
  assign n11755 = x117 & n11384 ;
  assign n11756 = ( ~n11389 & n11754 ) | ( ~n11389 & n11755 ) | ( n11754 & n11755 ) ;
  assign n11757 = ( n11389 & n11754 ) | ( n11389 & n11755 ) | ( n11754 & n11755 ) ;
  assign n11758 = ( n11389 & n11756 ) | ( n11389 & ~n11757 ) | ( n11756 & ~n11757 ) ;
  assign n11759 = ( x118 & n11753 ) | ( x118 & ~n11758 ) | ( n11753 & ~n11758 ) ;
  assign n11760 = ( x118 & n11390 ) | ( x118 & ~n11437 ) | ( n11390 & ~n11437 ) ;
  assign n11761 = x118 & n11390 ;
  assign n11762 = ( n11395 & n11760 ) | ( n11395 & n11761 ) | ( n11760 & n11761 ) ;
  assign n11763 = ( ~n11395 & n11760 ) | ( ~n11395 & n11761 ) | ( n11760 & n11761 ) ;
  assign n11764 = ( n11395 & ~n11762 ) | ( n11395 & n11763 ) | ( ~n11762 & n11763 ) ;
  assign n11765 = ( x119 & n11759 ) | ( x119 & ~n11764 ) | ( n11759 & ~n11764 ) ;
  assign n11766 = ( x119 & n11396 ) | ( x119 & ~n11437 ) | ( n11396 & ~n11437 ) ;
  assign n11767 = x119 & n11396 ;
  assign n11768 = ( ~n11401 & n11766 ) | ( ~n11401 & n11767 ) | ( n11766 & n11767 ) ;
  assign n11769 = ( n11401 & n11766 ) | ( n11401 & n11767 ) | ( n11766 & n11767 ) ;
  assign n11770 = ( n11401 & n11768 ) | ( n11401 & ~n11769 ) | ( n11768 & ~n11769 ) ;
  assign n11771 = ( x120 & n11765 ) | ( x120 & ~n11770 ) | ( n11765 & ~n11770 ) ;
  assign n11772 = ( x120 & n11402 ) | ( x120 & ~n11437 ) | ( n11402 & ~n11437 ) ;
  assign n11773 = x120 & n11402 ;
  assign n11774 = ( n11407 & n11772 ) | ( n11407 & n11773 ) | ( n11772 & n11773 ) ;
  assign n11775 = ( ~n11407 & n11772 ) | ( ~n11407 & n11773 ) | ( n11772 & n11773 ) ;
  assign n11776 = ( n11407 & ~n11774 ) | ( n11407 & n11775 ) | ( ~n11774 & n11775 ) ;
  assign n11777 = ( x121 & n11771 ) | ( x121 & ~n11776 ) | ( n11771 & ~n11776 ) ;
  assign n11778 = ( x121 & n11408 ) | ( x121 & ~n11437 ) | ( n11408 & ~n11437 ) ;
  assign n11779 = x121 & n11408 ;
  assign n11780 = ( ~n11413 & n11778 ) | ( ~n11413 & n11779 ) | ( n11778 & n11779 ) ;
  assign n11781 = ( n11413 & n11778 ) | ( n11413 & n11779 ) | ( n11778 & n11779 ) ;
  assign n11782 = ( n11413 & n11780 ) | ( n11413 & ~n11781 ) | ( n11780 & ~n11781 ) ;
  assign n11783 = ( x122 & n11777 ) | ( x122 & ~n11782 ) | ( n11777 & ~n11782 ) ;
  assign n11784 = ( x122 & n11414 ) | ( x122 & ~n11437 ) | ( n11414 & ~n11437 ) ;
  assign n11785 = x122 & n11414 ;
  assign n11786 = ( n11419 & n11784 ) | ( n11419 & n11785 ) | ( n11784 & n11785 ) ;
  assign n11787 = ( ~n11419 & n11784 ) | ( ~n11419 & n11785 ) | ( n11784 & n11785 ) ;
  assign n11788 = ( n11419 & ~n11786 ) | ( n11419 & n11787 ) | ( ~n11786 & n11787 ) ;
  assign n11789 = ( x123 & n11783 ) | ( x123 & ~n11788 ) | ( n11783 & ~n11788 ) ;
  assign n11790 = ( x123 & n11420 ) | ( x123 & ~n11437 ) | ( n11420 & ~n11437 ) ;
  assign n11791 = x123 & n11420 ;
  assign n11792 = ( ~n11425 & n11790 ) | ( ~n11425 & n11791 ) | ( n11790 & n11791 ) ;
  assign n11793 = ( n11425 & n11790 ) | ( n11425 & n11791 ) | ( n11790 & n11791 ) ;
  assign n11794 = ( n11425 & n11792 ) | ( n11425 & ~n11793 ) | ( n11792 & ~n11793 ) ;
  assign n11795 = ( x124 & n11789 ) | ( x124 & ~n11794 ) | ( n11789 & ~n11794 ) ;
  assign n11796 = ( x124 & n11426 ) | ( x124 & ~n11437 ) | ( n11426 & ~n11437 ) ;
  assign n11797 = x124 & n11426 ;
  assign n11798 = ( ~n11431 & n11796 ) | ( ~n11431 & n11797 ) | ( n11796 & n11797 ) ;
  assign n11799 = ( n11431 & n11796 ) | ( n11431 & n11797 ) | ( n11796 & n11797 ) ;
  assign n11800 = ( n11431 & n11798 ) | ( n11431 & ~n11799 ) | ( n11798 & ~n11799 ) ;
  assign n11801 = ( x125 & n11795 ) | ( x125 & ~n11800 ) | ( n11795 & ~n11800 ) ;
  assign n11802 = ( x126 & ~n11435 ) | ( x126 & n11801 ) | ( ~n11435 & n11801 ) ;
  assign n11803 = x127 | n11802 ;
  assign n11804 = ( x1 & ~x64 ) | ( x1 & n11803 ) | ( ~x64 & n11803 ) ;
  assign n11805 = ~x1 & n11803 ;
  assign n11806 = ( n129 & n11804 ) | ( n129 & ~n11805 ) | ( n11804 & ~n11805 ) ;
  assign n11807 = ~x0 & x64 ;
  assign n11808 = ( x65 & ~n11806 ) | ( x65 & n11807 ) | ( ~n11806 & n11807 ) ;
  assign n11809 = ( x65 & n129 ) | ( x65 & ~n11803 ) | ( n129 & ~n11803 ) ;
  assign n11810 = x65 & n129 ;
  assign n11811 = ( n11440 & n11809 ) | ( n11440 & n11810 ) | ( n11809 & n11810 ) ;
  assign n11812 = ( ~n11440 & n11809 ) | ( ~n11440 & n11810 ) | ( n11809 & n11810 ) ;
  assign n11813 = ( n11440 & ~n11811 ) | ( n11440 & n11812 ) | ( ~n11811 & n11812 ) ;
  assign n11814 = ( x66 & n11808 ) | ( x66 & ~n11813 ) | ( n11808 & ~n11813 ) ;
  assign n11815 = ( x66 & n11441 ) | ( x66 & ~n11803 ) | ( n11441 & ~n11803 ) ;
  assign n11816 = x66 & n11441 ;
  assign n11817 = ( n11446 & n11815 ) | ( n11446 & n11816 ) | ( n11815 & n11816 ) ;
  assign n11818 = ( ~n11446 & n11815 ) | ( ~n11446 & n11816 ) | ( n11815 & n11816 ) ;
  assign n11819 = ( n11446 & ~n11817 ) | ( n11446 & n11818 ) | ( ~n11817 & n11818 ) ;
  assign n11820 = ( x67 & n11814 ) | ( x67 & ~n11819 ) | ( n11814 & ~n11819 ) ;
  assign n11821 = ( x67 & n11447 ) | ( x67 & ~n11803 ) | ( n11447 & ~n11803 ) ;
  assign n11822 = x67 & n11447 ;
  assign n11823 = ( ~n11452 & n11821 ) | ( ~n11452 & n11822 ) | ( n11821 & n11822 ) ;
  assign n11824 = ( n11452 & n11821 ) | ( n11452 & n11822 ) | ( n11821 & n11822 ) ;
  assign n11825 = ( n11452 & n11823 ) | ( n11452 & ~n11824 ) | ( n11823 & ~n11824 ) ;
  assign n11826 = ( x68 & n11820 ) | ( x68 & ~n11825 ) | ( n11820 & ~n11825 ) ;
  assign n11827 = ( x68 & n11453 ) | ( x68 & ~n11803 ) | ( n11453 & ~n11803 ) ;
  assign n11828 = x68 & n11453 ;
  assign n11829 = ( n11458 & n11827 ) | ( n11458 & n11828 ) | ( n11827 & n11828 ) ;
  assign n11830 = ( ~n11458 & n11827 ) | ( ~n11458 & n11828 ) | ( n11827 & n11828 ) ;
  assign n11831 = ( n11458 & ~n11829 ) | ( n11458 & n11830 ) | ( ~n11829 & n11830 ) ;
  assign n11832 = ( x69 & n11826 ) | ( x69 & ~n11831 ) | ( n11826 & ~n11831 ) ;
  assign n11833 = ( x69 & n11459 ) | ( x69 & ~n11803 ) | ( n11459 & ~n11803 ) ;
  assign n11834 = x69 & n11459 ;
  assign n11835 = ( ~n11464 & n11833 ) | ( ~n11464 & n11834 ) | ( n11833 & n11834 ) ;
  assign n11836 = ( n11464 & n11833 ) | ( n11464 & n11834 ) | ( n11833 & n11834 ) ;
  assign n11837 = ( n11464 & n11835 ) | ( n11464 & ~n11836 ) | ( n11835 & ~n11836 ) ;
  assign n11838 = ( x70 & n11832 ) | ( x70 & ~n11837 ) | ( n11832 & ~n11837 ) ;
  assign n11839 = ( x70 & n11465 ) | ( x70 & ~n11803 ) | ( n11465 & ~n11803 ) ;
  assign n11840 = x70 & n11465 ;
  assign n11841 = ( n11470 & n11839 ) | ( n11470 & n11840 ) | ( n11839 & n11840 ) ;
  assign n11842 = ( ~n11470 & n11839 ) | ( ~n11470 & n11840 ) | ( n11839 & n11840 ) ;
  assign n11843 = ( n11470 & ~n11841 ) | ( n11470 & n11842 ) | ( ~n11841 & n11842 ) ;
  assign n11844 = ( x71 & n11838 ) | ( x71 & ~n11843 ) | ( n11838 & ~n11843 ) ;
  assign n11845 = ( x71 & n11471 ) | ( x71 & ~n11803 ) | ( n11471 & ~n11803 ) ;
  assign n11846 = x71 & n11471 ;
  assign n11847 = ( ~n11476 & n11845 ) | ( ~n11476 & n11846 ) | ( n11845 & n11846 ) ;
  assign n11848 = ( n11476 & n11845 ) | ( n11476 & n11846 ) | ( n11845 & n11846 ) ;
  assign n11849 = ( n11476 & n11847 ) | ( n11476 & ~n11848 ) | ( n11847 & ~n11848 ) ;
  assign n11850 = ( x72 & n11844 ) | ( x72 & ~n11849 ) | ( n11844 & ~n11849 ) ;
  assign n11851 = ( x72 & n11477 ) | ( x72 & ~n11803 ) | ( n11477 & ~n11803 ) ;
  assign n11852 = x72 & n11477 ;
  assign n11853 = ( n11482 & n11851 ) | ( n11482 & n11852 ) | ( n11851 & n11852 ) ;
  assign n11854 = ( ~n11482 & n11851 ) | ( ~n11482 & n11852 ) | ( n11851 & n11852 ) ;
  assign n11855 = ( n11482 & ~n11853 ) | ( n11482 & n11854 ) | ( ~n11853 & n11854 ) ;
  assign n11856 = ( x73 & n11850 ) | ( x73 & ~n11855 ) | ( n11850 & ~n11855 ) ;
  assign n11857 = ( x73 & n11483 ) | ( x73 & ~n11803 ) | ( n11483 & ~n11803 ) ;
  assign n11858 = x73 & n11483 ;
  assign n11859 = ( ~n11488 & n11857 ) | ( ~n11488 & n11858 ) | ( n11857 & n11858 ) ;
  assign n11860 = ( n11488 & n11857 ) | ( n11488 & n11858 ) | ( n11857 & n11858 ) ;
  assign n11861 = ( n11488 & n11859 ) | ( n11488 & ~n11860 ) | ( n11859 & ~n11860 ) ;
  assign n11862 = ( x74 & n11856 ) | ( x74 & ~n11861 ) | ( n11856 & ~n11861 ) ;
  assign n11863 = ( x74 & n11489 ) | ( x74 & ~n11803 ) | ( n11489 & ~n11803 ) ;
  assign n11864 = x74 & n11489 ;
  assign n11865 = ( n11494 & n11863 ) | ( n11494 & n11864 ) | ( n11863 & n11864 ) ;
  assign n11866 = ( ~n11494 & n11863 ) | ( ~n11494 & n11864 ) | ( n11863 & n11864 ) ;
  assign n11867 = ( n11494 & ~n11865 ) | ( n11494 & n11866 ) | ( ~n11865 & n11866 ) ;
  assign n11868 = ( x75 & n11862 ) | ( x75 & ~n11867 ) | ( n11862 & ~n11867 ) ;
  assign n11869 = ( x75 & n11495 ) | ( x75 & ~n11803 ) | ( n11495 & ~n11803 ) ;
  assign n11870 = x75 & n11495 ;
  assign n11871 = ( ~n11500 & n11869 ) | ( ~n11500 & n11870 ) | ( n11869 & n11870 ) ;
  assign n11872 = ( n11500 & n11869 ) | ( n11500 & n11870 ) | ( n11869 & n11870 ) ;
  assign n11873 = ( n11500 & n11871 ) | ( n11500 & ~n11872 ) | ( n11871 & ~n11872 ) ;
  assign n11874 = ( x76 & n11868 ) | ( x76 & ~n11873 ) | ( n11868 & ~n11873 ) ;
  assign n11875 = ( x76 & n11501 ) | ( x76 & ~n11803 ) | ( n11501 & ~n11803 ) ;
  assign n11876 = x76 & n11501 ;
  assign n11877 = ( n11506 & n11875 ) | ( n11506 & n11876 ) | ( n11875 & n11876 ) ;
  assign n11878 = ( ~n11506 & n11875 ) | ( ~n11506 & n11876 ) | ( n11875 & n11876 ) ;
  assign n11879 = ( n11506 & ~n11877 ) | ( n11506 & n11878 ) | ( ~n11877 & n11878 ) ;
  assign n11880 = ( x77 & n11874 ) | ( x77 & ~n11879 ) | ( n11874 & ~n11879 ) ;
  assign n11881 = ( x77 & n11507 ) | ( x77 & ~n11803 ) | ( n11507 & ~n11803 ) ;
  assign n11882 = x77 & n11507 ;
  assign n11883 = ( ~n11512 & n11881 ) | ( ~n11512 & n11882 ) | ( n11881 & n11882 ) ;
  assign n11884 = ( n11512 & n11881 ) | ( n11512 & n11882 ) | ( n11881 & n11882 ) ;
  assign n11885 = ( n11512 & n11883 ) | ( n11512 & ~n11884 ) | ( n11883 & ~n11884 ) ;
  assign n11886 = ( x78 & n11880 ) | ( x78 & ~n11885 ) | ( n11880 & ~n11885 ) ;
  assign n11887 = ( x78 & n11513 ) | ( x78 & ~n11803 ) | ( n11513 & ~n11803 ) ;
  assign n11888 = x78 & n11513 ;
  assign n11889 = ( n11518 & n11887 ) | ( n11518 & n11888 ) | ( n11887 & n11888 ) ;
  assign n11890 = ( ~n11518 & n11887 ) | ( ~n11518 & n11888 ) | ( n11887 & n11888 ) ;
  assign n11891 = ( n11518 & ~n11889 ) | ( n11518 & n11890 ) | ( ~n11889 & n11890 ) ;
  assign n11892 = ( x79 & n11886 ) | ( x79 & ~n11891 ) | ( n11886 & ~n11891 ) ;
  assign n11893 = ( x79 & n11519 ) | ( x79 & ~n11803 ) | ( n11519 & ~n11803 ) ;
  assign n11894 = x79 & n11519 ;
  assign n11895 = ( ~n11524 & n11893 ) | ( ~n11524 & n11894 ) | ( n11893 & n11894 ) ;
  assign n11896 = ( n11524 & n11893 ) | ( n11524 & n11894 ) | ( n11893 & n11894 ) ;
  assign n11897 = ( n11524 & n11895 ) | ( n11524 & ~n11896 ) | ( n11895 & ~n11896 ) ;
  assign n11898 = ( x80 & n11892 ) | ( x80 & ~n11897 ) | ( n11892 & ~n11897 ) ;
  assign n11899 = ( x80 & n11525 ) | ( x80 & ~n11803 ) | ( n11525 & ~n11803 ) ;
  assign n11900 = x80 & n11525 ;
  assign n11901 = ( n11530 & n11899 ) | ( n11530 & n11900 ) | ( n11899 & n11900 ) ;
  assign n11902 = ( ~n11530 & n11899 ) | ( ~n11530 & n11900 ) | ( n11899 & n11900 ) ;
  assign n11903 = ( n11530 & ~n11901 ) | ( n11530 & n11902 ) | ( ~n11901 & n11902 ) ;
  assign n11904 = ( x81 & n11898 ) | ( x81 & ~n11903 ) | ( n11898 & ~n11903 ) ;
  assign n11905 = ( x81 & n11531 ) | ( x81 & ~n11803 ) | ( n11531 & ~n11803 ) ;
  assign n11906 = x81 & n11531 ;
  assign n11907 = ( ~n11536 & n11905 ) | ( ~n11536 & n11906 ) | ( n11905 & n11906 ) ;
  assign n11908 = ( n11536 & n11905 ) | ( n11536 & n11906 ) | ( n11905 & n11906 ) ;
  assign n11909 = ( n11536 & n11907 ) | ( n11536 & ~n11908 ) | ( n11907 & ~n11908 ) ;
  assign n11910 = ( x82 & n11904 ) | ( x82 & ~n11909 ) | ( n11904 & ~n11909 ) ;
  assign n11911 = ( x82 & n11537 ) | ( x82 & ~n11803 ) | ( n11537 & ~n11803 ) ;
  assign n11912 = x82 & n11537 ;
  assign n11913 = ( n11542 & n11911 ) | ( n11542 & n11912 ) | ( n11911 & n11912 ) ;
  assign n11914 = ( ~n11542 & n11911 ) | ( ~n11542 & n11912 ) | ( n11911 & n11912 ) ;
  assign n11915 = ( n11542 & ~n11913 ) | ( n11542 & n11914 ) | ( ~n11913 & n11914 ) ;
  assign n11916 = ( x83 & n11910 ) | ( x83 & ~n11915 ) | ( n11910 & ~n11915 ) ;
  assign n11917 = ( x83 & n11543 ) | ( x83 & ~n11803 ) | ( n11543 & ~n11803 ) ;
  assign n11918 = x83 & n11543 ;
  assign n11919 = ( ~n11548 & n11917 ) | ( ~n11548 & n11918 ) | ( n11917 & n11918 ) ;
  assign n11920 = ( n11548 & n11917 ) | ( n11548 & n11918 ) | ( n11917 & n11918 ) ;
  assign n11921 = ( n11548 & n11919 ) | ( n11548 & ~n11920 ) | ( n11919 & ~n11920 ) ;
  assign n11922 = ( x84 & n11916 ) | ( x84 & ~n11921 ) | ( n11916 & ~n11921 ) ;
  assign n11923 = ( x84 & n11549 ) | ( x84 & ~n11803 ) | ( n11549 & ~n11803 ) ;
  assign n11924 = x84 & n11549 ;
  assign n11925 = ( n11554 & n11923 ) | ( n11554 & n11924 ) | ( n11923 & n11924 ) ;
  assign n11926 = ( ~n11554 & n11923 ) | ( ~n11554 & n11924 ) | ( n11923 & n11924 ) ;
  assign n11927 = ( n11554 & ~n11925 ) | ( n11554 & n11926 ) | ( ~n11925 & n11926 ) ;
  assign n11928 = ( x85 & n11922 ) | ( x85 & ~n11927 ) | ( n11922 & ~n11927 ) ;
  assign n11929 = ( x85 & n11555 ) | ( x85 & ~n11803 ) | ( n11555 & ~n11803 ) ;
  assign n11930 = x85 & n11555 ;
  assign n11931 = ( ~n11560 & n11929 ) | ( ~n11560 & n11930 ) | ( n11929 & n11930 ) ;
  assign n11932 = ( n11560 & n11929 ) | ( n11560 & n11930 ) | ( n11929 & n11930 ) ;
  assign n11933 = ( n11560 & n11931 ) | ( n11560 & ~n11932 ) | ( n11931 & ~n11932 ) ;
  assign n11934 = ( x86 & n11928 ) | ( x86 & ~n11933 ) | ( n11928 & ~n11933 ) ;
  assign n11935 = ( x86 & n11561 ) | ( x86 & ~n11803 ) | ( n11561 & ~n11803 ) ;
  assign n11936 = x86 & n11561 ;
  assign n11937 = ( n11566 & n11935 ) | ( n11566 & n11936 ) | ( n11935 & n11936 ) ;
  assign n11938 = ( ~n11566 & n11935 ) | ( ~n11566 & n11936 ) | ( n11935 & n11936 ) ;
  assign n11939 = ( n11566 & ~n11937 ) | ( n11566 & n11938 ) | ( ~n11937 & n11938 ) ;
  assign n11940 = ( x87 & n11934 ) | ( x87 & ~n11939 ) | ( n11934 & ~n11939 ) ;
  assign n11941 = ( x87 & n11567 ) | ( x87 & ~n11803 ) | ( n11567 & ~n11803 ) ;
  assign n11942 = x87 & n11567 ;
  assign n11943 = ( ~n11572 & n11941 ) | ( ~n11572 & n11942 ) | ( n11941 & n11942 ) ;
  assign n11944 = ( n11572 & n11941 ) | ( n11572 & n11942 ) | ( n11941 & n11942 ) ;
  assign n11945 = ( n11572 & n11943 ) | ( n11572 & ~n11944 ) | ( n11943 & ~n11944 ) ;
  assign n11946 = ( x88 & n11940 ) | ( x88 & ~n11945 ) | ( n11940 & ~n11945 ) ;
  assign n11947 = ( x88 & n11573 ) | ( x88 & ~n11803 ) | ( n11573 & ~n11803 ) ;
  assign n11948 = x88 & n11573 ;
  assign n11949 = ( n11578 & n11947 ) | ( n11578 & n11948 ) | ( n11947 & n11948 ) ;
  assign n11950 = ( ~n11578 & n11947 ) | ( ~n11578 & n11948 ) | ( n11947 & n11948 ) ;
  assign n11951 = ( n11578 & ~n11949 ) | ( n11578 & n11950 ) | ( ~n11949 & n11950 ) ;
  assign n11952 = ( x89 & n11946 ) | ( x89 & ~n11951 ) | ( n11946 & ~n11951 ) ;
  assign n11953 = ( x89 & n11579 ) | ( x89 & ~n11803 ) | ( n11579 & ~n11803 ) ;
  assign n11954 = x89 & n11579 ;
  assign n11955 = ( ~n11584 & n11953 ) | ( ~n11584 & n11954 ) | ( n11953 & n11954 ) ;
  assign n11956 = ( n11584 & n11953 ) | ( n11584 & n11954 ) | ( n11953 & n11954 ) ;
  assign n11957 = ( n11584 & n11955 ) | ( n11584 & ~n11956 ) | ( n11955 & ~n11956 ) ;
  assign n11958 = ( x90 & n11952 ) | ( x90 & ~n11957 ) | ( n11952 & ~n11957 ) ;
  assign n11959 = ( x90 & n11585 ) | ( x90 & ~n11803 ) | ( n11585 & ~n11803 ) ;
  assign n11960 = x90 & n11585 ;
  assign n11961 = ( n11590 & n11959 ) | ( n11590 & n11960 ) | ( n11959 & n11960 ) ;
  assign n11962 = ( ~n11590 & n11959 ) | ( ~n11590 & n11960 ) | ( n11959 & n11960 ) ;
  assign n11963 = ( n11590 & ~n11961 ) | ( n11590 & n11962 ) | ( ~n11961 & n11962 ) ;
  assign n11964 = ( x91 & n11958 ) | ( x91 & ~n11963 ) | ( n11958 & ~n11963 ) ;
  assign n11965 = ( x91 & n11591 ) | ( x91 & ~n11803 ) | ( n11591 & ~n11803 ) ;
  assign n11966 = x91 & n11591 ;
  assign n11967 = ( ~n11596 & n11965 ) | ( ~n11596 & n11966 ) | ( n11965 & n11966 ) ;
  assign n11968 = ( n11596 & n11965 ) | ( n11596 & n11966 ) | ( n11965 & n11966 ) ;
  assign n11969 = ( n11596 & n11967 ) | ( n11596 & ~n11968 ) | ( n11967 & ~n11968 ) ;
  assign n11970 = ( x92 & n11964 ) | ( x92 & ~n11969 ) | ( n11964 & ~n11969 ) ;
  assign n11971 = ( x92 & n11597 ) | ( x92 & ~n11803 ) | ( n11597 & ~n11803 ) ;
  assign n11972 = x92 & n11597 ;
  assign n11973 = ( n11602 & n11971 ) | ( n11602 & n11972 ) | ( n11971 & n11972 ) ;
  assign n11974 = ( ~n11602 & n11971 ) | ( ~n11602 & n11972 ) | ( n11971 & n11972 ) ;
  assign n11975 = ( n11602 & ~n11973 ) | ( n11602 & n11974 ) | ( ~n11973 & n11974 ) ;
  assign n11976 = ( x93 & n11970 ) | ( x93 & ~n11975 ) | ( n11970 & ~n11975 ) ;
  assign n11977 = ( x93 & n11603 ) | ( x93 & ~n11803 ) | ( n11603 & ~n11803 ) ;
  assign n11978 = x93 & n11603 ;
  assign n11979 = ( ~n11608 & n11977 ) | ( ~n11608 & n11978 ) | ( n11977 & n11978 ) ;
  assign n11980 = ( n11608 & n11977 ) | ( n11608 & n11978 ) | ( n11977 & n11978 ) ;
  assign n11981 = ( n11608 & n11979 ) | ( n11608 & ~n11980 ) | ( n11979 & ~n11980 ) ;
  assign n11982 = ( x94 & n11976 ) | ( x94 & ~n11981 ) | ( n11976 & ~n11981 ) ;
  assign n11983 = ( x94 & n11609 ) | ( x94 & ~n11803 ) | ( n11609 & ~n11803 ) ;
  assign n11984 = x94 & n11609 ;
  assign n11985 = ( n11614 & n11983 ) | ( n11614 & n11984 ) | ( n11983 & n11984 ) ;
  assign n11986 = ( ~n11614 & n11983 ) | ( ~n11614 & n11984 ) | ( n11983 & n11984 ) ;
  assign n11987 = ( n11614 & ~n11985 ) | ( n11614 & n11986 ) | ( ~n11985 & n11986 ) ;
  assign n11988 = ( x95 & n11982 ) | ( x95 & ~n11987 ) | ( n11982 & ~n11987 ) ;
  assign n11989 = ( x95 & n11615 ) | ( x95 & ~n11803 ) | ( n11615 & ~n11803 ) ;
  assign n11990 = x95 & n11615 ;
  assign n11991 = ( ~n11620 & n11989 ) | ( ~n11620 & n11990 ) | ( n11989 & n11990 ) ;
  assign n11992 = ( n11620 & n11989 ) | ( n11620 & n11990 ) | ( n11989 & n11990 ) ;
  assign n11993 = ( n11620 & n11991 ) | ( n11620 & ~n11992 ) | ( n11991 & ~n11992 ) ;
  assign n11994 = ( x96 & n11988 ) | ( x96 & ~n11993 ) | ( n11988 & ~n11993 ) ;
  assign n11995 = ( x96 & n11621 ) | ( x96 & ~n11803 ) | ( n11621 & ~n11803 ) ;
  assign n11996 = x96 & n11621 ;
  assign n11997 = ( n11626 & n11995 ) | ( n11626 & n11996 ) | ( n11995 & n11996 ) ;
  assign n11998 = ( ~n11626 & n11995 ) | ( ~n11626 & n11996 ) | ( n11995 & n11996 ) ;
  assign n11999 = ( n11626 & ~n11997 ) | ( n11626 & n11998 ) | ( ~n11997 & n11998 ) ;
  assign n12000 = ( x97 & n11994 ) | ( x97 & ~n11999 ) | ( n11994 & ~n11999 ) ;
  assign n12001 = ( x97 & n11627 ) | ( x97 & ~n11803 ) | ( n11627 & ~n11803 ) ;
  assign n12002 = x97 & n11627 ;
  assign n12003 = ( ~n11632 & n12001 ) | ( ~n11632 & n12002 ) | ( n12001 & n12002 ) ;
  assign n12004 = ( n11632 & n12001 ) | ( n11632 & n12002 ) | ( n12001 & n12002 ) ;
  assign n12005 = ( n11632 & n12003 ) | ( n11632 & ~n12004 ) | ( n12003 & ~n12004 ) ;
  assign n12006 = ( x98 & n12000 ) | ( x98 & ~n12005 ) | ( n12000 & ~n12005 ) ;
  assign n12007 = ( x98 & n11633 ) | ( x98 & ~n11803 ) | ( n11633 & ~n11803 ) ;
  assign n12008 = x98 & n11633 ;
  assign n12009 = ( n11638 & n12007 ) | ( n11638 & n12008 ) | ( n12007 & n12008 ) ;
  assign n12010 = ( ~n11638 & n12007 ) | ( ~n11638 & n12008 ) | ( n12007 & n12008 ) ;
  assign n12011 = ( n11638 & ~n12009 ) | ( n11638 & n12010 ) | ( ~n12009 & n12010 ) ;
  assign n12012 = ( x99 & n12006 ) | ( x99 & ~n12011 ) | ( n12006 & ~n12011 ) ;
  assign n12013 = ( x99 & n11639 ) | ( x99 & ~n11803 ) | ( n11639 & ~n11803 ) ;
  assign n12014 = x99 & n11639 ;
  assign n12015 = ( ~n11644 & n12013 ) | ( ~n11644 & n12014 ) | ( n12013 & n12014 ) ;
  assign n12016 = ( n11644 & n12013 ) | ( n11644 & n12014 ) | ( n12013 & n12014 ) ;
  assign n12017 = ( n11644 & n12015 ) | ( n11644 & ~n12016 ) | ( n12015 & ~n12016 ) ;
  assign n12018 = ( x100 & n12012 ) | ( x100 & ~n12017 ) | ( n12012 & ~n12017 ) ;
  assign n12019 = ( x100 & n11645 ) | ( x100 & ~n11803 ) | ( n11645 & ~n11803 ) ;
  assign n12020 = x100 & n11645 ;
  assign n12021 = ( n11650 & n12019 ) | ( n11650 & n12020 ) | ( n12019 & n12020 ) ;
  assign n12022 = ( ~n11650 & n12019 ) | ( ~n11650 & n12020 ) | ( n12019 & n12020 ) ;
  assign n12023 = ( n11650 & ~n12021 ) | ( n11650 & n12022 ) | ( ~n12021 & n12022 ) ;
  assign n12024 = ( x101 & n12018 ) | ( x101 & ~n12023 ) | ( n12018 & ~n12023 ) ;
  assign n12025 = ( x101 & n11651 ) | ( x101 & ~n11803 ) | ( n11651 & ~n11803 ) ;
  assign n12026 = x101 & n11651 ;
  assign n12027 = ( ~n11656 & n12025 ) | ( ~n11656 & n12026 ) | ( n12025 & n12026 ) ;
  assign n12028 = ( n11656 & n12025 ) | ( n11656 & n12026 ) | ( n12025 & n12026 ) ;
  assign n12029 = ( n11656 & n12027 ) | ( n11656 & ~n12028 ) | ( n12027 & ~n12028 ) ;
  assign n12030 = ( x102 & n12024 ) | ( x102 & ~n12029 ) | ( n12024 & ~n12029 ) ;
  assign n12031 = ( x102 & n11657 ) | ( x102 & ~n11803 ) | ( n11657 & ~n11803 ) ;
  assign n12032 = x102 & n11657 ;
  assign n12033 = ( n11662 & n12031 ) | ( n11662 & n12032 ) | ( n12031 & n12032 ) ;
  assign n12034 = ( ~n11662 & n12031 ) | ( ~n11662 & n12032 ) | ( n12031 & n12032 ) ;
  assign n12035 = ( n11662 & ~n12033 ) | ( n11662 & n12034 ) | ( ~n12033 & n12034 ) ;
  assign n12036 = ( x103 & n12030 ) | ( x103 & ~n12035 ) | ( n12030 & ~n12035 ) ;
  assign n12037 = ( x103 & n11663 ) | ( x103 & ~n11803 ) | ( n11663 & ~n11803 ) ;
  assign n12038 = x103 & n11663 ;
  assign n12039 = ( ~n11668 & n12037 ) | ( ~n11668 & n12038 ) | ( n12037 & n12038 ) ;
  assign n12040 = ( n11668 & n12037 ) | ( n11668 & n12038 ) | ( n12037 & n12038 ) ;
  assign n12041 = ( n11668 & n12039 ) | ( n11668 & ~n12040 ) | ( n12039 & ~n12040 ) ;
  assign n12042 = ( x104 & n12036 ) | ( x104 & ~n12041 ) | ( n12036 & ~n12041 ) ;
  assign n12043 = ( x104 & n11669 ) | ( x104 & ~n11803 ) | ( n11669 & ~n11803 ) ;
  assign n12044 = x104 & n11669 ;
  assign n12045 = ( n11674 & n12043 ) | ( n11674 & n12044 ) | ( n12043 & n12044 ) ;
  assign n12046 = ( ~n11674 & n12043 ) | ( ~n11674 & n12044 ) | ( n12043 & n12044 ) ;
  assign n12047 = ( n11674 & ~n12045 ) | ( n11674 & n12046 ) | ( ~n12045 & n12046 ) ;
  assign n12048 = ( x105 & n12042 ) | ( x105 & ~n12047 ) | ( n12042 & ~n12047 ) ;
  assign n12049 = ( x105 & n11675 ) | ( x105 & ~n11803 ) | ( n11675 & ~n11803 ) ;
  assign n12050 = x105 & n11675 ;
  assign n12051 = ( ~n11680 & n12049 ) | ( ~n11680 & n12050 ) | ( n12049 & n12050 ) ;
  assign n12052 = ( n11680 & n12049 ) | ( n11680 & n12050 ) | ( n12049 & n12050 ) ;
  assign n12053 = ( n11680 & n12051 ) | ( n11680 & ~n12052 ) | ( n12051 & ~n12052 ) ;
  assign n12054 = ( x106 & n12048 ) | ( x106 & ~n12053 ) | ( n12048 & ~n12053 ) ;
  assign n12055 = ( x106 & n11681 ) | ( x106 & ~n11803 ) | ( n11681 & ~n11803 ) ;
  assign n12056 = x106 & n11681 ;
  assign n12057 = ( n11686 & n12055 ) | ( n11686 & n12056 ) | ( n12055 & n12056 ) ;
  assign n12058 = ( ~n11686 & n12055 ) | ( ~n11686 & n12056 ) | ( n12055 & n12056 ) ;
  assign n12059 = ( n11686 & ~n12057 ) | ( n11686 & n12058 ) | ( ~n12057 & n12058 ) ;
  assign n12060 = ( x107 & n12054 ) | ( x107 & ~n12059 ) | ( n12054 & ~n12059 ) ;
  assign n12061 = ( x107 & n11687 ) | ( x107 & ~n11803 ) | ( n11687 & ~n11803 ) ;
  assign n12062 = x107 & n11687 ;
  assign n12063 = ( ~n11692 & n12061 ) | ( ~n11692 & n12062 ) | ( n12061 & n12062 ) ;
  assign n12064 = ( n11692 & n12061 ) | ( n11692 & n12062 ) | ( n12061 & n12062 ) ;
  assign n12065 = ( n11692 & n12063 ) | ( n11692 & ~n12064 ) | ( n12063 & ~n12064 ) ;
  assign n12066 = ( x108 & n12060 ) | ( x108 & ~n12065 ) | ( n12060 & ~n12065 ) ;
  assign n12067 = ( x108 & n11693 ) | ( x108 & ~n11803 ) | ( n11693 & ~n11803 ) ;
  assign n12068 = x108 & n11693 ;
  assign n12069 = ( n11698 & n12067 ) | ( n11698 & n12068 ) | ( n12067 & n12068 ) ;
  assign n12070 = ( ~n11698 & n12067 ) | ( ~n11698 & n12068 ) | ( n12067 & n12068 ) ;
  assign n12071 = ( n11698 & ~n12069 ) | ( n11698 & n12070 ) | ( ~n12069 & n12070 ) ;
  assign n12072 = ( x109 & n12066 ) | ( x109 & ~n12071 ) | ( n12066 & ~n12071 ) ;
  assign n12073 = ( x109 & n11699 ) | ( x109 & ~n11803 ) | ( n11699 & ~n11803 ) ;
  assign n12074 = x109 & n11699 ;
  assign n12075 = ( ~n11704 & n12073 ) | ( ~n11704 & n12074 ) | ( n12073 & n12074 ) ;
  assign n12076 = ( n11704 & n12073 ) | ( n11704 & n12074 ) | ( n12073 & n12074 ) ;
  assign n12077 = ( n11704 & n12075 ) | ( n11704 & ~n12076 ) | ( n12075 & ~n12076 ) ;
  assign n12078 = ( x110 & n12072 ) | ( x110 & ~n12077 ) | ( n12072 & ~n12077 ) ;
  assign n12079 = ( x110 & n11705 ) | ( x110 & ~n11803 ) | ( n11705 & ~n11803 ) ;
  assign n12080 = x110 & n11705 ;
  assign n12081 = ( n11710 & n12079 ) | ( n11710 & n12080 ) | ( n12079 & n12080 ) ;
  assign n12082 = ( ~n11710 & n12079 ) | ( ~n11710 & n12080 ) | ( n12079 & n12080 ) ;
  assign n12083 = ( n11710 & ~n12081 ) | ( n11710 & n12082 ) | ( ~n12081 & n12082 ) ;
  assign n12084 = ( x111 & n12078 ) | ( x111 & ~n12083 ) | ( n12078 & ~n12083 ) ;
  assign n12085 = ( x111 & n11711 ) | ( x111 & ~n11803 ) | ( n11711 & ~n11803 ) ;
  assign n12086 = x111 & n11711 ;
  assign n12087 = ( ~n11716 & n12085 ) | ( ~n11716 & n12086 ) | ( n12085 & n12086 ) ;
  assign n12088 = ( n11716 & n12085 ) | ( n11716 & n12086 ) | ( n12085 & n12086 ) ;
  assign n12089 = ( n11716 & n12087 ) | ( n11716 & ~n12088 ) | ( n12087 & ~n12088 ) ;
  assign n12090 = ( x112 & n12084 ) | ( x112 & ~n12089 ) | ( n12084 & ~n12089 ) ;
  assign n12091 = ( x112 & n11717 ) | ( x112 & ~n11803 ) | ( n11717 & ~n11803 ) ;
  assign n12092 = x112 & n11717 ;
  assign n12093 = ( n11722 & n12091 ) | ( n11722 & n12092 ) | ( n12091 & n12092 ) ;
  assign n12094 = ( ~n11722 & n12091 ) | ( ~n11722 & n12092 ) | ( n12091 & n12092 ) ;
  assign n12095 = ( n11722 & ~n12093 ) | ( n11722 & n12094 ) | ( ~n12093 & n12094 ) ;
  assign n12096 = ( x113 & n12090 ) | ( x113 & ~n12095 ) | ( n12090 & ~n12095 ) ;
  assign n12097 = ( x113 & n11723 ) | ( x113 & ~n11803 ) | ( n11723 & ~n11803 ) ;
  assign n12098 = x113 & n11723 ;
  assign n12099 = ( ~n11728 & n12097 ) | ( ~n11728 & n12098 ) | ( n12097 & n12098 ) ;
  assign n12100 = ( n11728 & n12097 ) | ( n11728 & n12098 ) | ( n12097 & n12098 ) ;
  assign n12101 = ( n11728 & n12099 ) | ( n11728 & ~n12100 ) | ( n12099 & ~n12100 ) ;
  assign n12102 = ( x114 & n12096 ) | ( x114 & ~n12101 ) | ( n12096 & ~n12101 ) ;
  assign n12103 = ( x114 & n11729 ) | ( x114 & ~n11803 ) | ( n11729 & ~n11803 ) ;
  assign n12104 = x114 & n11729 ;
  assign n12105 = ( n11734 & n12103 ) | ( n11734 & n12104 ) | ( n12103 & n12104 ) ;
  assign n12106 = ( ~n11734 & n12103 ) | ( ~n11734 & n12104 ) | ( n12103 & n12104 ) ;
  assign n12107 = ( n11734 & ~n12105 ) | ( n11734 & n12106 ) | ( ~n12105 & n12106 ) ;
  assign n12108 = ( x115 & n12102 ) | ( x115 & ~n12107 ) | ( n12102 & ~n12107 ) ;
  assign n12109 = ( x115 & n11735 ) | ( x115 & ~n11803 ) | ( n11735 & ~n11803 ) ;
  assign n12110 = x115 & n11735 ;
  assign n12111 = ( ~n11740 & n12109 ) | ( ~n11740 & n12110 ) | ( n12109 & n12110 ) ;
  assign n12112 = ( n11740 & n12109 ) | ( n11740 & n12110 ) | ( n12109 & n12110 ) ;
  assign n12113 = ( n11740 & n12111 ) | ( n11740 & ~n12112 ) | ( n12111 & ~n12112 ) ;
  assign n12114 = ( x116 & n12108 ) | ( x116 & ~n12113 ) | ( n12108 & ~n12113 ) ;
  assign n12115 = ( x116 & n11741 ) | ( x116 & ~n11803 ) | ( n11741 & ~n11803 ) ;
  assign n12116 = x116 & n11741 ;
  assign n12117 = ( n11746 & n12115 ) | ( n11746 & n12116 ) | ( n12115 & n12116 ) ;
  assign n12118 = ( ~n11746 & n12115 ) | ( ~n11746 & n12116 ) | ( n12115 & n12116 ) ;
  assign n12119 = ( n11746 & ~n12117 ) | ( n11746 & n12118 ) | ( ~n12117 & n12118 ) ;
  assign n12120 = ( x117 & n12114 ) | ( x117 & ~n12119 ) | ( n12114 & ~n12119 ) ;
  assign n12121 = ( x117 & n11747 ) | ( x117 & ~n11803 ) | ( n11747 & ~n11803 ) ;
  assign n12122 = x117 & n11747 ;
  assign n12123 = ( ~n11752 & n12121 ) | ( ~n11752 & n12122 ) | ( n12121 & n12122 ) ;
  assign n12124 = ( n11752 & n12121 ) | ( n11752 & n12122 ) | ( n12121 & n12122 ) ;
  assign n12125 = ( n11752 & n12123 ) | ( n11752 & ~n12124 ) | ( n12123 & ~n12124 ) ;
  assign n12126 = ( x118 & n12120 ) | ( x118 & ~n12125 ) | ( n12120 & ~n12125 ) ;
  assign n12127 = ( x118 & n11753 ) | ( x118 & ~n11803 ) | ( n11753 & ~n11803 ) ;
  assign n12128 = x118 & n11753 ;
  assign n12129 = ( n11758 & n12127 ) | ( n11758 & n12128 ) | ( n12127 & n12128 ) ;
  assign n12130 = ( ~n11758 & n12127 ) | ( ~n11758 & n12128 ) | ( n12127 & n12128 ) ;
  assign n12131 = ( n11758 & ~n12129 ) | ( n11758 & n12130 ) | ( ~n12129 & n12130 ) ;
  assign n12132 = ( x119 & n12126 ) | ( x119 & ~n12131 ) | ( n12126 & ~n12131 ) ;
  assign n12133 = ( x119 & n11759 ) | ( x119 & ~n11803 ) | ( n11759 & ~n11803 ) ;
  assign n12134 = x119 & n11759 ;
  assign n12135 = ( ~n11764 & n12133 ) | ( ~n11764 & n12134 ) | ( n12133 & n12134 ) ;
  assign n12136 = ( n11764 & n12133 ) | ( n11764 & n12134 ) | ( n12133 & n12134 ) ;
  assign n12137 = ( n11764 & n12135 ) | ( n11764 & ~n12136 ) | ( n12135 & ~n12136 ) ;
  assign n12138 = ( x120 & n12132 ) | ( x120 & ~n12137 ) | ( n12132 & ~n12137 ) ;
  assign n12139 = ( x120 & n11765 ) | ( x120 & ~n11803 ) | ( n11765 & ~n11803 ) ;
  assign n12140 = x120 & n11765 ;
  assign n12141 = ( n11770 & n12139 ) | ( n11770 & n12140 ) | ( n12139 & n12140 ) ;
  assign n12142 = ( ~n11770 & n12139 ) | ( ~n11770 & n12140 ) | ( n12139 & n12140 ) ;
  assign n12143 = ( n11770 & ~n12141 ) | ( n11770 & n12142 ) | ( ~n12141 & n12142 ) ;
  assign n12144 = ( x121 & n12138 ) | ( x121 & ~n12143 ) | ( n12138 & ~n12143 ) ;
  assign n12145 = ( x121 & n11771 ) | ( x121 & ~n11803 ) | ( n11771 & ~n11803 ) ;
  assign n12146 = x121 & n11771 ;
  assign n12147 = ( ~n11776 & n12145 ) | ( ~n11776 & n12146 ) | ( n12145 & n12146 ) ;
  assign n12148 = ( n11776 & n12145 ) | ( n11776 & n12146 ) | ( n12145 & n12146 ) ;
  assign n12149 = ( n11776 & n12147 ) | ( n11776 & ~n12148 ) | ( n12147 & ~n12148 ) ;
  assign n12150 = ( x122 & n12144 ) | ( x122 & ~n12149 ) | ( n12144 & ~n12149 ) ;
  assign n12151 = ( x122 & n11777 ) | ( x122 & ~n11803 ) | ( n11777 & ~n11803 ) ;
  assign n12152 = x122 & n11777 ;
  assign n12153 = ( n11782 & n12151 ) | ( n11782 & n12152 ) | ( n12151 & n12152 ) ;
  assign n12154 = ( ~n11782 & n12151 ) | ( ~n11782 & n12152 ) | ( n12151 & n12152 ) ;
  assign n12155 = ( n11782 & ~n12153 ) | ( n11782 & n12154 ) | ( ~n12153 & n12154 ) ;
  assign n12156 = ( x123 & n12150 ) | ( x123 & ~n12155 ) | ( n12150 & ~n12155 ) ;
  assign n12157 = ( x123 & n11783 ) | ( x123 & ~n11803 ) | ( n11783 & ~n11803 ) ;
  assign n12158 = x123 & n11783 ;
  assign n12159 = ( ~n11788 & n12157 ) | ( ~n11788 & n12158 ) | ( n12157 & n12158 ) ;
  assign n12160 = ( n11788 & n12157 ) | ( n11788 & n12158 ) | ( n12157 & n12158 ) ;
  assign n12161 = ( n11788 & n12159 ) | ( n11788 & ~n12160 ) | ( n12159 & ~n12160 ) ;
  assign n12162 = ( x124 & n12156 ) | ( x124 & ~n12161 ) | ( n12156 & ~n12161 ) ;
  assign n12163 = ( x124 & n11789 ) | ( x124 & ~n11803 ) | ( n11789 & ~n11803 ) ;
  assign n12164 = x124 & n11789 ;
  assign n12165 = ( n11794 & n12163 ) | ( n11794 & n12164 ) | ( n12163 & n12164 ) ;
  assign n12166 = ( ~n11794 & n12163 ) | ( ~n11794 & n12164 ) | ( n12163 & n12164 ) ;
  assign n12167 = ( n11794 & ~n12165 ) | ( n11794 & n12166 ) | ( ~n12165 & n12166 ) ;
  assign n12168 = ( x125 & n12162 ) | ( x125 & ~n12167 ) | ( n12162 & ~n12167 ) ;
  assign n12169 = ( x125 & n11795 ) | ( x125 & ~n11803 ) | ( n11795 & ~n11803 ) ;
  assign n12170 = x125 & n11795 ;
  assign n12171 = ( n11800 & n12169 ) | ( n11800 & n12170 ) | ( n12169 & n12170 ) ;
  assign n12172 = ( ~n11800 & n12169 ) | ( ~n11800 & n12170 ) | ( n12169 & n12170 ) ;
  assign n12173 = ( n11800 & ~n12171 ) | ( n11800 & n12172 ) | ( ~n12171 & n12172 ) ;
  assign n12174 = ( x126 & n12168 ) | ( x126 & ~n12173 ) | ( n12168 & ~n12173 ) ;
  assign n12175 = x126 | n11801 ;
  assign n12176 = ( x126 & x127 ) | ( x126 & n11801 ) | ( x127 & n11801 ) ;
  assign n12177 = ( n11435 & ~n12175 ) | ( n11435 & n12176 ) | ( ~n12175 & n12176 ) ;
  assign n12178 = ( x127 & n12174 ) | ( x127 & ~n12177 ) | ( n12174 & ~n12177 ) ;
  assign n12179 = ~x63 & x64 ;
  assign n12180 = n197 | n12179 ;
  assign n12181 = ( x0 & ~x64 ) | ( x0 & n12178 ) | ( ~x64 & n12178 ) ;
  assign n12182 = ~x0 & n12178 ;
  assign n12183 = ( n11807 & n12181 ) | ( n11807 & ~n12182 ) | ( n12181 & ~n12182 ) ;
  assign n12184 = ( x65 & n11807 ) | ( x65 & ~n12178 ) | ( n11807 & ~n12178 ) ;
  assign n12185 = x65 & n11807 ;
  assign n12186 = ( n11806 & n12184 ) | ( n11806 & n12185 ) | ( n12184 & n12185 ) ;
  assign n12187 = ( ~n11806 & n12184 ) | ( ~n11806 & n12185 ) | ( n12184 & n12185 ) ;
  assign n12188 = ( n11806 & ~n12186 ) | ( n11806 & n12187 ) | ( ~n12186 & n12187 ) ;
  assign n12189 = ( x66 & n11808 ) | ( x66 & ~n12178 ) | ( n11808 & ~n12178 ) ;
  assign n12190 = x66 & n11808 ;
  assign n12191 = ( n11813 & n12189 ) | ( n11813 & n12190 ) | ( n12189 & n12190 ) ;
  assign n12192 = ( ~n11813 & n12189 ) | ( ~n11813 & n12190 ) | ( n12189 & n12190 ) ;
  assign n12193 = ( n11813 & ~n12191 ) | ( n11813 & n12192 ) | ( ~n12191 & n12192 ) ;
  assign n12194 = ( x67 & n11814 ) | ( x67 & ~n12178 ) | ( n11814 & ~n12178 ) ;
  assign n12195 = x67 & n11814 ;
  assign n12196 = ( ~n11819 & n12194 ) | ( ~n11819 & n12195 ) | ( n12194 & n12195 ) ;
  assign n12197 = ( n11819 & n12194 ) | ( n11819 & n12195 ) | ( n12194 & n12195 ) ;
  assign n12198 = ( n11819 & n12196 ) | ( n11819 & ~n12197 ) | ( n12196 & ~n12197 ) ;
  assign n12199 = ( x68 & n11820 ) | ( x68 & ~n12178 ) | ( n11820 & ~n12178 ) ;
  assign n12200 = x68 & n11820 ;
  assign n12201 = ( n11825 & n12199 ) | ( n11825 & n12200 ) | ( n12199 & n12200 ) ;
  assign n12202 = ( ~n11825 & n12199 ) | ( ~n11825 & n12200 ) | ( n12199 & n12200 ) ;
  assign n12203 = ( n11825 & ~n12201 ) | ( n11825 & n12202 ) | ( ~n12201 & n12202 ) ;
  assign n12204 = ( x69 & n11826 ) | ( x69 & ~n12178 ) | ( n11826 & ~n12178 ) ;
  assign n12205 = x69 & n11826 ;
  assign n12206 = ( ~n11831 & n12204 ) | ( ~n11831 & n12205 ) | ( n12204 & n12205 ) ;
  assign n12207 = ( n11831 & n12204 ) | ( n11831 & n12205 ) | ( n12204 & n12205 ) ;
  assign n12208 = ( n11831 & n12206 ) | ( n11831 & ~n12207 ) | ( n12206 & ~n12207 ) ;
  assign n12209 = ( x70 & n11832 ) | ( x70 & ~n12178 ) | ( n11832 & ~n12178 ) ;
  assign n12210 = x70 & n11832 ;
  assign n12211 = ( n11837 & n12209 ) | ( n11837 & n12210 ) | ( n12209 & n12210 ) ;
  assign n12212 = ( ~n11837 & n12209 ) | ( ~n11837 & n12210 ) | ( n12209 & n12210 ) ;
  assign n12213 = ( n11837 & ~n12211 ) | ( n11837 & n12212 ) | ( ~n12211 & n12212 ) ;
  assign n12214 = ( x71 & n11838 ) | ( x71 & ~n12178 ) | ( n11838 & ~n12178 ) ;
  assign n12215 = x71 & n11838 ;
  assign n12216 = ( ~n11843 & n12214 ) | ( ~n11843 & n12215 ) | ( n12214 & n12215 ) ;
  assign n12217 = ( n11843 & n12214 ) | ( n11843 & n12215 ) | ( n12214 & n12215 ) ;
  assign n12218 = ( n11843 & n12216 ) | ( n11843 & ~n12217 ) | ( n12216 & ~n12217 ) ;
  assign n12219 = ( x72 & n11844 ) | ( x72 & ~n12178 ) | ( n11844 & ~n12178 ) ;
  assign n12220 = x72 & n11844 ;
  assign n12221 = ( n11849 & n12219 ) | ( n11849 & n12220 ) | ( n12219 & n12220 ) ;
  assign n12222 = ( ~n11849 & n12219 ) | ( ~n11849 & n12220 ) | ( n12219 & n12220 ) ;
  assign n12223 = ( n11849 & ~n12221 ) | ( n11849 & n12222 ) | ( ~n12221 & n12222 ) ;
  assign n12224 = ( x73 & n11850 ) | ( x73 & ~n12178 ) | ( n11850 & ~n12178 ) ;
  assign n12225 = x73 & n11850 ;
  assign n12226 = ( ~n11855 & n12224 ) | ( ~n11855 & n12225 ) | ( n12224 & n12225 ) ;
  assign n12227 = ( n11855 & n12224 ) | ( n11855 & n12225 ) | ( n12224 & n12225 ) ;
  assign n12228 = ( n11855 & n12226 ) | ( n11855 & ~n12227 ) | ( n12226 & ~n12227 ) ;
  assign n12229 = ( x74 & n11856 ) | ( x74 & ~n12178 ) | ( n11856 & ~n12178 ) ;
  assign n12230 = x74 & n11856 ;
  assign n12231 = ( n11861 & n12229 ) | ( n11861 & n12230 ) | ( n12229 & n12230 ) ;
  assign n12232 = ( ~n11861 & n12229 ) | ( ~n11861 & n12230 ) | ( n12229 & n12230 ) ;
  assign n12233 = ( n11861 & ~n12231 ) | ( n11861 & n12232 ) | ( ~n12231 & n12232 ) ;
  assign n12234 = ( x75 & n11862 ) | ( x75 & ~n12178 ) | ( n11862 & ~n12178 ) ;
  assign n12235 = x75 & n11862 ;
  assign n12236 = ( ~n11867 & n12234 ) | ( ~n11867 & n12235 ) | ( n12234 & n12235 ) ;
  assign n12237 = ( n11867 & n12234 ) | ( n11867 & n12235 ) | ( n12234 & n12235 ) ;
  assign n12238 = ( n11867 & n12236 ) | ( n11867 & ~n12237 ) | ( n12236 & ~n12237 ) ;
  assign n12239 = ( x76 & n11868 ) | ( x76 & ~n12178 ) | ( n11868 & ~n12178 ) ;
  assign n12240 = x76 & n11868 ;
  assign n12241 = ( n11873 & n12239 ) | ( n11873 & n12240 ) | ( n12239 & n12240 ) ;
  assign n12242 = ( ~n11873 & n12239 ) | ( ~n11873 & n12240 ) | ( n12239 & n12240 ) ;
  assign n12243 = ( n11873 & ~n12241 ) | ( n11873 & n12242 ) | ( ~n12241 & n12242 ) ;
  assign n12244 = ( x77 & n11874 ) | ( x77 & ~n12178 ) | ( n11874 & ~n12178 ) ;
  assign n12245 = x77 & n11874 ;
  assign n12246 = ( ~n11879 & n12244 ) | ( ~n11879 & n12245 ) | ( n12244 & n12245 ) ;
  assign n12247 = ( n11879 & n12244 ) | ( n11879 & n12245 ) | ( n12244 & n12245 ) ;
  assign n12248 = ( n11879 & n12246 ) | ( n11879 & ~n12247 ) | ( n12246 & ~n12247 ) ;
  assign n12249 = ( x78 & n11880 ) | ( x78 & ~n12178 ) | ( n11880 & ~n12178 ) ;
  assign n12250 = x78 & n11880 ;
  assign n12251 = ( n11885 & n12249 ) | ( n11885 & n12250 ) | ( n12249 & n12250 ) ;
  assign n12252 = ( ~n11885 & n12249 ) | ( ~n11885 & n12250 ) | ( n12249 & n12250 ) ;
  assign n12253 = ( n11885 & ~n12251 ) | ( n11885 & n12252 ) | ( ~n12251 & n12252 ) ;
  assign n12254 = ( x79 & n11886 ) | ( x79 & ~n12178 ) | ( n11886 & ~n12178 ) ;
  assign n12255 = x79 & n11886 ;
  assign n12256 = ( ~n11891 & n12254 ) | ( ~n11891 & n12255 ) | ( n12254 & n12255 ) ;
  assign n12257 = ( n11891 & n12254 ) | ( n11891 & n12255 ) | ( n12254 & n12255 ) ;
  assign n12258 = ( n11891 & n12256 ) | ( n11891 & ~n12257 ) | ( n12256 & ~n12257 ) ;
  assign n12259 = ( x80 & n11892 ) | ( x80 & ~n12178 ) | ( n11892 & ~n12178 ) ;
  assign n12260 = x80 & n11892 ;
  assign n12261 = ( n11897 & n12259 ) | ( n11897 & n12260 ) | ( n12259 & n12260 ) ;
  assign n12262 = ( ~n11897 & n12259 ) | ( ~n11897 & n12260 ) | ( n12259 & n12260 ) ;
  assign n12263 = ( n11897 & ~n12261 ) | ( n11897 & n12262 ) | ( ~n12261 & n12262 ) ;
  assign n12264 = ( x81 & n11898 ) | ( x81 & ~n12178 ) | ( n11898 & ~n12178 ) ;
  assign n12265 = x81 & n11898 ;
  assign n12266 = ( ~n11903 & n12264 ) | ( ~n11903 & n12265 ) | ( n12264 & n12265 ) ;
  assign n12267 = ( n11903 & n12264 ) | ( n11903 & n12265 ) | ( n12264 & n12265 ) ;
  assign n12268 = ( n11903 & n12266 ) | ( n11903 & ~n12267 ) | ( n12266 & ~n12267 ) ;
  assign n12269 = ( x82 & n11904 ) | ( x82 & ~n12178 ) | ( n11904 & ~n12178 ) ;
  assign n12270 = x82 & n11904 ;
  assign n12271 = ( n11909 & n12269 ) | ( n11909 & n12270 ) | ( n12269 & n12270 ) ;
  assign n12272 = ( ~n11909 & n12269 ) | ( ~n11909 & n12270 ) | ( n12269 & n12270 ) ;
  assign n12273 = ( n11909 & ~n12271 ) | ( n11909 & n12272 ) | ( ~n12271 & n12272 ) ;
  assign n12274 = ( x83 & n11910 ) | ( x83 & ~n12178 ) | ( n11910 & ~n12178 ) ;
  assign n12275 = x83 & n11910 ;
  assign n12276 = ( ~n11915 & n12274 ) | ( ~n11915 & n12275 ) | ( n12274 & n12275 ) ;
  assign n12277 = ( n11915 & n12274 ) | ( n11915 & n12275 ) | ( n12274 & n12275 ) ;
  assign n12278 = ( n11915 & n12276 ) | ( n11915 & ~n12277 ) | ( n12276 & ~n12277 ) ;
  assign n12279 = ( x84 & n11916 ) | ( x84 & ~n12178 ) | ( n11916 & ~n12178 ) ;
  assign n12280 = x84 & n11916 ;
  assign n12281 = ( n11921 & n12279 ) | ( n11921 & n12280 ) | ( n12279 & n12280 ) ;
  assign n12282 = ( ~n11921 & n12279 ) | ( ~n11921 & n12280 ) | ( n12279 & n12280 ) ;
  assign n12283 = ( n11921 & ~n12281 ) | ( n11921 & n12282 ) | ( ~n12281 & n12282 ) ;
  assign n12284 = ( x85 & n11922 ) | ( x85 & ~n12178 ) | ( n11922 & ~n12178 ) ;
  assign n12285 = x85 & n11922 ;
  assign n12286 = ( ~n11927 & n12284 ) | ( ~n11927 & n12285 ) | ( n12284 & n12285 ) ;
  assign n12287 = ( n11927 & n12284 ) | ( n11927 & n12285 ) | ( n12284 & n12285 ) ;
  assign n12288 = ( n11927 & n12286 ) | ( n11927 & ~n12287 ) | ( n12286 & ~n12287 ) ;
  assign n12289 = ( x86 & n11928 ) | ( x86 & ~n12178 ) | ( n11928 & ~n12178 ) ;
  assign n12290 = x86 & n11928 ;
  assign n12291 = ( n11933 & n12289 ) | ( n11933 & n12290 ) | ( n12289 & n12290 ) ;
  assign n12292 = ( ~n11933 & n12289 ) | ( ~n11933 & n12290 ) | ( n12289 & n12290 ) ;
  assign n12293 = ( n11933 & ~n12291 ) | ( n11933 & n12292 ) | ( ~n12291 & n12292 ) ;
  assign n12294 = ( x87 & n11934 ) | ( x87 & ~n12178 ) | ( n11934 & ~n12178 ) ;
  assign n12295 = x87 & n11934 ;
  assign n12296 = ( ~n11939 & n12294 ) | ( ~n11939 & n12295 ) | ( n12294 & n12295 ) ;
  assign n12297 = ( n11939 & n12294 ) | ( n11939 & n12295 ) | ( n12294 & n12295 ) ;
  assign n12298 = ( n11939 & n12296 ) | ( n11939 & ~n12297 ) | ( n12296 & ~n12297 ) ;
  assign n12299 = ( x88 & n11940 ) | ( x88 & ~n12178 ) | ( n11940 & ~n12178 ) ;
  assign n12300 = x88 & n11940 ;
  assign n12301 = ( n11945 & n12299 ) | ( n11945 & n12300 ) | ( n12299 & n12300 ) ;
  assign n12302 = ( ~n11945 & n12299 ) | ( ~n11945 & n12300 ) | ( n12299 & n12300 ) ;
  assign n12303 = ( n11945 & ~n12301 ) | ( n11945 & n12302 ) | ( ~n12301 & n12302 ) ;
  assign n12304 = ( x89 & n11946 ) | ( x89 & ~n12178 ) | ( n11946 & ~n12178 ) ;
  assign n12305 = x89 & n11946 ;
  assign n12306 = ( ~n11951 & n12304 ) | ( ~n11951 & n12305 ) | ( n12304 & n12305 ) ;
  assign n12307 = ( n11951 & n12304 ) | ( n11951 & n12305 ) | ( n12304 & n12305 ) ;
  assign n12308 = ( n11951 & n12306 ) | ( n11951 & ~n12307 ) | ( n12306 & ~n12307 ) ;
  assign n12309 = ( x90 & n11952 ) | ( x90 & ~n12178 ) | ( n11952 & ~n12178 ) ;
  assign n12310 = x90 & n11952 ;
  assign n12311 = ( n11957 & n12309 ) | ( n11957 & n12310 ) | ( n12309 & n12310 ) ;
  assign n12312 = ( ~n11957 & n12309 ) | ( ~n11957 & n12310 ) | ( n12309 & n12310 ) ;
  assign n12313 = ( n11957 & ~n12311 ) | ( n11957 & n12312 ) | ( ~n12311 & n12312 ) ;
  assign n12314 = ( x91 & n11958 ) | ( x91 & ~n12178 ) | ( n11958 & ~n12178 ) ;
  assign n12315 = x91 & n11958 ;
  assign n12316 = ( ~n11963 & n12314 ) | ( ~n11963 & n12315 ) | ( n12314 & n12315 ) ;
  assign n12317 = ( n11963 & n12314 ) | ( n11963 & n12315 ) | ( n12314 & n12315 ) ;
  assign n12318 = ( n11963 & n12316 ) | ( n11963 & ~n12317 ) | ( n12316 & ~n12317 ) ;
  assign n12319 = ( x92 & n11964 ) | ( x92 & ~n12178 ) | ( n11964 & ~n12178 ) ;
  assign n12320 = x92 & n11964 ;
  assign n12321 = ( n11969 & n12319 ) | ( n11969 & n12320 ) | ( n12319 & n12320 ) ;
  assign n12322 = ( ~n11969 & n12319 ) | ( ~n11969 & n12320 ) | ( n12319 & n12320 ) ;
  assign n12323 = ( n11969 & ~n12321 ) | ( n11969 & n12322 ) | ( ~n12321 & n12322 ) ;
  assign n12324 = ( x93 & n11970 ) | ( x93 & ~n12178 ) | ( n11970 & ~n12178 ) ;
  assign n12325 = x93 & n11970 ;
  assign n12326 = ( ~n11975 & n12324 ) | ( ~n11975 & n12325 ) | ( n12324 & n12325 ) ;
  assign n12327 = ( n11975 & n12324 ) | ( n11975 & n12325 ) | ( n12324 & n12325 ) ;
  assign n12328 = ( n11975 & n12326 ) | ( n11975 & ~n12327 ) | ( n12326 & ~n12327 ) ;
  assign n12329 = ( x94 & n11976 ) | ( x94 & ~n12178 ) | ( n11976 & ~n12178 ) ;
  assign n12330 = x94 & n11976 ;
  assign n12331 = ( n11981 & n12329 ) | ( n11981 & n12330 ) | ( n12329 & n12330 ) ;
  assign n12332 = ( ~n11981 & n12329 ) | ( ~n11981 & n12330 ) | ( n12329 & n12330 ) ;
  assign n12333 = ( n11981 & ~n12331 ) | ( n11981 & n12332 ) | ( ~n12331 & n12332 ) ;
  assign n12334 = ( x95 & n11982 ) | ( x95 & ~n12178 ) | ( n11982 & ~n12178 ) ;
  assign n12335 = x95 & n11982 ;
  assign n12336 = ( ~n11987 & n12334 ) | ( ~n11987 & n12335 ) | ( n12334 & n12335 ) ;
  assign n12337 = ( n11987 & n12334 ) | ( n11987 & n12335 ) | ( n12334 & n12335 ) ;
  assign n12338 = ( n11987 & n12336 ) | ( n11987 & ~n12337 ) | ( n12336 & ~n12337 ) ;
  assign n12339 = ( x96 & n11988 ) | ( x96 & ~n12178 ) | ( n11988 & ~n12178 ) ;
  assign n12340 = x96 & n11988 ;
  assign n12341 = ( n11993 & n12339 ) | ( n11993 & n12340 ) | ( n12339 & n12340 ) ;
  assign n12342 = ( ~n11993 & n12339 ) | ( ~n11993 & n12340 ) | ( n12339 & n12340 ) ;
  assign n12343 = ( n11993 & ~n12341 ) | ( n11993 & n12342 ) | ( ~n12341 & n12342 ) ;
  assign n12344 = ( x97 & n11994 ) | ( x97 & ~n12178 ) | ( n11994 & ~n12178 ) ;
  assign n12345 = x97 & n11994 ;
  assign n12346 = ( ~n11999 & n12344 ) | ( ~n11999 & n12345 ) | ( n12344 & n12345 ) ;
  assign n12347 = ( n11999 & n12344 ) | ( n11999 & n12345 ) | ( n12344 & n12345 ) ;
  assign n12348 = ( n11999 & n12346 ) | ( n11999 & ~n12347 ) | ( n12346 & ~n12347 ) ;
  assign n12349 = ( x98 & n12000 ) | ( x98 & ~n12178 ) | ( n12000 & ~n12178 ) ;
  assign n12350 = x98 & n12000 ;
  assign n12351 = ( n12005 & n12349 ) | ( n12005 & n12350 ) | ( n12349 & n12350 ) ;
  assign n12352 = ( ~n12005 & n12349 ) | ( ~n12005 & n12350 ) | ( n12349 & n12350 ) ;
  assign n12353 = ( n12005 & ~n12351 ) | ( n12005 & n12352 ) | ( ~n12351 & n12352 ) ;
  assign n12354 = ( x99 & n12006 ) | ( x99 & ~n12178 ) | ( n12006 & ~n12178 ) ;
  assign n12355 = x99 & n12006 ;
  assign n12356 = ( ~n12011 & n12354 ) | ( ~n12011 & n12355 ) | ( n12354 & n12355 ) ;
  assign n12357 = ( n12011 & n12354 ) | ( n12011 & n12355 ) | ( n12354 & n12355 ) ;
  assign n12358 = ( n12011 & n12356 ) | ( n12011 & ~n12357 ) | ( n12356 & ~n12357 ) ;
  assign n12359 = ( x100 & n12012 ) | ( x100 & ~n12178 ) | ( n12012 & ~n12178 ) ;
  assign n12360 = x100 & n12012 ;
  assign n12361 = ( n12017 & n12359 ) | ( n12017 & n12360 ) | ( n12359 & n12360 ) ;
  assign n12362 = ( ~n12017 & n12359 ) | ( ~n12017 & n12360 ) | ( n12359 & n12360 ) ;
  assign n12363 = ( n12017 & ~n12361 ) | ( n12017 & n12362 ) | ( ~n12361 & n12362 ) ;
  assign n12364 = ( x101 & n12018 ) | ( x101 & ~n12178 ) | ( n12018 & ~n12178 ) ;
  assign n12365 = x101 & n12018 ;
  assign n12366 = ( ~n12023 & n12364 ) | ( ~n12023 & n12365 ) | ( n12364 & n12365 ) ;
  assign n12367 = ( n12023 & n12364 ) | ( n12023 & n12365 ) | ( n12364 & n12365 ) ;
  assign n12368 = ( n12023 & n12366 ) | ( n12023 & ~n12367 ) | ( n12366 & ~n12367 ) ;
  assign n12369 = ( x102 & n12024 ) | ( x102 & ~n12178 ) | ( n12024 & ~n12178 ) ;
  assign n12370 = x102 & n12024 ;
  assign n12371 = ( n12029 & n12369 ) | ( n12029 & n12370 ) | ( n12369 & n12370 ) ;
  assign n12372 = ( ~n12029 & n12369 ) | ( ~n12029 & n12370 ) | ( n12369 & n12370 ) ;
  assign n12373 = ( n12029 & ~n12371 ) | ( n12029 & n12372 ) | ( ~n12371 & n12372 ) ;
  assign n12374 = ( x103 & n12030 ) | ( x103 & ~n12178 ) | ( n12030 & ~n12178 ) ;
  assign n12375 = x103 & n12030 ;
  assign n12376 = ( ~n12035 & n12374 ) | ( ~n12035 & n12375 ) | ( n12374 & n12375 ) ;
  assign n12377 = ( n12035 & n12374 ) | ( n12035 & n12375 ) | ( n12374 & n12375 ) ;
  assign n12378 = ( n12035 & n12376 ) | ( n12035 & ~n12377 ) | ( n12376 & ~n12377 ) ;
  assign n12379 = ( x104 & n12036 ) | ( x104 & ~n12178 ) | ( n12036 & ~n12178 ) ;
  assign n12380 = x104 & n12036 ;
  assign n12381 = ( n12041 & n12379 ) | ( n12041 & n12380 ) | ( n12379 & n12380 ) ;
  assign n12382 = ( ~n12041 & n12379 ) | ( ~n12041 & n12380 ) | ( n12379 & n12380 ) ;
  assign n12383 = ( n12041 & ~n12381 ) | ( n12041 & n12382 ) | ( ~n12381 & n12382 ) ;
  assign n12384 = ( x105 & n12042 ) | ( x105 & ~n12178 ) | ( n12042 & ~n12178 ) ;
  assign n12385 = x105 & n12042 ;
  assign n12386 = ( ~n12047 & n12384 ) | ( ~n12047 & n12385 ) | ( n12384 & n12385 ) ;
  assign n12387 = ( n12047 & n12384 ) | ( n12047 & n12385 ) | ( n12384 & n12385 ) ;
  assign n12388 = ( n12047 & n12386 ) | ( n12047 & ~n12387 ) | ( n12386 & ~n12387 ) ;
  assign n12389 = ( x106 & n12048 ) | ( x106 & ~n12178 ) | ( n12048 & ~n12178 ) ;
  assign n12390 = x106 & n12048 ;
  assign n12391 = ( n12053 & n12389 ) | ( n12053 & n12390 ) | ( n12389 & n12390 ) ;
  assign n12392 = ( ~n12053 & n12389 ) | ( ~n12053 & n12390 ) | ( n12389 & n12390 ) ;
  assign n12393 = ( n12053 & ~n12391 ) | ( n12053 & n12392 ) | ( ~n12391 & n12392 ) ;
  assign n12394 = ( x107 & n12054 ) | ( x107 & ~n12178 ) | ( n12054 & ~n12178 ) ;
  assign n12395 = x107 & n12054 ;
  assign n12396 = ( ~n12059 & n12394 ) | ( ~n12059 & n12395 ) | ( n12394 & n12395 ) ;
  assign n12397 = ( n12059 & n12394 ) | ( n12059 & n12395 ) | ( n12394 & n12395 ) ;
  assign n12398 = ( n12059 & n12396 ) | ( n12059 & ~n12397 ) | ( n12396 & ~n12397 ) ;
  assign n12399 = ( x108 & n12060 ) | ( x108 & ~n12178 ) | ( n12060 & ~n12178 ) ;
  assign n12400 = x108 & n12060 ;
  assign n12401 = ( n12065 & n12399 ) | ( n12065 & n12400 ) | ( n12399 & n12400 ) ;
  assign n12402 = ( ~n12065 & n12399 ) | ( ~n12065 & n12400 ) | ( n12399 & n12400 ) ;
  assign n12403 = ( n12065 & ~n12401 ) | ( n12065 & n12402 ) | ( ~n12401 & n12402 ) ;
  assign n12404 = ( x109 & n12066 ) | ( x109 & ~n12178 ) | ( n12066 & ~n12178 ) ;
  assign n12405 = x109 & n12066 ;
  assign n12406 = ( ~n12071 & n12404 ) | ( ~n12071 & n12405 ) | ( n12404 & n12405 ) ;
  assign n12407 = ( n12071 & n12404 ) | ( n12071 & n12405 ) | ( n12404 & n12405 ) ;
  assign n12408 = ( n12071 & n12406 ) | ( n12071 & ~n12407 ) | ( n12406 & ~n12407 ) ;
  assign n12409 = ( x110 & n12072 ) | ( x110 & ~n12178 ) | ( n12072 & ~n12178 ) ;
  assign n12410 = x110 & n12072 ;
  assign n12411 = ( n12077 & n12409 ) | ( n12077 & n12410 ) | ( n12409 & n12410 ) ;
  assign n12412 = ( ~n12077 & n12409 ) | ( ~n12077 & n12410 ) | ( n12409 & n12410 ) ;
  assign n12413 = ( n12077 & ~n12411 ) | ( n12077 & n12412 ) | ( ~n12411 & n12412 ) ;
  assign n12414 = ( x111 & n12078 ) | ( x111 & ~n12178 ) | ( n12078 & ~n12178 ) ;
  assign n12415 = x111 & n12078 ;
  assign n12416 = ( ~n12083 & n12414 ) | ( ~n12083 & n12415 ) | ( n12414 & n12415 ) ;
  assign n12417 = ( n12083 & n12414 ) | ( n12083 & n12415 ) | ( n12414 & n12415 ) ;
  assign n12418 = ( n12083 & n12416 ) | ( n12083 & ~n12417 ) | ( n12416 & ~n12417 ) ;
  assign n12419 = ( x112 & n12084 ) | ( x112 & ~n12178 ) | ( n12084 & ~n12178 ) ;
  assign n12420 = x112 & n12084 ;
  assign n12421 = ( n12089 & n12419 ) | ( n12089 & n12420 ) | ( n12419 & n12420 ) ;
  assign n12422 = ( ~n12089 & n12419 ) | ( ~n12089 & n12420 ) | ( n12419 & n12420 ) ;
  assign n12423 = ( n12089 & ~n12421 ) | ( n12089 & n12422 ) | ( ~n12421 & n12422 ) ;
  assign n12424 = ( x113 & n12090 ) | ( x113 & ~n12178 ) | ( n12090 & ~n12178 ) ;
  assign n12425 = x113 & n12090 ;
  assign n12426 = ( ~n12095 & n12424 ) | ( ~n12095 & n12425 ) | ( n12424 & n12425 ) ;
  assign n12427 = ( n12095 & n12424 ) | ( n12095 & n12425 ) | ( n12424 & n12425 ) ;
  assign n12428 = ( n12095 & n12426 ) | ( n12095 & ~n12427 ) | ( n12426 & ~n12427 ) ;
  assign n12429 = ( x114 & n12096 ) | ( x114 & ~n12178 ) | ( n12096 & ~n12178 ) ;
  assign n12430 = x114 & n12096 ;
  assign n12431 = ( n12101 & n12429 ) | ( n12101 & n12430 ) | ( n12429 & n12430 ) ;
  assign n12432 = ( ~n12101 & n12429 ) | ( ~n12101 & n12430 ) | ( n12429 & n12430 ) ;
  assign n12433 = ( n12101 & ~n12431 ) | ( n12101 & n12432 ) | ( ~n12431 & n12432 ) ;
  assign n12434 = ( x115 & n12102 ) | ( x115 & ~n12178 ) | ( n12102 & ~n12178 ) ;
  assign n12435 = x115 & n12102 ;
  assign n12436 = ( ~n12107 & n12434 ) | ( ~n12107 & n12435 ) | ( n12434 & n12435 ) ;
  assign n12437 = ( n12107 & n12434 ) | ( n12107 & n12435 ) | ( n12434 & n12435 ) ;
  assign n12438 = ( n12107 & n12436 ) | ( n12107 & ~n12437 ) | ( n12436 & ~n12437 ) ;
  assign n12439 = ( x116 & n12108 ) | ( x116 & ~n12178 ) | ( n12108 & ~n12178 ) ;
  assign n12440 = x116 & n12108 ;
  assign n12441 = ( n12113 & n12439 ) | ( n12113 & n12440 ) | ( n12439 & n12440 ) ;
  assign n12442 = ( ~n12113 & n12439 ) | ( ~n12113 & n12440 ) | ( n12439 & n12440 ) ;
  assign n12443 = ( n12113 & ~n12441 ) | ( n12113 & n12442 ) | ( ~n12441 & n12442 ) ;
  assign n12444 = ( x117 & n12114 ) | ( x117 & ~n12178 ) | ( n12114 & ~n12178 ) ;
  assign n12445 = x117 & n12114 ;
  assign n12446 = ( ~n12119 & n12444 ) | ( ~n12119 & n12445 ) | ( n12444 & n12445 ) ;
  assign n12447 = ( n12119 & n12444 ) | ( n12119 & n12445 ) | ( n12444 & n12445 ) ;
  assign n12448 = ( n12119 & n12446 ) | ( n12119 & ~n12447 ) | ( n12446 & ~n12447 ) ;
  assign n12449 = ( x118 & n12120 ) | ( x118 & ~n12178 ) | ( n12120 & ~n12178 ) ;
  assign n12450 = x118 & n12120 ;
  assign n12451 = ( n12125 & n12449 ) | ( n12125 & n12450 ) | ( n12449 & n12450 ) ;
  assign n12452 = ( ~n12125 & n12449 ) | ( ~n12125 & n12450 ) | ( n12449 & n12450 ) ;
  assign n12453 = ( n12125 & ~n12451 ) | ( n12125 & n12452 ) | ( ~n12451 & n12452 ) ;
  assign n12454 = ( x119 & n12126 ) | ( x119 & ~n12178 ) | ( n12126 & ~n12178 ) ;
  assign n12455 = x119 & n12126 ;
  assign n12456 = ( ~n12131 & n12454 ) | ( ~n12131 & n12455 ) | ( n12454 & n12455 ) ;
  assign n12457 = ( n12131 & n12454 ) | ( n12131 & n12455 ) | ( n12454 & n12455 ) ;
  assign n12458 = ( n12131 & n12456 ) | ( n12131 & ~n12457 ) | ( n12456 & ~n12457 ) ;
  assign n12459 = ( x120 & n12132 ) | ( x120 & ~n12178 ) | ( n12132 & ~n12178 ) ;
  assign n12460 = x120 & n12132 ;
  assign n12461 = ( n12137 & n12459 ) | ( n12137 & n12460 ) | ( n12459 & n12460 ) ;
  assign n12462 = ( ~n12137 & n12459 ) | ( ~n12137 & n12460 ) | ( n12459 & n12460 ) ;
  assign n12463 = ( n12137 & ~n12461 ) | ( n12137 & n12462 ) | ( ~n12461 & n12462 ) ;
  assign n12464 = ( x121 & n12138 ) | ( x121 & ~n12178 ) | ( n12138 & ~n12178 ) ;
  assign n12465 = x121 & n12138 ;
  assign n12466 = ( ~n12143 & n12464 ) | ( ~n12143 & n12465 ) | ( n12464 & n12465 ) ;
  assign n12467 = ( n12143 & n12464 ) | ( n12143 & n12465 ) | ( n12464 & n12465 ) ;
  assign n12468 = ( n12143 & n12466 ) | ( n12143 & ~n12467 ) | ( n12466 & ~n12467 ) ;
  assign n12469 = ( x122 & n12144 ) | ( x122 & ~n12178 ) | ( n12144 & ~n12178 ) ;
  assign n12470 = x122 & n12144 ;
  assign n12471 = ( n12149 & n12469 ) | ( n12149 & n12470 ) | ( n12469 & n12470 ) ;
  assign n12472 = ( ~n12149 & n12469 ) | ( ~n12149 & n12470 ) | ( n12469 & n12470 ) ;
  assign n12473 = ( n12149 & ~n12471 ) | ( n12149 & n12472 ) | ( ~n12471 & n12472 ) ;
  assign n12474 = ( x123 & n12150 ) | ( x123 & ~n12178 ) | ( n12150 & ~n12178 ) ;
  assign n12475 = x123 & n12150 ;
  assign n12476 = ( ~n12155 & n12474 ) | ( ~n12155 & n12475 ) | ( n12474 & n12475 ) ;
  assign n12477 = ( n12155 & n12474 ) | ( n12155 & n12475 ) | ( n12474 & n12475 ) ;
  assign n12478 = ( n12155 & n12476 ) | ( n12155 & ~n12477 ) | ( n12476 & ~n12477 ) ;
  assign n12479 = ( x124 & n12156 ) | ( x124 & ~n12178 ) | ( n12156 & ~n12178 ) ;
  assign n12480 = x124 & n12156 ;
  assign n12481 = ( n12161 & n12479 ) | ( n12161 & n12480 ) | ( n12479 & n12480 ) ;
  assign n12482 = ( ~n12161 & n12479 ) | ( ~n12161 & n12480 ) | ( n12479 & n12480 ) ;
  assign n12483 = ( n12161 & ~n12481 ) | ( n12161 & n12482 ) | ( ~n12481 & n12482 ) ;
  assign n12484 = ( x125 & n12162 ) | ( x125 & ~n12178 ) | ( n12162 & ~n12178 ) ;
  assign n12485 = x125 & n12162 ;
  assign n12486 = ( ~n12167 & n12484 ) | ( ~n12167 & n12485 ) | ( n12484 & n12485 ) ;
  assign n12487 = ( n12167 & n12484 ) | ( n12167 & n12485 ) | ( n12484 & n12485 ) ;
  assign n12488 = ( n12167 & n12486 ) | ( n12167 & ~n12487 ) | ( n12486 & ~n12487 ) ;
  assign n12489 = ( x126 & n12168 ) | ( x126 & ~n12178 ) | ( n12168 & ~n12178 ) ;
  assign n12490 = x126 & n12168 ;
  assign n12491 = ( ~n12173 & n12489 ) | ( ~n12173 & n12490 ) | ( n12489 & n12490 ) ;
  assign n12492 = ( n12173 & n12489 ) | ( n12173 & n12490 ) | ( n12489 & n12490 ) ;
  assign n12493 = ( n12173 & n12491 ) | ( n12173 & ~n12492 ) | ( n12491 & ~n12492 ) ;
  assign n12494 = ( x127 & ~n12174 ) | ( x127 & n12177 ) | ( ~n12174 & n12177 ) ;
  assign n12495 = ( ~x127 & n12174 ) | ( ~x127 & n12177 ) | ( n12174 & n12177 ) ;
  assign n12496 = n12494 & n12495 ;
  assign y0 = ~n12178 ;
  assign y1 = ~n11803 ;
  assign y2 = ~n11437 ;
  assign y3 = ~n11073 ;
  assign y4 = ~n10715 ;
  assign y5 = ~n10363 ;
  assign y6 = ~n10017 ;
  assign y7 = ~n9677 ;
  assign y8 = ~n9343 ;
  assign y9 = ~n9015 ;
  assign y10 = ~n8693 ;
  assign y11 = ~n8377 ;
  assign y12 = ~n8067 ;
  assign y13 = ~n7763 ;
  assign y14 = ~n7464 ;
  assign y15 = ~n7173 ;
  assign y16 = ~n6890 ;
  assign y17 = ~n6610 ;
  assign y18 = ~n6334 ;
  assign y19 = ~n6069 ;
  assign y20 = ~n5807 ;
  assign y21 = ~n5551 ;
  assign y22 = ~n5301 ;
  assign y23 = ~n5057 ;
  assign y24 = ~n4819 ;
  assign y25 = ~n4587 ;
  assign y26 = ~n4361 ;
  assign y27 = ~n4140 ;
  assign y28 = ~n3926 ;
  assign y29 = ~n3718 ;
  assign y30 = ~n3516 ;
  assign y31 = ~n3317 ;
  assign y32 = ~n3130 ;
  assign y33 = ~n2946 ;
  assign y34 = ~n2766 ;
  assign y35 = ~n2597 ;
  assign y36 = ~n2431 ;
  assign y37 = ~n2271 ;
  assign y38 = ~n2117 ;
  assign y39 = ~n1969 ;
  assign y40 = ~n1825 ;
  assign y41 = ~n1692 ;
  assign y42 = ~n1561 ;
  assign y43 = ~n1435 ;
  assign y44 = ~n1319 ;
  assign y45 = ~n1207 ;
  assign y46 = ~n1099 ;
  assign y47 = ~n1002 ;
  assign y48 = ~n905 ;
  assign y49 = ~n817 ;
  assign y50 = ~n734 ;
  assign y51 = ~n658 ;
  assign y52 = ~n585 ;
  assign y53 = ~n524 ;
  assign y54 = ~n465 ;
  assign y55 = ~n412 ;
  assign y56 = ~n369 ;
  assign y57 = ~n330 ;
  assign y58 = ~n285 ;
  assign y59 = ~n252 ;
  assign y60 = ~n233 ;
  assign y61 = ~n210 ;
  assign y62 = ~n200 ;
  assign y63 = ~n12180 ;
  assign y64 = n12183 ;
  assign y65 = n12188 ;
  assign y66 = n12193 ;
  assign y67 = n12198 ;
  assign y68 = n12203 ;
  assign y69 = n12208 ;
  assign y70 = n12213 ;
  assign y71 = n12218 ;
  assign y72 = n12223 ;
  assign y73 = n12228 ;
  assign y74 = n12233 ;
  assign y75 = n12238 ;
  assign y76 = n12243 ;
  assign y77 = n12248 ;
  assign y78 = n12253 ;
  assign y79 = n12258 ;
  assign y80 = n12263 ;
  assign y81 = n12268 ;
  assign y82 = n12273 ;
  assign y83 = n12278 ;
  assign y84 = n12283 ;
  assign y85 = n12288 ;
  assign y86 = n12293 ;
  assign y87 = n12298 ;
  assign y88 = n12303 ;
  assign y89 = n12308 ;
  assign y90 = n12313 ;
  assign y91 = n12318 ;
  assign y92 = n12323 ;
  assign y93 = n12328 ;
  assign y94 = n12333 ;
  assign y95 = n12338 ;
  assign y96 = n12343 ;
  assign y97 = n12348 ;
  assign y98 = n12353 ;
  assign y99 = n12358 ;
  assign y100 = n12363 ;
  assign y101 = n12368 ;
  assign y102 = n12373 ;
  assign y103 = n12378 ;
  assign y104 = n12383 ;
  assign y105 = n12388 ;
  assign y106 = n12393 ;
  assign y107 = n12398 ;
  assign y108 = n12403 ;
  assign y109 = n12408 ;
  assign y110 = n12413 ;
  assign y111 = n12418 ;
  assign y112 = n12423 ;
  assign y113 = n12428 ;
  assign y114 = n12433 ;
  assign y115 = n12438 ;
  assign y116 = n12443 ;
  assign y117 = n12448 ;
  assign y118 = n12453 ;
  assign y119 = n12458 ;
  assign y120 = n12463 ;
  assign y121 = n12468 ;
  assign y122 = n12473 ;
  assign y123 = n12478 ;
  assign y124 = n12483 ;
  assign y125 = n12488 ;
  assign y126 = n12493 ;
  assign y127 = n12496 ;
endmodule
