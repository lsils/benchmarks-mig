module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 ;
  assign n129 = x125 & ~x126 ;
  assign n130 = x121 & ~x122 ;
  assign n131 = x119 & ~x120 ;
  assign n132 = x117 & ~x118 ;
  assign n133 = x114 | x115 ;
  assign n134 = x112 | x113 ;
  assign n135 = x111 & ~n134 ;
  assign n136 = ( x113 & ~n133 ) | ( x113 & n135 ) | ( ~n133 & n135 ) ;
  assign n137 = ( x115 & ~x116 ) | ( x115 & n136 ) | ( ~x116 & n136 ) ;
  assign n138 = ( ~x118 & n132 ) | ( ~x118 & n137 ) | ( n132 & n137 ) ;
  assign n139 = ( ~x120 & n131 ) | ( ~x120 & n138 ) | ( n131 & n138 ) ;
  assign n140 = ( ~x122 & n130 ) | ( ~x122 & n139 ) | ( n130 & n139 ) ;
  assign n141 = x123 & ~x124 ;
  assign n142 = ( ~x124 & n140 ) | ( ~x124 & n141 ) | ( n140 & n141 ) ;
  assign n143 = ( ~x126 & n129 ) | ( ~x126 & n142 ) | ( n129 & n142 ) ;
  assign n144 = x110 | x112 ;
  assign n145 = x108 | x109 ;
  assign n146 = ( ~x109 & x114 ) | ( ~x109 & n145 ) | ( x114 & n145 ) ;
  assign n147 = x116 | n146 ;
  assign n148 = x118 | x120 ;
  assign n149 = x122 | x124 ;
  assign n150 = ( x126 & ~n148 ) | ( x126 & n149 ) | ( ~n148 & n149 ) ;
  assign n151 = n148 | n150 ;
  assign n152 = ( ~n144 & n147 ) | ( ~n144 & n151 ) | ( n147 & n151 ) ;
  assign n153 = n144 | n152 ;
  assign n154 = x107 | x109 ;
  assign n155 = x103 | x105 ;
  assign n156 = x104 & ~x105 ;
  assign n157 = x102 | x103 ;
  assign n158 = x99 | x101 ;
  assign n159 = x98 | x99 ;
  assign n160 = x96 | x97 ;
  assign n161 = ( ~x97 & n159 ) | ( ~x97 & n160 ) | ( n159 & n160 ) ;
  assign n162 = ~x101 & n161 ;
  assign n163 = ( x100 & ~n158 ) | ( x100 & n162 ) | ( ~n158 & n162 ) ;
  assign n164 = n157 | n163 ;
  assign n165 = ( ~n155 & n156 ) | ( ~n155 & n164 ) | ( n156 & n164 ) ;
  assign n166 = x106 | n165 ;
  assign n167 = x95 | x97 ;
  assign n168 = ( ~n155 & n158 ) | ( ~n155 & n167 ) | ( n158 & n167 ) ;
  assign n169 = x93 & ~x94 ;
  assign n170 = ( ~n155 & n168 ) | ( ~n155 & n169 ) | ( n168 & n169 ) ;
  assign n171 = n155 | n170 ;
  assign n172 = x88 | x89 ;
  assign n173 = x87 & ~n172 ;
  assign n174 = x84 | x85 ;
  assign n175 = x80 | x81 ;
  assign n176 = x76 | x77 ;
  assign n177 = x75 & ~n176 ;
  assign n178 = x70 | x71 ;
  assign n179 = x66 | x67 ;
  assign n180 = x64 | x65 ;
  assign n181 = x63 & ~n180 ;
  assign n182 = ( x65 & ~n179 ) | ( x65 & n181 ) | ( ~n179 & n181 ) ;
  assign n183 = ( x67 & ~x68 ) | ( x67 & n182 ) | ( ~x68 & n182 ) ;
  assign n184 = x69 & ~n178 ;
  assign n185 = ( ~n178 & n183 ) | ( ~n178 & n184 ) | ( n183 & n184 ) ;
  assign n186 = x72 | x73 ;
  assign n187 = ( x71 & n185 ) | ( x71 & ~n186 ) | ( n185 & ~n186 ) ;
  assign n188 = ( x73 & ~x74 ) | ( x73 & n187 ) | ( ~x74 & n187 ) ;
  assign n189 = ( ~n176 & n177 ) | ( ~n176 & n188 ) | ( n177 & n188 ) ;
  assign n190 = ( x77 & ~x78 ) | ( x77 & n189 ) | ( ~x78 & n189 ) ;
  assign n191 = x79 & ~n175 ;
  assign n192 = ( ~n175 & n190 ) | ( ~n175 & n191 ) | ( n190 & n191 ) ;
  assign n193 = ( x81 & ~x82 ) | ( x81 & n192 ) | ( ~x82 & n192 ) ;
  assign n194 = x83 & ~n174 ;
  assign n195 = ( ~n174 & n193 ) | ( ~n174 & n194 ) | ( n193 & n194 ) ;
  assign n196 = ( x85 & ~x86 ) | ( x85 & n195 ) | ( ~x86 & n195 ) ;
  assign n197 = ( ~n172 & n173 ) | ( ~n172 & n196 ) | ( n173 & n196 ) ;
  assign n198 = ( x89 & ~x90 ) | ( x89 & n197 ) | ( ~x90 & n197 ) ;
  assign n199 = x91 | n198 ;
  assign n200 = x92 | x93 ;
  assign n201 = x94 | x95 ;
  assign n202 = n200 | n201 ;
  assign n203 = ~n171 & n202 ;
  assign n204 = ( n171 & n199 ) | ( n171 & ~n203 ) | ( n199 & ~n203 ) ;
  assign n205 = ~n166 & n204 ;
  assign n206 = ~n154 & n205 ;
  assign n207 = ( ~n153 & n154 ) | ( ~n153 & n206 ) | ( n154 & n206 ) ;
  assign n208 = n143 | n207 ;
  assign n209 = x90 | x91 ;
  assign n210 = ( n172 & n202 ) | ( n172 & ~n209 ) | ( n202 & ~n209 ) ;
  assign n211 = n209 | n210 ;
  assign n212 = x86 | x87 ;
  assign n213 = n174 | n212 ;
  assign n214 = n211 | n213 ;
  assign n215 = x82 | x83 ;
  assign n216 = n175 | n215 ;
  assign n217 = n214 | n216 ;
  assign n218 = x78 | x79 ;
  assign n219 = n176 | n218 ;
  assign n220 = x74 | x75 ;
  assign n221 = n186 | n220 ;
  assign n222 = n219 | n221 ;
  assign n223 = n179 | n180 ;
  assign n224 = x68 | x69 ;
  assign n225 = n178 | n224 ;
  assign n226 = n223 | n225 ;
  assign n227 = n222 | n226 ;
  assign n228 = n217 | n227 ;
  assign n229 = x106 | x107 ;
  assign n230 = x110 | x111 ;
  assign n231 = n229 | n230 ;
  assign n232 = ( x105 & n156 ) | ( x105 & ~n229 ) | ( n156 & ~n229 ) ;
  assign n233 = n145 | n232 ;
  assign n234 = n231 | n233 ;
  assign n235 = x100 | x101 ;
  assign n236 = n157 | n235 ;
  assign n237 = n159 | n160 ;
  assign n238 = n236 | n237 ;
  assign n239 = n234 | n238 ;
  assign n240 = x120 | x121 ;
  assign n241 = x122 | x123 ;
  assign n242 = n240 | n241 ;
  assign n243 = x124 | x125 ;
  assign n244 = x126 | x127 ;
  assign n245 = n243 | n244 ;
  assign n246 = n242 | n245 ;
  assign n247 = x116 | x117 ;
  assign n248 = x118 | x119 ;
  assign n249 = n247 | n248 ;
  assign n250 = n133 | n134 ;
  assign n251 = n249 | n250 ;
  assign n252 = n246 | n251 ;
  assign n253 = n239 | n252 ;
  assign n254 = n228 | n253 ;
  assign n255 = x60 | x61 ;
  assign n256 = x54 | x55 ;
  assign n257 = ( ~x55 & x56 ) | ( ~x55 & n256 ) | ( x56 & n256 ) ;
  assign n258 = x58 | x59 ;
  assign n259 = x57 & ~n258 ;
  assign n260 = ( n257 & n258 ) | ( n257 & ~n259 ) | ( n258 & ~n259 ) ;
  assign n261 = ( ~x59 & n255 ) | ( ~x59 & n260 ) | ( n255 & n260 ) ;
  assign n262 = ( ~x61 & x62 ) | ( ~x61 & n261 ) | ( x62 & n261 ) ;
  assign n263 = n254 | n262 ;
  assign n264 = x51 & ~x52 ;
  assign n265 = x48 | x50 ;
  assign n266 = x46 | x47 ;
  assign n267 = x45 & ~n266 ;
  assign n268 = ( x47 & ~n265 ) | ( x47 & n267 ) | ( ~n265 & n267 ) ;
  assign n269 = ( x49 & ~x50 ) | ( x49 & n268 ) | ( ~x50 & n268 ) ;
  assign n270 = ( ~x52 & n264 ) | ( ~x52 & n269 ) | ( n264 & n269 ) ;
  assign n271 = x53 | x55 ;
  assign n272 = x57 | x59 ;
  assign n273 = ( x61 & ~n271 ) | ( x61 & n272 ) | ( ~n271 & n272 ) ;
  assign n274 = n271 | n273 ;
  assign n275 = ( x127 & ~n270 ) | ( x127 & n274 ) | ( ~n270 & n274 ) ;
  assign n276 = n270 | n275 ;
  assign n277 = ( x127 & ~n263 ) | ( x127 & n276 ) | ( ~n263 & n276 ) ;
  assign n278 = n208 | n277 ;
  assign n279 = x44 | x45 ;
  assign n280 = n266 | n279 ;
  assign n281 = ( ~x52 & n263 ) | ( ~x52 & n265 ) | ( n263 & n265 ) ;
  assign n282 = ( ~x52 & n280 ) | ( ~x52 & n281 ) | ( n280 & n281 ) ;
  assign n283 = x52 | n282 ;
  assign n284 = x42 | x43 ;
  assign n285 = x40 | x41 ;
  assign n286 = x32 | x34 ;
  assign n287 = x36 | n286 ;
  assign n288 = x30 | x31 ;
  assign n289 = x28 | x29 ;
  assign n290 = x26 | x27 ;
  assign n291 = x16 | x17 ;
  assign n292 = x12 | x13 ;
  assign n293 = x8 | x9 ;
  assign n294 = x7 & ~n293 ;
  assign n295 = x4 | x5 ;
  assign n296 = x2 | x3 ;
  assign n297 = x1 & ~n296 ;
  assign n298 = ( x3 & ~n295 ) | ( x3 & n297 ) | ( ~n295 & n297 ) ;
  assign n299 = ( x5 & ~x6 ) | ( x5 & n298 ) | ( ~x6 & n298 ) ;
  assign n300 = ( ~n293 & n294 ) | ( ~n293 & n299 ) | ( n294 & n299 ) ;
  assign n301 = ( x9 & ~x10 ) | ( x9 & n300 ) | ( ~x10 & n300 ) ;
  assign n302 = x11 & ~n292 ;
  assign n303 = ( ~n292 & n301 ) | ( ~n292 & n302 ) | ( n301 & n302 ) ;
  assign n304 = ( x13 & ~x14 ) | ( x13 & n303 ) | ( ~x14 & n303 ) ;
  assign n305 = x15 & ~n291 ;
  assign n306 = ( ~n291 & n304 ) | ( ~n291 & n305 ) | ( n304 & n305 ) ;
  assign n307 = ( x17 & ~x18 ) | ( x17 & n306 ) | ( ~x18 & n306 ) ;
  assign n308 = x19 | n307 ;
  assign n309 = x20 & ~x21 ;
  assign n310 = ( x21 & n308 ) | ( x21 & ~n309 ) | ( n308 & ~n309 ) ;
  assign n311 = x22 & ~x23 ;
  assign n312 = ( x23 & n310 ) | ( x23 & ~n311 ) | ( n310 & ~n311 ) ;
  assign n313 = x24 | x25 ;
  assign n314 = n312 & ~n313 ;
  assign n315 = ( x25 & ~n290 ) | ( x25 & n314 ) | ( ~n290 & n314 ) ;
  assign n316 = ( x27 & ~n289 ) | ( x27 & n315 ) | ( ~n289 & n315 ) ;
  assign n317 = ( x29 & ~n288 ) | ( x29 & n316 ) | ( ~n288 & n316 ) ;
  assign n318 = ( x31 & ~n287 ) | ( x31 & n317 ) | ( ~n287 & n317 ) ;
  assign n319 = x34 | x35 ;
  assign n320 = x33 & ~n319 ;
  assign n321 = x36 | x37 ;
  assign n322 = ( x35 & n320 ) | ( x35 & ~n321 ) | ( n320 & ~n321 ) ;
  assign n323 = ( x37 & ~x38 ) | ( x37 & n322 ) | ( ~x38 & n322 ) ;
  assign n324 = ( ~x38 & n318 ) | ( ~x38 & n323 ) | ( n318 & n323 ) ;
  assign n325 = x39 & ~n285 ;
  assign n326 = ( ~n285 & n324 ) | ( ~n285 & n325 ) | ( n324 & n325 ) ;
  assign n327 = ( x41 & ~n284 ) | ( x41 & n326 ) | ( ~n284 & n326 ) ;
  assign n328 = ( x43 & ~n283 ) | ( x43 & n327 ) | ( ~n283 & n327 ) ;
  assign n329 = n278 | n328 ;
  assign n330 = n133 & ~n249 ;
  assign n331 = ( ~n242 & n248 ) | ( ~n242 & n330 ) | ( n248 & n330 ) ;
  assign n332 = ( n241 & ~n243 ) | ( n241 & n331 ) | ( ~n243 & n331 ) ;
  assign n333 = n244 | n332 ;
  assign n334 = n252 & ~n333 ;
  assign n335 = n157 | n231 ;
  assign n336 = n235 & ~n335 ;
  assign n337 = ~n159 & n160 ;
  assign n338 = n201 | n212 ;
  assign n339 = ( n214 & ~n215 ) | ( n214 & n216 ) | ( ~n215 & n216 ) ;
  assign n340 = ( n211 & ~n338 ) | ( n211 & n339 ) | ( ~n338 & n339 ) ;
  assign n341 = ( n200 & ~n209 ) | ( n200 & n340 ) | ( ~n209 & n340 ) ;
  assign n342 = ~n201 & n341 ;
  assign n343 = ( ~n159 & n337 ) | ( ~n159 & n342 ) | ( n337 & n342 ) ;
  assign n344 = ( ~n335 & n336 ) | ( ~n335 & n343 ) | ( n336 & n343 ) ;
  assign n345 = ( ~n230 & n233 ) | ( ~n230 & n344 ) | ( n233 & n344 ) ;
  assign n346 = n159 | n215 ;
  assign n347 = ~n176 & n220 ;
  assign n348 = n209 | n218 ;
  assign n349 = ( ~n338 & n347 ) | ( ~n338 & n348 ) | ( n347 & n348 ) ;
  assign n350 = ( ~n338 & n346 ) | ( ~n338 & n349 ) | ( n346 & n349 ) ;
  assign n351 = n338 | n350 ;
  assign n352 = n335 | n351 ;
  assign n353 = x62 | x63 ;
  assign n354 = n255 | n353 ;
  assign n355 = x56 | x57 ;
  assign n356 = n256 & ~n355 ;
  assign n357 = n258 | n356 ;
  assign n358 = x52 | x53 ;
  assign n359 = n256 | n358 ;
  assign n360 = n355 | n359 ;
  assign n361 = x50 | x51 ;
  assign n362 = x48 | x49 ;
  assign n363 = n361 | n362 ;
  assign n364 = ( n280 & n284 ) | ( n280 & ~n285 ) | ( n284 & ~n285 ) ;
  assign n365 = n285 | n364 ;
  assign n366 = x38 | x39 ;
  assign n367 = n321 | n366 ;
  assign n368 = n319 & ~n367 ;
  assign n369 = ( ~n365 & n366 ) | ( ~n365 & n368 ) | ( n366 & n368 ) ;
  assign n370 = ( ~n279 & n284 ) | ( ~n279 & n369 ) | ( n284 & n369 ) ;
  assign n371 = n266 | n370 ;
  assign n372 = x22 | x23 ;
  assign n373 = n288 | n289 ;
  assign n374 = n290 | n313 ;
  assign n375 = n373 | n374 ;
  assign n376 = x20 | x21 ;
  assign n377 = n372 | n376 ;
  assign n378 = x18 | x19 ;
  assign n379 = x14 | x15 ;
  assign n380 = n292 | n379 ;
  assign n381 = x10 | x11 ;
  assign n382 = x6 | x7 ;
  assign n383 = n293 | n381 ;
  assign n384 = n295 | n382 ;
  assign n385 = n296 & ~n384 ;
  assign n386 = ( n382 & ~n383 ) | ( n382 & n385 ) | ( ~n383 & n385 ) ;
  assign n387 = ( ~n380 & n381 ) | ( ~n380 & n386 ) | ( n381 & n386 ) ;
  assign n388 = ( ~n291 & n379 ) | ( ~n291 & n387 ) | ( n379 & n387 ) ;
  assign n389 = n378 | n388 ;
  assign n390 = ~n377 & n389 ;
  assign n391 = ( n372 & ~n375 ) | ( n372 & n390 ) | ( ~n375 & n390 ) ;
  assign n392 = ( ~n289 & n290 ) | ( ~n289 & n391 ) | ( n290 & n391 ) ;
  assign n393 = n288 | n392 ;
  assign n394 = x32 | x33 ;
  assign n395 = ( n319 & n367 ) | ( n319 & ~n394 ) | ( n367 & ~n394 ) ;
  assign n396 = n394 | n395 ;
  assign n397 = n365 | n396 ;
  assign n398 = ~n371 & n397 ;
  assign n399 = ( n371 & n393 ) | ( n371 & ~n398 ) | ( n393 & ~n398 ) ;
  assign n400 = ~n363 & n399 ;
  assign n401 = ( ~n354 & n361 ) | ( ~n354 & n400 ) | ( n361 & n400 ) ;
  assign n402 = ~n360 & n401 ;
  assign n403 = ( ~n354 & n357 ) | ( ~n354 & n402 ) | ( n357 & n402 ) ;
  assign n404 = ( ~n227 & n353 ) | ( ~n227 & n403 ) | ( n353 & n403 ) ;
  assign n405 = n179 & ~n224 ;
  assign n406 = n178 | n405 ;
  assign n407 = ( ~n222 & n404 ) | ( ~n222 & n406 ) | ( n404 & n406 ) ;
  assign n408 = ~n345 & n407 ;
  assign n409 = ( ~n345 & n352 ) | ( ~n345 & n408 ) | ( n352 & n408 ) ;
  assign n410 = ( n333 & ~n334 ) | ( n333 & n409 ) | ( ~n334 & n409 ) ;
  assign n411 = n242 & ~n245 ;
  assign n412 = n145 | n230 ;
  assign n413 = ~n234 & n236 ;
  assign n414 = ( ~n250 & n412 ) | ( ~n250 & n413 ) | ( n412 & n413 ) ;
  assign n415 = n249 | n414 ;
  assign n416 = ( ~n202 & n211 ) | ( ~n202 & n253 ) | ( n211 & n253 ) ;
  assign n417 = ~n415 & n416 ;
  assign n418 = ( ~n245 & n411 ) | ( ~n245 & n417 ) | ( n411 & n417 ) ;
  assign n419 = n214 | n253 ;
  assign n420 = ( n291 & n377 ) | ( n291 & ~n378 ) | ( n377 & ~n378 ) ;
  assign n421 = n378 | n420 ;
  assign n422 = n380 | n383 ;
  assign n423 = n384 & ~n422 ;
  assign n424 = ( n380 & ~n421 ) | ( n380 & n423 ) | ( ~n421 & n423 ) ;
  assign n425 = ( ~n374 & n377 ) | ( ~n374 & n424 ) | ( n377 & n424 ) ;
  assign n426 = n373 & ~n396 ;
  assign n427 = ( ~n396 & n425 ) | ( ~n396 & n426 ) | ( n425 & n426 ) ;
  assign n428 = ( ~n365 & n367 ) | ( ~n365 & n427 ) | ( n367 & n427 ) ;
  assign n429 = ( n280 & ~n363 ) | ( n280 & n428 ) | ( ~n363 & n428 ) ;
  assign n430 = n359 | n429 ;
  assign n431 = n258 | n355 ;
  assign n432 = ~n354 & n431 ;
  assign n433 = ( n354 & n430 ) | ( n354 & ~n432 ) | ( n430 & ~n432 ) ;
  assign n434 = ~n226 & n433 ;
  assign n435 = ( ~n222 & n225 ) | ( ~n222 & n434 ) | ( n225 & n434 ) ;
  assign n436 = ( ~n216 & n219 ) | ( ~n216 & n435 ) | ( n219 & n435 ) ;
  assign n437 = ~n419 & n436 ;
  assign n438 = ( ~n418 & n419 ) | ( ~n418 & n437 ) | ( n419 & n437 ) ;
  assign n439 = ~n246 & n251 ;
  assign n440 = n354 | n431 ;
  assign n441 = n375 | n421 ;
  assign n442 = n422 & ~n441 ;
  assign n443 = ( n375 & ~n397 ) | ( n375 & n442 ) | ( ~n397 & n442 ) ;
  assign n444 = n359 | n363 ;
  assign n445 = n440 | n444 ;
  assign n446 = ( n365 & n443 ) | ( n365 & ~n445 ) | ( n443 & ~n445 ) ;
  assign n447 = ( ~n227 & n440 ) | ( ~n227 & n446 ) | ( n440 & n446 ) ;
  assign n448 = ( ~n217 & n222 ) | ( ~n217 & n447 ) | ( n222 & n447 ) ;
  assign n449 = ( n211 & ~n238 ) | ( n211 & n448 ) | ( ~n238 & n448 ) ;
  assign n450 = n234 | n449 ;
  assign n451 = ( n246 & ~n439 ) | ( n246 & n450 ) | ( ~n439 & n450 ) ;
  assign n452 = n397 | n445 ;
  assign n453 = n441 & ~n452 ;
  assign n454 = ( ~n228 & n445 ) | ( ~n228 & n453 ) | ( n445 & n453 ) ;
  assign n455 = ( n217 & ~n239 ) | ( n217 & n454 ) | ( ~n239 & n454 ) ;
  assign n456 = n252 | n455 ;
  assign n457 = n253 | n452 ;
  assign n458 = ( ~n228 & n253 ) | ( ~n228 & n457 ) | ( n253 & n457 ) ;
  assign n459 = x0 | x1 ;
  assign n460 = ( n296 & n384 ) | ( n296 & ~n459 ) | ( n384 & ~n459 ) ;
  assign n461 = n459 | n460 ;
  assign n462 = ( n422 & n441 ) | ( n422 & ~n461 ) | ( n441 & ~n461 ) ;
  assign n463 = n461 | n462 ;
  assign n464 = ( n254 & n452 ) | ( n254 & ~n463 ) | ( n452 & ~n463 ) ;
  assign n465 = n463 | n464 ;
  assign y0 = n329 ;
  assign y1 = n410 ;
  assign y2 = n438 ;
  assign y3 = n451 ;
  assign y4 = n456 ;
  assign y5 = n458 ;
  assign y6 = n254 ;
  assign y7 = n465 ;
endmodule
