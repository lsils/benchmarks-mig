module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 ;
  assign n148 = x11 | x22 ;
  assign n149 = x16 | x18 ;
  assign n150 = x19 | n149 ;
  assign n151 = x8 | x21 ;
  assign n152 = x10 | x14 ;
  assign n153 = n151 | n152 ;
  assign n154 = x4 | x7 ;
  assign n155 = x13 | n154 ;
  assign n156 = n153 | n155 ;
  assign n157 = n150 | n156 ;
  assign n158 = n148 | n157 ;
  assign n159 = x6 | x12 ;
  assign n160 = x5 | x9 ;
  assign n161 = n159 | n160 ;
  assign n162 = x17 | n161 ;
  assign n163 = n158 | n162 ;
  assign n164 = x54 & n163 ;
  assign n165 = x0 & ~n164 ;
  assign n166 = x3 | x129 ;
  assign n167 = x9 | x11 ;
  assign n168 = x5 | x22 ;
  assign n169 = n167 | n168 ;
  assign n170 = ( x56 & n167 ) | ( x56 & n168 ) | ( n167 & n168 ) ;
  assign n171 = ( x54 & ~n169 ) | ( x54 & n170 ) | ( ~n169 & n170 ) ;
  assign n172 = n166 | n171 ;
  assign n173 = x54 & ~n166 ;
  assign n174 = ~n162 & n173 ;
  assign n175 = ~n148 & n174 ;
  assign n176 = ( x10 & x14 ) | ( x10 & n151 ) | ( x14 & n151 ) ;
  assign n177 = n150 | n176 ;
  assign n178 = x8 & x21 ;
  assign n179 = ( x4 & ~n177 ) | ( x4 & n178 ) | ( ~n177 & n178 ) ;
  assign n180 = n177 | n179 ;
  assign n181 = n175 & ~n180 ;
  assign n182 = ( x7 & x13 ) | ( x7 & n153 ) | ( x13 & n153 ) ;
  assign n183 = n181 & ~n182 ;
  assign n184 = n172 & ~n183 ;
  assign n185 = n165 | n184 ;
  assign n186 = x1 & n181 ;
  assign n187 = x6 & x12 ;
  assign n188 = ~x17 & x54 ;
  assign n189 = x9 | n166 ;
  assign n190 = ( x5 & n159 ) | ( x5 & n189 ) | ( n159 & n189 ) ;
  assign n191 = ( n158 & n188 ) | ( n158 & n190 ) | ( n188 & n190 ) ;
  assign n192 = n188 & ~n191 ;
  assign n193 = ~n187 & n192 ;
  assign n194 = x1 | n188 ;
  assign n195 = ( n186 & ~n193 ) | ( n186 & n194 ) | ( ~n193 & n194 ) ;
  assign n196 = x7 | x13 ;
  assign n197 = ( n166 & n183 ) | ( n166 & ~n196 ) | ( n183 & ~n196 ) ;
  assign n198 = n183 & ~n197 ;
  assign n199 = ( n166 & n195 ) | ( n166 & ~n198 ) | ( n195 & ~n198 ) ;
  assign n200 = x122 & x127 ;
  assign n201 = x24 | x49 ;
  assign n202 = x42 | x44 ;
  assign n203 = x82 & ~n202 ;
  assign n204 = ~x40 & n203 ;
  assign n205 = ~x38 & n204 ;
  assign n206 = ~x50 & n205 ;
  assign n207 = ~x46 & n206 ;
  assign n208 = x41 | x43 ;
  assign n209 = n207 & ~n208 ;
  assign n210 = x45 | x47 ;
  assign n211 = x48 | n210 ;
  assign n212 = n209 & ~n211 ;
  assign n213 = ~n201 & n212 ;
  assign n214 = x2 | x15 ;
  assign n215 = x20 | n214 ;
  assign n216 = n213 & n215 ;
  assign n217 = ( x82 & ~n213 ) | ( x82 & n216 ) | ( ~n213 & n216 ) ;
  assign n218 = n200 | n217 ;
  assign n219 = x65 | n218 ;
  assign n220 = x82 | n200 ;
  assign n221 = ~x15 & n213 ;
  assign n222 = n220 & ~n221 ;
  assign n223 = x20 & n221 ;
  assign n224 = ( x2 & n222 ) | ( x2 & n223 ) | ( n222 & n223 ) ;
  assign n225 = ~x129 & n224 ;
  assign n226 = ( x129 & n219 ) | ( x129 & ~n225 ) | ( n219 & ~n225 ) ;
  assign n227 = x61 | x118 ;
  assign n228 = ( x129 & n163 ) | ( x129 & n227 ) | ( n163 & n227 ) ;
  assign n229 = x123 | x129 ;
  assign n230 = x0 & ~x113 ;
  assign n231 = ~n229 & n230 ;
  assign n232 = ( n163 & ~n228 ) | ( n163 & n231 ) | ( ~n228 & n231 ) ;
  assign n233 = x54 | n166 ;
  assign n234 = x4 & ~n233 ;
  assign n235 = x10 | n234 ;
  assign n236 = ( n183 & n234 ) | ( n183 & n235 ) | ( n234 & n235 ) ;
  assign n237 = x5 & ~n233 ;
  assign n238 = ~n156 & n175 ;
  assign n239 = x29 | n177 ;
  assign n240 = x59 | n239 ;
  assign n241 = n238 & ~n240 ;
  assign n242 = x25 | x28 ;
  assign n243 = ( ~x25 & n237 ) | ( ~x25 & n242 ) | ( n237 & n242 ) ;
  assign n244 = ( n237 & n241 ) | ( n237 & n243 ) | ( n241 & n243 ) ;
  assign n245 = x6 & ~n233 ;
  assign n246 = ( ~x28 & n242 ) | ( ~x28 & n245 ) | ( n242 & n245 ) ;
  assign n247 = ( n241 & n245 ) | ( n241 & n246 ) | ( n245 & n246 ) ;
  assign n248 = x7 & ~n233 ;
  assign n249 = x8 | n248 ;
  assign n250 = ( n183 & n248 ) | ( n183 & n249 ) | ( n248 & n249 ) ;
  assign n251 = x8 & ~n233 ;
  assign n252 = x21 | n251 ;
  assign n253 = ( n183 & n251 ) | ( n183 & n252 ) | ( n251 & n252 ) ;
  assign n254 = x9 & ~n233 ;
  assign n255 = x11 & ~x22 ;
  assign n256 = ~n157 & n174 ;
  assign n257 = n255 & ~n256 ;
  assign n258 = ( n254 & n255 ) | ( n254 & ~n257 ) | ( n255 & ~n257 ) ;
  assign n259 = x10 & ~n233 ;
  assign n260 = x14 | n259 ;
  assign n261 = ( n183 & n259 ) | ( n183 & n260 ) | ( n259 & n260 ) ;
  assign n262 = x11 & ~n233 ;
  assign n263 = ~x11 & n256 ;
  assign n264 = ( n148 & n262 ) | ( n148 & n263 ) | ( n262 & n263 ) ;
  assign n265 = ~x19 & n238 ;
  assign n266 = x12 & ~n233 ;
  assign n267 = ( ~x16 & n149 ) | ( ~x16 & n266 ) | ( n149 & n266 ) ;
  assign n268 = ( n265 & n266 ) | ( n265 & n267 ) | ( n266 & n267 ) ;
  assign n269 = x29 & x54 ;
  assign n270 = ( x59 & n242 ) | ( x59 & n269 ) | ( n242 & n269 ) ;
  assign n271 = n269 & ~n270 ;
  assign n272 = x13 & ~n166 ;
  assign n273 = ( ~n166 & n271 ) | ( ~n166 & n272 ) | ( n271 & n272 ) ;
  assign n274 = ~n164 & n273 ;
  assign n275 = x14 & ~n233 ;
  assign n276 = x13 | n275 ;
  assign n277 = ( n183 & n275 ) | ( n183 & n276 ) | ( n275 & n276 ) ;
  assign n278 = n215 & n220 ;
  assign n279 = n200 & ~n215 ;
  assign n280 = ( x70 & ~n278 ) | ( x70 & n279 ) | ( ~n278 & n279 ) ;
  assign n281 = x129 | n280 ;
  assign n282 = ( ~x15 & n213 ) | ( ~x15 & n220 ) | ( n213 & n220 ) ;
  assign n283 = ( ~n221 & n281 ) | ( ~n221 & n282 ) | ( n281 & n282 ) ;
  assign n284 = x16 & ~n233 ;
  assign n285 = ( x6 & ~n187 ) | ( x6 & n284 ) | ( ~n187 & n284 ) ;
  assign n286 = ( n192 & n284 ) | ( n192 & n285 ) | ( n284 & n285 ) ;
  assign n287 = x17 & ~n233 ;
  assign n288 = x59 & ~n242 ;
  assign n289 = ~n239 & n288 ;
  assign n290 = n287 | n289 ;
  assign n291 = ( n238 & n287 ) | ( n238 & n290 ) | ( n287 & n290 ) ;
  assign n292 = ~x18 & n265 ;
  assign n293 = x18 & ~n233 ;
  assign n294 = ( n149 & n292 ) | ( n149 & n293 ) | ( n292 & n293 ) ;
  assign n295 = x19 & ~n233 ;
  assign n296 = x17 & ~n161 ;
  assign n297 = n173 & n296 ;
  assign n298 = ~n158 & n297 ;
  assign n299 = n295 | n298 ;
  assign n300 = ~x20 & n222 ;
  assign n301 = ( x71 & ~n278 ) | ( x71 & n279 ) | ( ~n278 & n279 ) ;
  assign n302 = x129 | n301 ;
  assign n303 = n223 | n302 ;
  assign n304 = n300 | n303 ;
  assign n305 = x21 & ~n233 ;
  assign n306 = ( ~n149 & n150 ) | ( ~n149 & n305 ) | ( n150 & n305 ) ;
  assign n307 = ( n238 & n305 ) | ( n238 & n306 ) | ( n305 & n306 ) ;
  assign n308 = x22 & ~n233 ;
  assign n309 = x5 | n308 ;
  assign n310 = ( n192 & n308 ) | ( n192 & n309 ) | ( n308 & n309 ) ;
  assign n311 = ~x23 & x55 ;
  assign n312 = x61 & ~x129 ;
  assign n313 = ~n311 & n312 ;
  assign n314 = ~n212 & n220 ;
  assign n315 = x24 | n314 ;
  assign n316 = x24 & ~n212 ;
  assign n317 = x129 | n279 ;
  assign n318 = ( x129 & n213 ) | ( x129 & n317 ) | ( n213 & n317 ) ;
  assign n319 = ( n315 & ~n316 ) | ( n315 & n318 ) | ( ~n316 & n318 ) ;
  assign n320 = x63 & ~n218 ;
  assign n321 = n319 | n320 ;
  assign n322 = x53 | x58 ;
  assign n323 = x116 & ~n166 ;
  assign n324 = n322 & n323 ;
  assign n325 = ( x26 & x27 ) | ( x26 & n322 ) | ( x27 & n322 ) ;
  assign n326 = n166 | n325 ;
  assign n327 = x26 | x27 ;
  assign n328 = n322 | n327 ;
  assign n329 = x53 & x58 ;
  assign n330 = ( x85 & n328 ) | ( x85 & n329 ) | ( n328 & n329 ) ;
  assign n331 = n326 | n330 ;
  assign n332 = n324 | n331 ;
  assign n333 = x39 | x51 ;
  assign n334 = x52 | n333 ;
  assign n335 = ~x26 & n334 ;
  assign n336 = x85 & x116 ;
  assign n337 = x85 | x110 ;
  assign n338 = n328 | n337 ;
  assign n339 = x96 | n338 ;
  assign n340 = ( x100 & n336 ) | ( x100 & ~n339 ) | ( n336 & ~n339 ) ;
  assign n341 = x116 & n327 ;
  assign n342 = ( ~x26 & n334 ) | ( ~x26 & n341 ) | ( n334 & n341 ) ;
  assign n343 = ( ~n335 & n340 ) | ( ~n335 & n342 ) | ( n340 & n342 ) ;
  assign n344 = ~n332 & n343 ;
  assign n345 = x95 | x100 ;
  assign n346 = x97 | n345 ;
  assign n347 = ~n338 & n346 ;
  assign n348 = ( ~n166 & n336 ) | ( ~n166 & n347 ) | ( n336 & n347 ) ;
  assign n349 = n341 | n348 ;
  assign n350 = x25 & ~n349 ;
  assign n351 = ( ~n332 & n344 ) | ( ~n332 & n350 ) | ( n344 & n350 ) ;
  assign n352 = ~n334 & n341 ;
  assign n353 = ( x26 & n340 ) | ( x26 & ~n352 ) | ( n340 & ~n352 ) ;
  assign n354 = ~n331 & n353 ;
  assign n355 = x95 & ~n166 ;
  assign n356 = ~n339 & n355 ;
  assign n357 = ( ~n331 & n336 ) | ( ~n331 & n356 ) | ( n336 & n356 ) ;
  assign n358 = ( x27 & ~n331 ) | ( x27 & n357 ) | ( ~n331 & n357 ) ;
  assign n359 = ~n343 & n358 ;
  assign n360 = ( x28 & n341 ) | ( x28 & ~n347 ) | ( n341 & ~n347 ) ;
  assign n361 = ~n332 & n360 ;
  assign n362 = ~n343 & n357 ;
  assign n363 = ( ~n343 & n361 ) | ( ~n343 & n362 ) | ( n361 & n362 ) ;
  assign n364 = n339 | n345 ;
  assign n365 = n348 & ~n364 ;
  assign n366 = x58 & x116 ;
  assign n367 = x97 & n366 ;
  assign n368 = n331 & n367 ;
  assign n369 = ( n365 & n367 ) | ( n365 & ~n368 ) | ( n367 & ~n368 ) ;
  assign n370 = x29 & ~n332 ;
  assign n371 = n349 & n370 ;
  assign n372 = ( n369 & n370 ) | ( n369 & ~n371 ) | ( n370 & ~n371 ) ;
  assign n373 = ~x88 & x106 ;
  assign n374 = x129 | n373 ;
  assign n375 = ~x60 & x109 ;
  assign n376 = x30 | x109 ;
  assign n377 = ( x106 & ~n375 ) | ( x106 & n376 ) | ( ~n375 & n376 ) ;
  assign n378 = ~n374 & n377 ;
  assign n379 = ~x89 & x106 ;
  assign n380 = x129 | n379 ;
  assign n381 = ~x30 & x109 ;
  assign n382 = x31 | x109 ;
  assign n383 = ( x106 & ~n381 ) | ( x106 & n382 ) | ( ~n381 & n382 ) ;
  assign n384 = ~n380 & n383 ;
  assign n385 = ~x99 & x106 ;
  assign n386 = x129 | n385 ;
  assign n387 = ~x31 & x109 ;
  assign n388 = x32 | x109 ;
  assign n389 = ( x106 & ~n387 ) | ( x106 & n388 ) | ( ~n387 & n388 ) ;
  assign n390 = ~n386 & n389 ;
  assign n391 = ~x90 & x106 ;
  assign n392 = x129 | n391 ;
  assign n393 = ~x32 & x109 ;
  assign n394 = x33 | x109 ;
  assign n395 = ( x106 & ~n393 ) | ( x106 & n394 ) | ( ~n393 & n394 ) ;
  assign n396 = ~n392 & n395 ;
  assign n397 = ~x91 & x106 ;
  assign n398 = x129 | n397 ;
  assign n399 = ~x33 & x109 ;
  assign n400 = x34 | x109 ;
  assign n401 = ( x106 & ~n399 ) | ( x106 & n400 ) | ( ~n399 & n400 ) ;
  assign n402 = ~n398 & n401 ;
  assign n403 = ~x92 & x106 ;
  assign n404 = x129 | n403 ;
  assign n405 = ~x34 & x109 ;
  assign n406 = x35 | x109 ;
  assign n407 = ( x106 & ~n405 ) | ( x106 & n406 ) | ( ~n405 & n406 ) ;
  assign n408 = ~n404 & n407 ;
  assign n409 = ~x98 & x106 ;
  assign n410 = x129 | n409 ;
  assign n411 = ~x35 & x109 ;
  assign n412 = x36 | x109 ;
  assign n413 = ( x106 & ~n411 ) | ( x106 & n412 ) | ( ~n411 & n412 ) ;
  assign n414 = ~n410 & n413 ;
  assign n415 = ~x93 & x106 ;
  assign n416 = x129 | n415 ;
  assign n417 = ~x36 & x109 ;
  assign n418 = x37 | x109 ;
  assign n419 = ( x106 & ~n417 ) | ( x106 & n418 ) | ( ~n417 & n418 ) ;
  assign n420 = ~n416 & n419 ;
  assign n421 = ( ~n213 & n220 ) | ( ~n213 & n278 ) | ( n220 & n278 ) ;
  assign n422 = x38 & ~n204 ;
  assign n423 = ( n205 & ~n318 ) | ( n205 & n422 ) | ( ~n318 & n422 ) ;
  assign n424 = n421 & n423 ;
  assign n425 = x74 | n421 ;
  assign n426 = ( n318 & ~n424 ) | ( n318 & n425 ) | ( ~n424 & n425 ) ;
  assign n427 = ~x51 & x109 ;
  assign n428 = ~x52 & n427 ;
  assign n429 = ~x39 & n428 ;
  assign n430 = ( x39 & x106 ) | ( x39 & ~n428 ) | ( x106 & ~n428 ) ;
  assign n431 = ( ~x129 & n429 ) | ( ~x129 & n430 ) | ( n429 & n430 ) ;
  assign n432 = x73 | n218 ;
  assign n433 = x40 & ~n203 ;
  assign n434 = ( n204 & n218 ) | ( n204 & n433 ) | ( n218 & n433 ) ;
  assign n435 = ( n318 & n432 ) | ( n318 & ~n434 ) | ( n432 & ~n434 ) ;
  assign n436 = x76 | n218 ;
  assign n437 = ~x41 & n207 ;
  assign n438 = x41 & ~n207 ;
  assign n439 = ( n421 & n437 ) | ( n421 & n438 ) | ( n437 & n438 ) ;
  assign n440 = ( x129 & n436 ) | ( x129 & ~n439 ) | ( n436 & ~n439 ) ;
  assign n441 = x42 & n220 ;
  assign n442 = ~x44 & n217 ;
  assign n443 = x72 | n218 ;
  assign n444 = ( n441 & n442 ) | ( n441 & n443 ) | ( n442 & n443 ) ;
  assign n445 = ~n442 & n444 ;
  assign n446 = ( x129 & n443 ) | ( x129 & ~n444 ) | ( n443 & ~n444 ) ;
  assign n447 = ( n441 & ~n445 ) | ( n441 & n446 ) | ( ~n445 & n446 ) ;
  assign n448 = x43 & ~n437 ;
  assign n449 = ( n209 & n421 ) | ( n209 & n448 ) | ( n421 & n448 ) ;
  assign n450 = x77 | n218 ;
  assign n451 = ( x129 & ~n449 ) | ( x129 & n450 ) | ( ~n449 & n450 ) ;
  assign n452 = x67 | n200 ;
  assign n453 = x44 & n200 ;
  assign n454 = ( n217 & n452 ) | ( n217 & ~n453 ) | ( n452 & ~n453 ) ;
  assign n455 = ( x129 & ~n442 ) | ( x129 & n454 ) | ( ~n442 & n454 ) ;
  assign n456 = ~x47 & n209 ;
  assign n457 = ~x48 & n456 ;
  assign n458 = ~x45 & n314 ;
  assign n459 = ( n314 & n457 ) | ( n314 & n458 ) | ( n457 & n458 ) ;
  assign n460 = x68 & ~n421 ;
  assign n461 = n318 | n460 ;
  assign n462 = n459 | n461 ;
  assign n463 = x46 & ~n206 ;
  assign n464 = ( n207 & n421 ) | ( n207 & n463 ) | ( n421 & n463 ) ;
  assign n465 = x75 | n218 ;
  assign n466 = ( x129 & ~n464 ) | ( x129 & n465 ) | ( ~n464 & n465 ) ;
  assign n467 = x64 | n218 ;
  assign n468 = x47 & ~n209 ;
  assign n469 = ( n218 & n456 ) | ( n218 & n468 ) | ( n456 & n468 ) ;
  assign n470 = ( n318 & n467 ) | ( n318 & ~n469 ) | ( n467 & ~n469 ) ;
  assign n471 = x62 & ~n421 ;
  assign n472 = n318 | n471 ;
  assign n473 = ( ~x48 & n421 ) | ( ~x48 & n456 ) | ( n421 & n456 ) ;
  assign n474 = ( ~n457 & n472 ) | ( ~n457 & n473 ) | ( n472 & n473 ) ;
  assign n475 = x24 & n212 ;
  assign n476 = ( x49 & n314 ) | ( x49 & n475 ) | ( n314 & n475 ) ;
  assign n477 = ( n200 & ~n213 ) | ( n200 & n220 ) | ( ~n213 & n220 ) ;
  assign n478 = x69 | n477 ;
  assign n479 = ( ~n216 & n476 ) | ( ~n216 & n478 ) | ( n476 & n478 ) ;
  assign n480 = ( x129 & ~n476 ) | ( x129 & n479 ) | ( ~n476 & n479 ) ;
  assign n481 = x66 | n218 ;
  assign n482 = x50 & ~n205 ;
  assign n483 = ( n206 & n421 ) | ( n206 & n482 ) | ( n421 & n482 ) ;
  assign n484 = ( x129 & n481 ) | ( x129 & ~n483 ) | ( n481 & ~n483 ) ;
  assign n485 = ( x51 & x106 ) | ( x51 & ~x109 ) | ( x106 & ~x109 ) ;
  assign n486 = ( ~x129 & n427 ) | ( ~x129 & n485 ) | ( n427 & n485 ) ;
  assign n487 = ( x52 & x106 ) | ( x52 & ~n427 ) | ( x106 & ~n427 ) ;
  assign n488 = ( ~x129 & n428 ) | ( ~x129 & n487 ) | ( n428 & n487 ) ;
  assign n489 = x53 & ~n332 ;
  assign n490 = n369 | n489 ;
  assign n491 = ~x129 & n218 ;
  assign n492 = x114 & ~x122 ;
  assign n493 = ~n229 & n492 ;
  assign n494 = x37 | x116 ;
  assign n495 = ~x94 & x116 ;
  assign n496 = ( x26 & ~n494 ) | ( x26 & n495 ) | ( ~n494 & n495 ) ;
  assign n497 = x37 | x58 ;
  assign n498 = x94 | x116 ;
  assign n499 = x58 & ~n498 ;
  assign n500 = ( x26 & n497 ) | ( x26 & ~n499 ) | ( n497 & ~n499 ) ;
  assign n501 = ~n496 & n500 ;
  assign n502 = ~n331 & n501 ;
  assign n503 = x60 & n366 ;
  assign n504 = x57 & ~n366 ;
  assign n505 = ( ~n331 & n503 ) | ( ~n331 & n504 ) | ( n503 & n504 ) ;
  assign n506 = ( x58 & ~n324 ) | ( x58 & n352 ) | ( ~n324 & n352 ) ;
  assign n507 = ~n331 & n506 ;
  assign n508 = x96 & n347 ;
  assign n509 = x59 | n508 ;
  assign n510 = ( ~n349 & n508 ) | ( ~n349 & n509 ) | ( n508 & n509 ) ;
  assign n511 = ~n332 & n510 ;
  assign n512 = ~x117 & x123 ;
  assign n513 = ~x60 & x122 ;
  assign n514 = ( x60 & x117 ) | ( x60 & x122 ) | ( x117 & x122 ) ;
  assign n515 = ( n512 & ~n513 ) | ( n512 & n514 ) | ( ~n513 & n514 ) ;
  assign n516 = x114 | x122 ;
  assign n517 = x123 & ~x129 ;
  assign n518 = ~n516 & n517 ;
  assign n519 = x136 & ~x137 ;
  assign n520 = x132 & x133 ;
  assign n521 = x131 & n520 ;
  assign n522 = ~x138 & n521 ;
  assign n523 = n519 & n522 ;
  assign n524 = ~x140 & n523 ;
  assign n525 = x62 & ~n523 ;
  assign n526 = ( ~x129 & n524 ) | ( ~x129 & n525 ) | ( n524 & n525 ) ;
  assign n527 = x63 & ~n523 ;
  assign n528 = ~x142 & n523 ;
  assign n529 = ( ~x129 & n527 ) | ( ~x129 & n528 ) | ( n527 & n528 ) ;
  assign n530 = x64 & ~n523 ;
  assign n531 = ~x139 & n523 ;
  assign n532 = ( ~x129 & n530 ) | ( ~x129 & n531 ) | ( n530 & n531 ) ;
  assign n533 = x65 & ~n523 ;
  assign n534 = ~x146 & n523 ;
  assign n535 = ( ~x129 & n533 ) | ( ~x129 & n534 ) | ( n533 & n534 ) ;
  assign n536 = x136 | x137 ;
  assign n537 = n522 & ~n536 ;
  assign n538 = x66 & ~n537 ;
  assign n539 = ~x143 & n537 ;
  assign n540 = ( ~x129 & n538 ) | ( ~x129 & n539 ) | ( n538 & n539 ) ;
  assign n541 = x67 & ~n537 ;
  assign n542 = ~x139 & n537 ;
  assign n543 = ( ~x129 & n541 ) | ( ~x129 & n542 ) | ( n541 & n542 ) ;
  assign n544 = ~x141 & n523 ;
  assign n545 = x68 & ~n523 ;
  assign n546 = ( ~x129 & n544 ) | ( ~x129 & n545 ) | ( n544 & n545 ) ;
  assign n547 = ~x143 & n523 ;
  assign n548 = x69 & ~n523 ;
  assign n549 = ( ~x129 & n547 ) | ( ~x129 & n548 ) | ( n547 & n548 ) ;
  assign n550 = ~x144 & n523 ;
  assign n551 = x70 & ~n523 ;
  assign n552 = ( ~x129 & n550 ) | ( ~x129 & n551 ) | ( n550 & n551 ) ;
  assign n553 = ~x145 & n523 ;
  assign n554 = x71 & ~n523 ;
  assign n555 = ( ~x129 & n553 ) | ( ~x129 & n554 ) | ( n553 & n554 ) ;
  assign n556 = ~x140 & n537 ;
  assign n557 = x72 & ~n537 ;
  assign n558 = ( ~x129 & n556 ) | ( ~x129 & n557 ) | ( n556 & n557 ) ;
  assign n559 = x73 & ~n537 ;
  assign n560 = ~x141 & n537 ;
  assign n561 = ( ~x129 & n559 ) | ( ~x129 & n560 ) | ( n559 & n560 ) ;
  assign n562 = x74 & ~n537 ;
  assign n563 = ~x142 & n537 ;
  assign n564 = ( ~x129 & n562 ) | ( ~x129 & n563 ) | ( n562 & n563 ) ;
  assign n565 = x75 & ~n537 ;
  assign n566 = ~x144 & n537 ;
  assign n567 = ( ~x129 & n565 ) | ( ~x129 & n566 ) | ( n565 & n566 ) ;
  assign n568 = ~x145 & n537 ;
  assign n569 = x76 & ~n537 ;
  assign n570 = ( ~x129 & n568 ) | ( ~x129 & n569 ) | ( n568 & n569 ) ;
  assign n571 = x77 & ~n537 ;
  assign n572 = ~x146 & n537 ;
  assign n573 = ( ~x129 & n571 ) | ( ~x129 & n572 ) | ( n571 & n572 ) ;
  assign n574 = ~x136 & x137 ;
  assign n575 = n522 & n574 ;
  assign n576 = x142 & n575 ;
  assign n577 = x78 & ~n575 ;
  assign n578 = ( ~x129 & n576 ) | ( ~x129 & n577 ) | ( n576 & n577 ) ;
  assign n579 = x79 & ~n575 ;
  assign n580 = x143 & n575 ;
  assign n581 = ( ~x129 & n579 ) | ( ~x129 & n580 ) | ( n579 & n580 ) ;
  assign n582 = x80 & ~n575 ;
  assign n583 = x144 & n575 ;
  assign n584 = ( ~x129 & n582 ) | ( ~x129 & n583 ) | ( n582 & n583 ) ;
  assign n585 = x145 & n575 ;
  assign n586 = x81 & ~n575 ;
  assign n587 = ( ~x129 & n585 ) | ( ~x129 & n586 ) | ( n585 & n586 ) ;
  assign n588 = x146 & n575 ;
  assign n589 = x82 & ~n575 ;
  assign n590 = ( ~x129 & n588 ) | ( ~x129 & n589 ) | ( n588 & n589 ) ;
  assign n591 = x72 | x137 ;
  assign n592 = x87 & x137 ;
  assign n593 = ( x136 & n591 ) | ( x136 & ~n592 ) | ( n591 & ~n592 ) ;
  assign n594 = x119 | x136 ;
  assign n595 = ~x89 & x136 ;
  assign n596 = ( x137 & n594 ) | ( x137 & ~n595 ) | ( n594 & ~n595 ) ;
  assign n597 = x136 & x137 ;
  assign n598 = ( x115 & x137 ) | ( x115 & n597 ) | ( x137 & n597 ) ;
  assign n599 = ( x138 & ~n596 ) | ( x138 & n598 ) | ( ~n596 & n598 ) ;
  assign n600 = x62 | x137 ;
  assign n601 = x31 & x137 ;
  assign n602 = ( x136 & ~n600 ) | ( x136 & n601 ) | ( ~n600 & n601 ) ;
  assign n603 = ( x138 & n593 ) | ( x138 & n602 ) | ( n593 & n602 ) ;
  assign n604 = ( n593 & n599 ) | ( n593 & ~n603 ) | ( n599 & ~n603 ) ;
  assign n605 = x141 & n575 ;
  assign n606 = x84 & ~n575 ;
  assign n607 = ( ~x129 & n605 ) | ( ~x129 & n606 ) | ( n605 & n606 ) ;
  assign n608 = x85 & ~x116 ;
  assign n609 = ( ~n331 & n508 ) | ( ~n331 & n608 ) | ( n508 & n608 ) ;
  assign n610 = x86 & ~n575 ;
  assign n611 = x139 & n575 ;
  assign n612 = ( ~x129 & n610 ) | ( ~x129 & n611 ) | ( n610 & n611 ) ;
  assign n613 = x87 & ~n575 ;
  assign n614 = x140 & n575 ;
  assign n615 = ( ~x129 & n613 ) | ( ~x129 & n614 ) | ( n613 & n614 ) ;
  assign n616 = n522 & n597 ;
  assign n617 = x88 & ~n616 ;
  assign n618 = x139 & n616 ;
  assign n619 = ( ~x129 & n617 ) | ( ~x129 & n618 ) | ( n617 & n618 ) ;
  assign n620 = x140 & n616 ;
  assign n621 = x89 & ~n616 ;
  assign n622 = ( ~x129 & n620 ) | ( ~x129 & n621 ) | ( n620 & n621 ) ;
  assign n623 = x142 & n616 ;
  assign n624 = x90 & ~n616 ;
  assign n625 = ( ~x129 & n623 ) | ( ~x129 & n624 ) | ( n623 & n624 ) ;
  assign n626 = x143 & n616 ;
  assign n627 = x91 & ~n616 ;
  assign n628 = ( ~x129 & n626 ) | ( ~x129 & n627 ) | ( n626 & n627 ) ;
  assign n629 = x144 & n616 ;
  assign n630 = x92 & ~n616 ;
  assign n631 = ( ~x129 & n629 ) | ( ~x129 & n630 ) | ( n629 & n630 ) ;
  assign n632 = x93 & ~n616 ;
  assign n633 = x146 & n616 ;
  assign n634 = ( ~x129 & n632 ) | ( ~x129 & n633 ) | ( n632 & n633 ) ;
  assign n635 = x82 & x138 ;
  assign n636 = ~n536 & n635 ;
  assign n637 = n521 & n636 ;
  assign n638 = x142 & n637 ;
  assign n639 = x94 & ~n637 ;
  assign n640 = ( ~x129 & n638 ) | ( ~x129 & n639 ) | ( n638 & n639 ) ;
  assign n641 = x95 & ~n637 ;
  assign n642 = x143 & n637 ;
  assign n643 = x3 | x110 ;
  assign n644 = ~x129 & n521 ;
  assign n645 = ( x129 & n643 ) | ( x129 & ~n644 ) | ( n643 & ~n644 ) ;
  assign n646 = ( n641 & n642 ) | ( n641 & ~n645 ) | ( n642 & ~n645 ) ;
  assign n647 = x146 & n637 ;
  assign n648 = x96 & ~n637 ;
  assign n649 = ( ~n645 & n647 ) | ( ~n645 & n648 ) | ( n647 & n648 ) ;
  assign n650 = x145 & n637 ;
  assign n651 = x97 & ~n637 ;
  assign n652 = ( ~n645 & n650 ) | ( ~n645 & n651 ) | ( n650 & n651 ) ;
  assign n653 = x98 & ~n616 ;
  assign n654 = x145 & n616 ;
  assign n655 = ( ~x129 & n653 ) | ( ~x129 & n654 ) | ( n653 & n654 ) ;
  assign n656 = x99 & ~n616 ;
  assign n657 = x141 & n616 ;
  assign n658 = ( ~x129 & n656 ) | ( ~x129 & n657 ) | ( n656 & n657 ) ;
  assign n659 = x144 & n637 ;
  assign n660 = x100 & ~n637 ;
  assign n661 = ( ~n645 & n659 ) | ( ~n645 & n660 ) | ( n659 & n660 ) ;
  assign n662 = x77 & ~x138 ;
  assign n663 = ~x124 & x138 ;
  assign n664 = ( ~n536 & n662 ) | ( ~n536 & n663 ) | ( n662 & n663 ) ;
  assign n665 = ~x37 & x137 ;
  assign n666 = x136 & ~x138 ;
  assign n667 = ( x137 & n665 ) | ( x137 & ~n666 ) | ( n665 & ~n666 ) ;
  assign n668 = x96 & x138 ;
  assign n669 = x82 & ~x138 ;
  assign n670 = ( ~x136 & n668 ) | ( ~x136 & n669 ) | ( n668 & n669 ) ;
  assign n671 = x65 & ~x138 ;
  assign n672 = ~x93 & x138 ;
  assign n673 = ( n519 & n671 ) | ( n519 & n672 ) | ( n671 & n672 ) ;
  assign n674 = ( n667 & ~n670 ) | ( n667 & n673 ) | ( ~n670 & n673 ) ;
  assign n675 = n664 | n674 ;
  assign n676 = x91 & n519 ;
  assign n677 = x95 & n574 ;
  assign n678 = ( x138 & n676 ) | ( x138 & n677 ) | ( n676 & n677 ) ;
  assign n679 = x69 | x137 ;
  assign n680 = x34 & x137 ;
  assign n681 = ( x136 & ~n679 ) | ( x136 & n680 ) | ( ~n679 & n680 ) ;
  assign n682 = x66 | x137 ;
  assign n683 = x79 & x137 ;
  assign n684 = ( x136 & n682 ) | ( x136 & ~n683 ) | ( n682 & ~n683 ) ;
  assign n685 = ( x138 & ~n681 ) | ( x138 & n684 ) | ( ~n681 & n684 ) ;
  assign n686 = ~n678 & n685 ;
  assign n687 = x90 & n519 ;
  assign n688 = x94 & n574 ;
  assign n689 = ( x138 & n687 ) | ( x138 & n688 ) | ( n687 & n688 ) ;
  assign n690 = x74 | n536 ;
  assign n691 = x33 & n597 ;
  assign n692 = n690 & ~n691 ;
  assign n693 = ~x63 & n519 ;
  assign n694 = x78 & n574 ;
  assign n695 = n693 | n694 ;
  assign n696 = ( x138 & n692 ) | ( x138 & ~n695 ) | ( n692 & ~n695 ) ;
  assign n697 = ~n689 & n696 ;
  assign n698 = ~x112 & x138 ;
  assign n699 = n574 & n698 ;
  assign n700 = x99 & n519 ;
  assign n701 = ~x84 & n574 ;
  assign n702 = x73 | x138 ;
  assign n703 = ( x138 & ~n536 ) | ( x138 & n702 ) | ( ~n536 & n702 ) ;
  assign n704 = ( ~n700 & n701 ) | ( ~n700 & n703 ) | ( n701 & n703 ) ;
  assign n705 = x68 & ~x137 ;
  assign n706 = ~x32 & x137 ;
  assign n707 = ( n666 & n705 ) | ( n666 & n706 ) | ( n705 & n706 ) ;
  assign n708 = ( ~n699 & n704 ) | ( ~n699 & n707 ) | ( n704 & n707 ) ;
  assign n709 = x35 & n666 ;
  assign n710 = x100 & x138 ;
  assign n711 = x80 & ~x138 ;
  assign n712 = ( ~x136 & n710 ) | ( ~x136 & n711 ) | ( n710 & n711 ) ;
  assign n713 = ( x137 & n709 ) | ( x137 & n712 ) | ( n709 & n712 ) ;
  assign n714 = x125 | x136 ;
  assign n715 = ~x92 & x136 ;
  assign n716 = ( x138 & ~n714 ) | ( x138 & n715 ) | ( ~n714 & n715 ) ;
  assign n717 = x70 & x136 ;
  assign n718 = x75 & ~x136 ;
  assign n719 = ( ~x138 & n717 ) | ( ~x138 & n718 ) | ( n717 & n718 ) ;
  assign n720 = ( ~x137 & n716 ) | ( ~x137 & n719 ) | ( n716 & n719 ) ;
  assign n721 = ( x137 & ~n713 ) | ( x137 & n720 ) | ( ~n713 & n720 ) ;
  assign n722 = x23 & ~x136 ;
  assign n723 = x98 & x136 ;
  assign n724 = ( x138 & n722 ) | ( x138 & n723 ) | ( n722 & n723 ) ;
  assign n725 = x76 | x136 ;
  assign n726 = ~x71 & x136 ;
  assign n727 = ( x138 & n725 ) | ( x138 & ~n726 ) | ( n725 & ~n726 ) ;
  assign n728 = ( x137 & ~n724 ) | ( x137 & n727 ) | ( ~n724 & n727 ) ;
  assign n729 = x97 & ~x136 ;
  assign n730 = x138 & n729 ;
  assign n731 = x36 & x136 ;
  assign n732 = x81 & ~x136 ;
  assign n733 = ( ~x138 & n731 ) | ( ~x138 & n732 ) | ( n731 & n732 ) ;
  assign n734 = ( x137 & n730 ) | ( x137 & n733 ) | ( n730 & n733 ) ;
  assign n735 = n728 & ~n734 ;
  assign n736 = x67 | x138 ;
  assign n737 = x120 & x138 ;
  assign n738 = ( x136 & n736 ) | ( x136 & ~n737 ) | ( n736 & ~n737 ) ;
  assign n739 = x88 & x138 ;
  assign n740 = x64 | x138 ;
  assign n741 = ( x136 & n739 ) | ( x136 & ~n740 ) | ( n739 & ~n740 ) ;
  assign n742 = ( x137 & n738 ) | ( x137 & ~n741 ) | ( n738 & ~n741 ) ;
  assign n743 = x30 & n666 ;
  assign n744 = x86 & ~x138 ;
  assign n745 = x111 & x138 ;
  assign n746 = ( ~x136 & n744 ) | ( ~x136 & n745 ) | ( n744 & n745 ) ;
  assign n747 = ( x137 & n743 ) | ( x137 & n746 ) | ( n743 & n746 ) ;
  assign n748 = n742 & ~n747 ;
  assign n749 = ( x27 & n166 ) | ( x27 & ~n335 ) | ( n166 & ~n335 ) ;
  assign n750 = n341 & ~n749 ;
  assign n751 = n329 | n367 ;
  assign n752 = n324 & ~n751 ;
  assign n753 = x139 & n636 ;
  assign n754 = x111 & ~n636 ;
  assign n755 = ( n644 & n753 ) | ( n644 & n754 ) | ( n753 & n754 ) ;
  assign n756 = x141 & n636 ;
  assign n757 = x112 | n636 ;
  assign n758 = ( n644 & n756 ) | ( n644 & ~n757 ) | ( n756 & ~n757 ) ;
  assign n759 = x54 & n148 ;
  assign n760 = x54 | x113 ;
  assign n761 = ( n166 & ~n759 ) | ( n166 & n760 ) | ( ~n759 & n760 ) ;
  assign n762 = x115 | n636 ;
  assign n763 = x140 & n636 ;
  assign n764 = ( n644 & ~n762 ) | ( n644 & n763 ) | ( ~n762 & n763 ) ;
  assign n765 = x9 | x12 ;
  assign n766 = n154 & ~n765 ;
  assign n767 = ( n173 & n765 ) | ( n173 & n766 ) | ( n765 & n766 ) ;
  assign n768 = x122 & ~x129 ;
  assign n769 = ~x54 & x118 ;
  assign n770 = ( ~x129 & n271 ) | ( ~x129 & n769 ) | ( n271 & n769 ) ;
  assign n771 = ~x129 & n345 ;
  assign n772 = x120 | n643 ;
  assign n773 = x111 | x129 ;
  assign n774 = n772 & ~n773 ;
  assign n775 = x81 & x120 ;
  assign n776 = ~x129 & n775 ;
  assign n777 = x129 | x134 ;
  assign n778 = x129 | x135 ;
  assign n779 = x57 & ~x129 ;
  assign n780 = x3 & ~x129 ;
  assign n781 = ~x96 & x125 ;
  assign n782 = ( ~x129 & n780 ) | ( ~x129 & n781 ) | ( n780 & n781 ) ;
  assign n783 = ~x126 & n520 ;
  assign y0 = x108 ;
  assign y1 = x83 ;
  assign y2 = x104 ;
  assign y3 = x103 ;
  assign y4 = x102 ;
  assign y5 = x105 ;
  assign y6 = x107 ;
  assign y7 = x101 ;
  assign y8 = x126 ;
  assign y9 = x121 ;
  assign y10 = x1 ;
  assign y11 = x0 ;
  assign y12 = ~1'b0 ;
  assign y13 = x130 ;
  assign y14 = x128 ;
  assign y15 = n185 ;
  assign y16 = n199 ;
  assign y17 = ~n226 ;
  assign y18 = n232 ;
  assign y19 = n236 ;
  assign y20 = n244 ;
  assign y21 = n247 ;
  assign y22 = n250 ;
  assign y23 = n253 ;
  assign y24 = n258 ;
  assign y25 = n261 ;
  assign y26 = n264 ;
  assign y27 = n268 ;
  assign y28 = n274 ;
  assign y29 = n277 ;
  assign y30 = ~n283 ;
  assign y31 = n286 ;
  assign y32 = n291 ;
  assign y33 = n294 ;
  assign y34 = n299 ;
  assign y35 = ~n304 ;
  assign y36 = n307 ;
  assign y37 = n310 ;
  assign y38 = n313 ;
  assign y39 = ~n321 ;
  assign y40 = n351 ;
  assign y41 = n354 ;
  assign y42 = n359 ;
  assign y43 = n363 ;
  assign y44 = n372 ;
  assign y45 = n378 ;
  assign y46 = n384 ;
  assign y47 = n390 ;
  assign y48 = n396 ;
  assign y49 = n402 ;
  assign y50 = n408 ;
  assign y51 = n414 ;
  assign y52 = n420 ;
  assign y53 = ~n426 ;
  assign y54 = n431 ;
  assign y55 = ~n435 ;
  assign y56 = ~n440 ;
  assign y57 = ~n447 ;
  assign y58 = ~n451 ;
  assign y59 = ~n455 ;
  assign y60 = ~n462 ;
  assign y61 = ~n466 ;
  assign y62 = ~n470 ;
  assign y63 = ~n474 ;
  assign y64 = ~n480 ;
  assign y65 = ~n484 ;
  assign y66 = n486 ;
  assign y67 = n488 ;
  assign y68 = n490 ;
  assign y69 = ~n491 ;
  assign y70 = n493 ;
  assign y71 = n502 ;
  assign y72 = n505 ;
  assign y73 = n507 ;
  assign y74 = n511 ;
  assign y75 = n515 ;
  assign y76 = n518 ;
  assign y77 = ~n526 ;
  assign y78 = ~n529 ;
  assign y79 = ~n532 ;
  assign y80 = ~n535 ;
  assign y81 = ~n540 ;
  assign y82 = ~n543 ;
  assign y83 = ~n546 ;
  assign y84 = ~n549 ;
  assign y85 = ~n552 ;
  assign y86 = ~n555 ;
  assign y87 = ~n558 ;
  assign y88 = ~n561 ;
  assign y89 = ~n564 ;
  assign y90 = ~n567 ;
  assign y91 = ~n570 ;
  assign y92 = ~n573 ;
  assign y93 = n578 ;
  assign y94 = n581 ;
  assign y95 = n584 ;
  assign y96 = n587 ;
  assign y97 = n590 ;
  assign y98 = ~n604 ;
  assign y99 = n607 ;
  assign y100 = n609 ;
  assign y101 = n612 ;
  assign y102 = n615 ;
  assign y103 = n619 ;
  assign y104 = n622 ;
  assign y105 = n625 ;
  assign y106 = n628 ;
  assign y107 = n631 ;
  assign y108 = n634 ;
  assign y109 = n640 ;
  assign y110 = n646 ;
  assign y111 = n649 ;
  assign y112 = n652 ;
  assign y113 = n655 ;
  assign y114 = n658 ;
  assign y115 = n661 ;
  assign y116 = ~n675 ;
  assign y117 = ~n686 ;
  assign y118 = ~n697 ;
  assign y119 = ~n708 ;
  assign y120 = ~n721 ;
  assign y121 = n348 ;
  assign y122 = ~n735 ;
  assign y123 = ~n748 ;
  assign y124 = n750 ;
  assign y125 = n752 ;
  assign y126 = n755 ;
  assign y127 = n758 ;
  assign y128 = ~n761 ;
  assign y129 = n229 ;
  assign y130 = n764 ;
  assign y131 = n767 ;
  assign y132 = ~n768 ;
  assign y133 = n770 ;
  assign y134 = n771 ;
  assign y135 = n774 ;
  assign y136 = n776 ;
  assign y137 = n777 ;
  assign y138 = n778 ;
  assign y139 = n779 ;
  assign y140 = n782 ;
  assign y141 = n783 ;
endmodule
