module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 ;
  assign n12 = x2 & x3 ;
  assign n13 = x7 | x8 ;
  assign n14 = n12 | n13 ;
  assign n15 = x6 & ~x9 ;
  assign n16 = ( x2 & x3 ) | ( x2 & n15 ) | ( x3 & n15 ) ;
  assign n17 = ~n14 & n16 ;
  assign n18 = x1 & x4 ;
  assign n19 = x0 & ~n18 ;
  assign n20 = ( ~x0 & x5 ) | ( ~x0 & n18 ) | ( x5 & n18 ) ;
  assign n21 = x1 & ~x2 ;
  assign n22 = x6 | x7 ;
  assign n23 = ( x1 & ~x2 ) | ( x1 & x5 ) | ( ~x2 & x5 ) ;
  assign n24 = ( ~n21 & n22 ) | ( ~n21 & n23 ) | ( n22 & n23 ) ;
  assign n25 = ( n19 & n20 ) | ( n19 & ~n24 ) | ( n20 & ~n24 ) ;
  assign n26 = x3 & x4 ;
  assign n27 = ( x3 & x4 ) | ( x3 & x7 ) | ( x4 & x7 ) ;
  assign n28 = ( x8 & ~n26 ) | ( x8 & n27 ) | ( ~n26 & n27 ) ;
  assign n29 = n25 | n28 ;
  assign n30 = x4 & x5 ;
  assign n31 = x4 | x5 ;
  assign n32 = ( x8 & n30 ) | ( x8 & ~n31 ) | ( n30 & ~n31 ) ;
  assign n33 = x9 | n32 ;
  assign n34 = ( n17 & n29 ) | ( n17 & ~n33 ) | ( n29 & ~n33 ) ;
  assign n35 = x8 & x9 ;
  assign n36 = x6 & x7 ;
  assign n37 = ~n35 & n36 ;
  assign n38 = ( x10 & ~n22 ) | ( x10 & n37 ) | ( ~n22 & n37 ) ;
  assign n39 = x5 & x6 ;
  assign n40 = ( x5 & x6 ) | ( x5 & x9 ) | ( x6 & x9 ) ;
  assign n41 = ( x10 & ~n39 ) | ( x10 & n40 ) | ( ~n39 & n40 ) ;
  assign n42 = ~n38 & n41 ;
  assign n43 = ( n34 & ~n38 ) | ( n34 & n42 ) | ( ~n38 & n42 ) ;
  assign n44 = x8 | n36 ;
  assign n45 = x8 & n37 ;
  assign n46 = ( x10 & ~n44 ) | ( x10 & n45 ) | ( ~n44 & n45 ) ;
  assign n47 = x6 & n30 ;
  assign n48 = ( x6 & x8 ) | ( x6 & n30 ) | ( x8 & n30 ) ;
  assign n49 = ( x9 & ~n47 ) | ( x9 & n48 ) | ( ~n47 & n48 ) ;
  assign n50 = x5 | n26 ;
  assign n51 = x5 & n26 ;
  assign n52 = ( x7 & ~n50 ) | ( x7 & n51 ) | ( ~n50 & n51 ) ;
  assign n53 = ( ~x4 & x6 ) | ( ~x4 & n12 ) | ( x6 & n12 ) ;
  assign n54 = ( ~x4 & x7 ) | ( ~x4 & n12 ) | ( x7 & n12 ) ;
  assign n55 = n53 & ~n54 ;
  assign n56 = ( ~x8 & n52 ) | ( ~x8 & n55 ) | ( n52 & n55 ) ;
  assign n57 = ( x8 & ~n49 ) | ( x8 & n56 ) | ( ~n49 & n56 ) ;
  assign n58 = x5 & n36 ;
  assign n59 = x7 | n39 ;
  assign n60 = ( x9 & n58 ) | ( x9 & ~n59 ) | ( n58 & ~n59 ) ;
  assign n61 = x1 & x2 ;
  assign n62 = x3 & ~n61 ;
  assign n63 = ( ~x3 & x8 ) | ( ~x3 & n61 ) | ( x8 & n61 ) ;
  assign n64 = ( x5 & n62 ) | ( x5 & n63 ) | ( n62 & n63 ) ;
  assign n65 = n22 | n64 ;
  assign n66 = x2 & x4 ;
  assign n67 = ~x0 & x4 ;
  assign n68 = x1 & ~n67 ;
  assign n69 = n66 & n68 ;
  assign n70 = ( ~x5 & n66 ) | ( ~x5 & n68 ) | ( n66 & n68 ) ;
  assign n71 = ( n65 & ~n69 ) | ( n65 & n70 ) | ( ~n69 & n70 ) ;
  assign n72 = ( n57 & ~n60 ) | ( n57 & n71 ) | ( ~n60 & n71 ) ;
  assign n73 = ( x10 & ~n57 ) | ( x10 & n72 ) | ( ~n57 & n72 ) ;
  assign n74 = ~n46 & n73 ;
  assign n75 = ~x7 & x9 ;
  assign n76 = ( x7 & n22 ) | ( x7 & n30 ) | ( n22 & n30 ) ;
  assign n77 = ( ~x10 & n58 ) | ( ~x10 & n76 ) | ( n58 & n76 ) ;
  assign n78 = ( ~n58 & n75 ) | ( ~n58 & n77 ) | ( n75 & n77 ) ;
  assign n79 = x8 & n78 ;
  assign n80 = ( n37 & n45 ) | ( n37 & n60 ) | ( n45 & n60 ) ;
  assign n81 = ( x9 & x10 ) | ( x9 & n80 ) | ( x10 & n80 ) ;
  assign n82 = n79 | n81 ;
  assign n83 = x9 | x10 ;
  assign n84 = ( x7 & n26 ) | ( x7 & ~n61 ) | ( n26 & ~n61 ) ;
  assign n85 = x0 & ~x6 ;
  assign n86 = ( n26 & n51 ) | ( n26 & n85 ) | ( n51 & n85 ) ;
  assign n87 = ~n84 & n86 ;
  assign n88 = n83 | n87 ;
  assign n89 = x8 | n22 ;
  assign n90 = ( x3 & n26 ) | ( x3 & n61 ) | ( n26 & n61 ) ;
  assign n91 = x2 & ~n31 ;
  assign n92 = ( ~n69 & n90 ) | ( ~n69 & n91 ) | ( n90 & n91 ) ;
  assign n93 = ( n69 & ~n89 ) | ( n69 & n92 ) | ( ~n89 & n92 ) ;
  assign n94 = ~n14 & n30 ;
  assign n95 = x5 | x6 ;
  assign n96 = ( x6 & n26 ) | ( x6 & n95 ) | ( n26 & n95 ) ;
  assign n97 = x7 & ~n47 ;
  assign n98 = ( x2 & n26 ) | ( x2 & n51 ) | ( n26 & n51 ) ;
  assign n99 = ( x5 & ~x8 ) | ( x5 & n98 ) | ( ~x8 & n98 ) ;
  assign n100 = ( ~n51 & n97 ) | ( ~n51 & n99 ) | ( n97 & n99 ) ;
  assign n101 = ( n94 & n96 ) | ( n94 & n100 ) | ( n96 & n100 ) ;
  assign n102 = n93 | n101 ;
  assign n103 = ~n88 & n102 ;
  assign n104 = n82 | n103 ;
  assign n105 = n32 & n58 ;
  assign n106 = n31 | n89 ;
  assign n107 = x3 | n66 ;
  assign n108 = n83 | n107 ;
  assign n109 = ( ~n105 & n106 ) | ( ~n105 & n108 ) | ( n106 & n108 ) ;
  assign n110 = ( x4 & x6 ) | ( x4 & ~n30 ) | ( x6 & ~n30 ) ;
  assign n111 = ~x7 & n110 ;
  assign n112 = ( n47 & n52 ) | ( n47 & n55 ) | ( n52 & n55 ) ;
  assign n113 = n87 | n112 ;
  assign n114 = n111 & ~n113 ;
  assign n115 = ( x8 & ~n111 ) | ( x8 & n113 ) | ( ~n111 & n113 ) ;
  assign n116 = n105 & n107 ;
  assign n117 = x9 | n116 ;
  assign n118 = ( n114 & n115 ) | ( n114 & ~n117 ) | ( n115 & ~n117 ) ;
  assign n119 = x10 | n35 ;
  assign n120 = ( x10 & n58 ) | ( x10 & n119 ) | ( n58 & n119 ) ;
  assign n121 = n118 | n120 ;
  assign n122 = n88 | n95 ;
  assign n123 = n13 | n112 ;
  assign n124 = ~n116 & n123 ;
  assign n125 = ( n83 & n122 ) | ( n83 & ~n124 ) | ( n122 & ~n124 ) ;
  assign n126 = n83 | n123 ;
  assign y0 = n43 ;
  assign y1 = n74 ;
  assign y2 = n104 ;
  assign y3 = n109 ;
  assign y4 = n121 ;
  assign y5 = n125 ;
  assign y6 = n126 ;
endmodule
