module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 ;
  assign n65 = ~x0 & x1 ;
  assign n66 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n67 = x1 & x2 ;
  assign n68 = n66 & ~n67 ;
  assign n69 = x0 & x3 ;
  assign n70 = x2 & ~n69 ;
  assign n71 = ~x2 & n69 ;
  assign n72 = ( ~n65 & n70 ) | ( ~n65 & n71 ) | ( n70 & n71 ) ;
  assign n73 = x2 & x4 ;
  assign n74 = n69 & n73 ;
  assign n75 = x1 & x4 ;
  assign n76 = ( n69 & n74 ) | ( n69 & n75 ) | ( n74 & n75 ) ;
  assign n77 = x1 & x3 ;
  assign n78 = x0 & x4 ;
  assign n79 = n77 | n78 ;
  assign n80 = n67 & ~n79 ;
  assign n81 = x2 & x3 ;
  assign n82 = x0 & n81 ;
  assign n83 = ( ~n67 & n79 ) | ( ~n67 & n82 ) | ( n79 & n82 ) ;
  assign n84 = ( ~n76 & n80 ) | ( ~n76 & n83 ) | ( n80 & n83 ) ;
  assign n85 = x1 & x5 ;
  assign n86 = n78 & n85 ;
  assign n87 = x0 & x5 ;
  assign n88 = ( ~n69 & n75 ) | ( ~n69 & n87 ) | ( n75 & n87 ) ;
  assign n89 = n69 & n87 ;
  assign n90 = ( ~n86 & n88 ) | ( ~n86 & n89 ) | ( n88 & n89 ) ;
  assign n91 = ~x2 & x3 ;
  assign n92 = ( n67 & n74 ) | ( n67 & n79 ) | ( n74 & n79 ) ;
  assign n93 = ( n90 & n91 ) | ( n90 & n92 ) | ( n91 & n92 ) ;
  assign n94 = ( ~n90 & n91 ) | ( ~n90 & n92 ) | ( n91 & n92 ) ;
  assign n95 = ( n90 & ~n93 ) | ( n90 & n94 ) | ( ~n93 & n94 ) ;
  assign n96 = ( n69 & n75 ) | ( n69 & n86 ) | ( n75 & n86 ) ;
  assign n97 = n73 | n85 ;
  assign n98 = x2 & x5 ;
  assign n99 = n75 & n98 ;
  assign n100 = n97 & ~n99 ;
  assign n101 = x0 & x6 ;
  assign n102 = ( ~n81 & n100 ) | ( ~n81 & n101 ) | ( n100 & n101 ) ;
  assign n103 = ( n81 & n100 ) | ( n81 & n101 ) | ( n100 & n101 ) ;
  assign n104 = ( n81 & n102 ) | ( n81 & ~n103 ) | ( n102 & ~n103 ) ;
  assign n105 = ( ~n93 & n96 ) | ( ~n93 & n104 ) | ( n96 & n104 ) ;
  assign n106 = ( n93 & n96 ) | ( n93 & n104 ) | ( n96 & n104 ) ;
  assign n107 = ( n93 & n105 ) | ( n93 & ~n106 ) | ( n105 & ~n106 ) ;
  assign n108 = ~x6 & n99 ;
  assign n109 = x1 & x6 ;
  assign n110 = x4 | n109 ;
  assign n111 = x4 & n109 ;
  assign n112 = ( n99 & n110 ) | ( n99 & ~n111 ) | ( n110 & ~n111 ) ;
  assign n113 = ( n103 & n108 ) | ( n103 & n112 ) | ( n108 & n112 ) ;
  assign n114 = n103 | n112 ;
  assign n115 = ~n113 & n114 ;
  assign n116 = x0 & x7 ;
  assign n117 = x3 & x4 ;
  assign n118 = ( ~n98 & n116 ) | ( ~n98 & n117 ) | ( n116 & n117 ) ;
  assign n119 = ( n98 & n116 ) | ( n98 & n117 ) | ( n116 & n117 ) ;
  assign n120 = ( n98 & n118 ) | ( n98 & ~n119 ) | ( n118 & ~n119 ) ;
  assign n121 = ( n106 & n115 ) | ( n106 & n120 ) | ( n115 & n120 ) ;
  assign n122 = ( ~n106 & n115 ) | ( ~n106 & n120 ) | ( n115 & n120 ) ;
  assign n123 = ( n106 & ~n121 ) | ( n106 & n122 ) | ( ~n121 & n122 ) ;
  assign n124 = x2 & x8 ;
  assign n125 = n101 & n124 ;
  assign n126 = x2 & x6 ;
  assign n127 = x0 & x8 ;
  assign n128 = n126 | n127 ;
  assign n129 = ( n111 & n125 ) | ( n111 & n128 ) | ( n125 & n128 ) ;
  assign n130 = ( ~n111 & n125 ) | ( ~n111 & n128 ) | ( n125 & n128 ) ;
  assign n131 = ( n111 & ~n129 ) | ( n111 & n130 ) | ( ~n129 & n130 ) ;
  assign n132 = x3 & x5 ;
  assign n133 = x1 & x7 ;
  assign n134 = n132 & n133 ;
  assign n135 = n132 | n133 ;
  assign n136 = ~n134 & n135 ;
  assign n137 = ( n119 & n131 ) | ( n119 & n136 ) | ( n131 & n136 ) ;
  assign n138 = ( ~n119 & n131 ) | ( ~n119 & n136 ) | ( n131 & n136 ) ;
  assign n139 = ( n119 & ~n137 ) | ( n119 & n138 ) | ( ~n137 & n138 ) ;
  assign n140 = ( ~n113 & n121 ) | ( ~n113 & n139 ) | ( n121 & n139 ) ;
  assign n141 = ( n113 & n121 ) | ( n113 & n139 ) | ( n121 & n139 ) ;
  assign n142 = ( n113 & n140 ) | ( n113 & ~n141 ) | ( n140 & ~n141 ) ;
  assign n143 = ~x1 & x5 ;
  assign n144 = x5 & x8 ;
  assign n145 = ( x1 & x5 ) | ( x1 & x8 ) | ( x5 & x8 ) ;
  assign n146 = ( n143 & ~n144 ) | ( n143 & n145 ) | ( ~n144 & n145 ) ;
  assign n147 = x0 & x9 ;
  assign n148 = ( n134 & n146 ) | ( n134 & n147 ) | ( n146 & n147 ) ;
  assign n149 = ( ~n134 & n146 ) | ( ~n134 & n147 ) | ( n146 & n147 ) ;
  assign n150 = ( n134 & ~n148 ) | ( n134 & n149 ) | ( ~n148 & n149 ) ;
  assign n151 = x2 & x7 ;
  assign n152 = x4 & x5 ;
  assign n153 = x3 & x6 ;
  assign n154 = ( ~n151 & n152 ) | ( ~n151 & n153 ) | ( n152 & n153 ) ;
  assign n155 = ( n151 & n152 ) | ( n151 & n153 ) | ( n152 & n153 ) ;
  assign n156 = ( n151 & n154 ) | ( n151 & ~n155 ) | ( n154 & ~n155 ) ;
  assign n157 = ( ~n129 & n150 ) | ( ~n129 & n156 ) | ( n150 & n156 ) ;
  assign n158 = ( n129 & n150 ) | ( n129 & n156 ) | ( n150 & n156 ) ;
  assign n159 = ( n129 & n157 ) | ( n129 & ~n158 ) | ( n157 & ~n158 ) ;
  assign n160 = ( ~n137 & n141 ) | ( ~n137 & n159 ) | ( n141 & n159 ) ;
  assign n161 = ( n137 & n141 ) | ( n137 & n159 ) | ( n141 & n159 ) ;
  assign n162 = ( n137 & n160 ) | ( n137 & ~n161 ) | ( n160 & ~n161 ) ;
  assign n163 = x1 & n144 ;
  assign n164 = ~x1 & x9 ;
  assign n165 = x4 & x6 ;
  assign n166 = ( x9 & n164 ) | ( x9 & n165 ) | ( n164 & n165 ) ;
  assign n167 = ( x9 & ~n164 ) | ( x9 & n165 ) | ( ~n164 & n165 ) ;
  assign n168 = ( n164 & ~n166 ) | ( n164 & n167 ) | ( ~n166 & n167 ) ;
  assign n169 = ( n155 & n163 ) | ( n155 & n168 ) | ( n163 & n168 ) ;
  assign n170 = ( n155 & ~n163 ) | ( n155 & n168 ) | ( ~n163 & n168 ) ;
  assign n171 = ( n163 & ~n169 ) | ( n163 & n170 ) | ( ~n169 & n170 ) ;
  assign n172 = x3 & x7 ;
  assign n173 = x0 & x10 ;
  assign n174 = ( ~n124 & n172 ) | ( ~n124 & n173 ) | ( n172 & n173 ) ;
  assign n175 = ( n124 & n172 ) | ( n124 & n173 ) | ( n172 & n173 ) ;
  assign n176 = ( n124 & n174 ) | ( n124 & ~n175 ) | ( n174 & ~n175 ) ;
  assign n177 = ( ~n148 & n171 ) | ( ~n148 & n176 ) | ( n171 & n176 ) ;
  assign n178 = ( n148 & n171 ) | ( n148 & n176 ) | ( n171 & n176 ) ;
  assign n179 = ( n148 & n177 ) | ( n148 & ~n178 ) | ( n177 & ~n178 ) ;
  assign n180 = ( n158 & n161 ) | ( n158 & n179 ) | ( n161 & n179 ) ;
  assign n181 = ( ~n158 & n161 ) | ( ~n158 & n179 ) | ( n161 & n179 ) ;
  assign n182 = ( n158 & ~n180 ) | ( n158 & n181 ) | ( ~n180 & n181 ) ;
  assign n183 = x2 & x9 ;
  assign n184 = x3 & x8 ;
  assign n185 = n183 | n184 ;
  assign n186 = x4 & x9 ;
  assign n187 = n109 & n186 ;
  assign n188 = x3 & x9 ;
  assign n189 = n124 & n188 ;
  assign n190 = ( ~n185 & n187 ) | ( ~n185 & n189 ) | ( n187 & n189 ) ;
  assign n191 = ( n185 & n187 ) | ( n185 & n189 ) | ( n187 & n189 ) ;
  assign n192 = ( n185 & n190 ) | ( n185 & ~n191 ) | ( n190 & ~n191 ) ;
  assign n193 = ~x1 & x6 ;
  assign n194 = ( x1 & x6 ) | ( x1 & x10 ) | ( x6 & x10 ) ;
  assign n195 = x6 & x10 ;
  assign n196 = ( n193 & n194 ) | ( n193 & ~n195 ) | ( n194 & ~n195 ) ;
  assign n197 = ( ~n175 & n192 ) | ( ~n175 & n196 ) | ( n192 & n196 ) ;
  assign n198 = ( n175 & n192 ) | ( n175 & n196 ) | ( n192 & n196 ) ;
  assign n199 = ( n175 & n197 ) | ( n175 & ~n198 ) | ( n197 & ~n198 ) ;
  assign n200 = x0 & x11 ;
  assign n201 = x5 & x6 ;
  assign n202 = x4 & x7 ;
  assign n203 = ( ~n200 & n201 ) | ( ~n200 & n202 ) | ( n201 & n202 ) ;
  assign n204 = ( n200 & n201 ) | ( n200 & n202 ) | ( n201 & n202 ) ;
  assign n205 = ( n200 & n203 ) | ( n200 & ~n204 ) | ( n203 & ~n204 ) ;
  assign n206 = ( ~n169 & n199 ) | ( ~n169 & n205 ) | ( n199 & n205 ) ;
  assign n207 = ( n169 & n199 ) | ( n169 & n205 ) | ( n199 & n205 ) ;
  assign n208 = ( n169 & n206 ) | ( n169 & ~n207 ) | ( n206 & ~n207 ) ;
  assign n209 = ( n178 & n180 ) | ( n178 & n208 ) | ( n180 & n208 ) ;
  assign n210 = ( ~n178 & n180 ) | ( ~n178 & n208 ) | ( n180 & n208 ) ;
  assign n211 = ( n178 & ~n209 ) | ( n178 & n210 ) | ( ~n209 & n210 ) ;
  assign n212 = x10 & n109 ;
  assign n213 = x4 & x8 ;
  assign n214 = x5 & x11 ;
  assign n215 = n133 & n214 ;
  assign n216 = x1 & x11 ;
  assign n217 = ~x11 & n85 ;
  assign n218 = ( x7 & n143 ) | ( x7 & n217 ) | ( n143 & n217 ) ;
  assign n219 = ( ~n215 & n216 ) | ( ~n215 & n218 ) | ( n216 & n218 ) ;
  assign n220 = ( n212 & n213 ) | ( n212 & n219 ) | ( n213 & n219 ) ;
  assign n221 = ( ~n212 & n213 ) | ( ~n212 & n219 ) | ( n213 & n219 ) ;
  assign n222 = ( n212 & ~n220 ) | ( n212 & n221 ) | ( ~n220 & n221 ) ;
  assign n223 = x0 & x12 ;
  assign n224 = x2 & x10 ;
  assign n225 = ( ~n188 & n223 ) | ( ~n188 & n224 ) | ( n223 & n224 ) ;
  assign n226 = ( n188 & n223 ) | ( n188 & n224 ) | ( n223 & n224 ) ;
  assign n227 = ( n188 & n225 ) | ( n188 & ~n226 ) | ( n225 & ~n226 ) ;
  assign n228 = ( n191 & n204 ) | ( n191 & n227 ) | ( n204 & n227 ) ;
  assign n229 = ( n191 & ~n204 ) | ( n191 & n227 ) | ( ~n204 & n227 ) ;
  assign n230 = ( n204 & ~n228 ) | ( n204 & n229 ) | ( ~n228 & n229 ) ;
  assign n231 = ( ~n198 & n222 ) | ( ~n198 & n230 ) | ( n222 & n230 ) ;
  assign n232 = ( n198 & n222 ) | ( n198 & n230 ) | ( n222 & n230 ) ;
  assign n233 = ( n198 & n231 ) | ( n198 & ~n232 ) | ( n231 & ~n232 ) ;
  assign n234 = ( n207 & n209 ) | ( n207 & n233 ) | ( n209 & n233 ) ;
  assign n235 = ( ~n207 & n209 ) | ( ~n207 & n233 ) | ( n209 & n233 ) ;
  assign n236 = ( n207 & ~n234 ) | ( n207 & n235 ) | ( ~n234 & n235 ) ;
  assign n237 = x2 & x11 ;
  assign n238 = x6 & x7 ;
  assign n239 = ( ~n144 & n237 ) | ( ~n144 & n238 ) | ( n237 & n238 ) ;
  assign n240 = ( n144 & n237 ) | ( n144 & n238 ) | ( n237 & n238 ) ;
  assign n241 = ( n144 & n239 ) | ( n144 & ~n240 ) | ( n239 & ~n240 ) ;
  assign n242 = x3 & x10 ;
  assign n243 = x0 & x13 ;
  assign n244 = ( ~n186 & n242 ) | ( ~n186 & n243 ) | ( n242 & n243 ) ;
  assign n245 = ( n186 & n242 ) | ( n186 & n243 ) | ( n242 & n243 ) ;
  assign n246 = ( n186 & n244 ) | ( n186 & ~n245 ) | ( n244 & ~n245 ) ;
  assign n247 = ( n220 & n241 ) | ( n220 & n246 ) | ( n241 & n246 ) ;
  assign n248 = ( ~n220 & n241 ) | ( ~n220 & n246 ) | ( n241 & n246 ) ;
  assign n249 = ( n220 & ~n247 ) | ( n220 & n248 ) | ( ~n247 & n248 ) ;
  assign n250 = ~x12 & n215 ;
  assign n251 = x1 & x12 ;
  assign n252 = x7 | n251 ;
  assign n253 = x12 & n133 ;
  assign n254 = ( n215 & n252 ) | ( n215 & ~n253 ) | ( n252 & ~n253 ) ;
  assign n255 = ( n226 & n250 ) | ( n226 & n254 ) | ( n250 & n254 ) ;
  assign n256 = ( ~n226 & n250 ) | ( ~n226 & n254 ) | ( n250 & n254 ) ;
  assign n257 = ( n226 & ~n255 ) | ( n226 & n256 ) | ( ~n255 & n256 ) ;
  assign n258 = ( n228 & n232 ) | ( n228 & n257 ) | ( n232 & n257 ) ;
  assign n259 = ( ~n228 & n232 ) | ( ~n228 & n257 ) | ( n232 & n257 ) ;
  assign n260 = ( n228 & ~n258 ) | ( n228 & n259 ) | ( ~n258 & n259 ) ;
  assign n261 = ( ~n234 & n249 ) | ( ~n234 & n260 ) | ( n249 & n260 ) ;
  assign n262 = ( n234 & n249 ) | ( n234 & n260 ) | ( n249 & n260 ) ;
  assign n263 = ( n234 & n261 ) | ( n234 & ~n262 ) | ( n261 & ~n262 ) ;
  assign n264 = x6 & x8 ;
  assign n265 = x1 & x13 ;
  assign n266 = n264 & n265 ;
  assign n267 = n264 | n265 ;
  assign n268 = ~n266 & n267 ;
  assign n269 = ( n240 & n245 ) | ( n240 & n268 ) | ( n245 & n268 ) ;
  assign n270 = ( n240 & n245 ) | ( n240 & ~n268 ) | ( n245 & ~n268 ) ;
  assign n271 = ( n268 & ~n269 ) | ( n268 & n270 ) | ( ~n269 & n270 ) ;
  assign n272 = x4 & x10 ;
  assign n273 = x5 & x9 ;
  assign n274 = n272 | n273 ;
  assign n275 = x5 & x10 ;
  assign n276 = n186 & n275 ;
  assign n277 = ( n253 & n274 ) | ( n253 & n276 ) | ( n274 & n276 ) ;
  assign n278 = ( ~n253 & n274 ) | ( ~n253 & n276 ) | ( n274 & n276 ) ;
  assign n279 = ( n253 & ~n277 ) | ( n253 & n278 ) | ( ~n277 & n278 ) ;
  assign n280 = x0 & x14 ;
  assign n281 = x2 & x12 ;
  assign n282 = x3 & x11 ;
  assign n283 = ( ~n280 & n281 ) | ( ~n280 & n282 ) | ( n281 & n282 ) ;
  assign n284 = ( n280 & n281 ) | ( n280 & n282 ) | ( n281 & n282 ) ;
  assign n285 = ( n280 & n283 ) | ( n280 & ~n284 ) | ( n283 & ~n284 ) ;
  assign n286 = ( ~n255 & n279 ) | ( ~n255 & n285 ) | ( n279 & n285 ) ;
  assign n287 = ( n255 & n279 ) | ( n255 & n285 ) | ( n279 & n285 ) ;
  assign n288 = ( n255 & n286 ) | ( n255 & ~n287 ) | ( n286 & ~n287 ) ;
  assign n289 = ( n247 & n271 ) | ( n247 & n288 ) | ( n271 & n288 ) ;
  assign n290 = ( ~n247 & n271 ) | ( ~n247 & n288 ) | ( n271 & n288 ) ;
  assign n291 = ( n247 & ~n289 ) | ( n247 & n290 ) | ( ~n289 & n290 ) ;
  assign n292 = ( n258 & n262 ) | ( n258 & n291 ) | ( n262 & n291 ) ;
  assign n293 = ( ~n258 & n262 ) | ( ~n258 & n291 ) | ( n262 & n291 ) ;
  assign n294 = ( n258 & ~n292 ) | ( n258 & n293 ) | ( ~n292 & n293 ) ;
  assign n295 = x4 & x11 ;
  assign n296 = x1 & x14 ;
  assign n297 = x8 & n296 ;
  assign n298 = x8 | n296 ;
  assign n299 = ~n297 & n298 ;
  assign n300 = ( n266 & n295 ) | ( n266 & n299 ) | ( n295 & n299 ) ;
  assign n301 = ( ~n266 & n295 ) | ( ~n266 & n299 ) | ( n295 & n299 ) ;
  assign n302 = ( n266 & ~n300 ) | ( n266 & n301 ) | ( ~n300 & n301 ) ;
  assign n303 = x2 & x13 ;
  assign n304 = x7 & x8 ;
  assign n305 = x6 & x9 ;
  assign n306 = ( ~n303 & n304 ) | ( ~n303 & n305 ) | ( n304 & n305 ) ;
  assign n307 = ( n303 & n304 ) | ( n303 & n305 ) | ( n304 & n305 ) ;
  assign n308 = ( n303 & n306 ) | ( n303 & ~n307 ) | ( n306 & ~n307 ) ;
  assign n309 = ( ~n269 & n302 ) | ( ~n269 & n308 ) | ( n302 & n308 ) ;
  assign n310 = ( n269 & n302 ) | ( n269 & n308 ) | ( n302 & n308 ) ;
  assign n311 = ( n269 & n309 ) | ( n269 & ~n310 ) | ( n309 & ~n310 ) ;
  assign n312 = x3 & x12 ;
  assign n313 = x0 & x15 ;
  assign n314 = ( ~n275 & n312 ) | ( ~n275 & n313 ) | ( n312 & n313 ) ;
  assign n315 = ( n275 & n312 ) | ( n275 & n313 ) | ( n312 & n313 ) ;
  assign n316 = ( n275 & n314 ) | ( n275 & ~n315 ) | ( n314 & ~n315 ) ;
  assign n317 = ( n277 & n284 ) | ( n277 & n316 ) | ( n284 & n316 ) ;
  assign n318 = ( ~n277 & n284 ) | ( ~n277 & n316 ) | ( n284 & n316 ) ;
  assign n319 = ( n277 & ~n317 ) | ( n277 & n318 ) | ( ~n317 & n318 ) ;
  assign n320 = ( ~n287 & n311 ) | ( ~n287 & n319 ) | ( n311 & n319 ) ;
  assign n321 = ( n287 & n311 ) | ( n287 & n319 ) | ( n311 & n319 ) ;
  assign n322 = ( n287 & n320 ) | ( n287 & ~n321 ) | ( n320 & ~n321 ) ;
  assign n323 = ( ~n289 & n292 ) | ( ~n289 & n322 ) | ( n292 & n322 ) ;
  assign n324 = ( n289 & n292 ) | ( n289 & n322 ) | ( n292 & n322 ) ;
  assign n325 = ( n289 & n323 ) | ( n289 & ~n324 ) | ( n323 & ~n324 ) ;
  assign n326 = x4 & x12 ;
  assign n327 = x3 & x13 ;
  assign n328 = x2 & x14 ;
  assign n329 = ( ~n326 & n327 ) | ( ~n326 & n328 ) | ( n327 & n328 ) ;
  assign n330 = ( n326 & n327 ) | ( n326 & n328 ) | ( n327 & n328 ) ;
  assign n331 = ( n326 & n329 ) | ( n326 & ~n330 ) | ( n329 & ~n330 ) ;
  assign n332 = x7 & x9 ;
  assign n333 = x1 & x15 ;
  assign n334 = n332 & n333 ;
  assign n335 = n332 | n333 ;
  assign n336 = ~n334 & n335 ;
  assign n337 = ( ~n297 & n307 ) | ( ~n297 & n336 ) | ( n307 & n336 ) ;
  assign n338 = ( n297 & n307 ) | ( n297 & n336 ) | ( n307 & n336 ) ;
  assign n339 = ( n297 & n337 ) | ( n297 & ~n338 ) | ( n337 & ~n338 ) ;
  assign n340 = ( n317 & n331 ) | ( n317 & n339 ) | ( n331 & n339 ) ;
  assign n341 = ( ~n317 & n331 ) | ( ~n317 & n339 ) | ( n331 & n339 ) ;
  assign n342 = ( n317 & ~n340 ) | ( n317 & n341 ) | ( ~n340 & n341 ) ;
  assign n343 = x0 & x16 ;
  assign n344 = ( n195 & n214 ) | ( n195 & n343 ) | ( n214 & n343 ) ;
  assign n345 = ( ~n195 & n214 ) | ( ~n195 & n343 ) | ( n214 & n343 ) ;
  assign n346 = ( n195 & ~n344 ) | ( n195 & n345 ) | ( ~n344 & n345 ) ;
  assign n347 = ( n300 & n315 ) | ( n300 & n346 ) | ( n315 & n346 ) ;
  assign n348 = ( ~n300 & n315 ) | ( ~n300 & n346 ) | ( n315 & n346 ) ;
  assign n349 = ( n300 & ~n347 ) | ( n300 & n348 ) | ( ~n347 & n348 ) ;
  assign n350 = ( n310 & n342 ) | ( n310 & n349 ) | ( n342 & n349 ) ;
  assign n351 = ( ~n310 & n342 ) | ( ~n310 & n349 ) | ( n342 & n349 ) ;
  assign n352 = ( n310 & ~n350 ) | ( n310 & n351 ) | ( ~n350 & n351 ) ;
  assign n353 = ( n321 & n324 ) | ( n321 & n352 ) | ( n324 & n352 ) ;
  assign n354 = ( ~n321 & n324 ) | ( ~n321 & n352 ) | ( n324 & n352 ) ;
  assign n355 = ( n321 & ~n353 ) | ( n321 & n354 ) | ( ~n353 & n354 ) ;
  assign n356 = x9 & x16 ;
  assign n357 = ( x1 & x9 ) | ( x1 & x16 ) | ( x9 & x16 ) ;
  assign n358 = ( n164 & ~n356 ) | ( n164 & n357 ) | ( ~n356 & n357 ) ;
  assign n359 = ( n330 & n344 ) | ( n330 & n358 ) | ( n344 & n358 ) ;
  assign n360 = ( n330 & n344 ) | ( n330 & ~n358 ) | ( n344 & ~n358 ) ;
  assign n361 = ( n358 & ~n359 ) | ( n358 & n360 ) | ( ~n359 & n360 ) ;
  assign n362 = ( n338 & n347 ) | ( n338 & n361 ) | ( n347 & n361 ) ;
  assign n363 = ( ~n338 & n347 ) | ( ~n338 & n361 ) | ( n347 & n361 ) ;
  assign n364 = ( n338 & ~n362 ) | ( n338 & n363 ) | ( ~n362 & n363 ) ;
  assign n365 = x5 & x12 ;
  assign n366 = x0 & x17 ;
  assign n367 = ( ~n334 & n365 ) | ( ~n334 & n366 ) | ( n365 & n366 ) ;
  assign n368 = ( n334 & n365 ) | ( n334 & n366 ) | ( n365 & n366 ) ;
  assign n369 = ( n334 & n367 ) | ( n334 & ~n368 ) | ( n367 & ~n368 ) ;
  assign n370 = x3 & x14 ;
  assign n371 = x8 & x9 ;
  assign n372 = x7 & x10 ;
  assign n373 = ( ~n370 & n371 ) | ( ~n370 & n372 ) | ( n371 & n372 ) ;
  assign n374 = ( n370 & n371 ) | ( n370 & n372 ) | ( n371 & n372 ) ;
  assign n375 = ( n370 & n373 ) | ( n370 & ~n374 ) | ( n373 & ~n374 ) ;
  assign n376 = x6 & x11 ;
  assign n377 = x4 & x13 ;
  assign n378 = x2 & x15 ;
  assign n379 = ( ~n376 & n377 ) | ( ~n376 & n378 ) | ( n377 & n378 ) ;
  assign n380 = ( n376 & n377 ) | ( n376 & n378 ) | ( n377 & n378 ) ;
  assign n381 = ( n376 & n379 ) | ( n376 & ~n380 ) | ( n379 & ~n380 ) ;
  assign n382 = ( ~n369 & n375 ) | ( ~n369 & n381 ) | ( n375 & n381 ) ;
  assign n383 = ( n369 & n375 ) | ( n369 & n381 ) | ( n375 & n381 ) ;
  assign n384 = ( n369 & n382 ) | ( n369 & ~n383 ) | ( n382 & ~n383 ) ;
  assign n385 = ( ~n340 & n364 ) | ( ~n340 & n384 ) | ( n364 & n384 ) ;
  assign n386 = ( n340 & n364 ) | ( n340 & n384 ) | ( n364 & n384 ) ;
  assign n387 = ( n340 & n385 ) | ( n340 & ~n386 ) | ( n385 & ~n386 ) ;
  assign n388 = ( n350 & n353 ) | ( n350 & n387 ) | ( n353 & n387 ) ;
  assign n389 = ( ~n350 & n353 ) | ( ~n350 & n387 ) | ( n353 & n387 ) ;
  assign n390 = ( n350 & ~n388 ) | ( n350 & n389 ) | ( ~n388 & n389 ) ;
  assign n391 = ( ~n368 & n374 ) | ( ~n368 & n380 ) | ( n374 & n380 ) ;
  assign n392 = ( n368 & n374 ) | ( n368 & n380 ) | ( n374 & n380 ) ;
  assign n393 = ( n368 & n391 ) | ( n368 & ~n392 ) | ( n391 & ~n392 ) ;
  assign n394 = ( ~n359 & n383 ) | ( ~n359 & n393 ) | ( n383 & n393 ) ;
  assign n395 = ( n359 & n383 ) | ( n359 & n393 ) | ( n383 & n393 ) ;
  assign n396 = ( n359 & n394 ) | ( n359 & ~n395 ) | ( n394 & ~n395 ) ;
  assign n397 = x4 & x14 ;
  assign n398 = x3 & x15 ;
  assign n399 = x2 & x16 ;
  assign n400 = ( ~n397 & n398 ) | ( ~n397 & n399 ) | ( n398 & n399 ) ;
  assign n401 = ( n397 & n398 ) | ( n397 & n399 ) | ( n398 & n399 ) ;
  assign n402 = ( n397 & n400 ) | ( n397 & ~n401 ) | ( n400 & ~n401 ) ;
  assign n403 = x7 & x11 ;
  assign n404 = x0 & x18 ;
  assign n405 = x5 & x13 ;
  assign n406 = ( ~n403 & n404 ) | ( ~n403 & n405 ) | ( n404 & n405 ) ;
  assign n407 = ( n403 & n404 ) | ( n403 & n405 ) | ( n404 & n405 ) ;
  assign n408 = ( n403 & n406 ) | ( n403 & ~n407 ) | ( n406 & ~n407 ) ;
  assign n409 = x1 & n356 ;
  assign n410 = x8 & x10 ;
  assign n411 = x1 & x17 ;
  assign n412 = n410 & n411 ;
  assign n413 = n410 | n411 ;
  assign n414 = ~n412 & n413 ;
  assign n415 = x6 & x12 ;
  assign n416 = ( n409 & n414 ) | ( n409 & n415 ) | ( n414 & n415 ) ;
  assign n417 = ( ~n409 & n414 ) | ( ~n409 & n415 ) | ( n414 & n415 ) ;
  assign n418 = ( n409 & ~n416 ) | ( n409 & n417 ) | ( ~n416 & n417 ) ;
  assign n419 = ( ~n402 & n408 ) | ( ~n402 & n418 ) | ( n408 & n418 ) ;
  assign n420 = ( n402 & n408 ) | ( n402 & n418 ) | ( n408 & n418 ) ;
  assign n421 = ( n402 & n419 ) | ( n402 & ~n420 ) | ( n419 & ~n420 ) ;
  assign n422 = ( ~n362 & n396 ) | ( ~n362 & n421 ) | ( n396 & n421 ) ;
  assign n423 = ( n362 & n396 ) | ( n362 & n421 ) | ( n396 & n421 ) ;
  assign n424 = ( n362 & n422 ) | ( n362 & ~n423 ) | ( n422 & ~n423 ) ;
  assign n425 = ( ~n386 & n388 ) | ( ~n386 & n424 ) | ( n388 & n424 ) ;
  assign n426 = ( n386 & n388 ) | ( n386 & n424 ) | ( n388 & n424 ) ;
  assign n427 = ( n386 & n425 ) | ( n386 & ~n426 ) | ( n425 & ~n426 ) ;
  assign n428 = x3 & x16 ;
  assign n429 = x9 & x10 ;
  assign n430 = x8 & x11 ;
  assign n431 = ( ~n428 & n429 ) | ( ~n428 & n430 ) | ( n429 & n430 ) ;
  assign n432 = ( n428 & n429 ) | ( n428 & n430 ) | ( n429 & n430 ) ;
  assign n433 = ( n428 & n431 ) | ( n428 & ~n432 ) | ( n431 & ~n432 ) ;
  assign n434 = ( ~n407 & n416 ) | ( ~n407 & n433 ) | ( n416 & n433 ) ;
  assign n435 = ( n407 & n416 ) | ( n407 & n433 ) | ( n416 & n433 ) ;
  assign n436 = ( n407 & n434 ) | ( n407 & ~n435 ) | ( n434 & ~n435 ) ;
  assign n437 = ~x18 & n412 ;
  assign n438 = n401 & n437 ;
  assign n439 = x1 & x18 ;
  assign n440 = x10 | n439 ;
  assign n441 = x10 & n439 ;
  assign n442 = ( n412 & n440 ) | ( n412 & ~n441 ) | ( n440 & ~n441 ) ;
  assign n443 = ( n401 & n437 ) | ( n401 & n442 ) | ( n437 & n442 ) ;
  assign n444 = n401 | n442 ;
  assign n445 = ( n438 & ~n443 ) | ( n438 & n444 ) | ( ~n443 & n444 ) ;
  assign n446 = ( ~n420 & n436 ) | ( ~n420 & n445 ) | ( n436 & n445 ) ;
  assign n447 = ( n420 & n436 ) | ( n420 & n445 ) | ( n436 & n445 ) ;
  assign n448 = ( n420 & n446 ) | ( n420 & ~n447 ) | ( n446 & ~n447 ) ;
  assign n449 = x0 & x19 ;
  assign n450 = x4 & x15 ;
  assign n451 = x2 & x17 ;
  assign n452 = ( ~n449 & n450 ) | ( ~n449 & n451 ) | ( n450 & n451 ) ;
  assign n453 = ( n449 & n450 ) | ( n449 & n451 ) | ( n450 & n451 ) ;
  assign n454 = ( n449 & n452 ) | ( n449 & ~n453 ) | ( n452 & ~n453 ) ;
  assign n455 = x5 & x14 ;
  assign n456 = x7 & x12 ;
  assign n457 = x6 & x13 ;
  assign n458 = ( ~n455 & n456 ) | ( ~n455 & n457 ) | ( n456 & n457 ) ;
  assign n459 = ( n455 & n456 ) | ( n455 & n457 ) | ( n456 & n457 ) ;
  assign n460 = ( n455 & n458 ) | ( n455 & ~n459 ) | ( n458 & ~n459 ) ;
  assign n461 = ( n392 & n454 ) | ( n392 & n460 ) | ( n454 & n460 ) ;
  assign n462 = ( ~n392 & n454 ) | ( ~n392 & n460 ) | ( n454 & n460 ) ;
  assign n463 = ( n392 & ~n461 ) | ( n392 & n462 ) | ( ~n461 & n462 ) ;
  assign n464 = ( ~n395 & n448 ) | ( ~n395 & n463 ) | ( n448 & n463 ) ;
  assign n465 = ( n395 & n448 ) | ( n395 & n463 ) | ( n448 & n463 ) ;
  assign n466 = ( n395 & n464 ) | ( n395 & ~n465 ) | ( n464 & ~n465 ) ;
  assign n467 = ( ~n423 & n426 ) | ( ~n423 & n466 ) | ( n426 & n466 ) ;
  assign n468 = ( n423 & n426 ) | ( n423 & n466 ) | ( n426 & n466 ) ;
  assign n469 = ( n423 & n467 ) | ( n423 & ~n468 ) | ( n467 & ~n468 ) ;
  assign n470 = x9 & x11 ;
  assign n471 = x1 & x19 ;
  assign n472 = n470 & n471 ;
  assign n473 = n470 | n471 ;
  assign n474 = ~n472 & n473 ;
  assign n475 = ( n432 & n453 ) | ( n432 & n474 ) | ( n453 & n474 ) ;
  assign n476 = ( ~n432 & n453 ) | ( ~n432 & n474 ) | ( n453 & n474 ) ;
  assign n477 = ( n432 & ~n475 ) | ( n432 & n476 ) | ( ~n475 & n476 ) ;
  assign n478 = x7 & x13 ;
  assign n479 = x0 & x20 ;
  assign n480 = ( ~n441 & n478 ) | ( ~n441 & n479 ) | ( n478 & n479 ) ;
  assign n481 = ( n441 & n478 ) | ( n441 & n479 ) | ( n478 & n479 ) ;
  assign n482 = ( n441 & n480 ) | ( n441 & ~n481 ) | ( n480 & ~n481 ) ;
  assign n483 = x8 & x12 ;
  assign n484 = x5 & x15 ;
  assign n485 = x6 & x14 ;
  assign n486 = ( ~n483 & n484 ) | ( ~n483 & n485 ) | ( n484 & n485 ) ;
  assign n487 = ( n483 & n484 ) | ( n483 & n485 ) | ( n484 & n485 ) ;
  assign n488 = ( n483 & n486 ) | ( n483 & ~n487 ) | ( n486 & ~n487 ) ;
  assign n489 = ( n459 & n482 ) | ( n459 & n488 ) | ( n482 & n488 ) ;
  assign n490 = ( ~n459 & n482 ) | ( ~n459 & n488 ) | ( n482 & n488 ) ;
  assign n491 = ( n459 & ~n489 ) | ( n459 & n490 ) | ( ~n489 & n490 ) ;
  assign n492 = ( ~n461 & n477 ) | ( ~n461 & n491 ) | ( n477 & n491 ) ;
  assign n493 = ( n461 & n477 ) | ( n461 & n491 ) | ( n477 & n491 ) ;
  assign n494 = ( n461 & n492 ) | ( n461 & ~n493 ) | ( n492 & ~n493 ) ;
  assign n495 = x2 & x18 ;
  assign n496 = x3 & x17 ;
  assign n497 = x4 & x16 ;
  assign n498 = ( ~n495 & n496 ) | ( ~n495 & n497 ) | ( n496 & n497 ) ;
  assign n499 = ( n495 & n496 ) | ( n495 & n497 ) | ( n496 & n497 ) ;
  assign n500 = ( n495 & n498 ) | ( n495 & ~n499 ) | ( n498 & ~n499 ) ;
  assign n501 = ( n435 & n443 ) | ( n435 & n500 ) | ( n443 & n500 ) ;
  assign n502 = ( ~n435 & n443 ) | ( ~n435 & n500 ) | ( n443 & n500 ) ;
  assign n503 = ( n435 & ~n501 ) | ( n435 & n502 ) | ( ~n501 & n502 ) ;
  assign n504 = ( n447 & n494 ) | ( n447 & n503 ) | ( n494 & n503 ) ;
  assign n505 = ( ~n447 & n494 ) | ( ~n447 & n503 ) | ( n494 & n503 ) ;
  assign n506 = ( n447 & ~n504 ) | ( n447 & n505 ) | ( ~n504 & n505 ) ;
  assign n507 = ( n465 & n468 ) | ( n465 & n506 ) | ( n468 & n506 ) ;
  assign n508 = ( ~n465 & n468 ) | ( ~n465 & n506 ) | ( n468 & n506 ) ;
  assign n509 = ( n465 & ~n507 ) | ( n465 & n508 ) | ( ~n507 & n508 ) ;
  assign n510 = ( ~n481 & n487 ) | ( ~n481 & n499 ) | ( n487 & n499 ) ;
  assign n511 = ( n481 & n487 ) | ( n481 & n499 ) | ( n487 & n499 ) ;
  assign n512 = ( n481 & n510 ) | ( n481 & ~n511 ) | ( n510 & ~n511 ) ;
  assign n513 = x5 & x16 ;
  assign n514 = x2 & x19 ;
  assign n515 = x3 & x18 ;
  assign n516 = ( ~n513 & n514 ) | ( ~n513 & n515 ) | ( n514 & n515 ) ;
  assign n517 = ( n513 & n514 ) | ( n513 & n515 ) | ( n514 & n515 ) ;
  assign n518 = ( n513 & n516 ) | ( n513 & ~n517 ) | ( n516 & ~n517 ) ;
  assign n519 = x4 & x17 ;
  assign n520 = x10 & x11 ;
  assign n521 = x9 & x12 ;
  assign n522 = ( ~n519 & n520 ) | ( ~n519 & n521 ) | ( n520 & n521 ) ;
  assign n523 = ( n519 & n520 ) | ( n519 & n521 ) | ( n520 & n521 ) ;
  assign n524 = ( n519 & n522 ) | ( n519 & ~n523 ) | ( n522 & ~n523 ) ;
  assign n525 = x6 & x15 ;
  assign n526 = x8 & x13 ;
  assign n527 = x7 & x14 ;
  assign n528 = ( ~n525 & n526 ) | ( ~n525 & n527 ) | ( n526 & n527 ) ;
  assign n529 = ( n525 & n526 ) | ( n525 & n527 ) | ( n526 & n527 ) ;
  assign n530 = ( n525 & n528 ) | ( n525 & ~n529 ) | ( n528 & ~n529 ) ;
  assign n531 = ( ~n518 & n524 ) | ( ~n518 & n530 ) | ( n524 & n530 ) ;
  assign n532 = ( n518 & n524 ) | ( n518 & n530 ) | ( n524 & n530 ) ;
  assign n533 = ( n518 & n531 ) | ( n518 & ~n532 ) | ( n531 & ~n532 ) ;
  assign n534 = ( ~n501 & n512 ) | ( ~n501 & n533 ) | ( n512 & n533 ) ;
  assign n535 = ( n501 & n512 ) | ( n501 & n533 ) | ( n512 & n533 ) ;
  assign n536 = ( n501 & n534 ) | ( n501 & ~n535 ) | ( n534 & ~n535 ) ;
  assign n537 = x0 & x21 ;
  assign n538 = x1 & x20 ;
  assign n539 = x11 & n538 ;
  assign n540 = x11 | n538 ;
  assign n541 = ~n539 & n540 ;
  assign n542 = ( n472 & n537 ) | ( n472 & n541 ) | ( n537 & n541 ) ;
  assign n543 = ( ~n472 & n537 ) | ( ~n472 & n541 ) | ( n537 & n541 ) ;
  assign n544 = ( n472 & ~n542 ) | ( n472 & n543 ) | ( ~n542 & n543 ) ;
  assign n545 = ( n475 & n489 ) | ( n475 & n544 ) | ( n489 & n544 ) ;
  assign n546 = ( ~n475 & n489 ) | ( ~n475 & n544 ) | ( n489 & n544 ) ;
  assign n547 = ( n475 & ~n545 ) | ( n475 & n546 ) | ( ~n545 & n546 ) ;
  assign n548 = ( ~n493 & n536 ) | ( ~n493 & n547 ) | ( n536 & n547 ) ;
  assign n549 = ( n493 & n536 ) | ( n493 & n547 ) | ( n536 & n547 ) ;
  assign n550 = ( n493 & n548 ) | ( n493 & ~n549 ) | ( n548 & ~n549 ) ;
  assign n551 = ( n504 & n507 ) | ( n504 & n550 ) | ( n507 & n550 ) ;
  assign n552 = ( ~n504 & n507 ) | ( ~n504 & n550 ) | ( n507 & n550 ) ;
  assign n553 = ( n504 & ~n551 ) | ( n504 & n552 ) | ( ~n551 & n552 ) ;
  assign n554 = ( n517 & n529 ) | ( n517 & ~n542 ) | ( n529 & ~n542 ) ;
  assign n555 = ( n517 & n529 ) | ( n517 & n542 ) | ( n529 & n542 ) ;
  assign n556 = ( n542 & n554 ) | ( n542 & ~n555 ) | ( n554 & ~n555 ) ;
  assign n557 = x3 & x19 ;
  assign n558 = x5 & x17 ;
  assign n559 = x4 & x18 ;
  assign n560 = ( ~n557 & n558 ) | ( ~n557 & n559 ) | ( n558 & n559 ) ;
  assign n561 = ( n557 & n558 ) | ( n557 & n559 ) | ( n558 & n559 ) ;
  assign n562 = ( n557 & n560 ) | ( n557 & ~n561 ) | ( n560 & ~n561 ) ;
  assign n563 = x6 & x16 ;
  assign n564 = x9 & x13 ;
  assign n565 = x2 & x20 ;
  assign n566 = ( ~n563 & n564 ) | ( ~n563 & n565 ) | ( n564 & n565 ) ;
  assign n567 = ( n563 & n564 ) | ( n563 & n565 ) | ( n564 & n565 ) ;
  assign n568 = ( n563 & n566 ) | ( n563 & ~n567 ) | ( n566 & ~n567 ) ;
  assign n569 = x0 & x22 ;
  assign n570 = x8 & x14 ;
  assign n571 = x7 & x15 ;
  assign n572 = ( ~n569 & n570 ) | ( ~n569 & n571 ) | ( n570 & n571 ) ;
  assign n573 = ( n569 & n570 ) | ( n569 & n571 ) | ( n570 & n571 ) ;
  assign n574 = ( n569 & n572 ) | ( n569 & ~n573 ) | ( n572 & ~n573 ) ;
  assign n575 = ( ~n562 & n568 ) | ( ~n562 & n574 ) | ( n568 & n574 ) ;
  assign n576 = ( n562 & n568 ) | ( n562 & n574 ) | ( n568 & n574 ) ;
  assign n577 = ( n562 & n575 ) | ( n562 & ~n576 ) | ( n575 & ~n576 ) ;
  assign n578 = ( ~n545 & n556 ) | ( ~n545 & n577 ) | ( n556 & n577 ) ;
  assign n579 = ( n545 & n556 ) | ( n545 & n577 ) | ( n556 & n577 ) ;
  assign n580 = ( n545 & n578 ) | ( n545 & ~n579 ) | ( n578 & ~n579 ) ;
  assign n581 = x10 & x12 ;
  assign n582 = x1 & x21 ;
  assign n583 = n581 & n582 ;
  assign n584 = n581 | n582 ;
  assign n585 = ~n583 & n584 ;
  assign n586 = ( ~n523 & n539 ) | ( ~n523 & n585 ) | ( n539 & n585 ) ;
  assign n587 = ( n523 & n539 ) | ( n523 & n585 ) | ( n539 & n585 ) ;
  assign n588 = ( n523 & n586 ) | ( n523 & ~n587 ) | ( n586 & ~n587 ) ;
  assign n589 = ( ~n511 & n532 ) | ( ~n511 & n588 ) | ( n532 & n588 ) ;
  assign n590 = ( n511 & n532 ) | ( n511 & n588 ) | ( n532 & n588 ) ;
  assign n591 = ( n511 & n589 ) | ( n511 & ~n590 ) | ( n589 & ~n590 ) ;
  assign n592 = ( n535 & n580 ) | ( n535 & n591 ) | ( n580 & n591 ) ;
  assign n593 = ( ~n535 & n580 ) | ( ~n535 & n591 ) | ( n580 & n591 ) ;
  assign n594 = ( n535 & ~n592 ) | ( n535 & n593 ) | ( ~n592 & n593 ) ;
  assign n595 = ( n549 & n551 ) | ( n549 & n594 ) | ( n551 & n594 ) ;
  assign n596 = ( ~n549 & n551 ) | ( ~n549 & n594 ) | ( n551 & n594 ) ;
  assign n597 = ( n549 & ~n595 ) | ( n549 & n596 ) | ( ~n595 & n596 ) ;
  assign n598 = x4 & x19 ;
  assign n599 = x11 & x12 ;
  assign n600 = x10 & x13 ;
  assign n601 = ( ~n598 & n599 ) | ( ~n598 & n600 ) | ( n599 & n600 ) ;
  assign n602 = ( n598 & n599 ) | ( n598 & n600 ) | ( n599 & n600 ) ;
  assign n603 = ( n598 & n601 ) | ( n598 & ~n602 ) | ( n601 & ~n602 ) ;
  assign n604 = x6 & x17 ;
  assign n605 = x5 & x18 ;
  assign n606 = x3 & x20 ;
  assign n607 = ( ~n604 & n605 ) | ( ~n604 & n606 ) | ( n605 & n606 ) ;
  assign n608 = ( n604 & n605 ) | ( n604 & n606 ) | ( n605 & n606 ) ;
  assign n609 = ( n604 & n607 ) | ( n604 & ~n608 ) | ( n607 & ~n608 ) ;
  assign n610 = ( n587 & n603 ) | ( n587 & n609 ) | ( n603 & n609 ) ;
  assign n611 = ( ~n587 & n603 ) | ( ~n587 & n609 ) | ( n603 & n609 ) ;
  assign n612 = ( n587 & ~n610 ) | ( n587 & n611 ) | ( ~n610 & n611 ) ;
  assign n613 = x7 & x16 ;
  assign n614 = x8 & x15 ;
  assign n615 = x9 & x14 ;
  assign n616 = ( ~n613 & n614 ) | ( ~n613 & n615 ) | ( n614 & n615 ) ;
  assign n617 = ( n613 & n614 ) | ( n613 & n615 ) | ( n614 & n615 ) ;
  assign n618 = ( n613 & n616 ) | ( n613 & ~n617 ) | ( n616 & ~n617 ) ;
  assign n619 = x2 & x23 ;
  assign n620 = n537 & n619 ;
  assign n621 = x0 & x23 ;
  assign n622 = x2 & x21 ;
  assign n623 = n621 | n622 ;
  assign n624 = ( n583 & n620 ) | ( n583 & n623 ) | ( n620 & n623 ) ;
  assign n625 = ( ~n583 & n620 ) | ( ~n583 & n623 ) | ( n620 & n623 ) ;
  assign n626 = ( n583 & ~n624 ) | ( n583 & n625 ) | ( ~n624 & n625 ) ;
  assign n627 = ( ~n573 & n618 ) | ( ~n573 & n626 ) | ( n618 & n626 ) ;
  assign n628 = ( n573 & n618 ) | ( n573 & n626 ) | ( n618 & n626 ) ;
  assign n629 = ( n573 & n627 ) | ( n573 & ~n628 ) | ( n627 & ~n628 ) ;
  assign n630 = ( ~n590 & n612 ) | ( ~n590 & n629 ) | ( n612 & n629 ) ;
  assign n631 = ( n590 & n612 ) | ( n590 & n629 ) | ( n612 & n629 ) ;
  assign n632 = ( n590 & n630 ) | ( n590 & ~n631 ) | ( n630 & ~n631 ) ;
  assign n633 = x1 & x22 ;
  assign n634 = x12 & n633 ;
  assign n635 = x12 | n633 ;
  assign n636 = ~n634 & n635 ;
  assign n637 = ( ~n561 & n567 ) | ( ~n561 & n636 ) | ( n567 & n636 ) ;
  assign n638 = ( n561 & n567 ) | ( n561 & n636 ) | ( n567 & n636 ) ;
  assign n639 = ( n561 & n637 ) | ( n561 & ~n638 ) | ( n637 & ~n638 ) ;
  assign n640 = ( ~n555 & n576 ) | ( ~n555 & n639 ) | ( n576 & n639 ) ;
  assign n641 = ( n555 & n576 ) | ( n555 & n639 ) | ( n576 & n639 ) ;
  assign n642 = ( n555 & n640 ) | ( n555 & ~n641 ) | ( n640 & ~n641 ) ;
  assign n643 = ( ~n579 & n632 ) | ( ~n579 & n642 ) | ( n632 & n642 ) ;
  assign n644 = ( n579 & n632 ) | ( n579 & n642 ) | ( n632 & n642 ) ;
  assign n645 = ( n579 & n643 ) | ( n579 & ~n644 ) | ( n643 & ~n644 ) ;
  assign n646 = ( n592 & n595 ) | ( n592 & n645 ) | ( n595 & n645 ) ;
  assign n647 = ( ~n592 & n595 ) | ( ~n592 & n645 ) | ( n595 & n645 ) ;
  assign n648 = ( n592 & ~n646 ) | ( n592 & n647 ) | ( ~n646 & n647 ) ;
  assign n649 = x0 & x24 ;
  assign n650 = x11 & x13 ;
  assign n651 = x1 & x23 ;
  assign n652 = n650 & n651 ;
  assign n653 = n650 | n651 ;
  assign n654 = ~n652 & n653 ;
  assign n655 = ( n634 & n649 ) | ( n634 & n654 ) | ( n649 & n654 ) ;
  assign n656 = ( ~n634 & n649 ) | ( ~n634 & n654 ) | ( n649 & n654 ) ;
  assign n657 = ( n634 & ~n655 ) | ( n634 & n656 ) | ( ~n655 & n656 ) ;
  assign n658 = x7 & x17 ;
  assign n659 = x2 & x22 ;
  assign n660 = x6 & x18 ;
  assign n661 = ( ~n658 & n659 ) | ( ~n658 & n660 ) | ( n659 & n660 ) ;
  assign n662 = ( n658 & n659 ) | ( n658 & n660 ) | ( n659 & n660 ) ;
  assign n663 = ( n658 & n661 ) | ( n658 & ~n662 ) | ( n661 & ~n662 ) ;
  assign n664 = ( ~n638 & n657 ) | ( ~n638 & n663 ) | ( n657 & n663 ) ;
  assign n665 = ( n638 & n657 ) | ( n638 & n663 ) | ( n657 & n663 ) ;
  assign n666 = ( n638 & n664 ) | ( n638 & ~n665 ) | ( n664 & ~n665 ) ;
  assign n667 = x8 & x16 ;
  assign n668 = x9 & x15 ;
  assign n669 = x10 & x14 ;
  assign n670 = ( ~n667 & n668 ) | ( ~n667 & n669 ) | ( n668 & n669 ) ;
  assign n671 = ( n667 & n668 ) | ( n667 & n669 ) | ( n668 & n669 ) ;
  assign n672 = ( n667 & n670 ) | ( n667 & ~n671 ) | ( n670 & ~n671 ) ;
  assign n673 = x3 & x21 ;
  assign n674 = x4 & x20 ;
  assign n675 = x5 & x19 ;
  assign n676 = ( ~n673 & n674 ) | ( ~n673 & n675 ) | ( n674 & n675 ) ;
  assign n677 = ( n673 & n674 ) | ( n673 & n675 ) | ( n674 & n675 ) ;
  assign n678 = ( n673 & n676 ) | ( n673 & ~n677 ) | ( n676 & ~n677 ) ;
  assign n679 = ( ~n624 & n672 ) | ( ~n624 & n678 ) | ( n672 & n678 ) ;
  assign n680 = ( n624 & n672 ) | ( n624 & n678 ) | ( n672 & n678 ) ;
  assign n681 = ( n624 & n679 ) | ( n624 & ~n680 ) | ( n679 & ~n680 ) ;
  assign n682 = ( n641 & n666 ) | ( n641 & n681 ) | ( n666 & n681 ) ;
  assign n683 = ( ~n641 & n666 ) | ( ~n641 & n681 ) | ( n666 & n681 ) ;
  assign n684 = ( n641 & ~n682 ) | ( n641 & n683 ) | ( ~n682 & n683 ) ;
  assign n685 = ( n602 & ~n608 ) | ( n602 & n617 ) | ( ~n608 & n617 ) ;
  assign n686 = ( n602 & n608 ) | ( n602 & n617 ) | ( n608 & n617 ) ;
  assign n687 = ( n608 & n685 ) | ( n608 & ~n686 ) | ( n685 & ~n686 ) ;
  assign n688 = ( ~n610 & n628 ) | ( ~n610 & n687 ) | ( n628 & n687 ) ;
  assign n689 = ( n610 & n628 ) | ( n610 & n687 ) | ( n628 & n687 ) ;
  assign n690 = ( n610 & n688 ) | ( n610 & ~n689 ) | ( n688 & ~n689 ) ;
  assign n691 = ( n631 & n684 ) | ( n631 & n690 ) | ( n684 & n690 ) ;
  assign n692 = ( ~n631 & n684 ) | ( ~n631 & n690 ) | ( n684 & n690 ) ;
  assign n693 = ( n631 & ~n691 ) | ( n631 & n692 ) | ( ~n691 & n692 ) ;
  assign n694 = ( ~n644 & n646 ) | ( ~n644 & n693 ) | ( n646 & n693 ) ;
  assign n695 = ( n644 & n646 ) | ( n644 & n693 ) | ( n646 & n693 ) ;
  assign n696 = ( n644 & n694 ) | ( n644 & ~n695 ) | ( n694 & ~n695 ) ;
  assign n697 = x7 & x18 ;
  assign n698 = x8 & x17 ;
  assign n699 = ( ~n356 & n697 ) | ( ~n356 & n698 ) | ( n697 & n698 ) ;
  assign n700 = ( n356 & n697 ) | ( n356 & n698 ) | ( n697 & n698 ) ;
  assign n701 = ( n356 & n699 ) | ( n356 & ~n700 ) | ( n699 & ~n700 ) ;
  assign n702 = x10 & x15 ;
  assign n703 = x0 & x25 ;
  assign n704 = ( ~n619 & n702 ) | ( ~n619 & n703 ) | ( n702 & n703 ) ;
  assign n705 = ( n619 & n702 ) | ( n619 & n703 ) | ( n702 & n703 ) ;
  assign n706 = ( n619 & n704 ) | ( n619 & ~n705 ) | ( n704 & ~n705 ) ;
  assign n707 = x6 & x19 ;
  assign n708 = x3 & x22 ;
  assign n709 = x4 & x21 ;
  assign n710 = ( ~n707 & n708 ) | ( ~n707 & n709 ) | ( n708 & n709 ) ;
  assign n711 = ( n707 & n708 ) | ( n707 & n709 ) | ( n708 & n709 ) ;
  assign n712 = ( n707 & n710 ) | ( n707 & ~n711 ) | ( n710 & ~n711 ) ;
  assign n713 = ( n701 & n706 ) | ( n701 & n712 ) | ( n706 & n712 ) ;
  assign n714 = ( ~n701 & n706 ) | ( ~n701 & n712 ) | ( n706 & n712 ) ;
  assign n715 = ( n701 & ~n713 ) | ( n701 & n714 ) | ( ~n713 & n714 ) ;
  assign n716 = x1 & x24 ;
  assign n717 = x13 & ~n652 ;
  assign n718 = ( ~n677 & n716 ) | ( ~n677 & n717 ) | ( n716 & n717 ) ;
  assign n719 = ( n677 & n716 ) | ( n677 & n717 ) | ( n716 & n717 ) ;
  assign n720 = ( n677 & n718 ) | ( n677 & ~n719 ) | ( n718 & ~n719 ) ;
  assign n721 = x5 & x20 ;
  assign n722 = x12 & x13 ;
  assign n723 = x11 & x14 ;
  assign n724 = ( ~n721 & n722 ) | ( ~n721 & n723 ) | ( n722 & n723 ) ;
  assign n725 = ( n721 & n722 ) | ( n721 & n723 ) | ( n722 & n723 ) ;
  assign n726 = ( n721 & n724 ) | ( n721 & ~n725 ) | ( n724 & ~n725 ) ;
  assign n727 = ( ~n686 & n720 ) | ( ~n686 & n726 ) | ( n720 & n726 ) ;
  assign n728 = ( n686 & n720 ) | ( n686 & n726 ) | ( n720 & n726 ) ;
  assign n729 = ( n686 & n727 ) | ( n686 & ~n728 ) | ( n727 & ~n728 ) ;
  assign n730 = ( ~n689 & n715 ) | ( ~n689 & n729 ) | ( n715 & n729 ) ;
  assign n731 = ( n689 & n715 ) | ( n689 & n729 ) | ( n715 & n729 ) ;
  assign n732 = ( n689 & n730 ) | ( n689 & ~n731 ) | ( n730 & ~n731 ) ;
  assign n733 = ( ~n655 & n662 ) | ( ~n655 & n671 ) | ( n662 & n671 ) ;
  assign n734 = ( n655 & n662 ) | ( n655 & n671 ) | ( n662 & n671 ) ;
  assign n735 = ( n655 & n733 ) | ( n655 & ~n734 ) | ( n733 & ~n734 ) ;
  assign n736 = ( n665 & n680 ) | ( n665 & n735 ) | ( n680 & n735 ) ;
  assign n737 = ( n665 & ~n680 ) | ( n665 & n735 ) | ( ~n680 & n735 ) ;
  assign n738 = ( n680 & ~n736 ) | ( n680 & n737 ) | ( ~n736 & n737 ) ;
  assign n739 = ( n682 & n732 ) | ( n682 & n738 ) | ( n732 & n738 ) ;
  assign n740 = ( n682 & ~n732 ) | ( n682 & n738 ) | ( ~n732 & n738 ) ;
  assign n741 = ( n732 & ~n739 ) | ( n732 & n740 ) | ( ~n739 & n740 ) ;
  assign n742 = ( ~n691 & n695 ) | ( ~n691 & n741 ) | ( n695 & n741 ) ;
  assign n743 = ( n691 & n695 ) | ( n691 & n741 ) | ( n695 & n741 ) ;
  assign n744 = ( n691 & n742 ) | ( n691 & ~n743 ) | ( n742 & ~n743 ) ;
  assign n745 = ( n652 & ~n718 ) | ( n652 & n719 ) | ( ~n718 & n719 ) ;
  assign n746 = x13 & n716 ;
  assign n747 = x0 & x26 ;
  assign n748 = x8 & x18 ;
  assign n749 = ( ~n746 & n747 ) | ( ~n746 & n748 ) | ( n747 & n748 ) ;
  assign n750 = ( n746 & n747 ) | ( n746 & n748 ) | ( n747 & n748 ) ;
  assign n751 = ( n746 & n749 ) | ( n746 & ~n750 ) | ( n749 & ~n750 ) ;
  assign n752 = ( ~n700 & n705 ) | ( ~n700 & n751 ) | ( n705 & n751 ) ;
  assign n753 = ( n700 & n705 ) | ( n700 & n751 ) | ( n705 & n751 ) ;
  assign n754 = ( n700 & n752 ) | ( n700 & ~n753 ) | ( n752 & ~n753 ) ;
  assign n755 = ( ~n734 & n745 ) | ( ~n734 & n754 ) | ( n745 & n754 ) ;
  assign n756 = ( n734 & n745 ) | ( n734 & n754 ) | ( n745 & n754 ) ;
  assign n757 = ( n734 & n755 ) | ( n734 & ~n756 ) | ( n755 & ~n756 ) ;
  assign n758 = x2 & x24 ;
  assign n759 = x3 & x23 ;
  assign n760 = x7 & x19 ;
  assign n761 = ( ~n758 & n759 ) | ( ~n758 & n760 ) | ( n759 & n760 ) ;
  assign n762 = ( n758 & n759 ) | ( n758 & n760 ) | ( n759 & n760 ) ;
  assign n763 = ( n758 & n761 ) | ( n758 & ~n762 ) | ( n761 & ~n762 ) ;
  assign n764 = x4 & x22 ;
  assign n765 = x6 & x20 ;
  assign n766 = x5 & x21 ;
  assign n767 = ( ~n764 & n765 ) | ( ~n764 & n766 ) | ( n765 & n766 ) ;
  assign n768 = ( n764 & n765 ) | ( n764 & n766 ) | ( n765 & n766 ) ;
  assign n769 = ( n764 & n767 ) | ( n764 & ~n768 ) | ( n767 & ~n768 ) ;
  assign n770 = x9 & x17 ;
  assign n771 = x11 & x15 ;
  assign n772 = x10 & x16 ;
  assign n773 = ( ~n770 & n771 ) | ( ~n770 & n772 ) | ( n771 & n772 ) ;
  assign n774 = ( n770 & n771 ) | ( n770 & n772 ) | ( n771 & n772 ) ;
  assign n775 = ( n770 & n773 ) | ( n770 & ~n774 ) | ( n773 & ~n774 ) ;
  assign n776 = ( ~n763 & n769 ) | ( ~n763 & n775 ) | ( n769 & n775 ) ;
  assign n777 = ( n763 & n769 ) | ( n763 & n775 ) | ( n769 & n775 ) ;
  assign n778 = ( n763 & n776 ) | ( n763 & ~n777 ) | ( n776 & ~n777 ) ;
  assign n779 = ( ~n736 & n757 ) | ( ~n736 & n778 ) | ( n757 & n778 ) ;
  assign n780 = ( n736 & n757 ) | ( n736 & n778 ) | ( n757 & n778 ) ;
  assign n781 = ( n736 & n779 ) | ( n736 & ~n780 ) | ( n779 & ~n780 ) ;
  assign n782 = x12 & x14 ;
  assign n783 = x1 & x25 ;
  assign n784 = n782 & n783 ;
  assign n785 = n782 | n783 ;
  assign n786 = ~n784 & n785 ;
  assign n787 = ( n711 & n725 ) | ( n711 & n786 ) | ( n725 & n786 ) ;
  assign n788 = ( ~n711 & n725 ) | ( ~n711 & n786 ) | ( n725 & n786 ) ;
  assign n789 = ( n711 & ~n787 ) | ( n711 & n788 ) | ( ~n787 & n788 ) ;
  assign n790 = ( ~n713 & n728 ) | ( ~n713 & n789 ) | ( n728 & n789 ) ;
  assign n791 = ( n713 & n728 ) | ( n713 & n789 ) | ( n728 & n789 ) ;
  assign n792 = ( n713 & n790 ) | ( n713 & ~n791 ) | ( n790 & ~n791 ) ;
  assign n793 = ( n731 & n781 ) | ( n731 & n792 ) | ( n781 & n792 ) ;
  assign n794 = ( ~n731 & n781 ) | ( ~n731 & n792 ) | ( n781 & n792 ) ;
  assign n795 = ( n731 & ~n793 ) | ( n731 & n794 ) | ( ~n793 & n794 ) ;
  assign n796 = ( n739 & n743 ) | ( n739 & n795 ) | ( n743 & n795 ) ;
  assign n797 = ( ~n739 & n743 ) | ( ~n739 & n795 ) | ( n743 & n795 ) ;
  assign n798 = ( n739 & ~n796 ) | ( n739 & n797 ) | ( ~n796 & n797 ) ;
  assign n799 = x11 & x16 ;
  assign n800 = x2 & x25 ;
  assign n801 = x7 & x20 ;
  assign n802 = ( ~n799 & n800 ) | ( ~n799 & n801 ) | ( n800 & n801 ) ;
  assign n803 = ( n799 & n800 ) | ( n799 & n801 ) | ( n800 & n801 ) ;
  assign n804 = ( n799 & n802 ) | ( n799 & ~n803 ) | ( n802 & ~n803 ) ;
  assign n805 = x8 & x19 ;
  assign n806 = x10 & x17 ;
  assign n807 = x9 & x18 ;
  assign n808 = ( ~n805 & n806 ) | ( ~n805 & n807 ) | ( n806 & n807 ) ;
  assign n809 = ( n805 & n806 ) | ( n805 & n807 ) | ( n806 & n807 ) ;
  assign n810 = ( n805 & n808 ) | ( n805 & ~n809 ) | ( n808 & ~n809 ) ;
  assign n811 = ( n750 & n804 ) | ( n750 & n810 ) | ( n804 & n810 ) ;
  assign n812 = ( ~n750 & n804 ) | ( ~n750 & n810 ) | ( n804 & n810 ) ;
  assign n813 = ( n750 & ~n811 ) | ( n750 & n812 ) | ( ~n811 & n812 ) ;
  assign n814 = ( n753 & n777 ) | ( n753 & ~n787 ) | ( n777 & ~n787 ) ;
  assign n815 = ( n753 & n777 ) | ( n753 & n787 ) | ( n777 & n787 ) ;
  assign n816 = ( n787 & n814 ) | ( n787 & ~n815 ) | ( n814 & ~n815 ) ;
  assign n817 = ( ~n791 & n813 ) | ( ~n791 & n816 ) | ( n813 & n816 ) ;
  assign n818 = ( n791 & n813 ) | ( n791 & n816 ) | ( n813 & n816 ) ;
  assign n819 = ( n791 & n817 ) | ( n791 & ~n818 ) | ( n817 & ~n818 ) ;
  assign n820 = ( ~n762 & n768 ) | ( ~n762 & n774 ) | ( n768 & n774 ) ;
  assign n821 = ( n762 & n768 ) | ( n762 & n774 ) | ( n768 & n774 ) ;
  assign n822 = ( n762 & n820 ) | ( n762 & ~n821 ) | ( n820 & ~n821 ) ;
  assign n823 = ~x1 & x14 ;
  assign n824 = ( x1 & x14 ) | ( x1 & x26 ) | ( x14 & x26 ) ;
  assign n825 = x14 & x26 ;
  assign n826 = ( n823 & n824 ) | ( n823 & ~n825 ) | ( n824 & ~n825 ) ;
  assign n827 = x0 & x27 ;
  assign n828 = ( n784 & n826 ) | ( n784 & n827 ) | ( n826 & n827 ) ;
  assign n829 = ( ~n784 & n826 ) | ( ~n784 & n827 ) | ( n826 & n827 ) ;
  assign n830 = ( n784 & ~n828 ) | ( n784 & n829 ) | ( ~n828 & n829 ) ;
  assign n831 = x6 & x21 ;
  assign n832 = x3 & x24 ;
  assign n833 = x4 & x23 ;
  assign n834 = ( ~n831 & n832 ) | ( ~n831 & n833 ) | ( n832 & n833 ) ;
  assign n835 = ( n831 & n832 ) | ( n831 & n833 ) | ( n832 & n833 ) ;
  assign n836 = ( n831 & n834 ) | ( n831 & ~n835 ) | ( n834 & ~n835 ) ;
  assign n837 = x5 & x22 ;
  assign n838 = x13 & x14 ;
  assign n839 = x12 & x15 ;
  assign n840 = ( ~n837 & n838 ) | ( ~n837 & n839 ) | ( n838 & n839 ) ;
  assign n841 = ( n837 & n838 ) | ( n837 & n839 ) | ( n838 & n839 ) ;
  assign n842 = ( n837 & n840 ) | ( n837 & ~n841 ) | ( n840 & ~n841 ) ;
  assign n843 = ( ~n830 & n836 ) | ( ~n830 & n842 ) | ( n836 & n842 ) ;
  assign n844 = ( n830 & n836 ) | ( n830 & n842 ) | ( n836 & n842 ) ;
  assign n845 = ( n830 & n843 ) | ( n830 & ~n844 ) | ( n843 & ~n844 ) ;
  assign n846 = ( ~n756 & n822 ) | ( ~n756 & n845 ) | ( n822 & n845 ) ;
  assign n847 = ( n756 & n822 ) | ( n756 & n845 ) | ( n822 & n845 ) ;
  assign n848 = ( n756 & n846 ) | ( n756 & ~n847 ) | ( n846 & ~n847 ) ;
  assign n849 = ( ~n780 & n819 ) | ( ~n780 & n848 ) | ( n819 & n848 ) ;
  assign n850 = ( n780 & n819 ) | ( n780 & n848 ) | ( n819 & n848 ) ;
  assign n851 = ( n780 & n849 ) | ( n780 & ~n850 ) | ( n849 & ~n850 ) ;
  assign n852 = ( ~n793 & n796 ) | ( ~n793 & n851 ) | ( n796 & n851 ) ;
  assign n853 = ( n793 & n796 ) | ( n793 & n851 ) | ( n796 & n851 ) ;
  assign n854 = ( n793 & n852 ) | ( n793 & ~n853 ) | ( n852 & ~n853 ) ;
  assign n855 = x7 & x21 ;
  assign n856 = x6 & x22 ;
  assign n857 = x5 & x23 ;
  assign n858 = ( ~n855 & n856 ) | ( ~n855 & n857 ) | ( n856 & n857 ) ;
  assign n859 = ( n855 & n856 ) | ( n855 & n857 ) | ( n856 & n857 ) ;
  assign n860 = ( n855 & n858 ) | ( n855 & ~n859 ) | ( n858 & ~n859 ) ;
  assign n861 = x8 & x20 ;
  assign n862 = x3 & x25 ;
  assign n863 = x4 & x24 ;
  assign n864 = ( ~n861 & n862 ) | ( ~n861 & n863 ) | ( n862 & n863 ) ;
  assign n865 = ( n861 & n862 ) | ( n861 & n863 ) | ( n862 & n863 ) ;
  assign n866 = ( n861 & n864 ) | ( n861 & ~n865 ) | ( n864 & ~n865 ) ;
  assign n867 = ( n828 & n860 ) | ( n828 & n866 ) | ( n860 & n866 ) ;
  assign n868 = ( ~n828 & n860 ) | ( ~n828 & n866 ) | ( n860 & n866 ) ;
  assign n869 = ( n828 & ~n867 ) | ( n828 & n868 ) | ( ~n867 & n868 ) ;
  assign n870 = x26 & n296 ;
  assign n871 = x13 & x15 ;
  assign n872 = x1 & x27 ;
  assign n873 = n871 & n872 ;
  assign n874 = n871 | n872 ;
  assign n875 = ~n873 & n874 ;
  assign n876 = ( n841 & n870 ) | ( n841 & n875 ) | ( n870 & n875 ) ;
  assign n877 = ( n841 & ~n870 ) | ( n841 & n875 ) | ( ~n870 & n875 ) ;
  assign n878 = ( n870 & ~n876 ) | ( n870 & n877 ) | ( ~n876 & n877 ) ;
  assign n879 = ( ~n811 & n844 ) | ( ~n811 & n878 ) | ( n844 & n878 ) ;
  assign n880 = ( n811 & n844 ) | ( n811 & n878 ) | ( n844 & n878 ) ;
  assign n881 = ( n811 & n879 ) | ( n811 & ~n880 ) | ( n879 & ~n880 ) ;
  assign n882 = ( ~n847 & n869 ) | ( ~n847 & n881 ) | ( n869 & n881 ) ;
  assign n883 = ( n847 & n869 ) | ( n847 & n881 ) | ( n869 & n881 ) ;
  assign n884 = ( n847 & n882 ) | ( n847 & ~n883 ) | ( n882 & ~n883 ) ;
  assign n885 = ( ~n803 & n809 ) | ( ~n803 & n835 ) | ( n809 & n835 ) ;
  assign n886 = ( n803 & n809 ) | ( n803 & n835 ) | ( n809 & n835 ) ;
  assign n887 = ( n803 & n885 ) | ( n803 & ~n886 ) | ( n885 & ~n886 ) ;
  assign n888 = x11 & x17 ;
  assign n889 = x0 & x28 ;
  assign n890 = x12 & x16 ;
  assign n891 = ( ~n888 & n889 ) | ( ~n888 & n890 ) | ( n889 & n890 ) ;
  assign n892 = ( n888 & n889 ) | ( n888 & n890 ) | ( n889 & n890 ) ;
  assign n893 = ( n888 & n891 ) | ( n888 & ~n892 ) | ( n891 & ~n892 ) ;
  assign n894 = x2 & x26 ;
  assign n895 = x10 & x18 ;
  assign n896 = x9 & x19 ;
  assign n897 = ( ~n894 & n895 ) | ( ~n894 & n896 ) | ( n895 & n896 ) ;
  assign n898 = ( n894 & n895 ) | ( n894 & n896 ) | ( n895 & n896 ) ;
  assign n899 = ( n894 & n897 ) | ( n894 & ~n898 ) | ( n897 & ~n898 ) ;
  assign n900 = ( n821 & n893 ) | ( n821 & n899 ) | ( n893 & n899 ) ;
  assign n901 = ( ~n821 & n893 ) | ( ~n821 & n899 ) | ( n893 & n899 ) ;
  assign n902 = ( n821 & ~n900 ) | ( n821 & n901 ) | ( ~n900 & n901 ) ;
  assign n903 = ( n815 & n887 ) | ( n815 & n902 ) | ( n887 & n902 ) ;
  assign n904 = ( ~n815 & n887 ) | ( ~n815 & n902 ) | ( n887 & n902 ) ;
  assign n905 = ( n815 & ~n903 ) | ( n815 & n904 ) | ( ~n903 & n904 ) ;
  assign n906 = ( n818 & n850 ) | ( n818 & n905 ) | ( n850 & n905 ) ;
  assign n907 = ( ~n818 & n850 ) | ( ~n818 & n905 ) | ( n850 & n905 ) ;
  assign n908 = ( n818 & ~n906 ) | ( n818 & n907 ) | ( ~n906 & n907 ) ;
  assign n909 = ( ~n853 & n884 ) | ( ~n853 & n908 ) | ( n884 & n908 ) ;
  assign n910 = ( n853 & n884 ) | ( n853 & n908 ) | ( n884 & n908 ) ;
  assign n911 = ( n853 & n909 ) | ( n853 & ~n910 ) | ( n909 & ~n910 ) ;
  assign n912 = x6 & x23 ;
  assign n913 = x14 & x15 ;
  assign n914 = x13 & x16 ;
  assign n915 = ( ~n912 & n913 ) | ( ~n912 & n914 ) | ( n913 & n914 ) ;
  assign n916 = ( n912 & n913 ) | ( n912 & n914 ) | ( n913 & n914 ) ;
  assign n917 = ( n912 & n915 ) | ( n912 & ~n916 ) | ( n915 & ~n916 ) ;
  assign n918 = ( ~n876 & n886 ) | ( ~n876 & n917 ) | ( n886 & n917 ) ;
  assign n919 = ( n876 & n886 ) | ( n876 & n917 ) | ( n886 & n917 ) ;
  assign n920 = ( n876 & n918 ) | ( n876 & ~n919 ) | ( n918 & ~n919 ) ;
  assign n921 = ~x1 & x15 ;
  assign n922 = ( x1 & x15 ) | ( x1 & x28 ) | ( x15 & x28 ) ;
  assign n923 = x15 & x28 ;
  assign n924 = ( n921 & n922 ) | ( n921 & ~n923 ) | ( n922 & ~n923 ) ;
  assign n925 = ( ~n859 & n865 ) | ( ~n859 & n924 ) | ( n865 & n924 ) ;
  assign n926 = ( n859 & n865 ) | ( n859 & n924 ) | ( n865 & n924 ) ;
  assign n927 = ( n859 & n925 ) | ( n859 & ~n926 ) | ( n925 & ~n926 ) ;
  assign n928 = x4 & x25 ;
  assign n929 = x7 & x22 ;
  assign n930 = x5 & x24 ;
  assign n931 = ( ~n928 & n929 ) | ( ~n928 & n930 ) | ( n929 & n930 ) ;
  assign n932 = ( n928 & n929 ) | ( n928 & n930 ) | ( n929 & n930 ) ;
  assign n933 = ( n928 & n931 ) | ( n928 & ~n932 ) | ( n931 & ~n932 ) ;
  assign n934 = x9 & x20 ;
  assign n935 = x10 & x19 ;
  assign n936 = x11 & x18 ;
  assign n937 = ( ~n934 & n935 ) | ( ~n934 & n936 ) | ( n935 & n936 ) ;
  assign n938 = ( n934 & n935 ) | ( n934 & n936 ) | ( n935 & n936 ) ;
  assign n939 = ( n934 & n937 ) | ( n934 & ~n938 ) | ( n937 & ~n938 ) ;
  assign n940 = x12 & x17 ;
  assign n941 = x3 & x26 ;
  assign n942 = x8 & x21 ;
  assign n943 = ( ~n940 & n941 ) | ( ~n940 & n942 ) | ( n941 & n942 ) ;
  assign n944 = ( n940 & n941 ) | ( n940 & n942 ) | ( n941 & n942 ) ;
  assign n945 = ( n940 & n943 ) | ( n940 & ~n944 ) | ( n943 & ~n944 ) ;
  assign n946 = ( ~n933 & n939 ) | ( ~n933 & n945 ) | ( n939 & n945 ) ;
  assign n947 = ( n933 & n939 ) | ( n933 & n945 ) | ( n939 & n945 ) ;
  assign n948 = ( n933 & n946 ) | ( n933 & ~n947 ) | ( n946 & ~n947 ) ;
  assign n949 = ( ~n920 & n927 ) | ( ~n920 & n948 ) | ( n927 & n948 ) ;
  assign n950 = ( n920 & n927 ) | ( n920 & n948 ) | ( n927 & n948 ) ;
  assign n951 = ( n920 & n949 ) | ( n920 & ~n950 ) | ( n949 & ~n950 ) ;
  assign n952 = x0 & x29 ;
  assign n953 = x2 & x27 ;
  assign n954 = n952 | n953 ;
  assign n955 = x2 & x29 ;
  assign n956 = n827 & n955 ;
  assign n957 = ( n873 & n954 ) | ( n873 & n956 ) | ( n954 & n956 ) ;
  assign n958 = ( ~n873 & n954 ) | ( ~n873 & n956 ) | ( n954 & n956 ) ;
  assign n959 = ( n873 & ~n957 ) | ( n873 & n958 ) | ( ~n957 & n958 ) ;
  assign n960 = ( n892 & n898 ) | ( n892 & n959 ) | ( n898 & n959 ) ;
  assign n961 = ( ~n892 & n898 ) | ( ~n892 & n959 ) | ( n898 & n959 ) ;
  assign n962 = ( n892 & ~n960 ) | ( n892 & n961 ) | ( ~n960 & n961 ) ;
  assign n963 = ( n867 & n900 ) | ( n867 & n962 ) | ( n900 & n962 ) ;
  assign n964 = ( ~n867 & n900 ) | ( ~n867 & n962 ) | ( n900 & n962 ) ;
  assign n965 = ( n867 & ~n963 ) | ( n867 & n964 ) | ( ~n963 & n964 ) ;
  assign n966 = ( n880 & n903 ) | ( n880 & n965 ) | ( n903 & n965 ) ;
  assign n967 = ( ~n880 & n903 ) | ( ~n880 & n965 ) | ( n903 & n965 ) ;
  assign n968 = ( n880 & ~n966 ) | ( n880 & n967 ) | ( ~n966 & n967 ) ;
  assign n969 = ( ~n883 & n951 ) | ( ~n883 & n968 ) | ( n951 & n968 ) ;
  assign n970 = ( n883 & n951 ) | ( n883 & n968 ) | ( n951 & n968 ) ;
  assign n971 = ( n883 & n969 ) | ( n883 & ~n970 ) | ( n969 & ~n970 ) ;
  assign n972 = ( n906 & n910 ) | ( n906 & n971 ) | ( n910 & n971 ) ;
  assign n973 = ( ~n906 & n910 ) | ( ~n906 & n971 ) | ( n910 & n971 ) ;
  assign n974 = ( n906 & ~n972 ) | ( n906 & n973 ) | ( ~n972 & n973 ) ;
  assign n975 = x28 & n333 ;
  assign n976 = x14 & x16 ;
  assign n977 = x1 & x29 ;
  assign n978 = n976 & n977 ;
  assign n979 = n976 | n977 ;
  assign n980 = ~n978 & n979 ;
  assign n981 = x0 & x30 ;
  assign n982 = ( n975 & n980 ) | ( n975 & n981 ) | ( n980 & n981 ) ;
  assign n983 = ( ~n975 & n980 ) | ( ~n975 & n981 ) | ( n980 & n981 ) ;
  assign n984 = ( n975 & ~n982 ) | ( n975 & n983 ) | ( ~n982 & n983 ) ;
  assign n985 = ( n926 & n960 ) | ( n926 & n984 ) | ( n960 & n984 ) ;
  assign n986 = ( ~n926 & n960 ) | ( ~n926 & n984 ) | ( n960 & n984 ) ;
  assign n987 = ( n926 & ~n985 ) | ( n926 & n986 ) | ( ~n985 & n986 ) ;
  assign n988 = ( ~n938 & n944 ) | ( ~n938 & n957 ) | ( n944 & n957 ) ;
  assign n989 = ( n938 & n944 ) | ( n938 & n957 ) | ( n944 & n957 ) ;
  assign n990 = ( n938 & n988 ) | ( n938 & ~n989 ) | ( n988 & ~n989 ) ;
  assign n991 = x13 & x17 ;
  assign n992 = x2 & x28 ;
  assign n993 = x9 & x21 ;
  assign n994 = ( ~n991 & n992 ) | ( ~n991 & n993 ) | ( n992 & n993 ) ;
  assign n995 = ( n991 & n992 ) | ( n991 & n993 ) | ( n992 & n993 ) ;
  assign n996 = ( n991 & n994 ) | ( n991 & ~n995 ) | ( n994 & ~n995 ) ;
  assign n997 = ( ~n916 & n932 ) | ( ~n916 & n996 ) | ( n932 & n996 ) ;
  assign n998 = ( n916 & n932 ) | ( n916 & n996 ) | ( n932 & n996 ) ;
  assign n999 = ( n916 & n997 ) | ( n916 & ~n998 ) | ( n997 & ~n998 ) ;
  assign n1000 = ( ~n947 & n990 ) | ( ~n947 & n999 ) | ( n990 & n999 ) ;
  assign n1001 = ( n947 & n990 ) | ( n947 & n999 ) | ( n990 & n999 ) ;
  assign n1002 = ( n947 & n1000 ) | ( n947 & ~n1001 ) | ( n1000 & ~n1001 ) ;
  assign n1003 = ( ~n950 & n987 ) | ( ~n950 & n1002 ) | ( n987 & n1002 ) ;
  assign n1004 = ( n950 & n987 ) | ( n950 & n1002 ) | ( n987 & n1002 ) ;
  assign n1005 = ( n950 & n1003 ) | ( n950 & ~n1004 ) | ( n1003 & ~n1004 ) ;
  assign n1006 = x10 & x20 ;
  assign n1007 = x11 & x19 ;
  assign n1008 = x12 & x18 ;
  assign n1009 = ( ~n1006 & n1007 ) | ( ~n1006 & n1008 ) | ( n1007 & n1008 ) ;
  assign n1010 = ( n1006 & n1007 ) | ( n1006 & n1008 ) | ( n1007 & n1008 ) ;
  assign n1011 = ( n1006 & n1009 ) | ( n1006 & ~n1010 ) | ( n1009 & ~n1010 ) ;
  assign n1012 = x3 & x27 ;
  assign n1013 = x4 & x26 ;
  assign n1014 = x8 & x22 ;
  assign n1015 = ( ~n1012 & n1013 ) | ( ~n1012 & n1014 ) | ( n1013 & n1014 ) ;
  assign n1016 = ( n1012 & n1013 ) | ( n1012 & n1014 ) | ( n1013 & n1014 ) ;
  assign n1017 = ( n1012 & n1015 ) | ( n1012 & ~n1016 ) | ( n1015 & ~n1016 ) ;
  assign n1018 = x5 & x25 ;
  assign n1019 = x7 & x23 ;
  assign n1020 = x6 & x24 ;
  assign n1021 = ( ~n1018 & n1019 ) | ( ~n1018 & n1020 ) | ( n1019 & n1020 ) ;
  assign n1022 = ( n1018 & n1019 ) | ( n1018 & n1020 ) | ( n1019 & n1020 ) ;
  assign n1023 = ( n1018 & n1021 ) | ( n1018 & ~n1022 ) | ( n1021 & ~n1022 ) ;
  assign n1024 = ( ~n1011 & n1017 ) | ( ~n1011 & n1023 ) | ( n1017 & n1023 ) ;
  assign n1025 = ( n1011 & n1017 ) | ( n1011 & n1023 ) | ( n1017 & n1023 ) ;
  assign n1026 = ( n1011 & n1024 ) | ( n1011 & ~n1025 ) | ( n1024 & ~n1025 ) ;
  assign n1027 = ( n919 & n963 ) | ( n919 & n1026 ) | ( n963 & n1026 ) ;
  assign n1028 = ( ~n919 & n963 ) | ( ~n919 & n1026 ) | ( n963 & n1026 ) ;
  assign n1029 = ( n919 & ~n1027 ) | ( n919 & n1028 ) | ( ~n1027 & n1028 ) ;
  assign n1030 = ( ~n966 & n1005 ) | ( ~n966 & n1029 ) | ( n1005 & n1029 ) ;
  assign n1031 = ( n966 & n1005 ) | ( n966 & n1029 ) | ( n1005 & n1029 ) ;
  assign n1032 = ( n966 & n1030 ) | ( n966 & ~n1031 ) | ( n1030 & ~n1031 ) ;
  assign n1033 = ( ~n970 & n972 ) | ( ~n970 & n1032 ) | ( n972 & n1032 ) ;
  assign n1034 = ( n970 & n972 ) | ( n970 & n1032 ) | ( n972 & n1032 ) ;
  assign n1035 = ( n970 & n1033 ) | ( n970 & ~n1034 ) | ( n1033 & ~n1034 ) ;
  assign n1036 = x1 & x30 ;
  assign n1037 = x16 & ~n978 ;
  assign n1038 = ( ~n1022 & n1036 ) | ( ~n1022 & n1037 ) | ( n1036 & n1037 ) ;
  assign n1039 = ( n1022 & n1036 ) | ( n1022 & n1037 ) | ( n1036 & n1037 ) ;
  assign n1040 = ( n1022 & n1038 ) | ( n1022 & ~n1039 ) | ( n1038 & ~n1039 ) ;
  assign n1041 = ( ~n989 & n998 ) | ( ~n989 & n1040 ) | ( n998 & n1040 ) ;
  assign n1042 = ( n989 & n998 ) | ( n989 & n1040 ) | ( n998 & n1040 ) ;
  assign n1043 = ( n989 & n1041 ) | ( n989 & ~n1042 ) | ( n1041 & ~n1042 ) ;
  assign n1044 = ( n995 & ~n1010 ) | ( n995 & n1016 ) | ( ~n1010 & n1016 ) ;
  assign n1045 = ( n995 & n1010 ) | ( n995 & n1016 ) | ( n1010 & n1016 ) ;
  assign n1046 = ( n1010 & n1044 ) | ( n1010 & ~n1045 ) | ( n1044 & ~n1045 ) ;
  assign n1047 = ( ~n985 & n1025 ) | ( ~n985 & n1046 ) | ( n1025 & n1046 ) ;
  assign n1048 = ( n985 & n1025 ) | ( n985 & n1046 ) | ( n1025 & n1046 ) ;
  assign n1049 = ( n985 & n1047 ) | ( n985 & ~n1048 ) | ( n1047 & ~n1048 ) ;
  assign n1050 = ( ~n1027 & n1043 ) | ( ~n1027 & n1049 ) | ( n1043 & n1049 ) ;
  assign n1051 = ( n1027 & n1043 ) | ( n1027 & n1049 ) | ( n1043 & n1049 ) ;
  assign n1052 = ( n1027 & n1050 ) | ( n1027 & ~n1051 ) | ( n1050 & ~n1051 ) ;
  assign n1053 = x11 & x20 ;
  assign n1054 = x12 & x19 ;
  assign n1055 = x13 & x18 ;
  assign n1056 = ( ~n1053 & n1054 ) | ( ~n1053 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1057 = ( n1053 & n1054 ) | ( n1053 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1058 = ( n1053 & n1056 ) | ( n1053 & ~n1057 ) | ( n1056 & ~n1057 ) ;
  assign n1059 = x10 & x21 ;
  assign n1060 = x0 & x31 ;
  assign n1061 = x9 & x22 ;
  assign n1062 = ( ~n1059 & n1060 ) | ( ~n1059 & n1061 ) | ( n1060 & n1061 ) ;
  assign n1063 = ( n1059 & n1060 ) | ( n1059 & n1061 ) | ( n1060 & n1061 ) ;
  assign n1064 = ( n1059 & n1062 ) | ( n1059 & ~n1063 ) | ( n1062 & ~n1063 ) ;
  assign n1065 = ( n982 & n1058 ) | ( n982 & n1064 ) | ( n1058 & n1064 ) ;
  assign n1066 = ( ~n982 & n1058 ) | ( ~n982 & n1064 ) | ( n1058 & n1064 ) ;
  assign n1067 = ( n982 & ~n1065 ) | ( n982 & n1066 ) | ( ~n1065 & n1066 ) ;
  assign n1068 = x3 & x28 ;
  assign n1069 = x4 & x27 ;
  assign n1070 = ( ~n955 & n1068 ) | ( ~n955 & n1069 ) | ( n1068 & n1069 ) ;
  assign n1071 = ( n955 & n1068 ) | ( n955 & n1069 ) | ( n1068 & n1069 ) ;
  assign n1072 = ( n955 & n1070 ) | ( n955 & ~n1071 ) | ( n1070 & ~n1071 ) ;
  assign n1073 = x6 & x25 ;
  assign n1074 = x15 & x16 ;
  assign n1075 = x14 & x17 ;
  assign n1076 = ( ~n1073 & n1074 ) | ( ~n1073 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1077 = ( n1073 & n1074 ) | ( n1073 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1078 = ( n1073 & n1076 ) | ( n1073 & ~n1077 ) | ( n1076 & ~n1077 ) ;
  assign n1079 = x8 & x23 ;
  assign n1080 = x7 & x24 ;
  assign n1081 = x5 & x26 ;
  assign n1082 = ( ~n1079 & n1080 ) | ( ~n1079 & n1081 ) | ( n1080 & n1081 ) ;
  assign n1083 = ( n1079 & n1080 ) | ( n1079 & n1081 ) | ( n1080 & n1081 ) ;
  assign n1084 = ( n1079 & n1082 ) | ( n1079 & ~n1083 ) | ( n1082 & ~n1083 ) ;
  assign n1085 = ( ~n1072 & n1078 ) | ( ~n1072 & n1084 ) | ( n1078 & n1084 ) ;
  assign n1086 = ( n1072 & n1078 ) | ( n1072 & n1084 ) | ( n1078 & n1084 ) ;
  assign n1087 = ( n1072 & n1085 ) | ( n1072 & ~n1086 ) | ( n1085 & ~n1086 ) ;
  assign n1088 = ( ~n1001 & n1067 ) | ( ~n1001 & n1087 ) | ( n1067 & n1087 ) ;
  assign n1089 = ( n1001 & n1067 ) | ( n1001 & n1087 ) | ( n1067 & n1087 ) ;
  assign n1090 = ( n1001 & n1088 ) | ( n1001 & ~n1089 ) | ( n1088 & ~n1089 ) ;
  assign n1091 = ( ~n1004 & n1052 ) | ( ~n1004 & n1090 ) | ( n1052 & n1090 ) ;
  assign n1092 = ( n1004 & n1052 ) | ( n1004 & n1090 ) | ( n1052 & n1090 ) ;
  assign n1093 = ( n1004 & n1091 ) | ( n1004 & ~n1092 ) | ( n1091 & ~n1092 ) ;
  assign n1094 = ( n1031 & n1034 ) | ( n1031 & n1093 ) | ( n1034 & n1093 ) ;
  assign n1095 = ( ~n1031 & n1034 ) | ( ~n1031 & n1093 ) | ( n1034 & n1093 ) ;
  assign n1096 = ( n1031 & ~n1094 ) | ( n1031 & n1095 ) | ( ~n1094 & n1095 ) ;
  assign n1097 = ( n978 & ~n1038 ) | ( n978 & n1039 ) | ( ~n1038 & n1039 ) ;
  assign n1098 = x8 & x24 ;
  assign n1099 = x7 & x25 ;
  assign n1100 = x6 & x26 ;
  assign n1101 = ( ~n1098 & n1099 ) | ( ~n1098 & n1100 ) | ( n1099 & n1100 ) ;
  assign n1102 = ( n1098 & n1099 ) | ( n1098 & n1100 ) | ( n1099 & n1100 ) ;
  assign n1103 = ( n1098 & n1101 ) | ( n1098 & ~n1102 ) | ( n1101 & ~n1102 ) ;
  assign n1104 = x9 & x23 ;
  assign n1105 = x4 & x28 ;
  assign n1106 = x5 & x27 ;
  assign n1107 = ( ~n1104 & n1105 ) | ( ~n1104 & n1106 ) | ( n1105 & n1106 ) ;
  assign n1108 = ( n1104 & n1105 ) | ( n1104 & n1106 ) | ( n1105 & n1106 ) ;
  assign n1109 = ( n1104 & n1107 ) | ( n1104 & ~n1108 ) | ( n1107 & ~n1108 ) ;
  assign n1110 = ( n1097 & n1103 ) | ( n1097 & n1109 ) | ( n1103 & n1109 ) ;
  assign n1111 = ( ~n1097 & n1103 ) | ( ~n1097 & n1109 ) | ( n1103 & n1109 ) ;
  assign n1112 = ( n1097 & ~n1110 ) | ( n1097 & n1111 ) | ( ~n1110 & n1111 ) ;
  assign n1113 = x16 & n1036 ;
  assign n1114 = x0 & x32 ;
  assign n1115 = x2 & x30 ;
  assign n1116 = ( ~n1113 & n1114 ) | ( ~n1113 & n1115 ) | ( n1114 & n1115 ) ;
  assign n1117 = ( n1113 & n1114 ) | ( n1113 & n1115 ) | ( n1114 & n1115 ) ;
  assign n1118 = ( n1113 & n1116 ) | ( n1113 & ~n1117 ) | ( n1116 & ~n1117 ) ;
  assign n1119 = x11 & x21 ;
  assign n1120 = x13 & x19 ;
  assign n1121 = x12 & x20 ;
  assign n1122 = ( ~n1119 & n1120 ) | ( ~n1119 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1123 = ( n1119 & n1120 ) | ( n1119 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1124 = ( n1119 & n1122 ) | ( n1119 & ~n1123 ) | ( n1122 & ~n1123 ) ;
  assign n1125 = x14 & x18 ;
  assign n1126 = x3 & x29 ;
  assign n1127 = x10 & x22 ;
  assign n1128 = ( ~n1125 & n1126 ) | ( ~n1125 & n1127 ) | ( n1126 & n1127 ) ;
  assign n1129 = ( n1125 & n1126 ) | ( n1125 & n1127 ) | ( n1126 & n1127 ) ;
  assign n1130 = ( n1125 & n1128 ) | ( n1125 & ~n1129 ) | ( n1128 & ~n1129 ) ;
  assign n1131 = ( ~n1118 & n1124 ) | ( ~n1118 & n1130 ) | ( n1124 & n1130 ) ;
  assign n1132 = ( n1118 & n1124 ) | ( n1118 & n1130 ) | ( n1124 & n1130 ) ;
  assign n1133 = ( n1118 & n1131 ) | ( n1118 & ~n1132 ) | ( n1131 & ~n1132 ) ;
  assign n1134 = ( n1048 & n1112 ) | ( n1048 & n1133 ) | ( n1112 & n1133 ) ;
  assign n1135 = ( ~n1048 & n1112 ) | ( ~n1048 & n1133 ) | ( n1112 & n1133 ) ;
  assign n1136 = ( n1048 & ~n1134 ) | ( n1048 & n1135 ) | ( ~n1134 & n1135 ) ;
  assign n1137 = ( n1057 & ~n1063 ) | ( n1057 & n1071 ) | ( ~n1063 & n1071 ) ;
  assign n1138 = ( n1057 & n1063 ) | ( n1057 & n1071 ) | ( n1063 & n1071 ) ;
  assign n1139 = ( n1063 & n1137 ) | ( n1063 & ~n1138 ) | ( n1137 & ~n1138 ) ;
  assign n1140 = x15 & x17 ;
  assign n1141 = x1 & x31 ;
  assign n1142 = n1140 & n1141 ;
  assign n1143 = n1140 | n1141 ;
  assign n1144 = ~n1142 & n1143 ;
  assign n1145 = ( n1077 & n1083 ) | ( n1077 & n1144 ) | ( n1083 & n1144 ) ;
  assign n1146 = ( ~n1077 & n1083 ) | ( ~n1077 & n1144 ) | ( n1083 & n1144 ) ;
  assign n1147 = ( n1077 & ~n1145 ) | ( n1077 & n1146 ) | ( ~n1145 & n1146 ) ;
  assign n1148 = ( ~n1042 & n1139 ) | ( ~n1042 & n1147 ) | ( n1139 & n1147 ) ;
  assign n1149 = ( n1042 & n1139 ) | ( n1042 & n1147 ) | ( n1139 & n1147 ) ;
  assign n1150 = ( n1042 & n1148 ) | ( n1042 & ~n1149 ) | ( n1148 & ~n1149 ) ;
  assign n1151 = ( n1045 & ~n1065 ) | ( n1045 & n1086 ) | ( ~n1065 & n1086 ) ;
  assign n1152 = ( n1045 & n1065 ) | ( n1045 & n1086 ) | ( n1065 & n1086 ) ;
  assign n1153 = ( n1065 & n1151 ) | ( n1065 & ~n1152 ) | ( n1151 & ~n1152 ) ;
  assign n1154 = ( n1089 & n1150 ) | ( n1089 & n1153 ) | ( n1150 & n1153 ) ;
  assign n1155 = ( ~n1089 & n1150 ) | ( ~n1089 & n1153 ) | ( n1150 & n1153 ) ;
  assign n1156 = ( n1089 & ~n1154 ) | ( n1089 & n1155 ) | ( ~n1154 & n1155 ) ;
  assign n1157 = ( ~n1051 & n1136 ) | ( ~n1051 & n1156 ) | ( n1136 & n1156 ) ;
  assign n1158 = ( n1051 & n1136 ) | ( n1051 & n1156 ) | ( n1136 & n1156 ) ;
  assign n1159 = ( n1051 & n1157 ) | ( n1051 & ~n1158 ) | ( n1157 & ~n1158 ) ;
  assign n1160 = ( n1092 & n1094 ) | ( n1092 & n1159 ) | ( n1094 & n1159 ) ;
  assign n1161 = ( ~n1092 & n1094 ) | ( ~n1092 & n1159 ) | ( n1094 & n1159 ) ;
  assign n1162 = ( n1092 & ~n1160 ) | ( n1092 & n1161 ) | ( ~n1160 & n1161 ) ;
  assign n1163 = ( ~n1117 & n1123 ) | ( ~n1117 & n1129 ) | ( n1123 & n1129 ) ;
  assign n1164 = ( n1117 & n1123 ) | ( n1117 & n1129 ) | ( n1123 & n1129 ) ;
  assign n1165 = ( n1117 & n1163 ) | ( n1117 & ~n1164 ) | ( n1163 & ~n1164 ) ;
  assign n1166 = x2 & x31 ;
  assign n1167 = x0 & x33 ;
  assign n1168 = x11 & x22 ;
  assign n1169 = ( ~n1166 & n1167 ) | ( ~n1166 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1170 = ( n1166 & n1167 ) | ( n1166 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1171 = ( n1166 & n1169 ) | ( n1166 & ~n1170 ) | ( n1169 & ~n1170 ) ;
  assign n1172 = ( ~n1102 & n1108 ) | ( ~n1102 & n1171 ) | ( n1108 & n1171 ) ;
  assign n1173 = ( n1102 & n1108 ) | ( n1102 & n1171 ) | ( n1108 & n1171 ) ;
  assign n1174 = ( n1102 & n1172 ) | ( n1102 & ~n1173 ) | ( n1172 & ~n1173 ) ;
  assign n1175 = x3 & x30 ;
  assign n1176 = x4 & x29 ;
  assign n1177 = x9 & x24 ;
  assign n1178 = ( ~n1175 & n1176 ) | ( ~n1175 & n1177 ) | ( n1176 & n1177 ) ;
  assign n1179 = ( n1175 & n1176 ) | ( n1175 & n1177 ) | ( n1176 & n1177 ) ;
  assign n1180 = ( n1175 & n1178 ) | ( n1175 & ~n1179 ) | ( n1178 & ~n1179 ) ;
  assign n1181 = x7 & x26 ;
  assign n1182 = x16 & x17 ;
  assign n1183 = x15 & x18 ;
  assign n1184 = ( ~n1181 & n1182 ) | ( ~n1181 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1185 = ( n1181 & n1182 ) | ( n1181 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1186 = ( n1181 & n1184 ) | ( n1181 & ~n1185 ) | ( n1184 & ~n1185 ) ;
  assign n1187 = x5 & x28 ;
  assign n1188 = x8 & x25 ;
  assign n1189 = x6 & x27 ;
  assign n1190 = ( ~n1187 & n1188 ) | ( ~n1187 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1191 = ( n1187 & n1188 ) | ( n1187 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1192 = ( n1187 & n1190 ) | ( n1187 & ~n1191 ) | ( n1190 & ~n1191 ) ;
  assign n1193 = ( ~n1180 & n1186 ) | ( ~n1180 & n1192 ) | ( n1186 & n1192 ) ;
  assign n1194 = ( n1180 & n1186 ) | ( n1180 & n1192 ) | ( n1186 & n1192 ) ;
  assign n1195 = ( n1180 & n1193 ) | ( n1180 & ~n1194 ) | ( n1193 & ~n1194 ) ;
  assign n1196 = ( n1165 & n1174 ) | ( n1165 & n1195 ) | ( n1174 & n1195 ) ;
  assign n1197 = ( ~n1165 & n1174 ) | ( ~n1165 & n1195 ) | ( n1174 & n1195 ) ;
  assign n1198 = ( n1165 & ~n1196 ) | ( n1165 & n1197 ) | ( ~n1196 & n1197 ) ;
  assign n1199 = ( ~n1110 & n1132 ) | ( ~n1110 & n1138 ) | ( n1132 & n1138 ) ;
  assign n1200 = ( n1110 & n1132 ) | ( n1110 & n1138 ) | ( n1132 & n1138 ) ;
  assign n1201 = ( n1110 & n1199 ) | ( n1110 & ~n1200 ) | ( n1199 & ~n1200 ) ;
  assign n1202 = ( ~n1134 & n1198 ) | ( ~n1134 & n1201 ) | ( n1198 & n1201 ) ;
  assign n1203 = ( n1134 & n1198 ) | ( n1134 & n1201 ) | ( n1198 & n1201 ) ;
  assign n1204 = ( n1134 & n1202 ) | ( n1134 & ~n1203 ) | ( n1202 & ~n1203 ) ;
  assign n1205 = x10 & x23 ;
  assign n1206 = x1 & x32 ;
  assign n1207 = x17 & n1206 ;
  assign n1208 = x17 | n1206 ;
  assign n1209 = ~n1207 & n1208 ;
  assign n1210 = ( n1142 & n1205 ) | ( n1142 & n1209 ) | ( n1205 & n1209 ) ;
  assign n1211 = ( ~n1142 & n1205 ) | ( ~n1142 & n1209 ) | ( n1205 & n1209 ) ;
  assign n1212 = ( n1142 & ~n1210 ) | ( n1142 & n1211 ) | ( ~n1210 & n1211 ) ;
  assign n1213 = x12 & x21 ;
  assign n1214 = x13 & x20 ;
  assign n1215 = x14 & x19 ;
  assign n1216 = ( ~n1213 & n1214 ) | ( ~n1213 & n1215 ) | ( n1214 & n1215 ) ;
  assign n1217 = ( n1213 & n1214 ) | ( n1213 & n1215 ) | ( n1214 & n1215 ) ;
  assign n1218 = ( n1213 & n1216 ) | ( n1213 & ~n1217 ) | ( n1216 & ~n1217 ) ;
  assign n1219 = ( ~n1145 & n1212 ) | ( ~n1145 & n1218 ) | ( n1212 & n1218 ) ;
  assign n1220 = ( n1145 & n1212 ) | ( n1145 & n1218 ) | ( n1212 & n1218 ) ;
  assign n1221 = ( n1145 & n1219 ) | ( n1145 & ~n1220 ) | ( n1219 & ~n1220 ) ;
  assign n1222 = ( ~n1149 & n1152 ) | ( ~n1149 & n1221 ) | ( n1152 & n1221 ) ;
  assign n1223 = ( n1149 & n1152 ) | ( n1149 & n1221 ) | ( n1152 & n1221 ) ;
  assign n1224 = ( n1149 & n1222 ) | ( n1149 & ~n1223 ) | ( n1222 & ~n1223 ) ;
  assign n1225 = ( ~n1154 & n1204 ) | ( ~n1154 & n1224 ) | ( n1204 & n1224 ) ;
  assign n1226 = ( n1154 & n1204 ) | ( n1154 & n1224 ) | ( n1204 & n1224 ) ;
  assign n1227 = ( n1154 & n1225 ) | ( n1154 & ~n1226 ) | ( n1225 & ~n1226 ) ;
  assign n1228 = ( ~n1158 & n1160 ) | ( ~n1158 & n1227 ) | ( n1160 & n1227 ) ;
  assign n1229 = ( n1158 & n1160 ) | ( n1158 & n1227 ) | ( n1160 & n1227 ) ;
  assign n1230 = ( n1158 & n1228 ) | ( n1158 & ~n1229 ) | ( n1228 & ~n1229 ) ;
  assign n1231 = ( n1170 & ~n1179 ) | ( n1170 & n1191 ) | ( ~n1179 & n1191 ) ;
  assign n1232 = ( n1170 & n1179 ) | ( n1170 & n1191 ) | ( n1179 & n1191 ) ;
  assign n1233 = ( n1179 & n1231 ) | ( n1179 & ~n1232 ) | ( n1231 & ~n1232 ) ;
  assign n1234 = x16 & x18 ;
  assign n1235 = x1 & x33 ;
  assign n1236 = n1234 & n1235 ;
  assign n1237 = n1234 | n1235 ;
  assign n1238 = ~n1236 & n1237 ;
  assign n1239 = ( ~n1185 & n1207 ) | ( ~n1185 & n1238 ) | ( n1207 & n1238 ) ;
  assign n1240 = ( n1185 & n1207 ) | ( n1185 & n1238 ) | ( n1207 & n1238 ) ;
  assign n1241 = ( n1185 & n1239 ) | ( n1185 & ~n1240 ) | ( n1239 & ~n1240 ) ;
  assign n1242 = ( ~n1194 & n1233 ) | ( ~n1194 & n1241 ) | ( n1233 & n1241 ) ;
  assign n1243 = ( n1194 & n1233 ) | ( n1194 & n1241 ) | ( n1233 & n1241 ) ;
  assign n1244 = ( n1194 & n1242 ) | ( n1194 & ~n1243 ) | ( n1242 & ~n1243 ) ;
  assign n1245 = x2 & x32 ;
  assign n1246 = x12 & x22 ;
  assign n1247 = x11 & x23 ;
  assign n1248 = ( ~n1245 & n1246 ) | ( ~n1245 & n1247 ) | ( n1246 & n1247 ) ;
  assign n1249 = ( n1245 & n1246 ) | ( n1245 & n1247 ) | ( n1246 & n1247 ) ;
  assign n1250 = ( n1245 & n1248 ) | ( n1245 & ~n1249 ) | ( n1248 & ~n1249 ) ;
  assign n1251 = ( n1210 & n1217 ) | ( n1210 & n1250 ) | ( n1217 & n1250 ) ;
  assign n1252 = ( ~n1210 & n1217 ) | ( ~n1210 & n1250 ) | ( n1217 & n1250 ) ;
  assign n1253 = ( n1210 & ~n1251 ) | ( n1210 & n1252 ) | ( ~n1251 & n1252 ) ;
  assign n1254 = x6 & x28 ;
  assign n1255 = x8 & x26 ;
  assign n1256 = x7 & x27 ;
  assign n1257 = ( ~n1254 & n1255 ) | ( ~n1254 & n1256 ) | ( n1255 & n1256 ) ;
  assign n1258 = ( n1254 & n1255 ) | ( n1254 & n1256 ) | ( n1255 & n1256 ) ;
  assign n1259 = ( n1254 & n1257 ) | ( n1254 & ~n1258 ) | ( n1257 & ~n1258 ) ;
  assign n1260 = x10 & x24 ;
  assign n1261 = x5 & x29 ;
  assign n1262 = x9 & x25 ;
  assign n1263 = ( ~n1260 & n1261 ) | ( ~n1260 & n1262 ) | ( n1261 & n1262 ) ;
  assign n1264 = ( n1260 & n1261 ) | ( n1260 & n1262 ) | ( n1261 & n1262 ) ;
  assign n1265 = ( n1260 & n1263 ) | ( n1260 & ~n1264 ) | ( n1263 & ~n1264 ) ;
  assign n1266 = x13 & x21 ;
  assign n1267 = x14 & x20 ;
  assign n1268 = x15 & x19 ;
  assign n1269 = ( ~n1266 & n1267 ) | ( ~n1266 & n1268 ) | ( n1267 & n1268 ) ;
  assign n1270 = ( n1266 & n1267 ) | ( n1266 & n1268 ) | ( n1267 & n1268 ) ;
  assign n1271 = ( n1266 & n1269 ) | ( n1266 & ~n1270 ) | ( n1269 & ~n1270 ) ;
  assign n1272 = ( ~n1259 & n1265 ) | ( ~n1259 & n1271 ) | ( n1265 & n1271 ) ;
  assign n1273 = ( n1259 & n1265 ) | ( n1259 & n1271 ) | ( n1265 & n1271 ) ;
  assign n1274 = ( n1259 & n1272 ) | ( n1259 & ~n1273 ) | ( n1272 & ~n1273 ) ;
  assign n1275 = ( n1220 & n1253 ) | ( n1220 & n1274 ) | ( n1253 & n1274 ) ;
  assign n1276 = ( ~n1220 & n1253 ) | ( ~n1220 & n1274 ) | ( n1253 & n1274 ) ;
  assign n1277 = ( n1220 & ~n1275 ) | ( n1220 & n1276 ) | ( ~n1275 & n1276 ) ;
  assign n1278 = ( ~n1223 & n1244 ) | ( ~n1223 & n1277 ) | ( n1244 & n1277 ) ;
  assign n1279 = ( n1223 & n1244 ) | ( n1223 & n1277 ) | ( n1244 & n1277 ) ;
  assign n1280 = ( n1223 & n1278 ) | ( n1223 & ~n1279 ) | ( n1278 & ~n1279 ) ;
  assign n1281 = x0 & x34 ;
  assign n1282 = x3 & x31 ;
  assign n1283 = x4 & x30 ;
  assign n1284 = ( ~n1281 & n1282 ) | ( ~n1281 & n1283 ) | ( n1282 & n1283 ) ;
  assign n1285 = ( n1281 & n1282 ) | ( n1281 & n1283 ) | ( n1282 & n1283 ) ;
  assign n1286 = ( n1281 & n1284 ) | ( n1281 & ~n1285 ) | ( n1284 & ~n1285 ) ;
  assign n1287 = ( ~n1164 & n1173 ) | ( ~n1164 & n1286 ) | ( n1173 & n1286 ) ;
  assign n1288 = ( n1164 & n1173 ) | ( n1164 & n1286 ) | ( n1173 & n1286 ) ;
  assign n1289 = ( n1164 & n1287 ) | ( n1164 & ~n1288 ) | ( n1287 & ~n1288 ) ;
  assign n1290 = ( ~n1196 & n1200 ) | ( ~n1196 & n1289 ) | ( n1200 & n1289 ) ;
  assign n1291 = ( n1196 & n1200 ) | ( n1196 & n1289 ) | ( n1200 & n1289 ) ;
  assign n1292 = ( n1196 & n1290 ) | ( n1196 & ~n1291 ) | ( n1290 & ~n1291 ) ;
  assign n1293 = ( n1203 & n1280 ) | ( n1203 & n1292 ) | ( n1280 & n1292 ) ;
  assign n1294 = ( n1203 & ~n1280 ) | ( n1203 & n1292 ) | ( ~n1280 & n1292 ) ;
  assign n1295 = ( n1280 & ~n1293 ) | ( n1280 & n1294 ) | ( ~n1293 & n1294 ) ;
  assign n1296 = ( n1226 & n1229 ) | ( n1226 & n1295 ) | ( n1229 & n1295 ) ;
  assign n1297 = ( ~n1226 & n1229 ) | ( ~n1226 & n1295 ) | ( n1229 & n1295 ) ;
  assign n1298 = ( n1226 & ~n1296 ) | ( n1226 & n1297 ) | ( ~n1296 & n1297 ) ;
  assign n1299 = ( n1232 & n1240 ) | ( n1232 & ~n1251 ) | ( n1240 & ~n1251 ) ;
  assign n1300 = ( n1232 & n1240 ) | ( n1232 & n1251 ) | ( n1240 & n1251 ) ;
  assign n1301 = ( n1251 & n1299 ) | ( n1251 & ~n1300 ) | ( n1299 & ~n1300 ) ;
  assign n1302 = ( n1243 & n1275 ) | ( n1243 & n1301 ) | ( n1275 & n1301 ) ;
  assign n1303 = ( n1243 & n1275 ) | ( n1243 & ~n1301 ) | ( n1275 & ~n1301 ) ;
  assign n1304 = ( n1301 & ~n1302 ) | ( n1301 & n1303 ) | ( ~n1302 & n1303 ) ;
  assign n1305 = ( n1249 & ~n1270 ) | ( n1249 & n1285 ) | ( ~n1270 & n1285 ) ;
  assign n1306 = ( n1249 & n1270 ) | ( n1249 & n1285 ) | ( n1270 & n1285 ) ;
  assign n1307 = ( n1270 & n1305 ) | ( n1270 & ~n1306 ) | ( n1305 & ~n1306 ) ;
  assign n1308 = ~x1 & x18 ;
  assign n1309 = ( x1 & x18 ) | ( x1 & x34 ) | ( x18 & x34 ) ;
  assign n1310 = x18 & x34 ;
  assign n1311 = ( n1308 & n1309 ) | ( n1308 & ~n1310 ) | ( n1309 & ~n1310 ) ;
  assign n1312 = ( ~n1258 & n1264 ) | ( ~n1258 & n1311 ) | ( n1264 & n1311 ) ;
  assign n1313 = ( n1258 & n1264 ) | ( n1258 & n1311 ) | ( n1264 & n1311 ) ;
  assign n1314 = ( n1258 & n1312 ) | ( n1258 & ~n1313 ) | ( n1312 & ~n1313 ) ;
  assign n1315 = ( ~n1273 & n1307 ) | ( ~n1273 & n1314 ) | ( n1307 & n1314 ) ;
  assign n1316 = ( n1273 & n1307 ) | ( n1273 & n1314 ) | ( n1307 & n1314 ) ;
  assign n1317 = ( n1273 & n1315 ) | ( n1273 & ~n1316 ) | ( n1315 & ~n1316 ) ;
  assign n1318 = x7 & x28 ;
  assign n1319 = x17 & x18 ;
  assign n1320 = x16 & x19 ;
  assign n1321 = ( ~n1318 & n1319 ) | ( ~n1318 & n1320 ) | ( n1319 & n1320 ) ;
  assign n1322 = ( n1318 & n1319 ) | ( n1318 & n1320 ) | ( n1319 & n1320 ) ;
  assign n1323 = ( n1318 & n1321 ) | ( n1318 & ~n1322 ) | ( n1321 & ~n1322 ) ;
  assign n1324 = x4 & x31 ;
  assign n1325 = x9 & x26 ;
  assign n1326 = x10 & x25 ;
  assign n1327 = ( ~n1324 & n1325 ) | ( ~n1324 & n1326 ) | ( n1325 & n1326 ) ;
  assign n1328 = ( n1324 & n1325 ) | ( n1324 & n1326 ) | ( n1325 & n1326 ) ;
  assign n1329 = ( n1324 & n1327 ) | ( n1324 & ~n1328 ) | ( n1327 & ~n1328 ) ;
  assign n1330 = x5 & x30 ;
  assign n1331 = x8 & x27 ;
  assign n1332 = x6 & x29 ;
  assign n1333 = ( ~n1330 & n1331 ) | ( ~n1330 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1334 = ( n1330 & n1331 ) | ( n1330 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1335 = ( n1330 & n1333 ) | ( n1330 & ~n1334 ) | ( n1333 & ~n1334 ) ;
  assign n1336 = ( ~n1323 & n1329 ) | ( ~n1323 & n1335 ) | ( n1329 & n1335 ) ;
  assign n1337 = ( n1323 & n1329 ) | ( n1323 & n1335 ) | ( n1329 & n1335 ) ;
  assign n1338 = ( n1323 & n1336 ) | ( n1323 & ~n1337 ) | ( n1336 & ~n1337 ) ;
  assign n1339 = x0 & x35 ;
  assign n1340 = x2 & x33 ;
  assign n1341 = ( ~n1236 & n1339 ) | ( ~n1236 & n1340 ) | ( n1339 & n1340 ) ;
  assign n1342 = ( n1236 & n1339 ) | ( n1236 & n1340 ) | ( n1339 & n1340 ) ;
  assign n1343 = ( n1236 & n1341 ) | ( n1236 & ~n1342 ) | ( n1341 & ~n1342 ) ;
  assign n1344 = x13 & x22 ;
  assign n1345 = x15 & x20 ;
  assign n1346 = x14 & x21 ;
  assign n1347 = ( ~n1344 & n1345 ) | ( ~n1344 & n1346 ) | ( n1345 & n1346 ) ;
  assign n1348 = ( n1344 & n1345 ) | ( n1344 & n1346 ) | ( n1345 & n1346 ) ;
  assign n1349 = ( n1344 & n1347 ) | ( n1344 & ~n1348 ) | ( n1347 & ~n1348 ) ;
  assign n1350 = x3 & x32 ;
  assign n1351 = x12 & x23 ;
  assign n1352 = x11 & x24 ;
  assign n1353 = ( ~n1350 & n1351 ) | ( ~n1350 & n1352 ) | ( n1351 & n1352 ) ;
  assign n1354 = ( n1350 & n1351 ) | ( n1350 & n1352 ) | ( n1351 & n1352 ) ;
  assign n1355 = ( n1350 & n1353 ) | ( n1350 & ~n1354 ) | ( n1353 & ~n1354 ) ;
  assign n1356 = ( ~n1343 & n1349 ) | ( ~n1343 & n1355 ) | ( n1349 & n1355 ) ;
  assign n1357 = ( n1343 & n1349 ) | ( n1343 & n1355 ) | ( n1349 & n1355 ) ;
  assign n1358 = ( n1343 & n1356 ) | ( n1343 & ~n1357 ) | ( n1356 & ~n1357 ) ;
  assign n1359 = ( n1288 & n1338 ) | ( n1288 & n1358 ) | ( n1338 & n1358 ) ;
  assign n1360 = ( ~n1288 & n1338 ) | ( ~n1288 & n1358 ) | ( n1338 & n1358 ) ;
  assign n1361 = ( n1288 & ~n1359 ) | ( n1288 & n1360 ) | ( ~n1359 & n1360 ) ;
  assign n1362 = ( ~n1291 & n1317 ) | ( ~n1291 & n1361 ) | ( n1317 & n1361 ) ;
  assign n1363 = ( n1291 & n1317 ) | ( n1291 & n1361 ) | ( n1317 & n1361 ) ;
  assign n1364 = ( n1291 & n1362 ) | ( n1291 & ~n1363 ) | ( n1362 & ~n1363 ) ;
  assign n1365 = ( ~n1279 & n1304 ) | ( ~n1279 & n1364 ) | ( n1304 & n1364 ) ;
  assign n1366 = ( n1279 & n1304 ) | ( n1279 & n1364 ) | ( n1304 & n1364 ) ;
  assign n1367 = ( n1279 & n1365 ) | ( n1279 & ~n1366 ) | ( n1365 & ~n1366 ) ;
  assign n1368 = ( ~n1293 & n1296 ) | ( ~n1293 & n1367 ) | ( n1296 & n1367 ) ;
  assign n1369 = ( n1293 & n1296 ) | ( n1293 & n1367 ) | ( n1296 & n1367 ) ;
  assign n1370 = ( n1293 & n1368 ) | ( n1293 & ~n1369 ) | ( n1368 & ~n1369 ) ;
  assign n1371 = ( n1322 & n1328 ) | ( n1322 & n1334 ) | ( n1328 & n1334 ) ;
  assign n1372 = ( ~n1322 & n1328 ) | ( ~n1322 & n1334 ) | ( n1328 & n1334 ) ;
  assign n1373 = ( n1322 & ~n1371 ) | ( n1322 & n1372 ) | ( ~n1371 & n1372 ) ;
  assign n1374 = ( n1342 & n1348 ) | ( n1342 & n1354 ) | ( n1348 & n1354 ) ;
  assign n1375 = ( ~n1342 & n1348 ) | ( ~n1342 & n1354 ) | ( n1348 & n1354 ) ;
  assign n1376 = ( n1342 & ~n1374 ) | ( n1342 & n1375 ) | ( ~n1374 & n1375 ) ;
  assign n1377 = ( ~n1337 & n1373 ) | ( ~n1337 & n1376 ) | ( n1373 & n1376 ) ;
  assign n1378 = ( n1337 & n1373 ) | ( n1337 & n1376 ) | ( n1373 & n1376 ) ;
  assign n1379 = ( n1337 & n1377 ) | ( n1337 & ~n1378 ) | ( n1377 & ~n1378 ) ;
  assign n1380 = x6 & x30 ;
  assign n1381 = x7 & x29 ;
  assign n1382 = x8 & x28 ;
  assign n1383 = ( ~n1380 & n1381 ) | ( ~n1380 & n1382 ) | ( n1381 & n1382 ) ;
  assign n1384 = ( n1380 & n1381 ) | ( n1380 & n1382 ) | ( n1381 & n1382 ) ;
  assign n1385 = ( n1380 & n1383 ) | ( n1380 & ~n1384 ) | ( n1383 & ~n1384 ) ;
  assign n1386 = x10 & x26 ;
  assign n1387 = x5 & x31 ;
  assign n1388 = x9 & x27 ;
  assign n1389 = ( ~n1386 & n1387 ) | ( ~n1386 & n1388 ) | ( n1387 & n1388 ) ;
  assign n1390 = ( n1386 & n1387 ) | ( n1386 & n1388 ) | ( n1387 & n1388 ) ;
  assign n1391 = ( n1386 & n1389 ) | ( n1386 & ~n1390 ) | ( n1389 & ~n1390 ) ;
  assign n1392 = x2 & x34 ;
  assign n1393 = x12 & x24 ;
  assign n1394 = x13 & x23 ;
  assign n1395 = ( ~n1392 & n1393 ) | ( ~n1392 & n1394 ) | ( n1393 & n1394 ) ;
  assign n1396 = ( n1392 & n1393 ) | ( n1392 & n1394 ) | ( n1393 & n1394 ) ;
  assign n1397 = ( n1392 & n1395 ) | ( n1392 & ~n1396 ) | ( n1395 & ~n1396 ) ;
  assign n1398 = ( ~n1385 & n1391 ) | ( ~n1385 & n1397 ) | ( n1391 & n1397 ) ;
  assign n1399 = ( n1385 & n1391 ) | ( n1385 & n1397 ) | ( n1391 & n1397 ) ;
  assign n1400 = ( n1385 & n1398 ) | ( n1385 & ~n1399 ) | ( n1398 & ~n1399 ) ;
  assign n1401 = x14 & x22 ;
  assign n1402 = x15 & x21 ;
  assign n1403 = x16 & x20 ;
  assign n1404 = ( ~n1401 & n1402 ) | ( ~n1401 & n1403 ) | ( n1402 & n1403 ) ;
  assign n1405 = ( n1401 & n1402 ) | ( n1401 & n1403 ) | ( n1402 & n1403 ) ;
  assign n1406 = ( n1401 & n1404 ) | ( n1401 & ~n1405 ) | ( n1404 & ~n1405 ) ;
  assign n1407 = x3 & x33 ;
  assign n1408 = x11 & x25 ;
  assign n1409 = x4 & x32 ;
  assign n1410 = ( ~n1407 & n1408 ) | ( ~n1407 & n1409 ) | ( n1408 & n1409 ) ;
  assign n1411 = ( n1407 & n1408 ) | ( n1407 & n1409 ) | ( n1408 & n1409 ) ;
  assign n1412 = ( n1407 & n1410 ) | ( n1407 & ~n1411 ) | ( n1410 & ~n1411 ) ;
  assign n1413 = x34 & n439 ;
  assign n1414 = x0 & x36 ;
  assign n1415 = x17 & x19 ;
  assign n1416 = x1 & x35 ;
  assign n1417 = n1415 & n1416 ;
  assign n1418 = n1415 | n1416 ;
  assign n1419 = ~n1417 & n1418 ;
  assign n1420 = ( n1413 & n1414 ) | ( n1413 & n1419 ) | ( n1414 & n1419 ) ;
  assign n1421 = ( ~n1413 & n1414 ) | ( ~n1413 & n1419 ) | ( n1414 & n1419 ) ;
  assign n1422 = ( n1413 & ~n1420 ) | ( n1413 & n1421 ) | ( ~n1420 & n1421 ) ;
  assign n1423 = ( ~n1406 & n1412 ) | ( ~n1406 & n1422 ) | ( n1412 & n1422 ) ;
  assign n1424 = ( n1406 & n1412 ) | ( n1406 & n1422 ) | ( n1412 & n1422 ) ;
  assign n1425 = ( n1406 & n1423 ) | ( n1406 & ~n1424 ) | ( n1423 & ~n1424 ) ;
  assign n1426 = ( ~n1300 & n1400 ) | ( ~n1300 & n1425 ) | ( n1400 & n1425 ) ;
  assign n1427 = ( n1300 & n1400 ) | ( n1300 & n1425 ) | ( n1400 & n1425 ) ;
  assign n1428 = ( n1300 & n1426 ) | ( n1300 & ~n1427 ) | ( n1426 & ~n1427 ) ;
  assign n1429 = ( ~n1302 & n1379 ) | ( ~n1302 & n1428 ) | ( n1379 & n1428 ) ;
  assign n1430 = ( n1302 & n1379 ) | ( n1302 & n1428 ) | ( n1379 & n1428 ) ;
  assign n1431 = ( n1302 & n1429 ) | ( n1302 & ~n1430 ) | ( n1429 & ~n1430 ) ;
  assign n1432 = ( n1306 & ~n1313 ) | ( n1306 & n1357 ) | ( ~n1313 & n1357 ) ;
  assign n1433 = ( n1306 & n1313 ) | ( n1306 & n1357 ) | ( n1313 & n1357 ) ;
  assign n1434 = ( n1313 & n1432 ) | ( n1313 & ~n1433 ) | ( n1432 & ~n1433 ) ;
  assign n1435 = ( n1316 & n1359 ) | ( n1316 & n1434 ) | ( n1359 & n1434 ) ;
  assign n1436 = ( n1316 & n1359 ) | ( n1316 & ~n1434 ) | ( n1359 & ~n1434 ) ;
  assign n1437 = ( n1434 & ~n1435 ) | ( n1434 & n1436 ) | ( ~n1435 & n1436 ) ;
  assign n1438 = ( n1363 & n1431 ) | ( n1363 & n1437 ) | ( n1431 & n1437 ) ;
  assign n1439 = ( ~n1363 & n1431 ) | ( ~n1363 & n1437 ) | ( n1431 & n1437 ) ;
  assign n1440 = ( n1363 & ~n1438 ) | ( n1363 & n1439 ) | ( ~n1438 & n1439 ) ;
  assign n1441 = ( n1366 & n1369 ) | ( n1366 & n1440 ) | ( n1369 & n1440 ) ;
  assign n1442 = ( ~n1366 & n1369 ) | ( ~n1366 & n1440 ) | ( n1369 & n1440 ) ;
  assign n1443 = ( n1366 & ~n1441 ) | ( n1366 & n1442 ) | ( ~n1441 & n1442 ) ;
  assign n1444 = x8 & x29 ;
  assign n1445 = x18 & x19 ;
  assign n1446 = x17 & x20 ;
  assign n1447 = ( ~n1444 & n1445 ) | ( ~n1444 & n1446 ) | ( n1445 & n1446 ) ;
  assign n1448 = ( n1444 & n1445 ) | ( n1444 & n1446 ) | ( n1445 & n1446 ) ;
  assign n1449 = ( n1444 & n1447 ) | ( n1444 & ~n1448 ) | ( n1447 & ~n1448 ) ;
  assign n1450 = x11 & x26 ;
  assign n1451 = x5 & x32 ;
  assign n1452 = x10 & x27 ;
  assign n1453 = ( ~n1450 & n1451 ) | ( ~n1450 & n1452 ) | ( n1451 & n1452 ) ;
  assign n1454 = ( n1450 & n1451 ) | ( n1450 & n1452 ) | ( n1451 & n1452 ) ;
  assign n1455 = ( n1450 & n1453 ) | ( n1450 & ~n1454 ) | ( n1453 & ~n1454 ) ;
  assign n1456 = ( ~n1374 & n1449 ) | ( ~n1374 & n1455 ) | ( n1449 & n1455 ) ;
  assign n1457 = ( n1374 & n1449 ) | ( n1374 & n1455 ) | ( n1449 & n1455 ) ;
  assign n1458 = ( n1374 & n1456 ) | ( n1374 & ~n1457 ) | ( n1456 & ~n1457 ) ;
  assign n1459 = x16 & x21 ;
  assign n1460 = x2 & x35 ;
  assign n1461 = x3 & x34 ;
  assign n1462 = ( ~n1459 & n1460 ) | ( ~n1459 & n1461 ) | ( n1460 & n1461 ) ;
  assign n1463 = ( n1459 & n1460 ) | ( n1459 & n1461 ) | ( n1460 & n1461 ) ;
  assign n1464 = ( n1459 & n1462 ) | ( n1459 & ~n1463 ) | ( n1462 & ~n1463 ) ;
  assign n1465 = x9 & x28 ;
  assign n1466 = x6 & x31 ;
  assign n1467 = x7 & x30 ;
  assign n1468 = ( ~n1465 & n1466 ) | ( ~n1465 & n1467 ) | ( n1466 & n1467 ) ;
  assign n1469 = ( n1465 & n1466 ) | ( n1465 & n1467 ) | ( n1466 & n1467 ) ;
  assign n1470 = ( n1465 & n1468 ) | ( n1465 & ~n1469 ) | ( n1468 & ~n1469 ) ;
  assign n1471 = x0 & x37 ;
  assign n1472 = x12 & x25 ;
  assign n1473 = x4 & x33 ;
  assign n1474 = ( ~n1471 & n1472 ) | ( ~n1471 & n1473 ) | ( n1472 & n1473 ) ;
  assign n1475 = ( n1471 & n1472 ) | ( n1471 & n1473 ) | ( n1472 & n1473 ) ;
  assign n1476 = ( n1471 & n1474 ) | ( n1471 & ~n1475 ) | ( n1474 & ~n1475 ) ;
  assign n1477 = ( ~n1464 & n1470 ) | ( ~n1464 & n1476 ) | ( n1470 & n1476 ) ;
  assign n1478 = ( n1464 & n1470 ) | ( n1464 & n1476 ) | ( n1470 & n1476 ) ;
  assign n1479 = ( n1464 & n1477 ) | ( n1464 & ~n1478 ) | ( n1477 & ~n1478 ) ;
  assign n1480 = ( n1433 & n1458 ) | ( n1433 & n1479 ) | ( n1458 & n1479 ) ;
  assign n1481 = ( ~n1433 & n1458 ) | ( ~n1433 & n1479 ) | ( n1458 & n1479 ) ;
  assign n1482 = ( n1433 & ~n1480 ) | ( n1433 & n1481 ) | ( ~n1480 & n1481 ) ;
  assign n1483 = x13 & x24 ;
  assign n1484 = x14 & x23 ;
  assign n1485 = x15 & x22 ;
  assign n1486 = ( ~n1483 & n1484 ) | ( ~n1483 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1487 = ( n1483 & n1484 ) | ( n1483 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1488 = ( n1483 & n1486 ) | ( n1483 & ~n1487 ) | ( n1486 & ~n1487 ) ;
  assign n1489 = ( ~n1390 & n1420 ) | ( ~n1390 & n1488 ) | ( n1420 & n1488 ) ;
  assign n1490 = ( n1390 & n1420 ) | ( n1390 & n1488 ) | ( n1420 & n1488 ) ;
  assign n1491 = ( n1390 & n1489 ) | ( n1390 & ~n1490 ) | ( n1489 & ~n1490 ) ;
  assign n1492 = ( n1396 & n1405 ) | ( n1396 & ~n1411 ) | ( n1405 & ~n1411 ) ;
  assign n1493 = ( n1396 & n1405 ) | ( n1396 & n1411 ) | ( n1405 & n1411 ) ;
  assign n1494 = ( n1411 & n1492 ) | ( n1411 & ~n1493 ) | ( n1492 & ~n1493 ) ;
  assign n1495 = ( ~n1424 & n1491 ) | ( ~n1424 & n1494 ) | ( n1491 & n1494 ) ;
  assign n1496 = ( n1424 & n1491 ) | ( n1424 & n1494 ) | ( n1491 & n1494 ) ;
  assign n1497 = ( n1424 & n1495 ) | ( n1424 & ~n1496 ) | ( n1495 & ~n1496 ) ;
  assign n1498 = ( ~n1435 & n1482 ) | ( ~n1435 & n1497 ) | ( n1482 & n1497 ) ;
  assign n1499 = ( n1435 & n1482 ) | ( n1435 & n1497 ) | ( n1482 & n1497 ) ;
  assign n1500 = ( n1435 & n1498 ) | ( n1435 & ~n1499 ) | ( n1498 & ~n1499 ) ;
  assign n1501 = ~x36 & n1417 ;
  assign n1502 = x1 & x36 ;
  assign n1503 = x19 | n1502 ;
  assign n1504 = x36 & n471 ;
  assign n1505 = ( n1417 & n1503 ) | ( n1417 & ~n1504 ) | ( n1503 & ~n1504 ) ;
  assign n1506 = ( n1384 & n1501 ) | ( n1384 & n1505 ) | ( n1501 & n1505 ) ;
  assign n1507 = ( n1384 & ~n1501 ) | ( n1384 & n1505 ) | ( ~n1501 & n1505 ) ;
  assign n1508 = ( n1501 & ~n1506 ) | ( n1501 & n1507 ) | ( ~n1506 & n1507 ) ;
  assign n1509 = ( n1371 & n1399 ) | ( n1371 & n1508 ) | ( n1399 & n1508 ) ;
  assign n1510 = ( ~n1371 & n1399 ) | ( ~n1371 & n1508 ) | ( n1399 & n1508 ) ;
  assign n1511 = ( n1371 & ~n1509 ) | ( n1371 & n1510 ) | ( ~n1509 & n1510 ) ;
  assign n1512 = ( n1378 & n1427 ) | ( n1378 & n1511 ) | ( n1427 & n1511 ) ;
  assign n1513 = ( ~n1378 & n1427 ) | ( ~n1378 & n1511 ) | ( n1427 & n1511 ) ;
  assign n1514 = ( n1378 & ~n1512 ) | ( n1378 & n1513 ) | ( ~n1512 & n1513 ) ;
  assign n1515 = ( ~n1430 & n1500 ) | ( ~n1430 & n1514 ) | ( n1500 & n1514 ) ;
  assign n1516 = ( n1430 & n1500 ) | ( n1430 & n1514 ) | ( n1500 & n1514 ) ;
  assign n1517 = ( n1430 & n1515 ) | ( n1430 & ~n1516 ) | ( n1515 & ~n1516 ) ;
  assign n1518 = ( ~n1438 & n1441 ) | ( ~n1438 & n1517 ) | ( n1441 & n1517 ) ;
  assign n1519 = ( n1438 & n1441 ) | ( n1438 & n1517 ) | ( n1441 & n1517 ) ;
  assign n1520 = ( n1438 & n1518 ) | ( n1438 & ~n1519 ) | ( n1518 & ~n1519 ) ;
  assign n1521 = ( n1463 & ~n1475 ) | ( n1463 & n1487 ) | ( ~n1475 & n1487 ) ;
  assign n1522 = ( n1463 & n1475 ) | ( n1463 & n1487 ) | ( n1475 & n1487 ) ;
  assign n1523 = ( n1475 & n1521 ) | ( n1475 & ~n1522 ) | ( n1521 & ~n1522 ) ;
  assign n1524 = x9 & x29 ;
  assign n1525 = x7 & x31 ;
  assign n1526 = x8 & x30 ;
  assign n1527 = ( ~n1524 & n1525 ) | ( ~n1524 & n1526 ) | ( n1525 & n1526 ) ;
  assign n1528 = ( n1524 & n1525 ) | ( n1524 & n1526 ) | ( n1525 & n1526 ) ;
  assign n1529 = ( n1524 & n1527 ) | ( n1524 & ~n1528 ) | ( n1527 & ~n1528 ) ;
  assign n1530 = x5 & x33 ;
  assign n1531 = x6 & x32 ;
  assign n1532 = x10 & x28 ;
  assign n1533 = ( ~n1530 & n1531 ) | ( ~n1530 & n1532 ) | ( n1531 & n1532 ) ;
  assign n1534 = ( n1530 & n1531 ) | ( n1530 & n1532 ) | ( n1531 & n1532 ) ;
  assign n1535 = ( n1530 & n1533 ) | ( n1530 & ~n1534 ) | ( n1533 & ~n1534 ) ;
  assign n1536 = x15 & x23 ;
  assign n1537 = x16 & x22 ;
  assign n1538 = x17 & x21 ;
  assign n1539 = ( ~n1536 & n1537 ) | ( ~n1536 & n1538 ) | ( n1537 & n1538 ) ;
  assign n1540 = ( n1536 & n1537 ) | ( n1536 & n1538 ) | ( n1537 & n1538 ) ;
  assign n1541 = ( n1536 & n1539 ) | ( n1536 & ~n1540 ) | ( n1539 & ~n1540 ) ;
  assign n1542 = ( ~n1529 & n1535 ) | ( ~n1529 & n1541 ) | ( n1535 & n1541 ) ;
  assign n1543 = ( n1529 & n1535 ) | ( n1529 & n1541 ) | ( n1535 & n1541 ) ;
  assign n1544 = ( n1529 & n1542 ) | ( n1529 & ~n1543 ) | ( n1542 & ~n1543 ) ;
  assign n1545 = ( ~n1457 & n1523 ) | ( ~n1457 & n1544 ) | ( n1523 & n1544 ) ;
  assign n1546 = ( n1457 & n1523 ) | ( n1457 & n1544 ) | ( n1523 & n1544 ) ;
  assign n1547 = ( n1457 & n1545 ) | ( n1457 & ~n1546 ) | ( n1545 & ~n1546 ) ;
  assign n1548 = ( ~n1480 & n1496 ) | ( ~n1480 & n1547 ) | ( n1496 & n1547 ) ;
  assign n1549 = ( n1480 & n1496 ) | ( n1480 & n1547 ) | ( n1496 & n1547 ) ;
  assign n1550 = ( n1480 & n1548 ) | ( n1480 & ~n1549 ) | ( n1548 & ~n1549 ) ;
  assign n1551 = x18 & x20 ;
  assign n1552 = x1 & x37 ;
  assign n1553 = n1551 & n1552 ;
  assign n1554 = n1551 | n1552 ;
  assign n1555 = ~n1553 & n1554 ;
  assign n1556 = ( n1448 & n1469 ) | ( n1448 & n1555 ) | ( n1469 & n1555 ) ;
  assign n1557 = ( ~n1448 & n1469 ) | ( ~n1448 & n1555 ) | ( n1469 & n1555 ) ;
  assign n1558 = ( n1448 & ~n1556 ) | ( n1448 & n1557 ) | ( ~n1556 & n1557 ) ;
  assign n1559 = ( n1478 & n1490 ) | ( n1478 & n1558 ) | ( n1490 & n1558 ) ;
  assign n1560 = ( ~n1478 & n1490 ) | ( ~n1478 & n1558 ) | ( n1490 & n1558 ) ;
  assign n1561 = ( n1478 & ~n1559 ) | ( n1478 & n1560 ) | ( ~n1559 & n1560 ) ;
  assign n1562 = x12 & x26 ;
  assign n1563 = x4 & x34 ;
  assign n1564 = x11 & x27 ;
  assign n1565 = ( ~n1562 & n1563 ) | ( ~n1562 & n1564 ) | ( n1563 & n1564 ) ;
  assign n1566 = ( n1562 & n1563 ) | ( n1562 & n1564 ) | ( n1563 & n1564 ) ;
  assign n1567 = ( n1562 & n1565 ) | ( n1562 & ~n1566 ) | ( n1565 & ~n1566 ) ;
  assign n1568 = ( ~n1493 & n1506 ) | ( ~n1493 & n1567 ) | ( n1506 & n1567 ) ;
  assign n1569 = ( n1493 & n1506 ) | ( n1493 & n1567 ) | ( n1506 & n1567 ) ;
  assign n1570 = ( n1493 & n1568 ) | ( n1493 & ~n1569 ) | ( n1568 & ~n1569 ) ;
  assign n1571 = x3 & x35 ;
  assign n1572 = x13 & x25 ;
  assign n1573 = x14 & x24 ;
  assign n1574 = ( ~n1571 & n1572 ) | ( ~n1571 & n1573 ) | ( n1572 & n1573 ) ;
  assign n1575 = ( n1571 & n1572 ) | ( n1571 & n1573 ) | ( n1572 & n1573 ) ;
  assign n1576 = ( n1571 & n1574 ) | ( n1571 & ~n1575 ) | ( n1574 & ~n1575 ) ;
  assign n1577 = x2 & x38 ;
  assign n1578 = n1414 & n1577 ;
  assign n1579 = x0 & x38 ;
  assign n1580 = x2 & x36 ;
  assign n1581 = n1579 | n1580 ;
  assign n1582 = ( n1504 & n1578 ) | ( n1504 & n1581 ) | ( n1578 & n1581 ) ;
  assign n1583 = ( ~n1504 & n1578 ) | ( ~n1504 & n1581 ) | ( n1578 & n1581 ) ;
  assign n1584 = ( n1504 & ~n1582 ) | ( n1504 & n1583 ) | ( ~n1582 & n1583 ) ;
  assign n1585 = ( ~n1454 & n1576 ) | ( ~n1454 & n1584 ) | ( n1576 & n1584 ) ;
  assign n1586 = ( n1454 & n1576 ) | ( n1454 & n1584 ) | ( n1576 & n1584 ) ;
  assign n1587 = ( n1454 & n1585 ) | ( n1454 & ~n1586 ) | ( n1585 & ~n1586 ) ;
  assign n1588 = ( n1509 & n1570 ) | ( n1509 & n1587 ) | ( n1570 & n1587 ) ;
  assign n1589 = ( ~n1509 & n1570 ) | ( ~n1509 & n1587 ) | ( n1570 & n1587 ) ;
  assign n1590 = ( n1509 & ~n1588 ) | ( n1509 & n1589 ) | ( ~n1588 & n1589 ) ;
  assign n1591 = ( ~n1512 & n1561 ) | ( ~n1512 & n1590 ) | ( n1561 & n1590 ) ;
  assign n1592 = ( n1512 & n1561 ) | ( n1512 & n1590 ) | ( n1561 & n1590 ) ;
  assign n1593 = ( n1512 & n1591 ) | ( n1512 & ~n1592 ) | ( n1591 & ~n1592 ) ;
  assign n1594 = ( ~n1499 & n1550 ) | ( ~n1499 & n1593 ) | ( n1550 & n1593 ) ;
  assign n1595 = ( n1499 & n1550 ) | ( n1499 & n1593 ) | ( n1550 & n1593 ) ;
  assign n1596 = ( n1499 & n1594 ) | ( n1499 & ~n1595 ) | ( n1594 & ~n1595 ) ;
  assign n1597 = ( n1516 & n1519 ) | ( n1516 & n1596 ) | ( n1519 & n1596 ) ;
  assign n1598 = ( ~n1516 & n1519 ) | ( ~n1516 & n1596 ) | ( n1519 & n1596 ) ;
  assign n1599 = ( n1516 & ~n1597 ) | ( n1516 & n1598 ) | ( ~n1597 & n1598 ) ;
  assign n1600 = ~x1 & x20 ;
  assign n1601 = ( x1 & x20 ) | ( x1 & x38 ) | ( x20 & x38 ) ;
  assign n1602 = x20 & x38 ;
  assign n1603 = ( n1600 & n1601 ) | ( n1600 & ~n1602 ) | ( n1601 & ~n1602 ) ;
  assign n1604 = x0 & x39 ;
  assign n1605 = ( n1553 & n1603 ) | ( n1553 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1606 = ( ~n1553 & n1603 ) | ( ~n1553 & n1604 ) | ( n1603 & n1604 ) ;
  assign n1607 = ( n1553 & ~n1605 ) | ( n1553 & n1606 ) | ( ~n1605 & n1606 ) ;
  assign n1608 = ( ~n1522 & n1556 ) | ( ~n1522 & n1607 ) | ( n1556 & n1607 ) ;
  assign n1609 = ( n1522 & n1556 ) | ( n1522 & n1607 ) | ( n1556 & n1607 ) ;
  assign n1610 = ( n1522 & n1608 ) | ( n1522 & ~n1609 ) | ( n1608 & ~n1609 ) ;
  assign n1611 = ( ~n1540 & n1575 ) | ( ~n1540 & n1582 ) | ( n1575 & n1582 ) ;
  assign n1612 = ( n1540 & n1575 ) | ( n1540 & n1582 ) | ( n1575 & n1582 ) ;
  assign n1613 = ( n1540 & n1611 ) | ( n1540 & ~n1612 ) | ( n1611 & ~n1612 ) ;
  assign n1614 = ( n1543 & n1586 ) | ( n1543 & n1613 ) | ( n1586 & n1613 ) ;
  assign n1615 = ( n1543 & n1586 ) | ( n1543 & ~n1613 ) | ( n1586 & ~n1613 ) ;
  assign n1616 = ( n1613 & ~n1614 ) | ( n1613 & n1615 ) | ( ~n1614 & n1615 ) ;
  assign n1617 = ( n1588 & n1610 ) | ( n1588 & n1616 ) | ( n1610 & n1616 ) ;
  assign n1618 = ( ~n1588 & n1610 ) | ( ~n1588 & n1616 ) | ( n1610 & n1616 ) ;
  assign n1619 = ( n1588 & ~n1617 ) | ( n1588 & n1618 ) | ( ~n1617 & n1618 ) ;
  assign n1620 = x2 & x37 ;
  assign n1621 = x3 & x36 ;
  assign n1622 = x13 & x26 ;
  assign n1623 = ( ~n1620 & n1621 ) | ( ~n1620 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1624 = ( n1620 & n1621 ) | ( n1620 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1625 = ( n1620 & n1623 ) | ( n1620 & ~n1624 ) | ( n1623 & ~n1624 ) ;
  assign n1626 = x6 & x33 ;
  assign n1627 = x9 & x30 ;
  assign n1628 = x7 & x32 ;
  assign n1629 = ( ~n1626 & n1627 ) | ( ~n1626 & n1628 ) | ( n1627 & n1628 ) ;
  assign n1630 = ( n1626 & n1627 ) | ( n1626 & n1628 ) | ( n1627 & n1628 ) ;
  assign n1631 = ( n1626 & n1629 ) | ( n1626 & ~n1630 ) | ( n1629 & ~n1630 ) ;
  assign n1632 = x14 & x25 ;
  assign n1633 = x15 & x24 ;
  assign n1634 = x16 & x23 ;
  assign n1635 = ( ~n1632 & n1633 ) | ( ~n1632 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1636 = ( n1632 & n1633 ) | ( n1632 & n1634 ) | ( n1633 & n1634 ) ;
  assign n1637 = ( n1632 & n1635 ) | ( n1632 & ~n1636 ) | ( n1635 & ~n1636 ) ;
  assign n1638 = ( ~n1625 & n1631 ) | ( ~n1625 & n1637 ) | ( n1631 & n1637 ) ;
  assign n1639 = ( n1625 & n1631 ) | ( n1625 & n1637 ) | ( n1631 & n1637 ) ;
  assign n1640 = ( n1625 & n1638 ) | ( n1625 & ~n1639 ) | ( n1638 & ~n1639 ) ;
  assign n1641 = ( n1546 & n1559 ) | ( n1546 & n1640 ) | ( n1559 & n1640 ) ;
  assign n1642 = ( ~n1546 & n1559 ) | ( ~n1546 & n1640 ) | ( n1559 & n1640 ) ;
  assign n1643 = ( n1546 & ~n1641 ) | ( n1546 & n1642 ) | ( ~n1641 & n1642 ) ;
  assign n1644 = ( ~n1528 & n1534 ) | ( ~n1528 & n1566 ) | ( n1534 & n1566 ) ;
  assign n1645 = ( n1528 & n1534 ) | ( n1528 & n1566 ) | ( n1534 & n1566 ) ;
  assign n1646 = ( n1528 & n1644 ) | ( n1528 & ~n1645 ) | ( n1644 & ~n1645 ) ;
  assign n1647 = x8 & x31 ;
  assign n1648 = x19 & x20 ;
  assign n1649 = x18 & x21 ;
  assign n1650 = ( ~n1647 & n1648 ) | ( ~n1647 & n1649 ) | ( n1648 & n1649 ) ;
  assign n1651 = ( n1647 & n1648 ) | ( n1647 & n1649 ) | ( n1648 & n1649 ) ;
  assign n1652 = ( n1647 & n1650 ) | ( n1647 & ~n1651 ) | ( n1650 & ~n1651 ) ;
  assign n1653 = x11 & x28 ;
  assign n1654 = x10 & x29 ;
  assign n1655 = x5 & x34 ;
  assign n1656 = ( ~n1653 & n1654 ) | ( ~n1653 & n1655 ) | ( n1654 & n1655 ) ;
  assign n1657 = ( n1653 & n1654 ) | ( n1653 & n1655 ) | ( n1654 & n1655 ) ;
  assign n1658 = ( n1653 & n1656 ) | ( n1653 & ~n1657 ) | ( n1656 & ~n1657 ) ;
  assign n1659 = x17 & x22 ;
  assign n1660 = x4 & x35 ;
  assign n1661 = x12 & x27 ;
  assign n1662 = ( ~n1659 & n1660 ) | ( ~n1659 & n1661 ) | ( n1660 & n1661 ) ;
  assign n1663 = ( n1659 & n1660 ) | ( n1659 & n1661 ) | ( n1660 & n1661 ) ;
  assign n1664 = ( n1659 & n1662 ) | ( n1659 & ~n1663 ) | ( n1662 & ~n1663 ) ;
  assign n1665 = ( ~n1652 & n1658 ) | ( ~n1652 & n1664 ) | ( n1658 & n1664 ) ;
  assign n1666 = ( n1652 & n1658 ) | ( n1652 & n1664 ) | ( n1658 & n1664 ) ;
  assign n1667 = ( n1652 & n1665 ) | ( n1652 & ~n1666 ) | ( n1665 & ~n1666 ) ;
  assign n1668 = ( ~n1569 & n1646 ) | ( ~n1569 & n1667 ) | ( n1646 & n1667 ) ;
  assign n1669 = ( n1569 & n1646 ) | ( n1569 & n1667 ) | ( n1646 & n1667 ) ;
  assign n1670 = ( n1569 & n1668 ) | ( n1569 & ~n1669 ) | ( n1668 & ~n1669 ) ;
  assign n1671 = ( n1549 & n1643 ) | ( n1549 & n1670 ) | ( n1643 & n1670 ) ;
  assign n1672 = ( ~n1549 & n1643 ) | ( ~n1549 & n1670 ) | ( n1643 & n1670 ) ;
  assign n1673 = ( n1549 & ~n1671 ) | ( n1549 & n1672 ) | ( ~n1671 & n1672 ) ;
  assign n1674 = ( n1592 & n1619 ) | ( n1592 & n1673 ) | ( n1619 & n1673 ) ;
  assign n1675 = ( ~n1592 & n1619 ) | ( ~n1592 & n1673 ) | ( n1619 & n1673 ) ;
  assign n1676 = ( n1592 & ~n1674 ) | ( n1592 & n1675 ) | ( ~n1674 & n1675 ) ;
  assign n1677 = ( n1595 & n1597 ) | ( n1595 & n1676 ) | ( n1597 & n1676 ) ;
  assign n1678 = ( ~n1595 & n1597 ) | ( ~n1595 & n1676 ) | ( n1597 & n1676 ) ;
  assign n1679 = ( n1595 & ~n1677 ) | ( n1595 & n1678 ) | ( ~n1677 & n1678 ) ;
  assign n1680 = ( n1624 & ~n1657 ) | ( n1624 & n1663 ) | ( ~n1657 & n1663 ) ;
  assign n1681 = ( n1624 & n1657 ) | ( n1624 & n1663 ) | ( n1657 & n1663 ) ;
  assign n1682 = ( n1657 & n1680 ) | ( n1657 & ~n1681 ) | ( n1680 & ~n1681 ) ;
  assign n1683 = ( n1639 & n1666 ) | ( n1639 & n1682 ) | ( n1666 & n1682 ) ;
  assign n1684 = ( ~n1639 & n1666 ) | ( ~n1639 & n1682 ) | ( n1666 & n1682 ) ;
  assign n1685 = ( n1639 & ~n1683 ) | ( n1639 & n1684 ) | ( ~n1683 & n1684 ) ;
  assign n1686 = ( ~n1641 & n1669 ) | ( ~n1641 & n1685 ) | ( n1669 & n1685 ) ;
  assign n1687 = ( n1641 & n1669 ) | ( n1641 & n1685 ) | ( n1669 & n1685 ) ;
  assign n1688 = ( n1641 & n1686 ) | ( n1641 & ~n1687 ) | ( n1686 & ~n1687 ) ;
  assign n1689 = ( ~n1605 & n1630 ) | ( ~n1605 & n1636 ) | ( n1630 & n1636 ) ;
  assign n1690 = ( n1605 & n1630 ) | ( n1605 & n1636 ) | ( n1630 & n1636 ) ;
  assign n1691 = ( n1605 & n1689 ) | ( n1605 & ~n1690 ) | ( n1689 & ~n1690 ) ;
  assign n1692 = x4 & x36 ;
  assign n1693 = x12 & x28 ;
  assign n1694 = x5 & x35 ;
  assign n1695 = ( ~n1692 & n1693 ) | ( ~n1692 & n1694 ) | ( n1693 & n1694 ) ;
  assign n1696 = ( n1692 & n1693 ) | ( n1692 & n1694 ) | ( n1693 & n1694 ) ;
  assign n1697 = ( n1692 & n1695 ) | ( n1692 & ~n1696 ) | ( n1695 & ~n1696 ) ;
  assign n1698 = x7 & x33 ;
  assign n1699 = x9 & x31 ;
  assign n1700 = x8 & x32 ;
  assign n1701 = ( ~n1698 & n1699 ) | ( ~n1698 & n1700 ) | ( n1699 & n1700 ) ;
  assign n1702 = ( n1698 & n1699 ) | ( n1698 & n1700 ) | ( n1699 & n1700 ) ;
  assign n1703 = ( n1698 & n1701 ) | ( n1698 & ~n1702 ) | ( n1701 & ~n1702 ) ;
  assign n1704 = x18 & x22 ;
  assign n1705 = x0 & x40 ;
  assign n1706 = ( ~n1577 & n1704 ) | ( ~n1577 & n1705 ) | ( n1704 & n1705 ) ;
  assign n1707 = ( n1577 & n1704 ) | ( n1577 & n1705 ) | ( n1704 & n1705 ) ;
  assign n1708 = ( n1577 & n1706 ) | ( n1577 & ~n1707 ) | ( n1706 & ~n1707 ) ;
  assign n1709 = ( ~n1697 & n1703 ) | ( ~n1697 & n1708 ) | ( n1703 & n1708 ) ;
  assign n1710 = ( n1697 & n1703 ) | ( n1697 & n1708 ) | ( n1703 & n1708 ) ;
  assign n1711 = ( n1697 & n1709 ) | ( n1697 & ~n1710 ) | ( n1709 & ~n1710 ) ;
  assign n1712 = ( ~n1609 & n1691 ) | ( ~n1609 & n1711 ) | ( n1691 & n1711 ) ;
  assign n1713 = ( n1609 & n1691 ) | ( n1609 & n1711 ) | ( n1691 & n1711 ) ;
  assign n1714 = ( n1609 & n1712 ) | ( n1609 & ~n1713 ) | ( n1712 & ~n1713 ) ;
  assign n1715 = x11 & x29 ;
  assign n1716 = x6 & x34 ;
  assign n1717 = x10 & x30 ;
  assign n1718 = ( ~n1715 & n1716 ) | ( ~n1715 & n1717 ) | ( n1716 & n1717 ) ;
  assign n1719 = ( n1715 & n1716 ) | ( n1715 & n1717 ) | ( n1716 & n1717 ) ;
  assign n1720 = ( n1715 & n1718 ) | ( n1715 & ~n1719 ) | ( n1718 & ~n1719 ) ;
  assign n1721 = x15 & x25 ;
  assign n1722 = x16 & x24 ;
  assign n1723 = x17 & x23 ;
  assign n1724 = ( ~n1721 & n1722 ) | ( ~n1721 & n1723 ) | ( n1722 & n1723 ) ;
  assign n1725 = ( n1721 & n1722 ) | ( n1721 & n1723 ) | ( n1722 & n1723 ) ;
  assign n1726 = ( n1721 & n1724 ) | ( n1721 & ~n1725 ) | ( n1724 & ~n1725 ) ;
  assign n1727 = x3 & x37 ;
  assign n1728 = x13 & x27 ;
  assign n1729 = ( ~n825 & n1727 ) | ( ~n825 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1730 = ( n825 & n1727 ) | ( n825 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1731 = ( n825 & n1729 ) | ( n825 & ~n1730 ) | ( n1729 & ~n1730 ) ;
  assign n1732 = ( ~n1720 & n1726 ) | ( ~n1720 & n1731 ) | ( n1726 & n1731 ) ;
  assign n1733 = ( n1720 & n1726 ) | ( n1720 & n1731 ) | ( n1726 & n1731 ) ;
  assign n1734 = ( n1720 & n1732 ) | ( n1720 & ~n1733 ) | ( n1732 & ~n1733 ) ;
  assign n1735 = x38 & n538 ;
  assign n1736 = x19 & x21 ;
  assign n1737 = x1 & x39 ;
  assign n1738 = n1736 & n1737 ;
  assign n1739 = n1736 | n1737 ;
  assign n1740 = ~n1738 & n1739 ;
  assign n1741 = ( n1651 & n1735 ) | ( n1651 & n1740 ) | ( n1735 & n1740 ) ;
  assign n1742 = ( n1651 & ~n1735 ) | ( n1651 & n1740 ) | ( ~n1735 & n1740 ) ;
  assign n1743 = ( n1735 & ~n1741 ) | ( n1735 & n1742 ) | ( ~n1741 & n1742 ) ;
  assign n1744 = ( ~n1612 & n1645 ) | ( ~n1612 & n1743 ) | ( n1645 & n1743 ) ;
  assign n1745 = ( n1612 & n1645 ) | ( n1612 & n1743 ) | ( n1645 & n1743 ) ;
  assign n1746 = ( n1612 & n1744 ) | ( n1612 & ~n1745 ) | ( n1744 & ~n1745 ) ;
  assign n1747 = ( ~n1614 & n1734 ) | ( ~n1614 & n1746 ) | ( n1734 & n1746 ) ;
  assign n1748 = ( n1614 & n1734 ) | ( n1614 & n1746 ) | ( n1734 & n1746 ) ;
  assign n1749 = ( n1614 & n1747 ) | ( n1614 & ~n1748 ) | ( n1747 & ~n1748 ) ;
  assign n1750 = ( n1617 & n1714 ) | ( n1617 & n1749 ) | ( n1714 & n1749 ) ;
  assign n1751 = ( ~n1617 & n1714 ) | ( ~n1617 & n1749 ) | ( n1714 & n1749 ) ;
  assign n1752 = ( n1617 & ~n1750 ) | ( n1617 & n1751 ) | ( ~n1750 & n1751 ) ;
  assign n1753 = ( n1671 & n1688 ) | ( n1671 & n1752 ) | ( n1688 & n1752 ) ;
  assign n1754 = ( n1671 & ~n1688 ) | ( n1671 & n1752 ) | ( ~n1688 & n1752 ) ;
  assign n1755 = ( n1688 & ~n1753 ) | ( n1688 & n1754 ) | ( ~n1753 & n1754 ) ;
  assign n1756 = ( ~n1674 & n1677 ) | ( ~n1674 & n1755 ) | ( n1677 & n1755 ) ;
  assign n1757 = ( n1674 & n1677 ) | ( n1674 & n1755 ) | ( n1677 & n1755 ) ;
  assign n1758 = ( n1674 & n1756 ) | ( n1674 & ~n1757 ) | ( n1756 & ~n1757 ) ;
  assign n1759 = ~x1 & x21 ;
  assign n1760 = ( x1 & x21 ) | ( x1 & x40 ) | ( x21 & x40 ) ;
  assign n1761 = x21 & x40 ;
  assign n1762 = ( n1759 & n1760 ) | ( n1759 & ~n1761 ) | ( n1760 & ~n1761 ) ;
  assign n1763 = ( ~n1702 & n1719 ) | ( ~n1702 & n1762 ) | ( n1719 & n1762 ) ;
  assign n1764 = ( n1702 & n1719 ) | ( n1702 & n1762 ) | ( n1719 & n1762 ) ;
  assign n1765 = ( n1702 & n1763 ) | ( n1702 & ~n1764 ) | ( n1763 & ~n1764 ) ;
  assign n1766 = ( n1707 & ~n1725 ) | ( n1707 & n1730 ) | ( ~n1725 & n1730 ) ;
  assign n1767 = ( n1707 & n1725 ) | ( n1707 & n1730 ) | ( n1725 & n1730 ) ;
  assign n1768 = ( n1725 & n1766 ) | ( n1725 & ~n1767 ) | ( n1766 & ~n1767 ) ;
  assign n1769 = ( n1710 & n1765 ) | ( n1710 & n1768 ) | ( n1765 & n1768 ) ;
  assign n1770 = ( n1710 & ~n1765 ) | ( n1710 & n1768 ) | ( ~n1765 & n1768 ) ;
  assign n1771 = ( n1765 & ~n1769 ) | ( n1765 & n1770 ) | ( ~n1769 & n1770 ) ;
  assign n1772 = ( n1713 & n1748 ) | ( n1713 & n1771 ) | ( n1748 & n1771 ) ;
  assign n1773 = ( ~n1713 & n1748 ) | ( ~n1713 & n1771 ) | ( n1748 & n1771 ) ;
  assign n1774 = ( n1713 & ~n1772 ) | ( n1713 & n1773 ) | ( ~n1772 & n1773 ) ;
  assign n1775 = ( n1681 & ~n1690 ) | ( n1681 & n1733 ) | ( ~n1690 & n1733 ) ;
  assign n1776 = ( n1681 & n1690 ) | ( n1681 & n1733 ) | ( n1690 & n1733 ) ;
  assign n1777 = ( n1690 & n1775 ) | ( n1690 & ~n1776 ) | ( n1775 & ~n1776 ) ;
  assign n1778 = x0 & x41 ;
  assign n1779 = x2 & x39 ;
  assign n1780 = n1778 | n1779 ;
  assign n1781 = x2 & x41 ;
  assign n1782 = n1604 & n1781 ;
  assign n1783 = ( n1738 & n1780 ) | ( n1738 & n1782 ) | ( n1780 & n1782 ) ;
  assign n1784 = ( ~n1738 & n1780 ) | ( ~n1738 & n1782 ) | ( n1780 & n1782 ) ;
  assign n1785 = ( n1738 & ~n1783 ) | ( n1738 & n1784 ) | ( ~n1783 & n1784 ) ;
  assign n1786 = x3 & x38 ;
  assign n1787 = x13 & x28 ;
  assign n1788 = x15 & x26 ;
  assign n1789 = ( ~n1786 & n1787 ) | ( ~n1786 & n1788 ) | ( n1787 & n1788 ) ;
  assign n1790 = ( n1786 & n1787 ) | ( n1786 & n1788 ) | ( n1787 & n1788 ) ;
  assign n1791 = ( n1786 & n1789 ) | ( n1786 & ~n1790 ) | ( n1789 & ~n1790 ) ;
  assign n1792 = ( ~n1696 & n1785 ) | ( ~n1696 & n1791 ) | ( n1785 & n1791 ) ;
  assign n1793 = ( n1696 & n1785 ) | ( n1696 & n1791 ) | ( n1785 & n1791 ) ;
  assign n1794 = ( n1696 & n1792 ) | ( n1696 & ~n1793 ) | ( n1792 & ~n1793 ) ;
  assign n1795 = ( ~n1683 & n1777 ) | ( ~n1683 & n1794 ) | ( n1777 & n1794 ) ;
  assign n1796 = ( n1683 & n1777 ) | ( n1683 & n1794 ) | ( n1777 & n1794 ) ;
  assign n1797 = ( n1683 & n1795 ) | ( n1683 & ~n1796 ) | ( n1795 & ~n1796 ) ;
  assign n1798 = x10 & x31 ;
  assign n1799 = x9 & x32 ;
  assign n1800 = x7 & x34 ;
  assign n1801 = ( ~n1798 & n1799 ) | ( ~n1798 & n1800 ) | ( n1799 & n1800 ) ;
  assign n1802 = ( n1798 & n1799 ) | ( n1798 & n1800 ) | ( n1799 & n1800 ) ;
  assign n1803 = ( n1798 & n1801 ) | ( n1798 & ~n1802 ) | ( n1801 & ~n1802 ) ;
  assign n1804 = x14 & x27 ;
  assign n1805 = x4 & x37 ;
  assign n1806 = x12 & x29 ;
  assign n1807 = ( ~n1804 & n1805 ) | ( ~n1804 & n1806 ) | ( n1805 & n1806 ) ;
  assign n1808 = ( n1804 & n1805 ) | ( n1804 & n1806 ) | ( n1805 & n1806 ) ;
  assign n1809 = ( n1804 & n1807 ) | ( n1804 & ~n1808 ) | ( n1807 & ~n1808 ) ;
  assign n1810 = x16 & x25 ;
  assign n1811 = x17 & x24 ;
  assign n1812 = x18 & x23 ;
  assign n1813 = ( ~n1810 & n1811 ) | ( ~n1810 & n1812 ) | ( n1811 & n1812 ) ;
  assign n1814 = ( n1810 & n1811 ) | ( n1810 & n1812 ) | ( n1811 & n1812 ) ;
  assign n1815 = ( n1810 & n1813 ) | ( n1810 & ~n1814 ) | ( n1813 & ~n1814 ) ;
  assign n1816 = ( ~n1803 & n1809 ) | ( ~n1803 & n1815 ) | ( n1809 & n1815 ) ;
  assign n1817 = ( n1803 & n1809 ) | ( n1803 & n1815 ) | ( n1809 & n1815 ) ;
  assign n1818 = ( n1803 & n1816 ) | ( n1803 & ~n1817 ) | ( n1816 & ~n1817 ) ;
  assign n1819 = x8 & x33 ;
  assign n1820 = x20 & x21 ;
  assign n1821 = x19 & x22 ;
  assign n1822 = ( ~n1819 & n1820 ) | ( ~n1819 & n1821 ) | ( n1820 & n1821 ) ;
  assign n1823 = ( n1819 & n1820 ) | ( n1819 & n1821 ) | ( n1820 & n1821 ) ;
  assign n1824 = ( n1819 & n1822 ) | ( n1819 & ~n1823 ) | ( n1822 & ~n1823 ) ;
  assign n1825 = x5 & x36 ;
  assign n1826 = x6 & x35 ;
  assign n1827 = x11 & x30 ;
  assign n1828 = ( ~n1825 & n1826 ) | ( ~n1825 & n1827 ) | ( n1826 & n1827 ) ;
  assign n1829 = ( n1825 & n1826 ) | ( n1825 & n1827 ) | ( n1826 & n1827 ) ;
  assign n1830 = ( n1825 & n1828 ) | ( n1825 & ~n1829 ) | ( n1828 & ~n1829 ) ;
  assign n1831 = ( n1741 & n1824 ) | ( n1741 & n1830 ) | ( n1824 & n1830 ) ;
  assign n1832 = ( ~n1741 & n1824 ) | ( ~n1741 & n1830 ) | ( n1824 & n1830 ) ;
  assign n1833 = ( n1741 & ~n1831 ) | ( n1741 & n1832 ) | ( ~n1831 & n1832 ) ;
  assign n1834 = ( n1745 & n1818 ) | ( n1745 & n1833 ) | ( n1818 & n1833 ) ;
  assign n1835 = ( n1745 & ~n1818 ) | ( n1745 & n1833 ) | ( ~n1818 & n1833 ) ;
  assign n1836 = ( n1818 & ~n1834 ) | ( n1818 & n1835 ) | ( ~n1834 & n1835 ) ;
  assign n1837 = ( ~n1687 & n1797 ) | ( ~n1687 & n1836 ) | ( n1797 & n1836 ) ;
  assign n1838 = ( n1687 & n1797 ) | ( n1687 & n1836 ) | ( n1797 & n1836 ) ;
  assign n1839 = ( n1687 & n1837 ) | ( n1687 & ~n1838 ) | ( n1837 & ~n1838 ) ;
  assign n1840 = ( n1750 & n1774 ) | ( n1750 & n1839 ) | ( n1774 & n1839 ) ;
  assign n1841 = ( ~n1750 & n1774 ) | ( ~n1750 & n1839 ) | ( n1774 & n1839 ) ;
  assign n1842 = ( n1750 & ~n1840 ) | ( n1750 & n1841 ) | ( ~n1840 & n1841 ) ;
  assign n1843 = ( ~n1753 & n1757 ) | ( ~n1753 & n1842 ) | ( n1757 & n1842 ) ;
  assign n1844 = ( n1753 & n1757 ) | ( n1753 & n1842 ) | ( n1757 & n1842 ) ;
  assign n1845 = ( n1753 & n1843 ) | ( n1753 & ~n1844 ) | ( n1843 & ~n1844 ) ;
  assign n1846 = ( ~n1767 & n1793 ) | ( ~n1767 & n1817 ) | ( n1793 & n1817 ) ;
  assign n1847 = ( n1767 & n1793 ) | ( n1767 & n1817 ) | ( n1793 & n1817 ) ;
  assign n1848 = ( n1767 & n1846 ) | ( n1767 & ~n1847 ) | ( n1846 & ~n1847 ) ;
  assign n1849 = ( n1796 & n1834 ) | ( n1796 & n1848 ) | ( n1834 & n1848 ) ;
  assign n1850 = ( ~n1796 & n1834 ) | ( ~n1796 & n1848 ) | ( n1834 & n1848 ) ;
  assign n1851 = ( n1796 & ~n1849 ) | ( n1796 & n1850 ) | ( ~n1849 & n1850 ) ;
  assign n1852 = ( n1808 & n1823 ) | ( n1808 & ~n1829 ) | ( n1823 & ~n1829 ) ;
  assign n1853 = ( n1808 & n1823 ) | ( n1808 & n1829 ) | ( n1823 & n1829 ) ;
  assign n1854 = ( n1829 & n1852 ) | ( n1829 & ~n1853 ) | ( n1852 & ~n1853 ) ;
  assign n1855 = ( n1783 & ~n1790 ) | ( n1783 & n1814 ) | ( ~n1790 & n1814 ) ;
  assign n1856 = ( n1783 & n1790 ) | ( n1783 & n1814 ) | ( n1790 & n1814 ) ;
  assign n1857 = ( n1790 & n1855 ) | ( n1790 & ~n1856 ) | ( n1855 & ~n1856 ) ;
  assign n1858 = ( ~n1831 & n1854 ) | ( ~n1831 & n1857 ) | ( n1854 & n1857 ) ;
  assign n1859 = ( n1831 & n1854 ) | ( n1831 & n1857 ) | ( n1854 & n1857 ) ;
  assign n1860 = ( n1831 & n1858 ) | ( n1831 & ~n1859 ) | ( n1858 & ~n1859 ) ;
  assign n1861 = x40 & n582 ;
  assign n1862 = x0 & x42 ;
  assign n1863 = x20 & x22 ;
  assign n1864 = x1 & x41 ;
  assign n1865 = n1863 & n1864 ;
  assign n1866 = n1863 | n1864 ;
  assign n1867 = ~n1865 & n1866 ;
  assign n1868 = ( n1861 & n1862 ) | ( n1861 & n1867 ) | ( n1862 & n1867 ) ;
  assign n1869 = ( ~n1861 & n1862 ) | ( ~n1861 & n1867 ) | ( n1862 & n1867 ) ;
  assign n1870 = ( n1861 & ~n1868 ) | ( n1861 & n1869 ) | ( ~n1868 & n1869 ) ;
  assign n1871 = x13 & x29 ;
  assign n1872 = x5 & x37 ;
  assign n1873 = x12 & x30 ;
  assign n1874 = ( ~n1871 & n1872 ) | ( ~n1871 & n1873 ) | ( n1872 & n1873 ) ;
  assign n1875 = ( n1871 & n1872 ) | ( n1871 & n1873 ) | ( n1872 & n1873 ) ;
  assign n1876 = ( n1871 & n1874 ) | ( n1871 & ~n1875 ) | ( n1874 & ~n1875 ) ;
  assign n1877 = ( ~n1764 & n1870 ) | ( ~n1764 & n1876 ) | ( n1870 & n1876 ) ;
  assign n1878 = ( n1764 & n1870 ) | ( n1764 & n1876 ) | ( n1870 & n1876 ) ;
  assign n1879 = ( n1764 & n1877 ) | ( n1764 & ~n1878 ) | ( n1877 & ~n1878 ) ;
  assign n1880 = ( ~n1769 & n1860 ) | ( ~n1769 & n1879 ) | ( n1860 & n1879 ) ;
  assign n1881 = ( n1769 & n1860 ) | ( n1769 & n1879 ) | ( n1860 & n1879 ) ;
  assign n1882 = ( n1769 & n1880 ) | ( n1769 & ~n1881 ) | ( n1880 & ~n1881 ) ;
  assign n1883 = x10 & x32 ;
  assign n1884 = x8 & x34 ;
  assign n1885 = x9 & x33 ;
  assign n1886 = ( ~n1883 & n1884 ) | ( ~n1883 & n1885 ) | ( n1884 & n1885 ) ;
  assign n1887 = ( n1883 & n1884 ) | ( n1883 & n1885 ) | ( n1884 & n1885 ) ;
  assign n1888 = ( n1883 & n1886 ) | ( n1883 & ~n1887 ) | ( n1886 & ~n1887 ) ;
  assign n1889 = x6 & x36 ;
  assign n1890 = x7 & x35 ;
  assign n1891 = x11 & x31 ;
  assign n1892 = ( ~n1889 & n1890 ) | ( ~n1889 & n1891 ) | ( n1890 & n1891 ) ;
  assign n1893 = ( n1889 & n1890 ) | ( n1889 & n1891 ) | ( n1890 & n1891 ) ;
  assign n1894 = ( n1889 & n1892 ) | ( n1889 & ~n1893 ) | ( n1892 & ~n1893 ) ;
  assign n1895 = ( n1802 & n1888 ) | ( n1802 & n1894 ) | ( n1888 & n1894 ) ;
  assign n1896 = ( ~n1802 & n1888 ) | ( ~n1802 & n1894 ) | ( n1888 & n1894 ) ;
  assign n1897 = ( n1802 & ~n1895 ) | ( n1802 & n1896 ) | ( ~n1895 & n1896 ) ;
  assign n1898 = x2 & x40 ;
  assign n1899 = x3 & x39 ;
  assign n1900 = x16 & x26 ;
  assign n1901 = ( ~n1898 & n1899 ) | ( ~n1898 & n1900 ) | ( n1899 & n1900 ) ;
  assign n1902 = ( n1898 & n1899 ) | ( n1898 & n1900 ) | ( n1899 & n1900 ) ;
  assign n1903 = ( n1898 & n1901 ) | ( n1898 & ~n1902 ) | ( n1901 & ~n1902 ) ;
  assign n1904 = x15 & x27 ;
  assign n1905 = x4 & x38 ;
  assign n1906 = x14 & x28 ;
  assign n1907 = ( ~n1904 & n1905 ) | ( ~n1904 & n1906 ) | ( n1905 & n1906 ) ;
  assign n1908 = ( n1904 & n1905 ) | ( n1904 & n1906 ) | ( n1905 & n1906 ) ;
  assign n1909 = ( n1904 & n1907 ) | ( n1904 & ~n1908 ) | ( n1907 & ~n1908 ) ;
  assign n1910 = x17 & x25 ;
  assign n1911 = x18 & x24 ;
  assign n1912 = x19 & x23 ;
  assign n1913 = ( ~n1910 & n1911 ) | ( ~n1910 & n1912 ) | ( n1911 & n1912 ) ;
  assign n1914 = ( n1910 & n1911 ) | ( n1910 & n1912 ) | ( n1911 & n1912 ) ;
  assign n1915 = ( n1910 & n1913 ) | ( n1910 & ~n1914 ) | ( n1913 & ~n1914 ) ;
  assign n1916 = ( ~n1903 & n1909 ) | ( ~n1903 & n1915 ) | ( n1909 & n1915 ) ;
  assign n1917 = ( n1903 & n1909 ) | ( n1903 & n1915 ) | ( n1909 & n1915 ) ;
  assign n1918 = ( n1903 & n1916 ) | ( n1903 & ~n1917 ) | ( n1916 & ~n1917 ) ;
  assign n1919 = ( ~n1776 & n1897 ) | ( ~n1776 & n1918 ) | ( n1897 & n1918 ) ;
  assign n1920 = ( n1776 & n1897 ) | ( n1776 & n1918 ) | ( n1897 & n1918 ) ;
  assign n1921 = ( n1776 & n1919 ) | ( n1776 & ~n1920 ) | ( n1919 & ~n1920 ) ;
  assign n1922 = ( n1772 & n1882 ) | ( n1772 & n1921 ) | ( n1882 & n1921 ) ;
  assign n1923 = ( ~n1772 & n1882 ) | ( ~n1772 & n1921 ) | ( n1882 & n1921 ) ;
  assign n1924 = ( n1772 & ~n1922 ) | ( n1772 & n1923 ) | ( ~n1922 & n1923 ) ;
  assign n1925 = ( ~n1838 & n1851 ) | ( ~n1838 & n1924 ) | ( n1851 & n1924 ) ;
  assign n1926 = ( n1838 & n1851 ) | ( n1838 & n1924 ) | ( n1851 & n1924 ) ;
  assign n1927 = ( n1838 & n1925 ) | ( n1838 & ~n1926 ) | ( n1925 & ~n1926 ) ;
  assign n1928 = ( ~n1840 & n1844 ) | ( ~n1840 & n1927 ) | ( n1844 & n1927 ) ;
  assign n1929 = ( n1840 & n1844 ) | ( n1840 & n1927 ) | ( n1844 & n1927 ) ;
  assign n1930 = ( n1840 & n1928 ) | ( n1840 & ~n1929 ) | ( n1928 & ~n1929 ) ;
  assign n1931 = x4 & x39 ;
  assign n1932 = x0 & x43 ;
  assign n1933 = x3 & x40 ;
  assign n1934 = ( ~n1931 & n1932 ) | ( ~n1931 & n1933 ) | ( n1932 & n1933 ) ;
  assign n1935 = ( n1931 & n1932 ) | ( n1931 & n1933 ) | ( n1932 & n1933 ) ;
  assign n1936 = ( n1931 & n1934 ) | ( n1931 & ~n1935 ) | ( n1934 & ~n1935 ) ;
  assign n1937 = x17 & x26 ;
  assign n1938 = x19 & x24 ;
  assign n1939 = x18 & x25 ;
  assign n1940 = ( ~n1937 & n1938 ) | ( ~n1937 & n1939 ) | ( n1938 & n1939 ) ;
  assign n1941 = ( n1937 & n1938 ) | ( n1937 & n1939 ) | ( n1938 & n1939 ) ;
  assign n1942 = ( n1937 & n1940 ) | ( n1937 & ~n1941 ) | ( n1940 & ~n1941 ) ;
  assign n1943 = x14 & x29 ;
  assign n1944 = x16 & x27 ;
  assign n1945 = ( ~n923 & n1943 ) | ( ~n923 & n1944 ) | ( n1943 & n1944 ) ;
  assign n1946 = ( n923 & n1943 ) | ( n923 & n1944 ) | ( n1943 & n1944 ) ;
  assign n1947 = ( n923 & n1945 ) | ( n923 & ~n1946 ) | ( n1945 & ~n1946 ) ;
  assign n1948 = ( ~n1936 & n1942 ) | ( ~n1936 & n1947 ) | ( n1942 & n1947 ) ;
  assign n1949 = ( n1936 & n1942 ) | ( n1936 & n1947 ) | ( n1942 & n1947 ) ;
  assign n1950 = ( n1936 & n1948 ) | ( n1936 & ~n1949 ) | ( n1948 & ~n1949 ) ;
  assign n1951 = x9 & x34 ;
  assign n1952 = x21 & x22 ;
  assign n1953 = x20 & x23 ;
  assign n1954 = ( ~n1951 & n1952 ) | ( ~n1951 & n1953 ) | ( n1952 & n1953 ) ;
  assign n1955 = ( n1951 & n1952 ) | ( n1951 & n1953 ) | ( n1952 & n1953 ) ;
  assign n1956 = ( n1951 & n1954 ) | ( n1951 & ~n1955 ) | ( n1954 & ~n1955 ) ;
  assign n1957 = x7 & x36 ;
  assign n1958 = x8 & x35 ;
  assign n1959 = x10 & x33 ;
  assign n1960 = ( ~n1957 & n1958 ) | ( ~n1957 & n1959 ) | ( n1958 & n1959 ) ;
  assign n1961 = ( n1957 & n1958 ) | ( n1957 & n1959 ) | ( n1958 & n1959 ) ;
  assign n1962 = ( n1957 & n1960 ) | ( n1957 & ~n1961 ) | ( n1960 & ~n1961 ) ;
  assign n1963 = x5 & x38 ;
  assign n1964 = x13 & x30 ;
  assign n1965 = ( ~n1781 & n1963 ) | ( ~n1781 & n1964 ) | ( n1963 & n1964 ) ;
  assign n1966 = ( n1781 & n1963 ) | ( n1781 & n1964 ) | ( n1963 & n1964 ) ;
  assign n1967 = ( n1781 & n1965 ) | ( n1781 & ~n1966 ) | ( n1965 & ~n1966 ) ;
  assign n1968 = ( ~n1956 & n1962 ) | ( ~n1956 & n1967 ) | ( n1962 & n1967 ) ;
  assign n1969 = ( n1956 & n1962 ) | ( n1956 & n1967 ) | ( n1962 & n1967 ) ;
  assign n1970 = ( n1956 & n1968 ) | ( n1956 & ~n1969 ) | ( n1968 & ~n1969 ) ;
  assign n1971 = ( n1847 & n1950 ) | ( n1847 & n1970 ) | ( n1950 & n1970 ) ;
  assign n1972 = ( ~n1847 & n1950 ) | ( ~n1847 & n1970 ) | ( n1950 & n1970 ) ;
  assign n1973 = ( n1847 & ~n1971 ) | ( n1847 & n1972 ) | ( ~n1971 & n1972 ) ;
  assign n1974 = ( n1893 & ~n1908 ) | ( n1893 & n1914 ) | ( ~n1908 & n1914 ) ;
  assign n1975 = ( n1893 & n1908 ) | ( n1893 & n1914 ) | ( n1908 & n1914 ) ;
  assign n1976 = ( n1908 & n1974 ) | ( n1908 & ~n1975 ) | ( n1974 & ~n1975 ) ;
  assign n1977 = ( n1868 & n1875 ) | ( n1868 & n1902 ) | ( n1875 & n1902 ) ;
  assign n1978 = ( ~n1868 & n1875 ) | ( ~n1868 & n1902 ) | ( n1875 & n1902 ) ;
  assign n1979 = ( n1868 & ~n1977 ) | ( n1868 & n1978 ) | ( ~n1977 & n1978 ) ;
  assign n1980 = ( ~n1878 & n1976 ) | ( ~n1878 & n1979 ) | ( n1976 & n1979 ) ;
  assign n1981 = ( n1878 & n1976 ) | ( n1878 & n1979 ) | ( n1976 & n1979 ) ;
  assign n1982 = ( n1878 & n1980 ) | ( n1878 & ~n1981 ) | ( n1980 & ~n1981 ) ;
  assign n1983 = x12 & x31 ;
  assign n1984 = x11 & x32 ;
  assign n1985 = x6 & x37 ;
  assign n1986 = ( ~n1983 & n1984 ) | ( ~n1983 & n1985 ) | ( n1984 & n1985 ) ;
  assign n1987 = ( n1983 & n1984 ) | ( n1983 & n1985 ) | ( n1984 & n1985 ) ;
  assign n1988 = ( n1983 & n1986 ) | ( n1983 & ~n1987 ) | ( n1986 & ~n1987 ) ;
  assign n1989 = ( ~n1853 & n1856 ) | ( ~n1853 & n1988 ) | ( n1856 & n1988 ) ;
  assign n1990 = ( n1853 & n1856 ) | ( n1853 & n1988 ) | ( n1856 & n1988 ) ;
  assign n1991 = ( n1853 & n1989 ) | ( n1853 & ~n1990 ) | ( n1989 & ~n1990 ) ;
  assign n1992 = ( n1859 & n1982 ) | ( n1859 & n1991 ) | ( n1982 & n1991 ) ;
  assign n1993 = ( ~n1859 & n1982 ) | ( ~n1859 & n1991 ) | ( n1982 & n1991 ) ;
  assign n1994 = ( n1859 & ~n1992 ) | ( n1859 & n1993 ) | ( ~n1992 & n1993 ) ;
  assign n1995 = ( n1849 & n1973 ) | ( n1849 & n1994 ) | ( n1973 & n1994 ) ;
  assign n1996 = ( ~n1849 & n1973 ) | ( ~n1849 & n1994 ) | ( n1973 & n1994 ) ;
  assign n1997 = ( n1849 & ~n1995 ) | ( n1849 & n1996 ) | ( ~n1995 & n1996 ) ;
  assign n1998 = ~x42 & n1865 ;
  assign n1999 = x1 & x42 ;
  assign n2000 = x22 | n1999 ;
  assign n2001 = x42 & n633 ;
  assign n2002 = ( n1865 & n2000 ) | ( n1865 & ~n2001 ) | ( n2000 & ~n2001 ) ;
  assign n2003 = ( n1887 & n1998 ) | ( n1887 & n2002 ) | ( n1998 & n2002 ) ;
  assign n2004 = ( n1887 & ~n1998 ) | ( n1887 & n2002 ) | ( ~n1998 & n2002 ) ;
  assign n2005 = ( n1998 & ~n2003 ) | ( n1998 & n2004 ) | ( ~n2003 & n2004 ) ;
  assign n2006 = ( n1895 & n1917 ) | ( n1895 & n2005 ) | ( n1917 & n2005 ) ;
  assign n2007 = ( ~n1895 & n1917 ) | ( ~n1895 & n2005 ) | ( n1917 & n2005 ) ;
  assign n2008 = ( n1895 & ~n2006 ) | ( n1895 & n2007 ) | ( ~n2006 & n2007 ) ;
  assign n2009 = ( n1881 & n1920 ) | ( n1881 & n2008 ) | ( n1920 & n2008 ) ;
  assign n2010 = ( ~n1881 & n1920 ) | ( ~n1881 & n2008 ) | ( n1920 & n2008 ) ;
  assign n2011 = ( n1881 & ~n2009 ) | ( n1881 & n2010 ) | ( ~n2009 & n2010 ) ;
  assign n2012 = ( n1922 & n1997 ) | ( n1922 & n2011 ) | ( n1997 & n2011 ) ;
  assign n2013 = ( ~n1922 & n1997 ) | ( ~n1922 & n2011 ) | ( n1997 & n2011 ) ;
  assign n2014 = ( n1922 & ~n2012 ) | ( n1922 & n2013 ) | ( ~n2012 & n2013 ) ;
  assign n2015 = ( n1926 & n1929 ) | ( n1926 & n2014 ) | ( n1929 & n2014 ) ;
  assign n2016 = ( ~n1926 & n1929 ) | ( ~n1926 & n2014 ) | ( n1929 & n2014 ) ;
  assign n2017 = ( n1926 & ~n2015 ) | ( n1926 & n2016 ) | ( ~n2015 & n2016 ) ;
  assign n2018 = ( ~n1935 & n1941 ) | ( ~n1935 & n1966 ) | ( n1941 & n1966 ) ;
  assign n2019 = ( n1935 & n1941 ) | ( n1935 & n1966 ) | ( n1941 & n1966 ) ;
  assign n2020 = ( n1935 & n2018 ) | ( n1935 & ~n2019 ) | ( n2018 & ~n2019 ) ;
  assign n2021 = ( n1949 & n1969 ) | ( n1949 & n2020 ) | ( n1969 & n2020 ) ;
  assign n2022 = ( ~n1949 & n1969 ) | ( ~n1949 & n2020 ) | ( n1969 & n2020 ) ;
  assign n2023 = ( n1949 & ~n2021 ) | ( n1949 & n2022 ) | ( ~n2021 & n2022 ) ;
  assign n2024 = ( n1971 & n1992 ) | ( n1971 & n2023 ) | ( n1992 & n2023 ) ;
  assign n2025 = ( ~n1971 & n1992 ) | ( ~n1971 & n2023 ) | ( n1992 & n2023 ) ;
  assign n2026 = ( n1971 & ~n2024 ) | ( n1971 & n2025 ) | ( ~n2024 & n2025 ) ;
  assign n2027 = x18 & x26 ;
  assign n2028 = x19 & x25 ;
  assign n2029 = x20 & x24 ;
  assign n2030 = ( ~n2027 & n2028 ) | ( ~n2027 & n2029 ) | ( n2028 & n2029 ) ;
  assign n2031 = ( n2027 & n2028 ) | ( n2027 & n2029 ) | ( n2028 & n2029 ) ;
  assign n2032 = ( n2027 & n2030 ) | ( n2027 & ~n2031 ) | ( n2030 & ~n2031 ) ;
  assign n2033 = x6 & x38 ;
  assign n2034 = x11 & x33 ;
  assign n2035 = x7 & x37 ;
  assign n2036 = ( ~n2033 & n2034 ) | ( ~n2033 & n2035 ) | ( n2034 & n2035 ) ;
  assign n2037 = ( n2033 & n2034 ) | ( n2033 & n2035 ) | ( n2034 & n2035 ) ;
  assign n2038 = ( n2033 & n2036 ) | ( n2033 & ~n2037 ) | ( n2036 & ~n2037 ) ;
  assign n2039 = x3 & x41 ;
  assign n2040 = x15 & x29 ;
  assign n2041 = x17 & x27 ;
  assign n2042 = ( ~n2039 & n2040 ) | ( ~n2039 & n2041 ) | ( n2040 & n2041 ) ;
  assign n2043 = ( n2039 & n2040 ) | ( n2039 & n2041 ) | ( n2040 & n2041 ) ;
  assign n2044 = ( n2039 & n2042 ) | ( n2039 & ~n2043 ) | ( n2042 & ~n2043 ) ;
  assign n2045 = ( ~n2032 & n2038 ) | ( ~n2032 & n2044 ) | ( n2038 & n2044 ) ;
  assign n2046 = ( n2032 & n2038 ) | ( n2032 & n2044 ) | ( n2038 & n2044 ) ;
  assign n2047 = ( n2032 & n2045 ) | ( n2032 & ~n2046 ) | ( n2045 & ~n2046 ) ;
  assign n2048 = x5 & x39 ;
  assign n2049 = x12 & x32 ;
  assign n2050 = x13 & x31 ;
  assign n2051 = ( ~n2048 & n2049 ) | ( ~n2048 & n2050 ) | ( n2049 & n2050 ) ;
  assign n2052 = ( n2048 & n2049 ) | ( n2048 & n2050 ) | ( n2049 & n2050 ) ;
  assign n2053 = ( n2048 & n2051 ) | ( n2048 & ~n2052 ) | ( n2051 & ~n2052 ) ;
  assign n2054 = x16 & x28 ;
  assign n2055 = x4 & x40 ;
  assign n2056 = x14 & x30 ;
  assign n2057 = ( ~n2054 & n2055 ) | ( ~n2054 & n2056 ) | ( n2055 & n2056 ) ;
  assign n2058 = ( n2054 & n2055 ) | ( n2054 & n2056 ) | ( n2055 & n2056 ) ;
  assign n2059 = ( n2054 & n2057 ) | ( n2054 & ~n2058 ) | ( n2057 & ~n2058 ) ;
  assign n2060 = x8 & x36 ;
  assign n2061 = x10 & x34 ;
  assign n2062 = x9 & x35 ;
  assign n2063 = ( ~n2060 & n2061 ) | ( ~n2060 & n2062 ) | ( n2061 & n2062 ) ;
  assign n2064 = ( n2060 & n2061 ) | ( n2060 & n2062 ) | ( n2061 & n2062 ) ;
  assign n2065 = ( n2060 & n2063 ) | ( n2060 & ~n2064 ) | ( n2063 & ~n2064 ) ;
  assign n2066 = ( ~n2053 & n2059 ) | ( ~n2053 & n2065 ) | ( n2059 & n2065 ) ;
  assign n2067 = ( n2053 & n2059 ) | ( n2053 & n2065 ) | ( n2059 & n2065 ) ;
  assign n2068 = ( n2053 & n2066 ) | ( n2053 & ~n2067 ) | ( n2066 & ~n2067 ) ;
  assign n2069 = ( n2006 & n2047 ) | ( n2006 & n2068 ) | ( n2047 & n2068 ) ;
  assign n2070 = ( ~n2006 & n2047 ) | ( ~n2006 & n2068 ) | ( n2047 & n2068 ) ;
  assign n2071 = ( n2006 & ~n2069 ) | ( n2006 & n2070 ) | ( ~n2069 & n2070 ) ;
  assign n2072 = x21 & x23 ;
  assign n2073 = x1 & x43 ;
  assign n2074 = n2072 & n2073 ;
  assign n2075 = n2072 | n2073 ;
  assign n2076 = ~n2074 & n2075 ;
  assign n2077 = ( ~n1955 & n1961 ) | ( ~n1955 & n2076 ) | ( n1961 & n2076 ) ;
  assign n2078 = ( n1955 & n1961 ) | ( n1955 & n2076 ) | ( n1961 & n2076 ) ;
  assign n2079 = ( n1955 & n2077 ) | ( n1955 & ~n2078 ) | ( n2077 & ~n2078 ) ;
  assign n2080 = x0 & x44 ;
  assign n2081 = x2 & x42 ;
  assign n2082 = n2080 | n2081 ;
  assign n2083 = x2 & x44 ;
  assign n2084 = n1862 & n2083 ;
  assign n2085 = ( n2001 & n2082 ) | ( n2001 & n2084 ) | ( n2082 & n2084 ) ;
  assign n2086 = ( n2001 & ~n2082 ) | ( n2001 & n2084 ) | ( ~n2082 & n2084 ) ;
  assign n2087 = ( n2082 & ~n2085 ) | ( n2082 & n2086 ) | ( ~n2085 & n2086 ) ;
  assign n2088 = ( n1946 & n1987 ) | ( n1946 & n2087 ) | ( n1987 & n2087 ) ;
  assign n2089 = ( ~n1946 & n1987 ) | ( ~n1946 & n2087 ) | ( n1987 & n2087 ) ;
  assign n2090 = ( n1946 & ~n2088 ) | ( n1946 & n2089 ) | ( ~n2088 & n2089 ) ;
  assign n2091 = ( ~n1990 & n2079 ) | ( ~n1990 & n2090 ) | ( n2079 & n2090 ) ;
  assign n2092 = ( n1990 & n2079 ) | ( n1990 & n2090 ) | ( n2079 & n2090 ) ;
  assign n2093 = ( n1990 & n2091 ) | ( n1990 & ~n2092 ) | ( n2091 & ~n2092 ) ;
  assign n2094 = ( n1975 & n1977 ) | ( n1975 & n2003 ) | ( n1977 & n2003 ) ;
  assign n2095 = ( n1975 & ~n1977 ) | ( n1975 & n2003 ) | ( ~n1977 & n2003 ) ;
  assign n2096 = ( n1977 & ~n2094 ) | ( n1977 & n2095 ) | ( ~n2094 & n2095 ) ;
  assign n2097 = ( ~n1981 & n2093 ) | ( ~n1981 & n2096 ) | ( n2093 & n2096 ) ;
  assign n2098 = ( n1981 & n2093 ) | ( n1981 & n2096 ) | ( n2093 & n2096 ) ;
  assign n2099 = ( n1981 & n2097 ) | ( n1981 & ~n2098 ) | ( n2097 & ~n2098 ) ;
  assign n2100 = ( ~n2009 & n2071 ) | ( ~n2009 & n2099 ) | ( n2071 & n2099 ) ;
  assign n2101 = ( n2009 & n2071 ) | ( n2009 & n2099 ) | ( n2071 & n2099 ) ;
  assign n2102 = ( n2009 & n2100 ) | ( n2009 & ~n2101 ) | ( n2100 & ~n2101 ) ;
  assign n2103 = ( ~n1995 & n2026 ) | ( ~n1995 & n2102 ) | ( n2026 & n2102 ) ;
  assign n2104 = ( n1995 & n2026 ) | ( n1995 & n2102 ) | ( n2026 & n2102 ) ;
  assign n2105 = ( n1995 & n2103 ) | ( n1995 & ~n2104 ) | ( n2103 & ~n2104 ) ;
  assign n2106 = ( ~n2012 & n2015 ) | ( ~n2012 & n2105 ) | ( n2015 & n2105 ) ;
  assign n2107 = ( n2012 & n2015 ) | ( n2012 & n2105 ) | ( n2015 & n2105 ) ;
  assign n2108 = ( n2012 & n2106 ) | ( n2012 & ~n2107 ) | ( n2106 & ~n2107 ) ;
  assign n2109 = ~x1 & x23 ;
  assign n2110 = ( x1 & x23 ) | ( x1 & x44 ) | ( x23 & x44 ) ;
  assign n2111 = x23 & x44 ;
  assign n2112 = ( n2109 & n2110 ) | ( n2109 & ~n2111 ) | ( n2110 & ~n2111 ) ;
  assign n2113 = x3 & x42 ;
  assign n2114 = ( n2074 & n2112 ) | ( n2074 & n2113 ) | ( n2112 & n2113 ) ;
  assign n2115 = ( ~n2074 & n2112 ) | ( ~n2074 & n2113 ) | ( n2112 & n2113 ) ;
  assign n2116 = ( n2074 & ~n2114 ) | ( n2074 & n2115 ) | ( ~n2114 & n2115 ) ;
  assign n2117 = x15 & x30 ;
  assign n2118 = x16 & x29 ;
  assign n2119 = x17 & x28 ;
  assign n2120 = ( ~n2117 & n2118 ) | ( ~n2117 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2121 = ( n2117 & n2118 ) | ( n2117 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2122 = ( n2117 & n2120 ) | ( n2117 & ~n2121 ) | ( n2120 & ~n2121 ) ;
  assign n2123 = x12 & x33 ;
  assign n2124 = x11 & x34 ;
  assign n2125 = x6 & x39 ;
  assign n2126 = ( ~n2123 & n2124 ) | ( ~n2123 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2127 = ( n2123 & n2124 ) | ( n2123 & n2125 ) | ( n2124 & n2125 ) ;
  assign n2128 = ( n2123 & n2126 ) | ( n2123 & ~n2127 ) | ( n2126 & ~n2127 ) ;
  assign n2129 = ( ~n2116 & n2122 ) | ( ~n2116 & n2128 ) | ( n2122 & n2128 ) ;
  assign n2130 = ( n2116 & n2122 ) | ( n2116 & n2128 ) | ( n2122 & n2128 ) ;
  assign n2131 = ( n2116 & n2129 ) | ( n2116 & ~n2130 ) | ( n2129 & ~n2130 ) ;
  assign n2132 = ( n2031 & n2043 ) | ( n2031 & n2085 ) | ( n2043 & n2085 ) ;
  assign n2133 = ( n2031 & n2043 ) | ( n2031 & ~n2085 ) | ( n2043 & ~n2085 ) ;
  assign n2134 = ( n2085 & ~n2132 ) | ( n2085 & n2133 ) | ( ~n2132 & n2133 ) ;
  assign n2135 = ( ~n2094 & n2131 ) | ( ~n2094 & n2134 ) | ( n2131 & n2134 ) ;
  assign n2136 = ( n2094 & n2131 ) | ( n2094 & n2134 ) | ( n2131 & n2134 ) ;
  assign n2137 = ( n2094 & n2135 ) | ( n2094 & ~n2136 ) | ( n2135 & ~n2136 ) ;
  assign n2138 = ( n2069 & n2098 ) | ( n2069 & n2137 ) | ( n2098 & n2137 ) ;
  assign n2139 = ( ~n2069 & n2098 ) | ( ~n2069 & n2137 ) | ( n2098 & n2137 ) ;
  assign n2140 = ( n2069 & ~n2138 ) | ( n2069 & n2139 ) | ( ~n2138 & n2139 ) ;
  assign n2141 = x13 & x32 ;
  assign n2142 = x14 & x31 ;
  assign n2143 = x5 & x40 ;
  assign n2144 = ( ~n2141 & n2142 ) | ( ~n2141 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2145 = ( n2141 & n2142 ) | ( n2141 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2146 = ( n2141 & n2144 ) | ( n2141 & ~n2145 ) | ( n2144 & ~n2145 ) ;
  assign n2147 = x18 & x27 ;
  assign n2148 = x20 & x25 ;
  assign n2149 = x19 & x26 ;
  assign n2150 = ( ~n2147 & n2148 ) | ( ~n2147 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2151 = ( n2147 & n2148 ) | ( n2147 & n2149 ) | ( n2148 & n2149 ) ;
  assign n2152 = ( n2147 & n2150 ) | ( n2147 & ~n2151 ) | ( n2150 & ~n2151 ) ;
  assign n2153 = ( n2064 & n2146 ) | ( n2064 & n2152 ) | ( n2146 & n2152 ) ;
  assign n2154 = ( ~n2064 & n2146 ) | ( ~n2064 & n2152 ) | ( n2146 & n2152 ) ;
  assign n2155 = ( n2064 & ~n2153 ) | ( n2064 & n2154 ) | ( ~n2153 & n2154 ) ;
  assign n2156 = x0 & x45 ;
  assign n2157 = x2 & x43 ;
  assign n2158 = x4 & x41 ;
  assign n2159 = ( ~n2156 & n2157 ) | ( ~n2156 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2160 = ( n2156 & n2157 ) | ( n2156 & n2158 ) | ( n2157 & n2158 ) ;
  assign n2161 = ( n2156 & n2159 ) | ( n2156 & ~n2160 ) | ( n2159 & ~n2160 ) ;
  assign n2162 = x10 & x35 ;
  assign n2163 = x22 & x23 ;
  assign n2164 = x21 & x24 ;
  assign n2165 = ( ~n2162 & n2163 ) | ( ~n2162 & n2164 ) | ( n2163 & n2164 ) ;
  assign n2166 = ( n2162 & n2163 ) | ( n2162 & n2164 ) | ( n2163 & n2164 ) ;
  assign n2167 = ( n2162 & n2165 ) | ( n2162 & ~n2166 ) | ( n2165 & ~n2166 ) ;
  assign n2168 = x7 & x38 ;
  assign n2169 = x8 & x37 ;
  assign n2170 = x9 & x36 ;
  assign n2171 = ( ~n2168 & n2169 ) | ( ~n2168 & n2170 ) | ( n2169 & n2170 ) ;
  assign n2172 = ( n2168 & n2169 ) | ( n2168 & n2170 ) | ( n2169 & n2170 ) ;
  assign n2173 = ( n2168 & n2171 ) | ( n2168 & ~n2172 ) | ( n2171 & ~n2172 ) ;
  assign n2174 = ( ~n2161 & n2167 ) | ( ~n2161 & n2173 ) | ( n2167 & n2173 ) ;
  assign n2175 = ( n2161 & n2167 ) | ( n2161 & n2173 ) | ( n2167 & n2173 ) ;
  assign n2176 = ( n2161 & n2174 ) | ( n2161 & ~n2175 ) | ( n2174 & ~n2175 ) ;
  assign n2177 = ( ~n2021 & n2155 ) | ( ~n2021 & n2176 ) | ( n2155 & n2176 ) ;
  assign n2178 = ( n2021 & n2155 ) | ( n2021 & n2176 ) | ( n2155 & n2176 ) ;
  assign n2179 = ( n2021 & n2177 ) | ( n2021 & ~n2178 ) | ( n2177 & ~n2178 ) ;
  assign n2180 = ( n2019 & n2078 ) | ( n2019 & n2088 ) | ( n2078 & n2088 ) ;
  assign n2181 = ( n2019 & n2078 ) | ( n2019 & ~n2088 ) | ( n2078 & ~n2088 ) ;
  assign n2182 = ( n2088 & ~n2180 ) | ( n2088 & n2181 ) | ( ~n2180 & n2181 ) ;
  assign n2183 = ( n2037 & ~n2052 ) | ( n2037 & n2058 ) | ( ~n2052 & n2058 ) ;
  assign n2184 = ( n2037 & n2052 ) | ( n2037 & n2058 ) | ( n2052 & n2058 ) ;
  assign n2185 = ( n2052 & n2183 ) | ( n2052 & ~n2184 ) | ( n2183 & ~n2184 ) ;
  assign n2186 = ( n2046 & n2067 ) | ( n2046 & n2185 ) | ( n2067 & n2185 ) ;
  assign n2187 = ( ~n2046 & n2067 ) | ( ~n2046 & n2185 ) | ( n2067 & n2185 ) ;
  assign n2188 = ( n2046 & ~n2186 ) | ( n2046 & n2187 ) | ( ~n2186 & n2187 ) ;
  assign n2189 = ( ~n2092 & n2182 ) | ( ~n2092 & n2188 ) | ( n2182 & n2188 ) ;
  assign n2190 = ( n2092 & n2182 ) | ( n2092 & n2188 ) | ( n2182 & n2188 ) ;
  assign n2191 = ( n2092 & n2189 ) | ( n2092 & ~n2190 ) | ( n2189 & ~n2190 ) ;
  assign n2192 = ( ~n2024 & n2179 ) | ( ~n2024 & n2191 ) | ( n2179 & n2191 ) ;
  assign n2193 = ( n2024 & n2179 ) | ( n2024 & n2191 ) | ( n2179 & n2191 ) ;
  assign n2194 = ( n2024 & n2192 ) | ( n2024 & ~n2193 ) | ( n2192 & ~n2193 ) ;
  assign n2195 = ( ~n2101 & n2140 ) | ( ~n2101 & n2194 ) | ( n2140 & n2194 ) ;
  assign n2196 = ( n2101 & n2140 ) | ( n2101 & n2194 ) | ( n2140 & n2194 ) ;
  assign n2197 = ( n2101 & n2195 ) | ( n2101 & ~n2196 ) | ( n2195 & ~n2196 ) ;
  assign n2198 = ( n2104 & n2107 ) | ( n2104 & n2197 ) | ( n2107 & n2197 ) ;
  assign n2199 = ( ~n2104 & n2107 ) | ( ~n2104 & n2197 ) | ( n2107 & n2197 ) ;
  assign n2200 = ( n2104 & ~n2198 ) | ( n2104 & n2199 ) | ( ~n2198 & n2199 ) ;
  assign n2201 = x14 & x32 ;
  assign n2202 = x6 & x40 ;
  assign n2203 = x13 & x33 ;
  assign n2204 = ( ~n2201 & n2202 ) | ( ~n2201 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2205 = ( n2201 & n2202 ) | ( n2201 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2206 = ( n2201 & n2204 ) | ( n2201 & ~n2205 ) | ( n2204 & ~n2205 ) ;
  assign n2207 = x15 & x31 ;
  assign n2208 = x5 & x41 ;
  assign n2209 = ( ~n2083 & n2207 ) | ( ~n2083 & n2208 ) | ( n2207 & n2208 ) ;
  assign n2210 = ( n2083 & n2207 ) | ( n2083 & n2208 ) | ( n2207 & n2208 ) ;
  assign n2211 = ( n2083 & n2209 ) | ( n2083 & ~n2210 ) | ( n2209 & ~n2210 ) ;
  assign n2212 = ( n2184 & n2206 ) | ( n2184 & n2211 ) | ( n2206 & n2211 ) ;
  assign n2213 = ( ~n2184 & n2206 ) | ( ~n2184 & n2211 ) | ( n2206 & n2211 ) ;
  assign n2214 = ( n2184 & ~n2212 ) | ( n2184 & n2213 ) | ( ~n2212 & n2213 ) ;
  assign n2215 = ( n2121 & ~n2127 ) | ( n2121 & n2151 ) | ( ~n2127 & n2151 ) ;
  assign n2216 = ( n2121 & n2127 ) | ( n2121 & n2151 ) | ( n2127 & n2151 ) ;
  assign n2217 = ( n2127 & n2215 ) | ( n2127 & ~n2216 ) | ( n2215 & ~n2216 ) ;
  assign n2218 = ( n2180 & n2214 ) | ( n2180 & n2217 ) | ( n2214 & n2217 ) ;
  assign n2219 = ( ~n2180 & n2214 ) | ( ~n2180 & n2217 ) | ( n2214 & n2217 ) ;
  assign n2220 = ( n2180 & ~n2218 ) | ( n2180 & n2219 ) | ( ~n2218 & n2219 ) ;
  assign n2221 = ( ~n2178 & n2190 ) | ( ~n2178 & n2220 ) | ( n2190 & n2220 ) ;
  assign n2222 = ( n2178 & n2190 ) | ( n2178 & n2220 ) | ( n2190 & n2220 ) ;
  assign n2223 = ( n2178 & n2221 ) | ( n2178 & ~n2222 ) | ( n2221 & ~n2222 ) ;
  assign n2224 = ( n2193 & n2196 ) | ( n2193 & n2223 ) | ( n2196 & n2223 ) ;
  assign n2225 = ( ~n2193 & n2196 ) | ( ~n2193 & n2223 ) | ( n2196 & n2223 ) ;
  assign n2226 = ( n2193 & ~n2224 ) | ( n2193 & n2225 ) | ( ~n2224 & n2225 ) ;
  assign n2227 = x12 & x34 ;
  assign n2228 = x7 & x39 ;
  assign n2229 = x8 & x38 ;
  assign n2230 = ( ~n2227 & n2228 ) | ( ~n2227 & n2229 ) | ( n2228 & n2229 ) ;
  assign n2231 = ( n2227 & n2228 ) | ( n2227 & n2229 ) | ( n2228 & n2229 ) ;
  assign n2232 = ( n2227 & n2230 ) | ( n2227 & ~n2231 ) | ( n2230 & ~n2231 ) ;
  assign n2233 = x16 & x30 ;
  assign n2234 = x17 & x29 ;
  assign n2235 = x18 & x28 ;
  assign n2236 = ( ~n2233 & n2234 ) | ( ~n2233 & n2235 ) | ( n2234 & n2235 ) ;
  assign n2237 = ( n2233 & n2234 ) | ( n2233 & n2235 ) | ( n2234 & n2235 ) ;
  assign n2238 = ( n2233 & n2236 ) | ( n2233 & ~n2237 ) | ( n2236 & ~n2237 ) ;
  assign n2239 = ( n2114 & n2232 ) | ( n2114 & n2238 ) | ( n2232 & n2238 ) ;
  assign n2240 = ( ~n2114 & n2232 ) | ( ~n2114 & n2238 ) | ( n2232 & n2238 ) ;
  assign n2241 = ( n2114 & ~n2239 ) | ( n2114 & n2240 ) | ( ~n2239 & n2240 ) ;
  assign n2242 = x3 & x43 ;
  assign n2243 = x0 & x46 ;
  assign n2244 = x4 & x42 ;
  assign n2245 = ( ~n2242 & n2243 ) | ( ~n2242 & n2244 ) | ( n2243 & n2244 ) ;
  assign n2246 = ( n2242 & n2243 ) | ( n2242 & n2244 ) | ( n2243 & n2244 ) ;
  assign n2247 = ( n2242 & n2245 ) | ( n2242 & ~n2246 ) | ( n2245 & ~n2246 ) ;
  assign n2248 = x19 & x27 ;
  assign n2249 = x20 & x26 ;
  assign n2250 = x21 & x25 ;
  assign n2251 = ( ~n2248 & n2249 ) | ( ~n2248 & n2250 ) | ( n2249 & n2250 ) ;
  assign n2252 = ( n2248 & n2249 ) | ( n2248 & n2250 ) | ( n2249 & n2250 ) ;
  assign n2253 = ( n2248 & n2251 ) | ( n2248 & ~n2252 ) | ( n2251 & ~n2252 ) ;
  assign n2254 = x9 & x37 ;
  assign n2255 = x11 & x35 ;
  assign n2256 = x10 & x36 ;
  assign n2257 = ( ~n2254 & n2255 ) | ( ~n2254 & n2256 ) | ( n2255 & n2256 ) ;
  assign n2258 = ( n2254 & n2255 ) | ( n2254 & n2256 ) | ( n2255 & n2256 ) ;
  assign n2259 = ( n2254 & n2257 ) | ( n2254 & ~n2258 ) | ( n2257 & ~n2258 ) ;
  assign n2260 = ( ~n2247 & n2253 ) | ( ~n2247 & n2259 ) | ( n2253 & n2259 ) ;
  assign n2261 = ( n2247 & n2253 ) | ( n2247 & n2259 ) | ( n2253 & n2259 ) ;
  assign n2262 = ( n2247 & n2260 ) | ( n2247 & ~n2261 ) | ( n2260 & ~n2261 ) ;
  assign n2263 = ( ~n2186 & n2241 ) | ( ~n2186 & n2262 ) | ( n2241 & n2262 ) ;
  assign n2264 = ( n2186 & n2241 ) | ( n2186 & n2262 ) | ( n2241 & n2262 ) ;
  assign n2265 = ( n2186 & n2263 ) | ( n2186 & ~n2264 ) | ( n2263 & ~n2264 ) ;
  assign n2266 = ( n2130 & n2153 ) | ( n2130 & n2175 ) | ( n2153 & n2175 ) ;
  assign n2267 = ( ~n2130 & n2153 ) | ( ~n2130 & n2175 ) | ( n2153 & n2175 ) ;
  assign n2268 = ( n2130 & ~n2266 ) | ( n2130 & n2267 ) | ( ~n2266 & n2267 ) ;
  assign n2269 = ( n2145 & n2160 ) | ( n2145 & n2172 ) | ( n2160 & n2172 ) ;
  assign n2270 = ( n2145 & n2160 ) | ( n2145 & ~n2172 ) | ( n2160 & ~n2172 ) ;
  assign n2271 = ( n2172 & ~n2269 ) | ( n2172 & n2270 ) | ( ~n2269 & n2270 ) ;
  assign n2272 = x44 & n651 ;
  assign n2273 = x22 & x24 ;
  assign n2274 = x1 & x45 ;
  assign n2275 = n2273 & n2274 ;
  assign n2276 = n2273 | n2274 ;
  assign n2277 = ~n2275 & n2276 ;
  assign n2278 = ( n2166 & n2272 ) | ( n2166 & n2277 ) | ( n2272 & n2277 ) ;
  assign n2279 = ( n2166 & ~n2272 ) | ( n2166 & n2277 ) | ( ~n2272 & n2277 ) ;
  assign n2280 = ( n2272 & ~n2278 ) | ( n2272 & n2279 ) | ( ~n2278 & n2279 ) ;
  assign n2281 = ( ~n2132 & n2271 ) | ( ~n2132 & n2280 ) | ( n2271 & n2280 ) ;
  assign n2282 = ( n2132 & n2271 ) | ( n2132 & n2280 ) | ( n2271 & n2280 ) ;
  assign n2283 = ( n2132 & n2281 ) | ( n2132 & ~n2282 ) | ( n2281 & ~n2282 ) ;
  assign n2284 = ( ~n2136 & n2268 ) | ( ~n2136 & n2283 ) | ( n2268 & n2283 ) ;
  assign n2285 = ( n2136 & n2268 ) | ( n2136 & n2283 ) | ( n2268 & n2283 ) ;
  assign n2286 = ( n2136 & n2284 ) | ( n2136 & ~n2285 ) | ( n2284 & ~n2285 ) ;
  assign n2287 = ( n2138 & n2265 ) | ( n2138 & n2286 ) | ( n2265 & n2286 ) ;
  assign n2288 = ( ~n2138 & n2265 ) | ( ~n2138 & n2286 ) | ( n2265 & n2286 ) ;
  assign n2289 = ( n2138 & ~n2287 ) | ( n2138 & n2288 ) | ( ~n2287 & n2288 ) ;
  assign n2290 = ( ~n2198 & n2226 ) | ( ~n2198 & n2289 ) | ( n2226 & n2289 ) ;
  assign n2291 = ( n2198 & n2226 ) | ( n2198 & n2289 ) | ( n2226 & n2289 ) ;
  assign n2292 = ( n2198 & n2290 ) | ( n2198 & ~n2291 ) | ( n2290 & ~n2291 ) ;
  assign n2293 = ( n2210 & n2246 ) | ( n2210 & ~n2252 ) | ( n2246 & ~n2252 ) ;
  assign n2294 = ( n2210 & n2246 ) | ( n2210 & n2252 ) | ( n2246 & n2252 ) ;
  assign n2295 = ( n2252 & n2293 ) | ( n2252 & ~n2294 ) | ( n2293 & ~n2294 ) ;
  assign n2296 = ( ~n2212 & n2261 ) | ( ~n2212 & n2295 ) | ( n2261 & n2295 ) ;
  assign n2297 = ( n2212 & n2261 ) | ( n2212 & n2295 ) | ( n2261 & n2295 ) ;
  assign n2298 = ( n2212 & n2296 ) | ( n2212 & ~n2297 ) | ( n2296 & ~n2297 ) ;
  assign n2299 = ( n2218 & n2264 ) | ( n2218 & n2298 ) | ( n2264 & n2298 ) ;
  assign n2300 = ( n2218 & n2264 ) | ( n2218 & ~n2298 ) | ( n2264 & ~n2298 ) ;
  assign n2301 = ( n2298 & ~n2299 ) | ( n2298 & n2300 ) | ( ~n2299 & n2300 ) ;
  assign n2302 = ( ~n2222 & n2285 ) | ( ~n2222 & n2301 ) | ( n2285 & n2301 ) ;
  assign n2303 = ( n2222 & n2285 ) | ( n2222 & n2301 ) | ( n2285 & n2301 ) ;
  assign n2304 = ( n2222 & n2302 ) | ( n2222 & ~n2303 ) | ( n2302 & ~n2303 ) ;
  assign n2305 = x13 & x34 ;
  assign n2306 = x12 & x35 ;
  assign n2307 = x7 & x40 ;
  assign n2308 = ( ~n2305 & n2306 ) | ( ~n2305 & n2307 ) | ( n2306 & n2307 ) ;
  assign n2309 = ( n2305 & n2306 ) | ( n2305 & n2307 ) | ( n2306 & n2307 ) ;
  assign n2310 = ( n2305 & n2308 ) | ( n2305 & ~n2309 ) | ( n2308 & ~n2309 ) ;
  assign n2311 = ( ~n2216 & n2278 ) | ( ~n2216 & n2310 ) | ( n2278 & n2310 ) ;
  assign n2312 = ( n2216 & n2278 ) | ( n2216 & n2310 ) | ( n2278 & n2310 ) ;
  assign n2313 = ( n2216 & n2311 ) | ( n2216 & ~n2312 ) | ( n2311 & ~n2312 ) ;
  assign n2314 = ( ~n2266 & n2282 ) | ( ~n2266 & n2313 ) | ( n2282 & n2313 ) ;
  assign n2315 = ( n2266 & n2282 ) | ( n2266 & n2313 ) | ( n2282 & n2313 ) ;
  assign n2316 = ( n2266 & n2314 ) | ( n2266 & ~n2315 ) | ( n2314 & ~n2315 ) ;
  assign n2317 = x3 & x44 ;
  assign n2318 = x4 & x43 ;
  assign n2319 = x15 & x32 ;
  assign n2320 = ( ~n2317 & n2318 ) | ( ~n2317 & n2319 ) | ( n2318 & n2319 ) ;
  assign n2321 = ( n2317 & n2318 ) | ( n2317 & n2319 ) | ( n2318 & n2319 ) ;
  assign n2322 = ( n2317 & n2320 ) | ( n2317 & ~n2321 ) | ( n2320 & ~n2321 ) ;
  assign n2323 = ( ~n2205 & n2237 ) | ( ~n2205 & n2322 ) | ( n2237 & n2322 ) ;
  assign n2324 = ( n2205 & n2237 ) | ( n2205 & n2322 ) | ( n2237 & n2322 ) ;
  assign n2325 = ( n2205 & n2323 ) | ( n2205 & ~n2324 ) | ( n2323 & ~n2324 ) ;
  assign n2326 = x5 & x42 ;
  assign n2327 = x6 & x41 ;
  assign n2328 = x14 & x33 ;
  assign n2329 = ( ~n2326 & n2327 ) | ( ~n2326 & n2328 ) | ( n2327 & n2328 ) ;
  assign n2330 = ( n2326 & n2327 ) | ( n2326 & n2328 ) | ( n2327 & n2328 ) ;
  assign n2331 = ( n2326 & n2329 ) | ( n2326 & ~n2330 ) | ( n2329 & ~n2330 ) ;
  assign n2332 = x10 & x37 ;
  assign n2333 = x23 & x24 ;
  assign n2334 = x22 & x25 ;
  assign n2335 = ( ~n2332 & n2333 ) | ( ~n2332 & n2334 ) | ( n2333 & n2334 ) ;
  assign n2336 = ( n2332 & n2333 ) | ( n2332 & n2334 ) | ( n2333 & n2334 ) ;
  assign n2337 = ( n2332 & n2335 ) | ( n2332 & ~n2336 ) | ( n2335 & ~n2336 ) ;
  assign n2338 = x8 & x39 ;
  assign n2339 = x11 & x36 ;
  assign n2340 = x9 & x38 ;
  assign n2341 = ( ~n2338 & n2339 ) | ( ~n2338 & n2340 ) | ( n2339 & n2340 ) ;
  assign n2342 = ( n2338 & n2339 ) | ( n2338 & n2340 ) | ( n2339 & n2340 ) ;
  assign n2343 = ( n2338 & n2341 ) | ( n2338 & ~n2342 ) | ( n2341 & ~n2342 ) ;
  assign n2344 = ( ~n2331 & n2337 ) | ( ~n2331 & n2343 ) | ( n2337 & n2343 ) ;
  assign n2345 = ( n2331 & n2337 ) | ( n2331 & n2343 ) | ( n2337 & n2343 ) ;
  assign n2346 = ( n2331 & n2344 ) | ( n2331 & ~n2345 ) | ( n2344 & ~n2345 ) ;
  assign n2347 = x0 & x47 ;
  assign n2348 = x2 & x45 ;
  assign n2349 = ( ~n2275 & n2347 ) | ( ~n2275 & n2348 ) | ( n2347 & n2348 ) ;
  assign n2350 = ( n2275 & n2347 ) | ( n2275 & n2348 ) | ( n2347 & n2348 ) ;
  assign n2351 = ( n2275 & n2349 ) | ( n2275 & ~n2350 ) | ( n2349 & ~n2350 ) ;
  assign n2352 = x16 & x31 ;
  assign n2353 = x18 & x29 ;
  assign n2354 = x17 & x30 ;
  assign n2355 = ( ~n2352 & n2353 ) | ( ~n2352 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2356 = ( n2352 & n2353 ) | ( n2352 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2357 = ( n2352 & n2355 ) | ( n2352 & ~n2356 ) | ( n2355 & ~n2356 ) ;
  assign n2358 = x19 & x28 ;
  assign n2359 = x21 & x26 ;
  assign n2360 = x20 & x27 ;
  assign n2361 = ( ~n2358 & n2359 ) | ( ~n2358 & n2360 ) | ( n2359 & n2360 ) ;
  assign n2362 = ( n2358 & n2359 ) | ( n2358 & n2360 ) | ( n2359 & n2360 ) ;
  assign n2363 = ( n2358 & n2361 ) | ( n2358 & ~n2362 ) | ( n2361 & ~n2362 ) ;
  assign n2364 = ( ~n2351 & n2357 ) | ( ~n2351 & n2363 ) | ( n2357 & n2363 ) ;
  assign n2365 = ( n2351 & n2357 ) | ( n2351 & n2363 ) | ( n2357 & n2363 ) ;
  assign n2366 = ( n2351 & n2364 ) | ( n2351 & ~n2365 ) | ( n2364 & ~n2365 ) ;
  assign n2367 = ( n2325 & n2346 ) | ( n2325 & n2366 ) | ( n2346 & n2366 ) ;
  assign n2368 = ( ~n2325 & n2346 ) | ( ~n2325 & n2366 ) | ( n2346 & n2366 ) ;
  assign n2369 = ( n2325 & ~n2367 ) | ( n2325 & n2368 ) | ( ~n2367 & n2368 ) ;
  assign n2370 = x24 & x46 ;
  assign n2371 = ( x1 & x24 ) | ( x1 & x46 ) | ( x24 & x46 ) ;
  assign n2372 = ~x1 & x24 ;
  assign n2373 = ( ~n2370 & n2371 ) | ( ~n2370 & n2372 ) | ( n2371 & n2372 ) ;
  assign n2374 = ( ~n2231 & n2258 ) | ( ~n2231 & n2373 ) | ( n2258 & n2373 ) ;
  assign n2375 = ( n2231 & n2258 ) | ( n2231 & n2373 ) | ( n2258 & n2373 ) ;
  assign n2376 = ( n2231 & n2374 ) | ( n2231 & ~n2375 ) | ( n2374 & ~n2375 ) ;
  assign n2377 = ( ~n2239 & n2269 ) | ( ~n2239 & n2376 ) | ( n2269 & n2376 ) ;
  assign n2378 = ( n2239 & n2269 ) | ( n2239 & n2376 ) | ( n2269 & n2376 ) ;
  assign n2379 = ( n2239 & n2377 ) | ( n2239 & ~n2378 ) | ( n2377 & ~n2378 ) ;
  assign n2380 = ( ~n2316 & n2369 ) | ( ~n2316 & n2379 ) | ( n2369 & n2379 ) ;
  assign n2381 = ( n2316 & n2369 ) | ( n2316 & n2379 ) | ( n2369 & n2379 ) ;
  assign n2382 = ( n2316 & n2380 ) | ( n2316 & ~n2381 ) | ( n2380 & ~n2381 ) ;
  assign n2383 = ( n2287 & n2304 ) | ( n2287 & n2382 ) | ( n2304 & n2382 ) ;
  assign n2384 = ( ~n2287 & n2304 ) | ( ~n2287 & n2382 ) | ( n2304 & n2382 ) ;
  assign n2385 = ( n2287 & ~n2383 ) | ( n2287 & n2384 ) | ( ~n2383 & n2384 ) ;
  assign n2386 = ( n2224 & n2291 ) | ( n2224 & n2385 ) | ( n2291 & n2385 ) ;
  assign n2387 = ( ~n2224 & n2291 ) | ( ~n2224 & n2385 ) | ( n2291 & n2385 ) ;
  assign n2388 = ( n2224 & ~n2386 ) | ( n2224 & n2387 ) | ( ~n2386 & n2387 ) ;
  assign n2389 = x9 & x39 ;
  assign n2390 = x11 & x37 ;
  assign n2391 = x10 & x38 ;
  assign n2392 = ( ~n2389 & n2390 ) | ( ~n2389 & n2391 ) | ( n2390 & n2391 ) ;
  assign n2393 = ( n2389 & n2390 ) | ( n2389 & n2391 ) | ( n2390 & n2391 ) ;
  assign n2394 = ( n2389 & n2392 ) | ( n2389 & ~n2393 ) | ( n2392 & ~n2393 ) ;
  assign n2395 = x14 & x34 ;
  assign n2396 = x6 & x42 ;
  assign n2397 = x13 & x35 ;
  assign n2398 = ( ~n2395 & n2396 ) | ( ~n2395 & n2397 ) | ( n2396 & n2397 ) ;
  assign n2399 = ( n2395 & n2396 ) | ( n2395 & n2397 ) | ( n2396 & n2397 ) ;
  assign n2400 = ( n2395 & n2398 ) | ( n2395 & ~n2399 ) | ( n2398 & ~n2399 ) ;
  assign n2401 = x7 & x41 ;
  assign n2402 = x12 & x36 ;
  assign n2403 = x8 & x40 ;
  assign n2404 = ( ~n2401 & n2402 ) | ( ~n2401 & n2403 ) | ( n2402 & n2403 ) ;
  assign n2405 = ( n2401 & n2402 ) | ( n2401 & n2403 ) | ( n2402 & n2403 ) ;
  assign n2406 = ( n2401 & n2404 ) | ( n2401 & ~n2405 ) | ( n2404 & ~n2405 ) ;
  assign n2407 = ( ~n2394 & n2400 ) | ( ~n2394 & n2406 ) | ( n2400 & n2406 ) ;
  assign n2408 = ( n2394 & n2400 ) | ( n2394 & n2406 ) | ( n2400 & n2406 ) ;
  assign n2409 = ( n2394 & n2407 ) | ( n2394 & ~n2408 ) | ( n2407 & ~n2408 ) ;
  assign n2410 = x17 & x31 ;
  assign n2411 = x18 & x30 ;
  assign n2412 = x19 & x29 ;
  assign n2413 = ( ~n2410 & n2411 ) | ( ~n2410 & n2412 ) | ( n2411 & n2412 ) ;
  assign n2414 = ( n2410 & n2411 ) | ( n2410 & n2412 ) | ( n2411 & n2412 ) ;
  assign n2415 = ( n2410 & n2413 ) | ( n2410 & ~n2414 ) | ( n2413 & ~n2414 ) ;
  assign n2416 = x20 & x28 ;
  assign n2417 = x21 & x27 ;
  assign n2418 = x22 & x26 ;
  assign n2419 = ( ~n2416 & n2417 ) | ( ~n2416 & n2418 ) | ( n2417 & n2418 ) ;
  assign n2420 = ( n2416 & n2417 ) | ( n2416 & n2418 ) | ( n2417 & n2418 ) ;
  assign n2421 = ( n2416 & n2419 ) | ( n2416 & ~n2420 ) | ( n2419 & ~n2420 ) ;
  assign n2422 = x4 & x44 ;
  assign n2423 = x5 & x43 ;
  assign n2424 = x15 & x33 ;
  assign n2425 = ( ~n2422 & n2423 ) | ( ~n2422 & n2424 ) | ( n2423 & n2424 ) ;
  assign n2426 = ( n2422 & n2423 ) | ( n2422 & n2424 ) | ( n2423 & n2424 ) ;
  assign n2427 = ( n2422 & n2425 ) | ( n2422 & ~n2426 ) | ( n2425 & ~n2426 ) ;
  assign n2428 = ( ~n2415 & n2421 ) | ( ~n2415 & n2427 ) | ( n2421 & n2427 ) ;
  assign n2429 = ( n2415 & n2421 ) | ( n2415 & n2427 ) | ( n2421 & n2427 ) ;
  assign n2430 = ( n2415 & n2428 ) | ( n2415 & ~n2429 ) | ( n2428 & ~n2429 ) ;
  assign n2431 = ( n2312 & n2409 ) | ( n2312 & n2430 ) | ( n2409 & n2430 ) ;
  assign n2432 = ( ~n2312 & n2409 ) | ( ~n2312 & n2430 ) | ( n2409 & n2430 ) ;
  assign n2433 = ( n2312 & ~n2431 ) | ( n2312 & n2432 ) | ( ~n2431 & n2432 ) ;
  assign n2434 = ( ~n2299 & n2315 ) | ( ~n2299 & n2433 ) | ( n2315 & n2433 ) ;
  assign n2435 = ( n2299 & n2315 ) | ( n2299 & n2433 ) | ( n2315 & n2433 ) ;
  assign n2436 = ( n2299 & n2434 ) | ( n2299 & ~n2435 ) | ( n2434 & ~n2435 ) ;
  assign n2437 = ( ~n2330 & n2342 ) | ( ~n2330 & n2362 ) | ( n2342 & n2362 ) ;
  assign n2438 = ( n2330 & n2342 ) | ( n2330 & n2362 ) | ( n2342 & n2362 ) ;
  assign n2439 = ( n2330 & n2437 ) | ( n2330 & ~n2438 ) | ( n2437 & ~n2438 ) ;
  assign n2440 = x2 & x46 ;
  assign n2441 = x3 & x45 ;
  assign n2442 = x16 & x32 ;
  assign n2443 = ( ~n2440 & n2441 ) | ( ~n2440 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2444 = ( n2440 & n2441 ) | ( n2440 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2445 = ( n2440 & n2443 ) | ( n2440 & ~n2444 ) | ( n2443 & ~n2444 ) ;
  assign n2446 = ( ~n2309 & n2336 ) | ( ~n2309 & n2445 ) | ( n2336 & n2445 ) ;
  assign n2447 = ( n2309 & n2336 ) | ( n2309 & n2445 ) | ( n2336 & n2445 ) ;
  assign n2448 = ( n2309 & n2446 ) | ( n2309 & ~n2447 ) | ( n2446 & ~n2447 ) ;
  assign n2449 = ( ~n2345 & n2439 ) | ( ~n2345 & n2448 ) | ( n2439 & n2448 ) ;
  assign n2450 = ( n2345 & n2439 ) | ( n2345 & n2448 ) | ( n2439 & n2448 ) ;
  assign n2451 = ( n2345 & n2449 ) | ( n2345 & ~n2450 ) | ( n2449 & ~n2450 ) ;
  assign n2452 = ( n2321 & ~n2350 ) | ( n2321 & n2356 ) | ( ~n2350 & n2356 ) ;
  assign n2453 = ( n2321 & n2350 ) | ( n2321 & n2356 ) | ( n2350 & n2356 ) ;
  assign n2454 = ( n2350 & n2452 ) | ( n2350 & ~n2453 ) | ( n2452 & ~n2453 ) ;
  assign n2455 = ( n2365 & n2375 ) | ( n2365 & n2454 ) | ( n2375 & n2454 ) ;
  assign n2456 = ( ~n2365 & n2375 ) | ( ~n2365 & n2454 ) | ( n2375 & n2454 ) ;
  assign n2457 = ( n2365 & ~n2455 ) | ( n2365 & n2456 ) | ( ~n2455 & n2456 ) ;
  assign n2458 = ( ~n2367 & n2451 ) | ( ~n2367 & n2457 ) | ( n2451 & n2457 ) ;
  assign n2459 = ( n2367 & n2451 ) | ( n2367 & n2457 ) | ( n2451 & n2457 ) ;
  assign n2460 = ( n2367 & n2458 ) | ( n2367 & ~n2459 ) | ( n2458 & ~n2459 ) ;
  assign n2461 = x1 & n2370 ;
  assign n2462 = x23 & x25 ;
  assign n2463 = x1 & x47 ;
  assign n2464 = n2462 & n2463 ;
  assign n2465 = n2462 | n2463 ;
  assign n2466 = ~n2464 & n2465 ;
  assign n2467 = x0 & x48 ;
  assign n2468 = ( n2461 & n2466 ) | ( n2461 & n2467 ) | ( n2466 & n2467 ) ;
  assign n2469 = ( ~n2461 & n2466 ) | ( ~n2461 & n2467 ) | ( n2466 & n2467 ) ;
  assign n2470 = ( n2461 & ~n2468 ) | ( n2461 & n2469 ) | ( ~n2468 & n2469 ) ;
  assign n2471 = ( ~n2294 & n2324 ) | ( ~n2294 & n2470 ) | ( n2324 & n2470 ) ;
  assign n2472 = ( n2294 & n2324 ) | ( n2294 & n2470 ) | ( n2324 & n2470 ) ;
  assign n2473 = ( n2294 & n2471 ) | ( n2294 & ~n2472 ) | ( n2471 & ~n2472 ) ;
  assign n2474 = ( ~n2297 & n2378 ) | ( ~n2297 & n2473 ) | ( n2378 & n2473 ) ;
  assign n2475 = ( n2297 & n2378 ) | ( n2297 & n2473 ) | ( n2378 & n2473 ) ;
  assign n2476 = ( n2297 & n2474 ) | ( n2297 & ~n2475 ) | ( n2474 & ~n2475 ) ;
  assign n2477 = ( ~n2381 & n2460 ) | ( ~n2381 & n2476 ) | ( n2460 & n2476 ) ;
  assign n2478 = ( n2381 & n2460 ) | ( n2381 & n2476 ) | ( n2460 & n2476 ) ;
  assign n2479 = ( n2381 & n2477 ) | ( n2381 & ~n2478 ) | ( n2477 & ~n2478 ) ;
  assign n2480 = ( n2303 & n2436 ) | ( n2303 & n2479 ) | ( n2436 & n2479 ) ;
  assign n2481 = ( ~n2303 & n2436 ) | ( ~n2303 & n2479 ) | ( n2436 & n2479 ) ;
  assign n2482 = ( n2303 & ~n2480 ) | ( n2303 & n2481 ) | ( ~n2480 & n2481 ) ;
  assign n2483 = ( ~n2383 & n2386 ) | ( ~n2383 & n2482 ) | ( n2386 & n2482 ) ;
  assign n2484 = ( n2383 & n2386 ) | ( n2383 & n2482 ) | ( n2386 & n2482 ) ;
  assign n2485 = ( n2383 & n2483 ) | ( n2383 & ~n2484 ) | ( n2483 & ~n2484 ) ;
  assign n2486 = x16 & x33 ;
  assign n2487 = x17 & x32 ;
  assign n2488 = x18 & x31 ;
  assign n2489 = ( ~n2486 & n2487 ) | ( ~n2486 & n2488 ) | ( n2487 & n2488 ) ;
  assign n2490 = ( n2486 & n2487 ) | ( n2486 & n2488 ) | ( n2487 & n2488 ) ;
  assign n2491 = ( n2486 & n2489 ) | ( n2486 & ~n2490 ) | ( n2489 & ~n2490 ) ;
  assign n2492 = x0 & x49 ;
  assign n2493 = x4 & x45 ;
  assign n2494 = x5 & x44 ;
  assign n2495 = ( ~n2492 & n2493 ) | ( ~n2492 & n2494 ) | ( n2493 & n2494 ) ;
  assign n2496 = ( n2492 & n2493 ) | ( n2492 & n2494 ) | ( n2493 & n2494 ) ;
  assign n2497 = ( n2492 & n2495 ) | ( n2492 & ~n2496 ) | ( n2495 & ~n2496 ) ;
  assign n2498 = ( n2468 & n2491 ) | ( n2468 & n2497 ) | ( n2491 & n2497 ) ;
  assign n2499 = ( ~n2468 & n2491 ) | ( ~n2468 & n2497 ) | ( n2491 & n2497 ) ;
  assign n2500 = ( n2468 & ~n2498 ) | ( n2468 & n2499 ) | ( ~n2498 & n2499 ) ;
  assign n2501 = x15 & x34 ;
  assign n2502 = x6 & x43 ;
  assign n2503 = x14 & x35 ;
  assign n2504 = ( ~n2501 & n2502 ) | ( ~n2501 & n2503 ) | ( n2502 & n2503 ) ;
  assign n2505 = ( n2501 & n2502 ) | ( n2501 & n2503 ) | ( n2502 & n2503 ) ;
  assign n2506 = ( n2501 & n2504 ) | ( n2501 & ~n2505 ) | ( n2504 & ~n2505 ) ;
  assign n2507 = x11 & x38 ;
  assign n2508 = x24 & x25 ;
  assign n2509 = x23 & x26 ;
  assign n2510 = ( ~n2507 & n2508 ) | ( ~n2507 & n2509 ) | ( n2508 & n2509 ) ;
  assign n2511 = ( n2507 & n2508 ) | ( n2507 & n2509 ) | ( n2508 & n2509 ) ;
  assign n2512 = ( n2507 & n2510 ) | ( n2507 & ~n2511 ) | ( n2510 & ~n2511 ) ;
  assign n2513 = x13 & x36 ;
  assign n2514 = x7 & x42 ;
  assign n2515 = x8 & x41 ;
  assign n2516 = ( ~n2513 & n2514 ) | ( ~n2513 & n2515 ) | ( n2514 & n2515 ) ;
  assign n2517 = ( n2513 & n2514 ) | ( n2513 & n2515 ) | ( n2514 & n2515 ) ;
  assign n2518 = ( n2513 & n2516 ) | ( n2513 & ~n2517 ) | ( n2516 & ~n2517 ) ;
  assign n2519 = ( ~n2506 & n2512 ) | ( ~n2506 & n2518 ) | ( n2512 & n2518 ) ;
  assign n2520 = ( n2506 & n2512 ) | ( n2506 & n2518 ) | ( n2512 & n2518 ) ;
  assign n2521 = ( n2506 & n2519 ) | ( n2506 & ~n2520 ) | ( n2519 & ~n2520 ) ;
  assign n2522 = x9 & x40 ;
  assign n2523 = x12 & x37 ;
  assign n2524 = x10 & x39 ;
  assign n2525 = ( ~n2522 & n2523 ) | ( ~n2522 & n2524 ) | ( n2523 & n2524 ) ;
  assign n2526 = ( n2522 & n2523 ) | ( n2522 & n2524 ) | ( n2523 & n2524 ) ;
  assign n2527 = ( n2522 & n2525 ) | ( n2522 & ~n2526 ) | ( n2525 & ~n2526 ) ;
  assign n2528 = x19 & x30 ;
  assign n2529 = x20 & x29 ;
  assign n2530 = x21 & x28 ;
  assign n2531 = ( ~n2528 & n2529 ) | ( ~n2528 & n2530 ) | ( n2529 & n2530 ) ;
  assign n2532 = ( n2528 & n2529 ) | ( n2528 & n2530 ) | ( n2529 & n2530 ) ;
  assign n2533 = ( n2528 & n2531 ) | ( n2528 & ~n2532 ) | ( n2531 & ~n2532 ) ;
  assign n2534 = x22 & x27 ;
  assign n2535 = x2 & x47 ;
  assign n2536 = x3 & x46 ;
  assign n2537 = ( ~n2534 & n2535 ) | ( ~n2534 & n2536 ) | ( n2535 & n2536 ) ;
  assign n2538 = ( n2534 & n2535 ) | ( n2534 & n2536 ) | ( n2535 & n2536 ) ;
  assign n2539 = ( n2534 & n2537 ) | ( n2534 & ~n2538 ) | ( n2537 & ~n2538 ) ;
  assign n2540 = ( ~n2527 & n2533 ) | ( ~n2527 & n2539 ) | ( n2533 & n2539 ) ;
  assign n2541 = ( n2527 & n2533 ) | ( n2527 & n2539 ) | ( n2533 & n2539 ) ;
  assign n2542 = ( n2527 & n2540 ) | ( n2527 & ~n2541 ) | ( n2540 & ~n2541 ) ;
  assign n2543 = ( n2500 & n2521 ) | ( n2500 & n2542 ) | ( n2521 & n2542 ) ;
  assign n2544 = ( ~n2500 & n2521 ) | ( ~n2500 & n2542 ) | ( n2521 & n2542 ) ;
  assign n2545 = ( n2500 & ~n2543 ) | ( n2500 & n2544 ) | ( ~n2543 & n2544 ) ;
  assign n2546 = ( n2459 & n2475 ) | ( n2459 & n2545 ) | ( n2475 & n2545 ) ;
  assign n2547 = ( ~n2459 & n2475 ) | ( ~n2459 & n2545 ) | ( n2475 & n2545 ) ;
  assign n2548 = ( n2459 & ~n2546 ) | ( n2459 & n2547 ) | ( ~n2546 & n2547 ) ;
  assign n2549 = ( n2399 & ~n2405 ) | ( n2399 & n2414 ) | ( ~n2405 & n2414 ) ;
  assign n2550 = ( n2399 & n2405 ) | ( n2399 & n2414 ) | ( n2405 & n2414 ) ;
  assign n2551 = ( n2405 & n2549 ) | ( n2405 & ~n2550 ) | ( n2549 & ~n2550 ) ;
  assign n2552 = ( n2429 & n2472 ) | ( n2429 & n2551 ) | ( n2472 & n2551 ) ;
  assign n2553 = ( n2429 & ~n2472 ) | ( n2429 & n2551 ) | ( ~n2472 & n2551 ) ;
  assign n2554 = ( n2472 & ~n2552 ) | ( n2472 & n2553 ) | ( ~n2552 & n2553 ) ;
  assign n2555 = ( n2420 & ~n2426 ) | ( n2420 & n2444 ) | ( ~n2426 & n2444 ) ;
  assign n2556 = ( n2420 & n2426 ) | ( n2420 & n2444 ) | ( n2426 & n2444 ) ;
  assign n2557 = ( n2426 & n2555 ) | ( n2426 & ~n2556 ) | ( n2555 & ~n2556 ) ;
  assign n2558 = ~x48 & n2464 ;
  assign n2559 = x1 & x48 ;
  assign n2560 = x25 | n2559 ;
  assign n2561 = x48 & n783 ;
  assign n2562 = ( n2464 & n2560 ) | ( n2464 & ~n2561 ) | ( n2560 & ~n2561 ) ;
  assign n2563 = ( n2393 & n2558 ) | ( n2393 & n2562 ) | ( n2558 & n2562 ) ;
  assign n2564 = ( n2393 & ~n2558 ) | ( n2393 & n2562 ) | ( ~n2558 & n2562 ) ;
  assign n2565 = ( n2558 & ~n2563 ) | ( n2558 & n2564 ) | ( ~n2563 & n2564 ) ;
  assign n2566 = ( n2408 & n2557 ) | ( n2408 & n2565 ) | ( n2557 & n2565 ) ;
  assign n2567 = ( ~n2408 & n2557 ) | ( ~n2408 & n2565 ) | ( n2557 & n2565 ) ;
  assign n2568 = ( n2408 & ~n2566 ) | ( n2408 & n2567 ) | ( ~n2566 & n2567 ) ;
  assign n2569 = ( ~n2431 & n2554 ) | ( ~n2431 & n2568 ) | ( n2554 & n2568 ) ;
  assign n2570 = ( n2431 & n2554 ) | ( n2431 & n2568 ) | ( n2554 & n2568 ) ;
  assign n2571 = ( n2431 & n2569 ) | ( n2431 & ~n2570 ) | ( n2569 & ~n2570 ) ;
  assign n2572 = ( n2438 & n2447 ) | ( n2438 & ~n2453 ) | ( n2447 & ~n2453 ) ;
  assign n2573 = ( n2438 & n2447 ) | ( n2438 & n2453 ) | ( n2447 & n2453 ) ;
  assign n2574 = ( n2453 & n2572 ) | ( n2453 & ~n2573 ) | ( n2572 & ~n2573 ) ;
  assign n2575 = ( n2450 & n2455 ) | ( n2450 & n2574 ) | ( n2455 & n2574 ) ;
  assign n2576 = ( ~n2450 & n2455 ) | ( ~n2450 & n2574 ) | ( n2455 & n2574 ) ;
  assign n2577 = ( n2450 & ~n2575 ) | ( n2450 & n2576 ) | ( ~n2575 & n2576 ) ;
  assign n2578 = ( ~n2435 & n2571 ) | ( ~n2435 & n2577 ) | ( n2571 & n2577 ) ;
  assign n2579 = ( n2435 & n2571 ) | ( n2435 & n2577 ) | ( n2571 & n2577 ) ;
  assign n2580 = ( n2435 & n2578 ) | ( n2435 & ~n2579 ) | ( n2578 & ~n2579 ) ;
  assign n2581 = ( ~n2478 & n2548 ) | ( ~n2478 & n2580 ) | ( n2548 & n2580 ) ;
  assign n2582 = ( n2478 & n2548 ) | ( n2478 & n2580 ) | ( n2548 & n2580 ) ;
  assign n2583 = ( n2478 & n2581 ) | ( n2478 & ~n2582 ) | ( n2581 & ~n2582 ) ;
  assign n2584 = ( ~n2480 & n2484 ) | ( ~n2480 & n2583 ) | ( n2484 & n2583 ) ;
  assign n2585 = ( n2480 & n2484 ) | ( n2480 & n2583 ) | ( n2484 & n2583 ) ;
  assign n2586 = ( n2480 & n2584 ) | ( n2480 & ~n2585 ) | ( n2584 & ~n2585 ) ;
  assign n2587 = ( n2496 & ~n2505 ) | ( n2496 & n2538 ) | ( ~n2505 & n2538 ) ;
  assign n2588 = ( n2496 & n2505 ) | ( n2496 & n2538 ) | ( n2505 & n2538 ) ;
  assign n2589 = ( n2505 & n2587 ) | ( n2505 & ~n2588 ) | ( n2587 & ~n2588 ) ;
  assign n2590 = ( n2550 & n2556 ) | ( n2550 & n2589 ) | ( n2556 & n2589 ) ;
  assign n2591 = ( ~n2550 & n2556 ) | ( ~n2550 & n2589 ) | ( n2556 & n2589 ) ;
  assign n2592 = ( n2550 & ~n2590 ) | ( n2550 & n2591 ) | ( ~n2590 & n2591 ) ;
  assign n2593 = ( ~n2552 & n2566 ) | ( ~n2552 & n2592 ) | ( n2566 & n2592 ) ;
  assign n2594 = ( n2552 & n2566 ) | ( n2552 & n2592 ) | ( n2566 & n2592 ) ;
  assign n2595 = ( n2552 & n2593 ) | ( n2552 & ~n2594 ) | ( n2593 & ~n2594 ) ;
  assign n2596 = ( n2490 & ~n2517 ) | ( n2490 & n2532 ) | ( ~n2517 & n2532 ) ;
  assign n2597 = ( n2490 & n2517 ) | ( n2490 & n2532 ) | ( n2517 & n2532 ) ;
  assign n2598 = ( n2517 & n2596 ) | ( n2517 & ~n2597 ) | ( n2596 & ~n2597 ) ;
  assign n2599 = ( n2520 & n2573 ) | ( n2520 & n2598 ) | ( n2573 & n2598 ) ;
  assign n2600 = ( ~n2520 & n2573 ) | ( ~n2520 & n2598 ) | ( n2573 & n2598 ) ;
  assign n2601 = ( n2520 & ~n2599 ) | ( n2520 & n2600 ) | ( ~n2599 & n2600 ) ;
  assign n2602 = x24 & x26 ;
  assign n2603 = x1 & x49 ;
  assign n2604 = n2602 & n2603 ;
  assign n2605 = n2602 | n2603 ;
  assign n2606 = ~n2604 & n2605 ;
  assign n2607 = ( n2511 & n2526 ) | ( n2511 & n2606 ) | ( n2526 & n2606 ) ;
  assign n2608 = ( ~n2511 & n2526 ) | ( ~n2511 & n2606 ) | ( n2526 & n2606 ) ;
  assign n2609 = ( n2511 & ~n2607 ) | ( n2511 & n2608 ) | ( ~n2607 & n2608 ) ;
  assign n2610 = ( ~n2498 & n2541 ) | ( ~n2498 & n2609 ) | ( n2541 & n2609 ) ;
  assign n2611 = ( n2498 & n2541 ) | ( n2498 & n2609 ) | ( n2541 & n2609 ) ;
  assign n2612 = ( n2498 & n2610 ) | ( n2498 & ~n2611 ) | ( n2610 & ~n2611 ) ;
  assign n2613 = ( n2543 & n2601 ) | ( n2543 & n2612 ) | ( n2601 & n2612 ) ;
  assign n2614 = ( ~n2543 & n2601 ) | ( ~n2543 & n2612 ) | ( n2601 & n2612 ) ;
  assign n2615 = ( n2543 & ~n2613 ) | ( n2543 & n2614 ) | ( ~n2613 & n2614 ) ;
  assign n2616 = ( n2546 & n2595 ) | ( n2546 & n2615 ) | ( n2595 & n2615 ) ;
  assign n2617 = ( ~n2546 & n2595 ) | ( ~n2546 & n2615 ) | ( n2595 & n2615 ) ;
  assign n2618 = ( n2546 & ~n2616 ) | ( n2546 & n2617 ) | ( ~n2616 & n2617 ) ;
  assign n2619 = x18 & x32 ;
  assign n2620 = x22 & x28 ;
  assign n2621 = x23 & x27 ;
  assign n2622 = ( ~n2619 & n2620 ) | ( ~n2619 & n2621 ) | ( n2620 & n2621 ) ;
  assign n2623 = ( n2619 & n2620 ) | ( n2619 & n2621 ) | ( n2620 & n2621 ) ;
  assign n2624 = ( n2619 & n2622 ) | ( n2619 & ~n2623 ) | ( n2622 & ~n2623 ) ;
  assign n2625 = x16 & x34 ;
  assign n2626 = x5 & x45 ;
  assign n2627 = x15 & x35 ;
  assign n2628 = ( ~n2625 & n2626 ) | ( ~n2625 & n2627 ) | ( n2626 & n2627 ) ;
  assign n2629 = ( n2625 & n2626 ) | ( n2625 & n2627 ) | ( n2626 & n2627 ) ;
  assign n2630 = ( n2625 & n2628 ) | ( n2625 & ~n2629 ) | ( n2628 & ~n2629 ) ;
  assign n2631 = ( n2563 & n2624 ) | ( n2563 & n2630 ) | ( n2624 & n2630 ) ;
  assign n2632 = ( ~n2563 & n2624 ) | ( ~n2563 & n2630 ) | ( n2624 & n2630 ) ;
  assign n2633 = ( n2563 & ~n2631 ) | ( n2563 & n2632 ) | ( ~n2631 & n2632 ) ;
  assign n2634 = x0 & x50 ;
  assign n2635 = x2 & x48 ;
  assign n2636 = ( ~n2561 & n2634 ) | ( ~n2561 & n2635 ) | ( n2634 & n2635 ) ;
  assign n2637 = ( n2561 & n2634 ) | ( n2561 & n2635 ) | ( n2634 & n2635 ) ;
  assign n2638 = ( n2561 & n2636 ) | ( n2561 & ~n2637 ) | ( n2636 & ~n2637 ) ;
  assign n2639 = x3 & x47 ;
  assign n2640 = x4 & x46 ;
  assign n2641 = x17 & x33 ;
  assign n2642 = ( ~n2639 & n2640 ) | ( ~n2639 & n2641 ) | ( n2640 & n2641 ) ;
  assign n2643 = ( n2639 & n2640 ) | ( n2639 & n2641 ) | ( n2640 & n2641 ) ;
  assign n2644 = ( n2639 & n2642 ) | ( n2639 & ~n2643 ) | ( n2642 & ~n2643 ) ;
  assign n2645 = x19 & x31 ;
  assign n2646 = x21 & x29 ;
  assign n2647 = x20 & x30 ;
  assign n2648 = ( ~n2645 & n2646 ) | ( ~n2645 & n2647 ) | ( n2646 & n2647 ) ;
  assign n2649 = ( n2645 & n2646 ) | ( n2645 & n2647 ) | ( n2646 & n2647 ) ;
  assign n2650 = ( n2645 & n2648 ) | ( n2645 & ~n2649 ) | ( n2648 & ~n2649 ) ;
  assign n2651 = ( ~n2638 & n2644 ) | ( ~n2638 & n2650 ) | ( n2644 & n2650 ) ;
  assign n2652 = ( n2638 & n2644 ) | ( n2638 & n2650 ) | ( n2644 & n2650 ) ;
  assign n2653 = ( n2638 & n2651 ) | ( n2638 & ~n2652 ) | ( n2651 & ~n2652 ) ;
  assign n2654 = x12 & x38 ;
  assign n2655 = x11 & x39 ;
  assign n2656 = x10 & x40 ;
  assign n2657 = ( ~n2654 & n2655 ) | ( ~n2654 & n2656 ) | ( n2655 & n2656 ) ;
  assign n2658 = ( n2654 & n2655 ) | ( n2654 & n2656 ) | ( n2655 & n2656 ) ;
  assign n2659 = ( n2654 & n2657 ) | ( n2654 & ~n2658 ) | ( n2657 & ~n2658 ) ;
  assign n2660 = x6 & x44 ;
  assign n2661 = x7 & x43 ;
  assign n2662 = x14 & x36 ;
  assign n2663 = ( ~n2660 & n2661 ) | ( ~n2660 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2664 = ( n2660 & n2661 ) | ( n2660 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2665 = ( n2660 & n2663 ) | ( n2660 & ~n2664 ) | ( n2663 & ~n2664 ) ;
  assign n2666 = x8 & x42 ;
  assign n2667 = x13 & x37 ;
  assign n2668 = x9 & x41 ;
  assign n2669 = ( ~n2666 & n2667 ) | ( ~n2666 & n2668 ) | ( n2667 & n2668 ) ;
  assign n2670 = ( n2666 & n2667 ) | ( n2666 & n2668 ) | ( n2667 & n2668 ) ;
  assign n2671 = ( n2666 & n2669 ) | ( n2666 & ~n2670 ) | ( n2669 & ~n2670 ) ;
  assign n2672 = ( ~n2659 & n2665 ) | ( ~n2659 & n2671 ) | ( n2665 & n2671 ) ;
  assign n2673 = ( n2659 & n2665 ) | ( n2659 & n2671 ) | ( n2665 & n2671 ) ;
  assign n2674 = ( n2659 & n2672 ) | ( n2659 & ~n2673 ) | ( n2672 & ~n2673 ) ;
  assign n2675 = ( n2633 & n2653 ) | ( n2633 & n2674 ) | ( n2653 & n2674 ) ;
  assign n2676 = ( ~n2633 & n2653 ) | ( ~n2633 & n2674 ) | ( n2653 & n2674 ) ;
  assign n2677 = ( n2633 & ~n2675 ) | ( n2633 & n2676 ) | ( ~n2675 & n2676 ) ;
  assign n2678 = ( n2570 & n2575 ) | ( n2570 & n2677 ) | ( n2575 & n2677 ) ;
  assign n2679 = ( n2570 & ~n2575 ) | ( n2570 & n2677 ) | ( ~n2575 & n2677 ) ;
  assign n2680 = ( n2575 & ~n2678 ) | ( n2575 & n2679 ) | ( ~n2678 & n2679 ) ;
  assign n2681 = ( n2579 & n2618 ) | ( n2579 & n2680 ) | ( n2618 & n2680 ) ;
  assign n2682 = ( ~n2579 & n2618 ) | ( ~n2579 & n2680 ) | ( n2618 & n2680 ) ;
  assign n2683 = ( n2579 & ~n2681 ) | ( n2579 & n2682 ) | ( ~n2681 & n2682 ) ;
  assign n2684 = ( ~n2582 & n2585 ) | ( ~n2582 & n2683 ) | ( n2585 & n2683 ) ;
  assign n2685 = ( n2582 & n2585 ) | ( n2582 & n2683 ) | ( n2585 & n2683 ) ;
  assign n2686 = ( n2582 & n2684 ) | ( n2582 & ~n2685 ) | ( n2684 & ~n2685 ) ;
  assign n2687 = x0 & x51 ;
  assign n2688 = x1 & x50 ;
  assign n2689 = x26 & n2688 ;
  assign n2690 = x26 | n2688 ;
  assign n2691 = ~n2689 & n2690 ;
  assign n2692 = ( n2604 & n2687 ) | ( n2604 & n2691 ) | ( n2687 & n2691 ) ;
  assign n2693 = ( ~n2604 & n2687 ) | ( ~n2604 & n2691 ) | ( n2687 & n2691 ) ;
  assign n2694 = ( n2604 & ~n2692 ) | ( n2604 & n2693 ) | ( ~n2692 & n2693 ) ;
  assign n2695 = x17 & x34 ;
  assign n2696 = x20 & x31 ;
  assign n2697 = x19 & x32 ;
  assign n2698 = ( ~n2695 & n2696 ) | ( ~n2695 & n2697 ) | ( n2696 & n2697 ) ;
  assign n2699 = ( n2695 & n2696 ) | ( n2695 & n2697 ) | ( n2696 & n2697 ) ;
  assign n2700 = ( n2695 & n2698 ) | ( n2695 & ~n2699 ) | ( n2698 & ~n2699 ) ;
  assign n2701 = ( ~n2597 & n2694 ) | ( ~n2597 & n2700 ) | ( n2694 & n2700 ) ;
  assign n2702 = ( n2597 & n2694 ) | ( n2597 & n2700 ) | ( n2694 & n2700 ) ;
  assign n2703 = ( n2597 & n2701 ) | ( n2597 & ~n2702 ) | ( n2701 & ~n2702 ) ;
  assign n2704 = x15 & x36 ;
  assign n2705 = x6 & x45 ;
  assign n2706 = x14 & x37 ;
  assign n2707 = ( ~n2704 & n2705 ) | ( ~n2704 & n2706 ) | ( n2705 & n2706 ) ;
  assign n2708 = ( n2704 & n2705 ) | ( n2704 & n2706 ) | ( n2705 & n2706 ) ;
  assign n2709 = ( n2704 & n2707 ) | ( n2704 & ~n2708 ) | ( n2707 & ~n2708 ) ;
  assign n2710 = x18 & x33 ;
  assign n2711 = x5 & x46 ;
  assign n2712 = x16 & x35 ;
  assign n2713 = ( ~n2710 & n2711 ) | ( ~n2710 & n2712 ) | ( n2711 & n2712 ) ;
  assign n2714 = ( n2710 & n2711 ) | ( n2710 & n2712 ) | ( n2711 & n2712 ) ;
  assign n2715 = ( n2710 & n2713 ) | ( n2710 & ~n2714 ) | ( n2713 & ~n2714 ) ;
  assign n2716 = x21 & x30 ;
  assign n2717 = x22 & x29 ;
  assign n2718 = x23 & x28 ;
  assign n2719 = ( ~n2716 & n2717 ) | ( ~n2716 & n2718 ) | ( n2717 & n2718 ) ;
  assign n2720 = ( n2716 & n2717 ) | ( n2716 & n2718 ) | ( n2717 & n2718 ) ;
  assign n2721 = ( n2716 & n2719 ) | ( n2716 & ~n2720 ) | ( n2719 & ~n2720 ) ;
  assign n2722 = ( ~n2709 & n2715 ) | ( ~n2709 & n2721 ) | ( n2715 & n2721 ) ;
  assign n2723 = ( n2709 & n2715 ) | ( n2709 & n2721 ) | ( n2715 & n2721 ) ;
  assign n2724 = ( n2709 & n2722 ) | ( n2709 & ~n2723 ) | ( n2722 & ~n2723 ) ;
  assign n2725 = x9 & x42 ;
  assign n2726 = x12 & x39 ;
  assign n2727 = x10 & x41 ;
  assign n2728 = ( ~n2725 & n2726 ) | ( ~n2725 & n2727 ) | ( n2726 & n2727 ) ;
  assign n2729 = ( n2725 & n2726 ) | ( n2725 & n2727 ) | ( n2726 & n2727 ) ;
  assign n2730 = ( n2725 & n2728 ) | ( n2725 & ~n2729 ) | ( n2728 & ~n2729 ) ;
  assign n2731 = x11 & x40 ;
  assign n2732 = x25 & x26 ;
  assign n2733 = x24 & x27 ;
  assign n2734 = ( ~n2731 & n2732 ) | ( ~n2731 & n2733 ) | ( n2732 & n2733 ) ;
  assign n2735 = ( n2731 & n2732 ) | ( n2731 & n2733 ) | ( n2732 & n2733 ) ;
  assign n2736 = ( n2731 & n2734 ) | ( n2731 & ~n2735 ) | ( n2734 & ~n2735 ) ;
  assign n2737 = x7 & x44 ;
  assign n2738 = x13 & x38 ;
  assign n2739 = x8 & x43 ;
  assign n2740 = ( ~n2737 & n2738 ) | ( ~n2737 & n2739 ) | ( n2738 & n2739 ) ;
  assign n2741 = ( n2737 & n2738 ) | ( n2737 & n2739 ) | ( n2738 & n2739 ) ;
  assign n2742 = ( n2737 & n2740 ) | ( n2737 & ~n2741 ) | ( n2740 & ~n2741 ) ;
  assign n2743 = ( ~n2730 & n2736 ) | ( ~n2730 & n2742 ) | ( n2736 & n2742 ) ;
  assign n2744 = ( n2730 & n2736 ) | ( n2730 & n2742 ) | ( n2736 & n2742 ) ;
  assign n2745 = ( n2730 & n2743 ) | ( n2730 & ~n2744 ) | ( n2743 & ~n2744 ) ;
  assign n2746 = ( ~n2703 & n2724 ) | ( ~n2703 & n2745 ) | ( n2724 & n2745 ) ;
  assign n2747 = ( n2703 & n2724 ) | ( n2703 & n2745 ) | ( n2724 & n2745 ) ;
  assign n2748 = ( n2703 & n2746 ) | ( n2703 & ~n2747 ) | ( n2746 & ~n2747 ) ;
  assign n2749 = ( ~n2594 & n2613 ) | ( ~n2594 & n2748 ) | ( n2613 & n2748 ) ;
  assign n2750 = ( n2594 & n2613 ) | ( n2594 & n2748 ) | ( n2613 & n2748 ) ;
  assign n2751 = ( n2594 & n2749 ) | ( n2594 & ~n2750 ) | ( n2749 & ~n2750 ) ;
  assign n2752 = ( n2588 & n2607 ) | ( n2588 & n2652 ) | ( n2607 & n2652 ) ;
  assign n2753 = ( ~n2588 & n2607 ) | ( ~n2588 & n2652 ) | ( n2607 & n2652 ) ;
  assign n2754 = ( n2588 & ~n2752 ) | ( n2588 & n2753 ) | ( ~n2752 & n2753 ) ;
  assign n2755 = ( ~n2599 & n2611 ) | ( ~n2599 & n2754 ) | ( n2611 & n2754 ) ;
  assign n2756 = ( n2599 & n2611 ) | ( n2599 & n2754 ) | ( n2611 & n2754 ) ;
  assign n2757 = ( n2599 & n2755 ) | ( n2599 & ~n2756 ) | ( n2755 & ~n2756 ) ;
  assign n2758 = x2 & x49 ;
  assign n2759 = x3 & x48 ;
  assign n2760 = x4 & x47 ;
  assign n2761 = ( ~n2758 & n2759 ) | ( ~n2758 & n2760 ) | ( n2759 & n2760 ) ;
  assign n2762 = ( n2758 & n2759 ) | ( n2758 & n2760 ) | ( n2759 & n2760 ) ;
  assign n2763 = ( n2758 & n2761 ) | ( n2758 & ~n2762 ) | ( n2761 & ~n2762 ) ;
  assign n2764 = ( ~n2629 & n2658 ) | ( ~n2629 & n2763 ) | ( n2658 & n2763 ) ;
  assign n2765 = ( n2629 & n2658 ) | ( n2629 & n2763 ) | ( n2658 & n2763 ) ;
  assign n2766 = ( n2629 & n2764 ) | ( n2629 & ~n2765 ) | ( n2764 & ~n2765 ) ;
  assign n2767 = ( ~n2590 & n2631 ) | ( ~n2590 & n2766 ) | ( n2631 & n2766 ) ;
  assign n2768 = ( n2590 & n2631 ) | ( n2590 & n2766 ) | ( n2631 & n2766 ) ;
  assign n2769 = ( n2590 & n2767 ) | ( n2590 & ~n2768 ) | ( n2767 & ~n2768 ) ;
  assign n2770 = ( ~n2637 & n2643 ) | ( ~n2637 & n2649 ) | ( n2643 & n2649 ) ;
  assign n2771 = ( n2637 & n2643 ) | ( n2637 & n2649 ) | ( n2643 & n2649 ) ;
  assign n2772 = ( n2637 & n2770 ) | ( n2637 & ~n2771 ) | ( n2770 & ~n2771 ) ;
  assign n2773 = ( n2623 & ~n2664 ) | ( n2623 & n2670 ) | ( ~n2664 & n2670 ) ;
  assign n2774 = ( n2623 & n2664 ) | ( n2623 & n2670 ) | ( n2664 & n2670 ) ;
  assign n2775 = ( n2664 & n2773 ) | ( n2664 & ~n2774 ) | ( n2773 & ~n2774 ) ;
  assign n2776 = ( n2673 & n2772 ) | ( n2673 & n2775 ) | ( n2772 & n2775 ) ;
  assign n2777 = ( ~n2673 & n2772 ) | ( ~n2673 & n2775 ) | ( n2772 & n2775 ) ;
  assign n2778 = ( n2673 & ~n2776 ) | ( n2673 & n2777 ) | ( ~n2776 & n2777 ) ;
  assign n2779 = ( n2675 & n2769 ) | ( n2675 & n2778 ) | ( n2769 & n2778 ) ;
  assign n2780 = ( n2675 & ~n2769 ) | ( n2675 & n2778 ) | ( ~n2769 & n2778 ) ;
  assign n2781 = ( n2769 & ~n2779 ) | ( n2769 & n2780 ) | ( ~n2779 & n2780 ) ;
  assign n2782 = ( n2678 & n2757 ) | ( n2678 & n2781 ) | ( n2757 & n2781 ) ;
  assign n2783 = ( ~n2678 & n2757 ) | ( ~n2678 & n2781 ) | ( n2757 & n2781 ) ;
  assign n2784 = ( n2678 & ~n2782 ) | ( n2678 & n2783 ) | ( ~n2782 & n2783 ) ;
  assign n2785 = ( ~n2616 & n2751 ) | ( ~n2616 & n2784 ) | ( n2751 & n2784 ) ;
  assign n2786 = ( n2616 & n2751 ) | ( n2616 & n2784 ) | ( n2751 & n2784 ) ;
  assign n2787 = ( n2616 & n2785 ) | ( n2616 & ~n2786 ) | ( n2785 & ~n2786 ) ;
  assign n2788 = ( n2681 & n2685 ) | ( n2681 & n2787 ) | ( n2685 & n2787 ) ;
  assign n2789 = ( ~n2681 & n2685 ) | ( ~n2681 & n2787 ) | ( n2685 & n2787 ) ;
  assign n2790 = ( n2681 & ~n2788 ) | ( n2681 & n2789 ) | ( ~n2788 & n2789 ) ;
  assign n2791 = x15 & x37 ;
  assign n2792 = x7 & x45 ;
  assign n2793 = x8 & x44 ;
  assign n2794 = ( ~n2791 & n2792 ) | ( ~n2791 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2795 = ( n2791 & n2792 ) | ( n2791 & n2793 ) | ( n2792 & n2793 ) ;
  assign n2796 = ( n2791 & n2794 ) | ( n2791 & ~n2795 ) | ( n2794 & ~n2795 ) ;
  assign n2797 = x10 & x42 ;
  assign n2798 = x12 & x40 ;
  assign n2799 = x11 & x41 ;
  assign n2800 = ( ~n2797 & n2798 ) | ( ~n2797 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2801 = ( n2797 & n2798 ) | ( n2797 & n2799 ) | ( n2798 & n2799 ) ;
  assign n2802 = ( n2797 & n2800 ) | ( n2797 & ~n2801 ) | ( n2800 & ~n2801 ) ;
  assign n2803 = x5 & x47 ;
  assign n2804 = x16 & x36 ;
  assign n2805 = x6 & x46 ;
  assign n2806 = ( ~n2803 & n2804 ) | ( ~n2803 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2807 = ( n2803 & n2804 ) | ( n2803 & n2805 ) | ( n2804 & n2805 ) ;
  assign n2808 = ( n2803 & n2806 ) | ( n2803 & ~n2807 ) | ( n2806 & ~n2807 ) ;
  assign n2809 = ( ~n2796 & n2802 ) | ( ~n2796 & n2808 ) | ( n2802 & n2808 ) ;
  assign n2810 = ( n2796 & n2802 ) | ( n2796 & n2808 ) | ( n2802 & n2808 ) ;
  assign n2811 = ( n2796 & n2809 ) | ( n2796 & ~n2810 ) | ( n2809 & ~n2810 ) ;
  assign n2812 = x14 & x38 ;
  assign n2813 = x9 & x43 ;
  assign n2814 = x13 & x39 ;
  assign n2815 = ( ~n2812 & n2813 ) | ( ~n2812 & n2814 ) | ( n2813 & n2814 ) ;
  assign n2816 = ( n2812 & n2813 ) | ( n2812 & n2814 ) | ( n2813 & n2814 ) ;
  assign n2817 = ( n2812 & n2815 ) | ( n2812 & ~n2816 ) | ( n2815 & ~n2816 ) ;
  assign n2818 = x22 & x30 ;
  assign n2819 = x23 & x29 ;
  assign n2820 = x24 & x28 ;
  assign n2821 = ( ~n2818 & n2819 ) | ( ~n2818 & n2820 ) | ( n2819 & n2820 ) ;
  assign n2822 = ( n2818 & n2819 ) | ( n2818 & n2820 ) | ( n2819 & n2820 ) ;
  assign n2823 = ( n2818 & n2821 ) | ( n2818 & ~n2822 ) | ( n2821 & ~n2822 ) ;
  assign n2824 = x20 & x32 ;
  assign n2825 = x21 & x31 ;
  assign n2826 = ( ~n1310 & n2824 ) | ( ~n1310 & n2825 ) | ( n2824 & n2825 ) ;
  assign n2827 = ( n1310 & n2824 ) | ( n1310 & n2825 ) | ( n2824 & n2825 ) ;
  assign n2828 = ( n1310 & n2826 ) | ( n1310 & ~n2827 ) | ( n2826 & ~n2827 ) ;
  assign n2829 = ( ~n2817 & n2823 ) | ( ~n2817 & n2828 ) | ( n2823 & n2828 ) ;
  assign n2830 = ( n2817 & n2823 ) | ( n2817 & n2828 ) | ( n2823 & n2828 ) ;
  assign n2831 = ( n2817 & n2829 ) | ( n2817 & ~n2830 ) | ( n2829 & ~n2830 ) ;
  assign n2832 = ( n2776 & n2811 ) | ( n2776 & n2831 ) | ( n2811 & n2831 ) ;
  assign n2833 = ( ~n2776 & n2811 ) | ( ~n2776 & n2831 ) | ( n2811 & n2831 ) ;
  assign n2834 = ( n2776 & ~n2832 ) | ( n2776 & n2833 ) | ( ~n2832 & n2833 ) ;
  assign n2835 = ( n2756 & n2779 ) | ( n2756 & n2834 ) | ( n2779 & n2834 ) ;
  assign n2836 = ( n2756 & ~n2779 ) | ( n2756 & n2834 ) | ( ~n2779 & n2834 ) ;
  assign n2837 = ( n2779 & ~n2835 ) | ( n2779 & n2836 ) | ( ~n2835 & n2836 ) ;
  assign n2838 = x19 & x33 ;
  assign n2839 = x2 & x50 ;
  assign n2840 = x3 & x49 ;
  assign n2841 = ( ~n2838 & n2839 ) | ( ~n2838 & n2840 ) | ( n2839 & n2840 ) ;
  assign n2842 = ( n2838 & n2839 ) | ( n2838 & n2840 ) | ( n2839 & n2840 ) ;
  assign n2843 = ( n2838 & n2841 ) | ( n2838 & ~n2842 ) | ( n2841 & ~n2842 ) ;
  assign n2844 = ( ~n2771 & n2774 ) | ( ~n2771 & n2843 ) | ( n2774 & n2843 ) ;
  assign n2845 = ( n2771 & n2774 ) | ( n2771 & n2843 ) | ( n2774 & n2843 ) ;
  assign n2846 = ( n2771 & n2844 ) | ( n2771 & ~n2845 ) | ( n2844 & ~n2845 ) ;
  assign n2847 = x25 & x27 ;
  assign n2848 = x1 & x51 ;
  assign n2849 = n2847 & n2848 ;
  assign n2850 = n2847 | n2848 ;
  assign n2851 = ~n2849 & n2850 ;
  assign n2852 = ( ~n2689 & n2735 ) | ( ~n2689 & n2851 ) | ( n2735 & n2851 ) ;
  assign n2853 = ( n2689 & n2735 ) | ( n2689 & n2851 ) | ( n2735 & n2851 ) ;
  assign n2854 = ( n2689 & n2852 ) | ( n2689 & ~n2853 ) | ( n2852 & ~n2853 ) ;
  assign n2855 = ( ~n2744 & n2765 ) | ( ~n2744 & n2854 ) | ( n2765 & n2854 ) ;
  assign n2856 = ( n2744 & n2765 ) | ( n2744 & n2854 ) | ( n2765 & n2854 ) ;
  assign n2857 = ( n2744 & n2855 ) | ( n2744 & ~n2856 ) | ( n2855 & ~n2856 ) ;
  assign n2858 = ( ~n2768 & n2846 ) | ( ~n2768 & n2857 ) | ( n2846 & n2857 ) ;
  assign n2859 = ( n2768 & n2846 ) | ( n2768 & n2857 ) | ( n2846 & n2857 ) ;
  assign n2860 = ( n2768 & n2858 ) | ( n2768 & ~n2859 ) | ( n2858 & ~n2859 ) ;
  assign n2861 = x4 & x48 ;
  assign n2862 = x0 & x52 ;
  assign n2863 = x17 & x35 ;
  assign n2864 = ( ~n2861 & n2862 ) | ( ~n2861 & n2863 ) | ( n2862 & n2863 ) ;
  assign n2865 = ( n2861 & n2862 ) | ( n2861 & n2863 ) | ( n2862 & n2863 ) ;
  assign n2866 = ( n2861 & n2864 ) | ( n2861 & ~n2865 ) | ( n2864 & ~n2865 ) ;
  assign n2867 = ( n2692 & n2729 ) | ( n2692 & n2866 ) | ( n2729 & n2866 ) ;
  assign n2868 = ( ~n2692 & n2729 ) | ( ~n2692 & n2866 ) | ( n2729 & n2866 ) ;
  assign n2869 = ( n2692 & ~n2867 ) | ( n2692 & n2868 ) | ( ~n2867 & n2868 ) ;
  assign n2870 = ( n2702 & n2752 ) | ( n2702 & n2869 ) | ( n2752 & n2869 ) ;
  assign n2871 = ( ~n2702 & n2752 ) | ( ~n2702 & n2869 ) | ( n2752 & n2869 ) ;
  assign n2872 = ( n2702 & ~n2870 ) | ( n2702 & n2871 ) | ( ~n2870 & n2871 ) ;
  assign n2873 = ( n2714 & ~n2720 ) | ( n2714 & n2741 ) | ( ~n2720 & n2741 ) ;
  assign n2874 = ( n2714 & n2720 ) | ( n2714 & n2741 ) | ( n2720 & n2741 ) ;
  assign n2875 = ( n2720 & n2873 ) | ( n2720 & ~n2874 ) | ( n2873 & ~n2874 ) ;
  assign n2876 = ( n2699 & ~n2708 ) | ( n2699 & n2762 ) | ( ~n2708 & n2762 ) ;
  assign n2877 = ( n2699 & n2708 ) | ( n2699 & n2762 ) | ( n2708 & n2762 ) ;
  assign n2878 = ( n2708 & n2876 ) | ( n2708 & ~n2877 ) | ( n2876 & ~n2877 ) ;
  assign n2879 = ( ~n2723 & n2875 ) | ( ~n2723 & n2878 ) | ( n2875 & n2878 ) ;
  assign n2880 = ( n2723 & n2875 ) | ( n2723 & n2878 ) | ( n2875 & n2878 ) ;
  assign n2881 = ( n2723 & n2879 ) | ( n2723 & ~n2880 ) | ( n2879 & ~n2880 ) ;
  assign n2882 = ( ~n2747 & n2872 ) | ( ~n2747 & n2881 ) | ( n2872 & n2881 ) ;
  assign n2883 = ( n2747 & n2872 ) | ( n2747 & n2881 ) | ( n2872 & n2881 ) ;
  assign n2884 = ( n2747 & n2882 ) | ( n2747 & ~n2883 ) | ( n2882 & ~n2883 ) ;
  assign n2885 = ( n2750 & n2860 ) | ( n2750 & n2884 ) | ( n2860 & n2884 ) ;
  assign n2886 = ( ~n2750 & n2860 ) | ( ~n2750 & n2884 ) | ( n2860 & n2884 ) ;
  assign n2887 = ( n2750 & ~n2885 ) | ( n2750 & n2886 ) | ( ~n2885 & n2886 ) ;
  assign n2888 = ( n2782 & n2837 ) | ( n2782 & n2887 ) | ( n2837 & n2887 ) ;
  assign n2889 = ( ~n2782 & n2837 ) | ( ~n2782 & n2887 ) | ( n2837 & n2887 ) ;
  assign n2890 = ( n2782 & ~n2888 ) | ( n2782 & n2889 ) | ( ~n2888 & n2889 ) ;
  assign n2891 = ( n2786 & n2788 ) | ( n2786 & n2890 ) | ( n2788 & n2890 ) ;
  assign n2892 = ( ~n2786 & n2788 ) | ( ~n2786 & n2890 ) | ( n2788 & n2890 ) ;
  assign n2893 = ( n2786 & ~n2891 ) | ( n2786 & n2892 ) | ( ~n2891 & n2892 ) ;
  assign n2894 = ( n2822 & ~n2842 ) | ( n2822 & n2865 ) | ( ~n2842 & n2865 ) ;
  assign n2895 = ( n2822 & n2842 ) | ( n2822 & n2865 ) | ( n2842 & n2865 ) ;
  assign n2896 = ( n2842 & n2894 ) | ( n2842 & ~n2895 ) | ( n2894 & ~n2895 ) ;
  assign n2897 = ( n2830 & n2867 ) | ( n2830 & n2896 ) | ( n2867 & n2896 ) ;
  assign n2898 = ( ~n2830 & n2867 ) | ( ~n2830 & n2896 ) | ( n2867 & n2896 ) ;
  assign n2899 = ( n2830 & ~n2897 ) | ( n2830 & n2898 ) | ( ~n2897 & n2898 ) ;
  assign n2900 = ( n2795 & ~n2807 ) | ( n2795 & n2827 ) | ( ~n2807 & n2827 ) ;
  assign n2901 = ( n2795 & n2807 ) | ( n2795 & n2827 ) | ( n2807 & n2827 ) ;
  assign n2902 = ( n2807 & n2900 ) | ( n2807 & ~n2901 ) | ( n2900 & ~n2901 ) ;
  assign n2903 = ~x1 & x27 ;
  assign n2904 = ( x1 & x27 ) | ( x1 & x52 ) | ( x27 & x52 ) ;
  assign n2905 = x27 & x52 ;
  assign n2906 = ( n2903 & n2904 ) | ( n2903 & ~n2905 ) | ( n2904 & ~n2905 ) ;
  assign n2907 = ( ~n2801 & n2816 ) | ( ~n2801 & n2906 ) | ( n2816 & n2906 ) ;
  assign n2908 = ( n2801 & n2816 ) | ( n2801 & n2906 ) | ( n2816 & n2906 ) ;
  assign n2909 = ( n2801 & n2907 ) | ( n2801 & ~n2908 ) | ( n2907 & ~n2908 ) ;
  assign n2910 = ( ~n2810 & n2902 ) | ( ~n2810 & n2909 ) | ( n2902 & n2909 ) ;
  assign n2911 = ( n2810 & n2902 ) | ( n2810 & n2909 ) | ( n2902 & n2909 ) ;
  assign n2912 = ( n2810 & n2910 ) | ( n2810 & ~n2911 ) | ( n2910 & ~n2911 ) ;
  assign n2913 = ( n2859 & n2899 ) | ( n2859 & n2912 ) | ( n2899 & n2912 ) ;
  assign n2914 = ( ~n2859 & n2899 ) | ( ~n2859 & n2912 ) | ( n2899 & n2912 ) ;
  assign n2915 = ( n2859 & ~n2913 ) | ( n2859 & n2914 ) | ( ~n2913 & n2914 ) ;
  assign n2916 = ( n2853 & ~n2874 ) | ( n2853 & n2877 ) | ( ~n2874 & n2877 ) ;
  assign n2917 = ( n2853 & n2874 ) | ( n2853 & n2877 ) | ( n2874 & n2877 ) ;
  assign n2918 = ( n2874 & n2916 ) | ( n2874 & ~n2917 ) | ( n2916 & ~n2917 ) ;
  assign n2919 = ( n2832 & n2870 ) | ( n2832 & n2918 ) | ( n2870 & n2918 ) ;
  assign n2920 = ( ~n2832 & n2870 ) | ( ~n2832 & n2918 ) | ( n2870 & n2918 ) ;
  assign n2921 = ( n2832 & ~n2919 ) | ( n2832 & n2920 ) | ( ~n2919 & n2920 ) ;
  assign n2922 = ( n2835 & n2915 ) | ( n2835 & n2921 ) | ( n2915 & n2921 ) ;
  assign n2923 = ( n2835 & ~n2915 ) | ( n2835 & n2921 ) | ( ~n2915 & n2921 ) ;
  assign n2924 = ( n2915 & ~n2922 ) | ( n2915 & n2923 ) | ( ~n2922 & n2923 ) ;
  assign n2925 = x3 & x50 ;
  assign n2926 = x2 & x51 ;
  assign n2927 = ( ~n2849 & n2925 ) | ( ~n2849 & n2926 ) | ( n2925 & n2926 ) ;
  assign n2928 = ( n2849 & n2925 ) | ( n2849 & n2926 ) | ( n2925 & n2926 ) ;
  assign n2929 = ( n2849 & n2927 ) | ( n2849 & ~n2928 ) | ( n2927 & ~n2928 ) ;
  assign n2930 = x19 & x34 ;
  assign n2931 = x21 & x32 ;
  assign n2932 = x20 & x33 ;
  assign n2933 = ( ~n2930 & n2931 ) | ( ~n2930 & n2932 ) | ( n2931 & n2932 ) ;
  assign n2934 = ( n2930 & n2931 ) | ( n2930 & n2932 ) | ( n2931 & n2932 ) ;
  assign n2935 = ( n2930 & n2933 ) | ( n2930 & ~n2934 ) | ( n2933 & ~n2934 ) ;
  assign n2936 = x4 & x49 ;
  assign n2937 = x17 & x36 ;
  assign n2938 = x18 & x35 ;
  assign n2939 = ( ~n2936 & n2937 ) | ( ~n2936 & n2938 ) | ( n2937 & n2938 ) ;
  assign n2940 = ( n2936 & n2937 ) | ( n2936 & n2938 ) | ( n2937 & n2938 ) ;
  assign n2941 = ( n2936 & n2939 ) | ( n2936 & ~n2940 ) | ( n2939 & ~n2940 ) ;
  assign n2942 = ( ~n2929 & n2935 ) | ( ~n2929 & n2941 ) | ( n2935 & n2941 ) ;
  assign n2943 = ( n2929 & n2935 ) | ( n2929 & n2941 ) | ( n2935 & n2941 ) ;
  assign n2944 = ( n2929 & n2942 ) | ( n2929 & ~n2943 ) | ( n2942 & ~n2943 ) ;
  assign n2945 = x8 & x45 ;
  assign n2946 = x14 & x39 ;
  assign n2947 = x9 & x44 ;
  assign n2948 = ( ~n2945 & n2946 ) | ( ~n2945 & n2947 ) | ( n2946 & n2947 ) ;
  assign n2949 = ( n2945 & n2946 ) | ( n2945 & n2947 ) | ( n2946 & n2947 ) ;
  assign n2950 = ( n2945 & n2948 ) | ( n2945 & ~n2949 ) | ( n2948 & ~n2949 ) ;
  assign n2951 = x6 & x47 ;
  assign n2952 = x15 & x38 ;
  assign n2953 = x7 & x46 ;
  assign n2954 = ( ~n2951 & n2952 ) | ( ~n2951 & n2953 ) | ( n2952 & n2953 ) ;
  assign n2955 = ( n2951 & n2952 ) | ( n2951 & n2953 ) | ( n2952 & n2953 ) ;
  assign n2956 = ( n2951 & n2954 ) | ( n2951 & ~n2955 ) | ( n2954 & ~n2955 ) ;
  assign n2957 = x0 & x53 ;
  assign n2958 = x5 & x48 ;
  assign n2959 = x16 & x37 ;
  assign n2960 = ( ~n2957 & n2958 ) | ( ~n2957 & n2959 ) | ( n2958 & n2959 ) ;
  assign n2961 = ( n2957 & n2958 ) | ( n2957 & n2959 ) | ( n2958 & n2959 ) ;
  assign n2962 = ( n2957 & n2960 ) | ( n2957 & ~n2961 ) | ( n2960 & ~n2961 ) ;
  assign n2963 = ( n2950 & n2956 ) | ( n2950 & n2962 ) | ( n2956 & n2962 ) ;
  assign n2964 = ( ~n2950 & n2956 ) | ( ~n2950 & n2962 ) | ( n2956 & n2962 ) ;
  assign n2965 = ( n2950 & ~n2963 ) | ( n2950 & n2964 ) | ( ~n2963 & n2964 ) ;
  assign n2966 = ( ~n2845 & n2944 ) | ( ~n2845 & n2965 ) | ( n2944 & n2965 ) ;
  assign n2967 = ( n2845 & n2944 ) | ( n2845 & n2965 ) | ( n2944 & n2965 ) ;
  assign n2968 = ( n2845 & n2966 ) | ( n2845 & ~n2967 ) | ( n2966 & ~n2967 ) ;
  assign n2969 = x11 & x42 ;
  assign n2970 = x26 & x27 ;
  assign n2971 = x25 & x28 ;
  assign n2972 = ( ~n2969 & n2970 ) | ( ~n2969 & n2971 ) | ( n2970 & n2971 ) ;
  assign n2973 = ( n2969 & n2970 ) | ( n2969 & n2971 ) | ( n2970 & n2971 ) ;
  assign n2974 = ( n2969 & n2972 ) | ( n2969 & ~n2973 ) | ( n2972 & ~n2973 ) ;
  assign n2975 = x22 & x31 ;
  assign n2976 = x24 & x29 ;
  assign n2977 = x23 & x30 ;
  assign n2978 = ( ~n2975 & n2976 ) | ( ~n2975 & n2977 ) | ( n2976 & n2977 ) ;
  assign n2979 = ( n2975 & n2976 ) | ( n2975 & n2977 ) | ( n2976 & n2977 ) ;
  assign n2980 = ( n2975 & n2978 ) | ( n2975 & ~n2979 ) | ( n2978 & ~n2979 ) ;
  assign n2981 = x13 & x40 ;
  assign n2982 = x12 & x41 ;
  assign n2983 = x10 & x43 ;
  assign n2984 = ( ~n2981 & n2982 ) | ( ~n2981 & n2983 ) | ( n2982 & n2983 ) ;
  assign n2985 = ( n2981 & n2982 ) | ( n2981 & n2983 ) | ( n2982 & n2983 ) ;
  assign n2986 = ( n2981 & n2984 ) | ( n2981 & ~n2985 ) | ( n2984 & ~n2985 ) ;
  assign n2987 = ( ~n2974 & n2980 ) | ( ~n2974 & n2986 ) | ( n2980 & n2986 ) ;
  assign n2988 = ( n2974 & n2980 ) | ( n2974 & n2986 ) | ( n2980 & n2986 ) ;
  assign n2989 = ( n2974 & n2987 ) | ( n2974 & ~n2988 ) | ( n2987 & ~n2988 ) ;
  assign n2990 = ( n2856 & n2880 ) | ( n2856 & n2989 ) | ( n2880 & n2989 ) ;
  assign n2991 = ( ~n2856 & n2880 ) | ( ~n2856 & n2989 ) | ( n2880 & n2989 ) ;
  assign n2992 = ( n2856 & ~n2990 ) | ( n2856 & n2991 ) | ( ~n2990 & n2991 ) ;
  assign n2993 = ( n2883 & n2968 ) | ( n2883 & n2992 ) | ( n2968 & n2992 ) ;
  assign n2994 = ( ~n2883 & n2968 ) | ( ~n2883 & n2992 ) | ( n2968 & n2992 ) ;
  assign n2995 = ( n2883 & ~n2993 ) | ( n2883 & n2994 ) | ( ~n2993 & n2994 ) ;
  assign n2996 = ( n2885 & n2924 ) | ( n2885 & n2995 ) | ( n2924 & n2995 ) ;
  assign n2997 = ( ~n2885 & n2924 ) | ( ~n2885 & n2995 ) | ( n2924 & n2995 ) ;
  assign n2998 = ( n2885 & ~n2996 ) | ( n2885 & n2997 ) | ( ~n2996 & n2997 ) ;
  assign n2999 = ( ~n2888 & n2891 ) | ( ~n2888 & n2998 ) | ( n2891 & n2998 ) ;
  assign n3000 = ( n2888 & n2891 ) | ( n2888 & n2998 ) | ( n2891 & n2998 ) ;
  assign n3001 = ( n2888 & n2999 ) | ( n2888 & ~n3000 ) | ( n2999 & ~n3000 ) ;
  assign n3002 = x52 & n872 ;
  assign n3003 = x26 & x28 ;
  assign n3004 = x1 & x53 ;
  assign n3005 = n3003 & n3004 ;
  assign n3006 = n3003 | n3004 ;
  assign n3007 = ~n3005 & n3006 ;
  assign n3008 = x0 & x54 ;
  assign n3009 = ( n3002 & n3007 ) | ( n3002 & n3008 ) | ( n3007 & n3008 ) ;
  assign n3010 = ( ~n3002 & n3007 ) | ( ~n3002 & n3008 ) | ( n3007 & n3008 ) ;
  assign n3011 = ( n3002 & ~n3009 ) | ( n3002 & n3010 ) | ( ~n3009 & n3010 ) ;
  assign n3012 = x23 & x31 ;
  assign n3013 = x24 & x30 ;
  assign n3014 = x25 & x29 ;
  assign n3015 = ( ~n3012 & n3013 ) | ( ~n3012 & n3014 ) | ( n3013 & n3014 ) ;
  assign n3016 = ( n3012 & n3013 ) | ( n3012 & n3014 ) | ( n3013 & n3014 ) ;
  assign n3017 = ( n3012 & n3015 ) | ( n3012 & ~n3016 ) | ( n3015 & ~n3016 ) ;
  assign n3018 = x19 & x35 ;
  assign n3019 = x21 & x33 ;
  assign n3020 = x22 & x32 ;
  assign n3021 = ( ~n3018 & n3019 ) | ( ~n3018 & n3020 ) | ( n3019 & n3020 ) ;
  assign n3022 = ( n3018 & n3019 ) | ( n3018 & n3020 ) | ( n3019 & n3020 ) ;
  assign n3023 = ( n3018 & n3021 ) | ( n3018 & ~n3022 ) | ( n3021 & ~n3022 ) ;
  assign n3024 = ( n3011 & n3017 ) | ( n3011 & n3023 ) | ( n3017 & n3023 ) ;
  assign n3025 = ( ~n3011 & n3017 ) | ( ~n3011 & n3023 ) | ( n3017 & n3023 ) ;
  assign n3026 = ( n3011 & ~n3024 ) | ( n3011 & n3025 ) | ( ~n3024 & n3025 ) ;
  assign n3027 = ( ~n2897 & n2911 ) | ( ~n2897 & n3026 ) | ( n2911 & n3026 ) ;
  assign n3028 = ( n2897 & n2911 ) | ( n2897 & n3026 ) | ( n2911 & n3026 ) ;
  assign n3029 = ( n2897 & n3027 ) | ( n2897 & ~n3028 ) | ( n3027 & ~n3028 ) ;
  assign n3030 = ( n2913 & n2919 ) | ( n2913 & n3029 ) | ( n2919 & n3029 ) ;
  assign n3031 = ( ~n2913 & n2919 ) | ( ~n2913 & n3029 ) | ( n2919 & n3029 ) ;
  assign n3032 = ( n2913 & ~n3030 ) | ( n2913 & n3031 ) | ( ~n3030 & n3031 ) ;
  assign n3033 = ( ~n2895 & n2901 ) | ( ~n2895 & n2908 ) | ( n2901 & n2908 ) ;
  assign n3034 = ( n2895 & n2901 ) | ( n2895 & n2908 ) | ( n2901 & n2908 ) ;
  assign n3035 = ( n2895 & n3033 ) | ( n2895 & ~n3034 ) | ( n3033 & ~n3034 ) ;
  assign n3036 = ( ~n2955 & n2961 ) | ( ~n2955 & n2973 ) | ( n2961 & n2973 ) ;
  assign n3037 = ( n2955 & n2961 ) | ( n2955 & n2973 ) | ( n2961 & n2973 ) ;
  assign n3038 = ( n2955 & n3036 ) | ( n2955 & ~n3037 ) | ( n3036 & ~n3037 ) ;
  assign n3039 = ( ~n2934 & n2940 ) | ( ~n2934 & n2979 ) | ( n2940 & n2979 ) ;
  assign n3040 = ( n2934 & n2940 ) | ( n2934 & n2979 ) | ( n2940 & n2979 ) ;
  assign n3041 = ( n2934 & n3039 ) | ( n2934 & ~n3040 ) | ( n3039 & ~n3040 ) ;
  assign n3042 = ( n2963 & n3038 ) | ( n2963 & n3041 ) | ( n3038 & n3041 ) ;
  assign n3043 = ( ~n2963 & n3038 ) | ( ~n2963 & n3041 ) | ( n3038 & n3041 ) ;
  assign n3044 = ( n2963 & ~n3042 ) | ( n2963 & n3043 ) | ( ~n3042 & n3043 ) ;
  assign n3045 = ( ~n2967 & n3035 ) | ( ~n2967 & n3044 ) | ( n3035 & n3044 ) ;
  assign n3046 = ( n2967 & n3035 ) | ( n2967 & n3044 ) | ( n3035 & n3044 ) ;
  assign n3047 = ( n2967 & n3045 ) | ( n2967 & ~n3046 ) | ( n3045 & ~n3046 ) ;
  assign n3048 = x17 & x37 ;
  assign n3049 = x6 & x48 ;
  assign n3050 = x16 & x38 ;
  assign n3051 = ( ~n3048 & n3049 ) | ( ~n3048 & n3050 ) | ( n3049 & n3050 ) ;
  assign n3052 = ( n3048 & n3049 ) | ( n3048 & n3050 ) | ( n3049 & n3050 ) ;
  assign n3053 = ( n3048 & n3051 ) | ( n3048 & ~n3052 ) | ( n3051 & ~n3052 ) ;
  assign n3054 = x18 & x36 ;
  assign n3055 = x20 & x34 ;
  assign n3056 = x5 & x49 ;
  assign n3057 = ( ~n3054 & n3055 ) | ( ~n3054 & n3056 ) | ( n3055 & n3056 ) ;
  assign n3058 = ( n3054 & n3055 ) | ( n3054 & n3056 ) | ( n3055 & n3056 ) ;
  assign n3059 = ( n3054 & n3057 ) | ( n3054 & ~n3058 ) | ( n3057 & ~n3058 ) ;
  assign n3060 = x13 & x41 ;
  assign n3061 = x11 & x43 ;
  assign n3062 = x12 & x42 ;
  assign n3063 = ( ~n3060 & n3061 ) | ( ~n3060 & n3062 ) | ( n3061 & n3062 ) ;
  assign n3064 = ( n3060 & n3061 ) | ( n3060 & n3062 ) | ( n3061 & n3062 ) ;
  assign n3065 = ( n3060 & n3063 ) | ( n3060 & ~n3064 ) | ( n3063 & ~n3064 ) ;
  assign n3066 = ( ~n3053 & n3059 ) | ( ~n3053 & n3065 ) | ( n3059 & n3065 ) ;
  assign n3067 = ( n3053 & n3059 ) | ( n3053 & n3065 ) | ( n3059 & n3065 ) ;
  assign n3068 = ( n3053 & n3066 ) | ( n3053 & ~n3067 ) | ( n3066 & ~n3067 ) ;
  assign n3069 = x9 & x45 ;
  assign n3070 = x14 & x40 ;
  assign n3071 = x10 & x44 ;
  assign n3072 = ( ~n3069 & n3070 ) | ( ~n3069 & n3071 ) | ( n3070 & n3071 ) ;
  assign n3073 = ( n3069 & n3070 ) | ( n3069 & n3071 ) | ( n3070 & n3071 ) ;
  assign n3074 = ( n3069 & n3072 ) | ( n3069 & ~n3073 ) | ( n3072 & ~n3073 ) ;
  assign n3075 = x7 & x47 ;
  assign n3076 = x15 & x39 ;
  assign n3077 = x8 & x46 ;
  assign n3078 = ( ~n3075 & n3076 ) | ( ~n3075 & n3077 ) | ( n3076 & n3077 ) ;
  assign n3079 = ( n3075 & n3076 ) | ( n3075 & n3077 ) | ( n3076 & n3077 ) ;
  assign n3080 = ( n3075 & n3078 ) | ( n3075 & ~n3079 ) | ( n3078 & ~n3079 ) ;
  assign n3081 = x2 & x52 ;
  assign n3082 = x3 & x51 ;
  assign n3083 = x4 & x50 ;
  assign n3084 = ( ~n3081 & n3082 ) | ( ~n3081 & n3083 ) | ( n3082 & n3083 ) ;
  assign n3085 = ( n3081 & n3082 ) | ( n3081 & n3083 ) | ( n3082 & n3083 ) ;
  assign n3086 = ( n3081 & n3084 ) | ( n3081 & ~n3085 ) | ( n3084 & ~n3085 ) ;
  assign n3087 = ( ~n3074 & n3080 ) | ( ~n3074 & n3086 ) | ( n3080 & n3086 ) ;
  assign n3088 = ( n3074 & n3080 ) | ( n3074 & n3086 ) | ( n3080 & n3086 ) ;
  assign n3089 = ( n3074 & n3087 ) | ( n3074 & ~n3088 ) | ( n3087 & ~n3088 ) ;
  assign n3090 = ( n2917 & n3068 ) | ( n2917 & n3089 ) | ( n3068 & n3089 ) ;
  assign n3091 = ( ~n2917 & n3068 ) | ( ~n2917 & n3089 ) | ( n3068 & n3089 ) ;
  assign n3092 = ( n2917 & ~n3090 ) | ( n2917 & n3091 ) | ( ~n3090 & n3091 ) ;
  assign n3093 = ( n2928 & n2949 ) | ( n2928 & n2985 ) | ( n2949 & n2985 ) ;
  assign n3094 = ( ~n2928 & n2949 ) | ( ~n2928 & n2985 ) | ( n2949 & n2985 ) ;
  assign n3095 = ( n2928 & ~n3093 ) | ( n2928 & n3094 ) | ( ~n3093 & n3094 ) ;
  assign n3096 = ( n2943 & n2988 ) | ( n2943 & n3095 ) | ( n2988 & n3095 ) ;
  assign n3097 = ( n2943 & n2988 ) | ( n2943 & ~n3095 ) | ( n2988 & ~n3095 ) ;
  assign n3098 = ( n3095 & ~n3096 ) | ( n3095 & n3097 ) | ( ~n3096 & n3097 ) ;
  assign n3099 = ( ~n2990 & n3092 ) | ( ~n2990 & n3098 ) | ( n3092 & n3098 ) ;
  assign n3100 = ( n2990 & n3092 ) | ( n2990 & n3098 ) | ( n3092 & n3098 ) ;
  assign n3101 = ( n2990 & n3099 ) | ( n2990 & ~n3100 ) | ( n3099 & ~n3100 ) ;
  assign n3102 = ( n2993 & n3047 ) | ( n2993 & n3101 ) | ( n3047 & n3101 ) ;
  assign n3103 = ( ~n2993 & n3047 ) | ( ~n2993 & n3101 ) | ( n3047 & n3101 ) ;
  assign n3104 = ( n2993 & ~n3102 ) | ( n2993 & n3103 ) | ( ~n3102 & n3103 ) ;
  assign n3105 = ( ~n2922 & n3032 ) | ( ~n2922 & n3104 ) | ( n3032 & n3104 ) ;
  assign n3106 = ( n2922 & n3032 ) | ( n2922 & n3104 ) | ( n3032 & n3104 ) ;
  assign n3107 = ( n2922 & n3105 ) | ( n2922 & ~n3106 ) | ( n3105 & ~n3106 ) ;
  assign n3108 = ( n2996 & n3000 ) | ( n2996 & n3107 ) | ( n3000 & n3107 ) ;
  assign n3109 = ( ~n2996 & n3000 ) | ( ~n2996 & n3107 ) | ( n3000 & n3107 ) ;
  assign n3110 = ( n2996 & ~n3108 ) | ( n2996 & n3109 ) | ( ~n3108 & n3109 ) ;
  assign n3111 = ~x54 & n3005 ;
  assign n3112 = n3064 & n3111 ;
  assign n3113 = x1 & x54 ;
  assign n3114 = x28 | n3113 ;
  assign n3115 = x28 & x54 ;
  assign n3116 = x1 & n3115 ;
  assign n3117 = ( n3005 & n3114 ) | ( n3005 & ~n3116 ) | ( n3114 & ~n3116 ) ;
  assign n3118 = ( n3064 & n3111 ) | ( n3064 & n3117 ) | ( n3111 & n3117 ) ;
  assign n3119 = n3064 | n3117 ;
  assign n3120 = ( n3112 & ~n3118 ) | ( n3112 & n3119 ) | ( ~n3118 & n3119 ) ;
  assign n3121 = ( n3037 & n3093 ) | ( n3037 & n3120 ) | ( n3093 & n3120 ) ;
  assign n3122 = ( n3037 & ~n3093 ) | ( n3037 & n3120 ) | ( ~n3093 & n3120 ) ;
  assign n3123 = ( n3093 & ~n3121 ) | ( n3093 & n3122 ) | ( ~n3121 & n3122 ) ;
  assign n3124 = ( n3058 & ~n3073 ) | ( n3058 & n3085 ) | ( ~n3073 & n3085 ) ;
  assign n3125 = ( n3058 & n3073 ) | ( n3058 & n3085 ) | ( n3073 & n3085 ) ;
  assign n3126 = ( n3073 & n3124 ) | ( n3073 & ~n3125 ) | ( n3124 & ~n3125 ) ;
  assign n3127 = x5 & x50 ;
  assign n3128 = x19 & x36 ;
  assign n3129 = x18 & x37 ;
  assign n3130 = ( ~n3127 & n3128 ) | ( ~n3127 & n3129 ) | ( n3128 & n3129 ) ;
  assign n3131 = ( n3127 & n3128 ) | ( n3127 & n3129 ) | ( n3128 & n3129 ) ;
  assign n3132 = ( n3127 & n3130 ) | ( n3127 & ~n3131 ) | ( n3130 & ~n3131 ) ;
  assign n3133 = ( n3009 & n3079 ) | ( n3009 & n3132 ) | ( n3079 & n3132 ) ;
  assign n3134 = ( ~n3009 & n3079 ) | ( ~n3009 & n3132 ) | ( n3079 & n3132 ) ;
  assign n3135 = ( n3009 & ~n3133 ) | ( n3009 & n3134 ) | ( ~n3133 & n3134 ) ;
  assign n3136 = ( ~n3024 & n3126 ) | ( ~n3024 & n3135 ) | ( n3126 & n3135 ) ;
  assign n3137 = ( n3024 & n3126 ) | ( n3024 & n3135 ) | ( n3126 & n3135 ) ;
  assign n3138 = ( n3024 & n3136 ) | ( n3024 & ~n3137 ) | ( n3136 & ~n3137 ) ;
  assign n3139 = ( n3090 & n3123 ) | ( n3090 & n3138 ) | ( n3123 & n3138 ) ;
  assign n3140 = ( ~n3090 & n3123 ) | ( ~n3090 & n3138 ) | ( n3123 & n3138 ) ;
  assign n3141 = ( n3090 & ~n3139 ) | ( n3090 & n3140 ) | ( ~n3139 & n3140 ) ;
  assign n3142 = x16 & x39 ;
  assign n3143 = x7 & x48 ;
  assign n3144 = x8 & x47 ;
  assign n3145 = ( ~n3142 & n3143 ) | ( ~n3142 & n3144 ) | ( n3143 & n3144 ) ;
  assign n3146 = ( n3142 & n3143 ) | ( n3142 & n3144 ) | ( n3143 & n3144 ) ;
  assign n3147 = ( n3142 & n3145 ) | ( n3142 & ~n3146 ) | ( n3145 & ~n3146 ) ;
  assign n3148 = x12 & x43 ;
  assign n3149 = x27 & x28 ;
  assign n3150 = x26 & x29 ;
  assign n3151 = ( ~n3148 & n3149 ) | ( ~n3148 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3152 = ( n3148 & n3149 ) | ( n3148 & n3150 ) | ( n3149 & n3150 ) ;
  assign n3153 = ( n3148 & n3151 ) | ( n3148 & ~n3152 ) | ( n3151 & ~n3152 ) ;
  assign n3154 = x10 & x45 ;
  assign n3155 = x13 & x42 ;
  assign n3156 = x11 & x44 ;
  assign n3157 = ( ~n3154 & n3155 ) | ( ~n3154 & n3156 ) | ( n3155 & n3156 ) ;
  assign n3158 = ( n3154 & n3155 ) | ( n3154 & n3156 ) | ( n3155 & n3156 ) ;
  assign n3159 = ( n3154 & n3157 ) | ( n3154 & ~n3158 ) | ( n3157 & ~n3158 ) ;
  assign n3160 = ( ~n3147 & n3153 ) | ( ~n3147 & n3159 ) | ( n3153 & n3159 ) ;
  assign n3161 = ( n3147 & n3153 ) | ( n3147 & n3159 ) | ( n3153 & n3159 ) ;
  assign n3162 = ( n3147 & n3160 ) | ( n3147 & ~n3161 ) | ( n3160 & ~n3161 ) ;
  assign n3163 = x0 & x55 ;
  assign n3164 = x4 & x51 ;
  assign n3165 = x2 & x53 ;
  assign n3166 = ( ~n3163 & n3164 ) | ( ~n3163 & n3165 ) | ( n3164 & n3165 ) ;
  assign n3167 = ( n3163 & n3164 ) | ( n3163 & n3165 ) | ( n3164 & n3165 ) ;
  assign n3168 = ( n3163 & n3166 ) | ( n3163 & ~n3167 ) | ( n3166 & ~n3167 ) ;
  assign n3169 = x23 & x32 ;
  assign n3170 = x25 & x30 ;
  assign n3171 = x24 & x31 ;
  assign n3172 = ( ~n3169 & n3170 ) | ( ~n3169 & n3171 ) | ( n3170 & n3171 ) ;
  assign n3173 = ( n3169 & n3170 ) | ( n3169 & n3171 ) | ( n3170 & n3171 ) ;
  assign n3174 = ( n3169 & n3172 ) | ( n3169 & ~n3173 ) | ( n3172 & ~n3173 ) ;
  assign n3175 = x20 & x35 ;
  assign n3176 = x22 & x33 ;
  assign n3177 = x21 & x34 ;
  assign n3178 = ( ~n3175 & n3176 ) | ( ~n3175 & n3177 ) | ( n3176 & n3177 ) ;
  assign n3179 = ( n3175 & n3176 ) | ( n3175 & n3177 ) | ( n3176 & n3177 ) ;
  assign n3180 = ( n3175 & n3178 ) | ( n3175 & ~n3179 ) | ( n3178 & ~n3179 ) ;
  assign n3181 = ( ~n3168 & n3174 ) | ( ~n3168 & n3180 ) | ( n3174 & n3180 ) ;
  assign n3182 = ( n3168 & n3174 ) | ( n3168 & n3180 ) | ( n3174 & n3180 ) ;
  assign n3183 = ( n3168 & n3181 ) | ( n3168 & ~n3182 ) | ( n3181 & ~n3182 ) ;
  assign n3184 = ( n3034 & n3162 ) | ( n3034 & n3183 ) | ( n3162 & n3183 ) ;
  assign n3185 = ( ~n3034 & n3162 ) | ( ~n3034 & n3183 ) | ( n3162 & n3183 ) ;
  assign n3186 = ( n3034 & ~n3184 ) | ( n3034 & n3185 ) | ( ~n3184 & n3185 ) ;
  assign n3187 = ( n3016 & ~n3022 ) | ( n3016 & n3052 ) | ( ~n3022 & n3052 ) ;
  assign n3188 = ( n3016 & n3022 ) | ( n3016 & n3052 ) | ( n3022 & n3052 ) ;
  assign n3189 = ( n3022 & n3187 ) | ( n3022 & ~n3188 ) | ( n3187 & ~n3188 ) ;
  assign n3190 = ( n3067 & n3088 ) | ( n3067 & n3189 ) | ( n3088 & n3189 ) ;
  assign n3191 = ( ~n3067 & n3088 ) | ( ~n3067 & n3189 ) | ( n3088 & n3189 ) ;
  assign n3192 = ( n3067 & ~n3190 ) | ( n3067 & n3191 ) | ( ~n3190 & n3191 ) ;
  assign n3193 = ( n3028 & n3186 ) | ( n3028 & n3192 ) | ( n3186 & n3192 ) ;
  assign n3194 = ( ~n3028 & n3186 ) | ( ~n3028 & n3192 ) | ( n3186 & n3192 ) ;
  assign n3195 = ( n3028 & ~n3193 ) | ( n3028 & n3194 ) | ( ~n3193 & n3194 ) ;
  assign n3196 = ( ~n3030 & n3141 ) | ( ~n3030 & n3195 ) | ( n3141 & n3195 ) ;
  assign n3197 = ( n3030 & n3141 ) | ( n3030 & n3195 ) | ( n3141 & n3195 ) ;
  assign n3198 = ( n3030 & n3196 ) | ( n3030 & ~n3197 ) | ( n3196 & ~n3197 ) ;
  assign n3199 = x14 & x41 ;
  assign n3200 = x15 & x40 ;
  assign n3201 = x9 & x46 ;
  assign n3202 = ( ~n3199 & n3200 ) | ( ~n3199 & n3201 ) | ( n3200 & n3201 ) ;
  assign n3203 = ( n3199 & n3200 ) | ( n3199 & n3201 ) | ( n3200 & n3201 ) ;
  assign n3204 = ( n3199 & n3202 ) | ( n3199 & ~n3203 ) | ( n3202 & ~n3203 ) ;
  assign n3205 = x3 & x52 ;
  assign n3206 = x6 & x49 ;
  assign n3207 = x17 & x38 ;
  assign n3208 = ( ~n3205 & n3206 ) | ( ~n3205 & n3207 ) | ( n3206 & n3207 ) ;
  assign n3209 = ( n3205 & n3206 ) | ( n3205 & n3207 ) | ( n3206 & n3207 ) ;
  assign n3210 = ( n3205 & n3208 ) | ( n3205 & ~n3209 ) | ( n3208 & ~n3209 ) ;
  assign n3211 = ( n3040 & n3204 ) | ( n3040 & n3210 ) | ( n3204 & n3210 ) ;
  assign n3212 = ( ~n3040 & n3204 ) | ( ~n3040 & n3210 ) | ( n3204 & n3210 ) ;
  assign n3213 = ( n3040 & ~n3211 ) | ( n3040 & n3212 ) | ( ~n3211 & n3212 ) ;
  assign n3214 = ( ~n3042 & n3096 ) | ( ~n3042 & n3213 ) | ( n3096 & n3213 ) ;
  assign n3215 = ( n3042 & n3096 ) | ( n3042 & n3213 ) | ( n3096 & n3213 ) ;
  assign n3216 = ( n3042 & n3214 ) | ( n3042 & ~n3215 ) | ( n3214 & ~n3215 ) ;
  assign n3217 = ( ~n3046 & n3100 ) | ( ~n3046 & n3216 ) | ( n3100 & n3216 ) ;
  assign n3218 = ( n3046 & n3100 ) | ( n3046 & n3216 ) | ( n3100 & n3216 ) ;
  assign n3219 = ( n3046 & n3217 ) | ( n3046 & ~n3218 ) | ( n3217 & ~n3218 ) ;
  assign n3220 = ( n3102 & n3198 ) | ( n3102 & n3219 ) | ( n3198 & n3219 ) ;
  assign n3221 = ( ~n3102 & n3198 ) | ( ~n3102 & n3219 ) | ( n3198 & n3219 ) ;
  assign n3222 = ( n3102 & ~n3220 ) | ( n3102 & n3221 ) | ( ~n3220 & n3221 ) ;
  assign n3223 = ( ~n3106 & n3108 ) | ( ~n3106 & n3222 ) | ( n3108 & n3222 ) ;
  assign n3224 = ( n3106 & n3108 ) | ( n3106 & n3222 ) | ( n3108 & n3222 ) ;
  assign n3225 = ( n3106 & n3223 ) | ( n3106 & ~n3224 ) | ( n3223 & ~n3224 ) ;
  assign n3226 = x11 & x45 ;
  assign n3227 = x13 & x43 ;
  assign n3228 = x12 & x44 ;
  assign n3229 = ( ~n3226 & n3227 ) | ( ~n3226 & n3228 ) | ( n3227 & n3228 ) ;
  assign n3230 = ( n3226 & n3227 ) | ( n3226 & n3228 ) | ( n3227 & n3228 ) ;
  assign n3231 = ( n3226 & n3229 ) | ( n3226 & ~n3230 ) | ( n3229 & ~n3230 ) ;
  assign n3232 = x6 & x50 ;
  assign n3233 = x7 & x49 ;
  assign n3234 = x17 & x39 ;
  assign n3235 = ( ~n3232 & n3233 ) | ( ~n3232 & n3234 ) | ( n3233 & n3234 ) ;
  assign n3236 = ( n3232 & n3233 ) | ( n3232 & n3234 ) | ( n3233 & n3234 ) ;
  assign n3237 = ( n3232 & n3235 ) | ( n3232 & ~n3236 ) | ( n3235 & ~n3236 ) ;
  assign n3238 = x16 & x40 ;
  assign n3239 = x15 & x41 ;
  assign n3240 = x8 & x48 ;
  assign n3241 = ( ~n3238 & n3239 ) | ( ~n3238 & n3240 ) | ( n3239 & n3240 ) ;
  assign n3242 = ( n3238 & n3239 ) | ( n3238 & n3240 ) | ( n3239 & n3240 ) ;
  assign n3243 = ( n3238 & n3241 ) | ( n3238 & ~n3242 ) | ( n3241 & ~n3242 ) ;
  assign n3244 = ( n3231 & n3237 ) | ( n3231 & n3243 ) | ( n3237 & n3243 ) ;
  assign n3245 = ( ~n3231 & n3237 ) | ( ~n3231 & n3243 ) | ( n3237 & n3243 ) ;
  assign n3246 = ( n3231 & ~n3244 ) | ( n3231 & n3245 ) | ( ~n3244 & n3245 ) ;
  assign n3247 = x24 & x32 ;
  assign n3248 = x25 & x31 ;
  assign n3249 = x26 & x30 ;
  assign n3250 = ( ~n3247 & n3248 ) | ( ~n3247 & n3249 ) | ( n3248 & n3249 ) ;
  assign n3251 = ( n3247 & n3248 ) | ( n3247 & n3249 ) | ( n3248 & n3249 ) ;
  assign n3252 = ( n3247 & n3250 ) | ( n3247 & ~n3251 ) | ( n3250 & ~n3251 ) ;
  assign n3253 = x9 & x47 ;
  assign n3254 = x14 & x42 ;
  assign n3255 = x10 & x46 ;
  assign n3256 = ( ~n3253 & n3254 ) | ( ~n3253 & n3255 ) | ( n3254 & n3255 ) ;
  assign n3257 = ( n3253 & n3254 ) | ( n3253 & n3255 ) | ( n3254 & n3255 ) ;
  assign n3258 = ( n3253 & n3256 ) | ( n3253 & ~n3257 ) | ( n3256 & ~n3257 ) ;
  assign n3259 = x20 & x36 ;
  assign n3260 = x22 & x34 ;
  assign n3261 = x23 & x33 ;
  assign n3262 = ( ~n3259 & n3260 ) | ( ~n3259 & n3261 ) | ( n3260 & n3261 ) ;
  assign n3263 = ( n3259 & n3260 ) | ( n3259 & n3261 ) | ( n3260 & n3261 ) ;
  assign n3264 = ( n3259 & n3262 ) | ( n3259 & ~n3263 ) | ( n3262 & ~n3263 ) ;
  assign n3265 = ( ~n3252 & n3258 ) | ( ~n3252 & n3264 ) | ( n3258 & n3264 ) ;
  assign n3266 = ( n3252 & n3258 ) | ( n3252 & n3264 ) | ( n3258 & n3264 ) ;
  assign n3267 = ( n3252 & n3265 ) | ( n3252 & ~n3266 ) | ( n3265 & ~n3266 ) ;
  assign n3268 = x0 & x56 ;
  assign n3269 = x2 & x54 ;
  assign n3270 = n3268 | n3269 ;
  assign n3271 = x2 & x56 ;
  assign n3272 = n3008 & n3271 ;
  assign n3273 = ( n3116 & n3270 ) | ( n3116 & n3272 ) | ( n3270 & n3272 ) ;
  assign n3274 = ( ~n3116 & n3270 ) | ( ~n3116 & n3272 ) | ( n3270 & n3272 ) ;
  assign n3275 = ( n3116 & ~n3273 ) | ( n3116 & n3274 ) | ( ~n3273 & n3274 ) ;
  assign n3276 = x19 & x37 ;
  assign n3277 = x3 & x53 ;
  assign n3278 = x4 & x52 ;
  assign n3279 = ( ~n3276 & n3277 ) | ( ~n3276 & n3278 ) | ( n3277 & n3278 ) ;
  assign n3280 = ( n3276 & n3277 ) | ( n3276 & n3278 ) | ( n3277 & n3278 ) ;
  assign n3281 = ( n3276 & n3279 ) | ( n3276 & ~n3280 ) | ( n3279 & ~n3280 ) ;
  assign n3282 = ( ~n3146 & n3275 ) | ( ~n3146 & n3281 ) | ( n3275 & n3281 ) ;
  assign n3283 = ( n3146 & n3275 ) | ( n3146 & n3281 ) | ( n3275 & n3281 ) ;
  assign n3284 = ( n3146 & n3282 ) | ( n3146 & ~n3283 ) | ( n3282 & ~n3283 ) ;
  assign n3285 = ( n3246 & n3267 ) | ( n3246 & n3284 ) | ( n3267 & n3284 ) ;
  assign n3286 = ( ~n3246 & n3267 ) | ( ~n3246 & n3284 ) | ( n3267 & n3284 ) ;
  assign n3287 = ( n3246 & ~n3285 ) | ( n3246 & n3286 ) | ( ~n3285 & n3286 ) ;
  assign n3288 = ( n3173 & n3179 ) | ( n3173 & n3209 ) | ( n3179 & n3209 ) ;
  assign n3289 = ( n3173 & ~n3179 ) | ( n3173 & n3209 ) | ( ~n3179 & n3209 ) ;
  assign n3290 = ( n3179 & ~n3288 ) | ( n3179 & n3289 ) | ( ~n3288 & n3289 ) ;
  assign n3291 = x27 & x29 ;
  assign n3292 = x1 & x55 ;
  assign n3293 = n3291 & n3292 ;
  assign n3294 = n3291 | n3292 ;
  assign n3295 = ~n3293 & n3294 ;
  assign n3296 = ( n3152 & n3158 ) | ( n3152 & n3295 ) | ( n3158 & n3295 ) ;
  assign n3297 = ( ~n3152 & n3158 ) | ( ~n3152 & n3295 ) | ( n3158 & n3295 ) ;
  assign n3298 = ( n3152 & ~n3296 ) | ( n3152 & n3297 ) | ( ~n3296 & n3297 ) ;
  assign n3299 = ( n3161 & n3290 ) | ( n3161 & n3298 ) | ( n3290 & n3298 ) ;
  assign n3300 = ( n3161 & ~n3290 ) | ( n3161 & n3298 ) | ( ~n3290 & n3298 ) ;
  assign n3301 = ( n3290 & ~n3299 ) | ( n3290 & n3300 ) | ( ~n3299 & n3300 ) ;
  assign n3302 = ( ~n3215 & n3287 ) | ( ~n3215 & n3301 ) | ( n3287 & n3301 ) ;
  assign n3303 = ( n3215 & n3287 ) | ( n3215 & n3301 ) | ( n3287 & n3301 ) ;
  assign n3304 = ( n3215 & n3302 ) | ( n3215 & ~n3303 ) | ( n3302 & ~n3303 ) ;
  assign n3305 = ( n3131 & ~n3167 ) | ( n3131 & n3203 ) | ( ~n3167 & n3203 ) ;
  assign n3306 = ( n3131 & n3167 ) | ( n3131 & n3203 ) | ( n3167 & n3203 ) ;
  assign n3307 = ( n3167 & n3305 ) | ( n3167 & ~n3306 ) | ( n3305 & ~n3306 ) ;
  assign n3308 = ( ~n3121 & n3211 ) | ( ~n3121 & n3307 ) | ( n3211 & n3307 ) ;
  assign n3309 = ( n3121 & n3211 ) | ( n3121 & n3307 ) | ( n3211 & n3307 ) ;
  assign n3310 = ( n3121 & n3308 ) | ( n3121 & ~n3309 ) | ( n3308 & ~n3309 ) ;
  assign n3311 = ( ~n3133 & n3182 ) | ( ~n3133 & n3188 ) | ( n3182 & n3188 ) ;
  assign n3312 = ( n3133 & n3182 ) | ( n3133 & n3188 ) | ( n3182 & n3188 ) ;
  assign n3313 = ( n3133 & n3311 ) | ( n3133 & ~n3312 ) | ( n3311 & ~n3312 ) ;
  assign n3314 = ( ~n3184 & n3310 ) | ( ~n3184 & n3313 ) | ( n3310 & n3313 ) ;
  assign n3315 = ( n3184 & n3310 ) | ( n3184 & n3313 ) | ( n3310 & n3313 ) ;
  assign n3316 = ( n3184 & n3314 ) | ( n3184 & ~n3315 ) | ( n3314 & ~n3315 ) ;
  assign n3317 = ( ~n3218 & n3304 ) | ( ~n3218 & n3316 ) | ( n3304 & n3316 ) ;
  assign n3318 = ( n3218 & n3304 ) | ( n3218 & n3316 ) | ( n3304 & n3316 ) ;
  assign n3319 = ( n3218 & n3317 ) | ( n3218 & ~n3318 ) | ( n3317 & ~n3318 ) ;
  assign n3320 = x21 & x35 ;
  assign n3321 = x5 & x51 ;
  assign n3322 = x18 & x38 ;
  assign n3323 = ( ~n3320 & n3321 ) | ( ~n3320 & n3322 ) | ( n3321 & n3322 ) ;
  assign n3324 = ( n3320 & n3321 ) | ( n3320 & n3322 ) | ( n3321 & n3322 ) ;
  assign n3325 = ( n3320 & n3323 ) | ( n3320 & ~n3324 ) | ( n3323 & ~n3324 ) ;
  assign n3326 = ( n3118 & n3125 ) | ( n3118 & n3325 ) | ( n3125 & n3325 ) ;
  assign n3327 = ( n3118 & ~n3125 ) | ( n3118 & n3325 ) | ( ~n3125 & n3325 ) ;
  assign n3328 = ( n3125 & ~n3326 ) | ( n3125 & n3327 ) | ( ~n3326 & n3327 ) ;
  assign n3329 = ( n3137 & n3190 ) | ( n3137 & n3328 ) | ( n3190 & n3328 ) ;
  assign n3330 = ( ~n3137 & n3190 ) | ( ~n3137 & n3328 ) | ( n3190 & n3328 ) ;
  assign n3331 = ( n3137 & ~n3329 ) | ( n3137 & n3330 ) | ( ~n3329 & n3330 ) ;
  assign n3332 = ( ~n3139 & n3193 ) | ( ~n3139 & n3331 ) | ( n3193 & n3331 ) ;
  assign n3333 = ( n3139 & n3193 ) | ( n3139 & n3331 ) | ( n3193 & n3331 ) ;
  assign n3334 = ( n3139 & n3332 ) | ( n3139 & ~n3333 ) | ( n3332 & ~n3333 ) ;
  assign n3335 = ( ~n3197 & n3319 ) | ( ~n3197 & n3334 ) | ( n3319 & n3334 ) ;
  assign n3336 = ( n3197 & n3319 ) | ( n3197 & n3334 ) | ( n3319 & n3334 ) ;
  assign n3337 = ( n3197 & n3335 ) | ( n3197 & ~n3336 ) | ( n3335 & ~n3336 ) ;
  assign n3338 = ( ~n3220 & n3224 ) | ( ~n3220 & n3337 ) | ( n3224 & n3337 ) ;
  assign n3339 = ( n3220 & n3224 ) | ( n3220 & n3337 ) | ( n3224 & n3337 ) ;
  assign n3340 = ( n3220 & n3338 ) | ( n3220 & ~n3339 ) | ( n3338 & ~n3339 ) ;
  assign n3341 = ( n3266 & ~n3283 ) | ( n3266 & n3296 ) | ( ~n3283 & n3296 ) ;
  assign n3342 = ( n3266 & n3283 ) | ( n3266 & n3296 ) | ( n3283 & n3296 ) ;
  assign n3343 = ( n3283 & n3341 ) | ( n3283 & ~n3342 ) | ( n3341 & ~n3342 ) ;
  assign n3344 = ( ~n3263 & n3273 ) | ( ~n3263 & n3280 ) | ( n3273 & n3280 ) ;
  assign n3345 = ( n3263 & n3273 ) | ( n3263 & n3280 ) | ( n3273 & n3280 ) ;
  assign n3346 = ( n3263 & n3344 ) | ( n3263 & ~n3345 ) | ( n3344 & ~n3345 ) ;
  assign n3347 = ( ~n3236 & n3242 ) | ( ~n3236 & n3251 ) | ( n3242 & n3251 ) ;
  assign n3348 = ( n3236 & n3242 ) | ( n3236 & n3251 ) | ( n3242 & n3251 ) ;
  assign n3349 = ( n3236 & n3347 ) | ( n3236 & ~n3348 ) | ( n3347 & ~n3348 ) ;
  assign n3350 = ( n3244 & n3346 ) | ( n3244 & n3349 ) | ( n3346 & n3349 ) ;
  assign n3351 = ( ~n3244 & n3346 ) | ( ~n3244 & n3349 ) | ( n3346 & n3349 ) ;
  assign n3352 = ( n3244 & ~n3350 ) | ( n3244 & n3351 ) | ( ~n3350 & n3351 ) ;
  assign n3353 = ( ~n3285 & n3343 ) | ( ~n3285 & n3352 ) | ( n3343 & n3352 ) ;
  assign n3354 = ( n3285 & n3343 ) | ( n3285 & n3352 ) | ( n3343 & n3352 ) ;
  assign n3355 = ( n3285 & n3353 ) | ( n3285 & ~n3354 ) | ( n3353 & ~n3354 ) ;
  assign n3356 = x15 & x42 ;
  assign n3357 = x9 & x48 ;
  assign n3358 = x10 & x47 ;
  assign n3359 = ( ~n3356 & n3357 ) | ( ~n3356 & n3358 ) | ( n3357 & n3358 ) ;
  assign n3360 = ( n3356 & n3357 ) | ( n3356 & n3358 ) | ( n3357 & n3358 ) ;
  assign n3361 = ( n3356 & n3359 ) | ( n3356 & ~n3360 ) | ( n3359 & ~n3360 ) ;
  assign n3362 = x5 & x52 ;
  assign n3363 = x19 & x38 ;
  assign n3364 = x20 & x37 ;
  assign n3365 = ( ~n3362 & n3363 ) | ( ~n3362 & n3364 ) | ( n3363 & n3364 ) ;
  assign n3366 = ( n3362 & n3363 ) | ( n3362 & n3364 ) | ( n3363 & n3364 ) ;
  assign n3367 = ( n3362 & n3365 ) | ( n3362 & ~n3366 ) | ( n3365 & ~n3366 ) ;
  assign n3368 = x3 & x54 ;
  assign n3369 = x4 & x53 ;
  assign n3370 = x2 & x55 ;
  assign n3371 = ( ~n3368 & n3369 ) | ( ~n3368 & n3370 ) | ( n3369 & n3370 ) ;
  assign n3372 = ( n3368 & n3369 ) | ( n3368 & n3370 ) | ( n3369 & n3370 ) ;
  assign n3373 = ( n3368 & n3371 ) | ( n3368 & ~n3372 ) | ( n3371 & ~n3372 ) ;
  assign n3374 = ( ~n3361 & n3367 ) | ( ~n3361 & n3373 ) | ( n3367 & n3373 ) ;
  assign n3375 = ( n3361 & n3367 ) | ( n3361 & n3373 ) | ( n3367 & n3373 ) ;
  assign n3376 = ( n3361 & n3374 ) | ( n3361 & ~n3375 ) | ( n3374 & ~n3375 ) ;
  assign n3377 = x12 & x45 ;
  assign n3378 = x28 & x29 ;
  assign n3379 = x27 & x30 ;
  assign n3380 = ( ~n3377 & n3378 ) | ( ~n3377 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3381 = ( n3377 & n3378 ) | ( n3377 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3382 = ( n3377 & n3380 ) | ( n3377 & ~n3381 ) | ( n3380 & ~n3381 ) ;
  assign n3383 = x18 & x39 ;
  assign n3384 = x6 & x51 ;
  assign n3385 = x17 & x40 ;
  assign n3386 = ( ~n3383 & n3384 ) | ( ~n3383 & n3385 ) | ( n3384 & n3385 ) ;
  assign n3387 = ( n3383 & n3384 ) | ( n3383 & n3385 ) | ( n3384 & n3385 ) ;
  assign n3388 = ( n3383 & n3386 ) | ( n3383 & ~n3387 ) | ( n3386 & ~n3387 ) ;
  assign n3389 = x14 & x43 ;
  assign n3390 = x13 & x44 ;
  assign n3391 = x11 & x46 ;
  assign n3392 = ( ~n3389 & n3390 ) | ( ~n3389 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3393 = ( n3389 & n3390 ) | ( n3389 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3394 = ( n3389 & n3392 ) | ( n3389 & ~n3393 ) | ( n3392 & ~n3393 ) ;
  assign n3395 = ( ~n3382 & n3388 ) | ( ~n3382 & n3394 ) | ( n3388 & n3394 ) ;
  assign n3396 = ( n3382 & n3388 ) | ( n3382 & n3394 ) | ( n3388 & n3394 ) ;
  assign n3397 = ( n3382 & n3395 ) | ( n3382 & ~n3396 ) | ( n3395 & ~n3396 ) ;
  assign n3398 = ( n3312 & n3376 ) | ( n3312 & n3397 ) | ( n3376 & n3397 ) ;
  assign n3399 = ( ~n3312 & n3376 ) | ( ~n3312 & n3397 ) | ( n3376 & n3397 ) ;
  assign n3400 = ( n3312 & ~n3398 ) | ( n3312 & n3399 ) | ( ~n3398 & n3399 ) ;
  assign n3401 = ( n3230 & ~n3257 ) | ( n3230 & n3324 ) | ( ~n3257 & n3324 ) ;
  assign n3402 = ( n3230 & n3257 ) | ( n3230 & n3324 ) | ( n3257 & n3324 ) ;
  assign n3403 = ( n3257 & n3401 ) | ( n3257 & ~n3402 ) | ( n3401 & ~n3402 ) ;
  assign n3404 = x24 & x33 ;
  assign n3405 = x26 & x31 ;
  assign n3406 = x25 & x32 ;
  assign n3407 = ( ~n3404 & n3405 ) | ( ~n3404 & n3406 ) | ( n3405 & n3406 ) ;
  assign n3408 = ( n3404 & n3405 ) | ( n3404 & n3406 ) | ( n3405 & n3406 ) ;
  assign n3409 = ( n3404 & n3407 ) | ( n3404 & ~n3408 ) | ( n3407 & ~n3408 ) ;
  assign n3410 = x21 & x36 ;
  assign n3411 = x23 & x34 ;
  assign n3412 = x22 & x35 ;
  assign n3413 = ( ~n3410 & n3411 ) | ( ~n3410 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3414 = ( n3410 & n3411 ) | ( n3410 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3415 = ( n3410 & n3413 ) | ( n3410 & ~n3414 ) | ( n3413 & ~n3414 ) ;
  assign n3416 = x7 & x50 ;
  assign n3417 = x8 & x49 ;
  assign n3418 = x16 & x41 ;
  assign n3419 = ( ~n3416 & n3417 ) | ( ~n3416 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3420 = ( n3416 & n3417 ) | ( n3416 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3421 = ( n3416 & n3419 ) | ( n3416 & ~n3420 ) | ( n3419 & ~n3420 ) ;
  assign n3422 = ( ~n3409 & n3415 ) | ( ~n3409 & n3421 ) | ( n3415 & n3421 ) ;
  assign n3423 = ( n3409 & n3415 ) | ( n3409 & n3421 ) | ( n3415 & n3421 ) ;
  assign n3424 = ( n3409 & n3422 ) | ( n3409 & ~n3423 ) | ( n3422 & ~n3423 ) ;
  assign n3425 = ( ~n3326 & n3403 ) | ( ~n3326 & n3424 ) | ( n3403 & n3424 ) ;
  assign n3426 = ( n3326 & n3403 ) | ( n3326 & n3424 ) | ( n3403 & n3424 ) ;
  assign n3427 = ( n3326 & n3425 ) | ( n3326 & ~n3426 ) | ( n3425 & ~n3426 ) ;
  assign n3428 = ( ~n3329 & n3400 ) | ( ~n3329 & n3427 ) | ( n3400 & n3427 ) ;
  assign n3429 = ( n3329 & n3400 ) | ( n3329 & n3427 ) | ( n3400 & n3427 ) ;
  assign n3430 = ( n3329 & n3428 ) | ( n3329 & ~n3429 ) | ( n3428 & ~n3429 ) ;
  assign n3431 = ( n3333 & n3355 ) | ( n3333 & n3430 ) | ( n3355 & n3430 ) ;
  assign n3432 = ( ~n3333 & n3355 ) | ( ~n3333 & n3430 ) | ( n3355 & n3430 ) ;
  assign n3433 = ( n3333 & ~n3431 ) | ( n3333 & n3432 ) | ( ~n3431 & n3432 ) ;
  assign n3434 = x0 & x57 ;
  assign n3435 = x1 & x56 ;
  assign n3436 = x29 & n3435 ;
  assign n3437 = x29 | n3435 ;
  assign n3438 = ~n3436 & n3437 ;
  assign n3439 = ( n3293 & n3434 ) | ( n3293 & n3438 ) | ( n3434 & n3438 ) ;
  assign n3440 = ( ~n3293 & n3434 ) | ( ~n3293 & n3438 ) | ( n3434 & n3438 ) ;
  assign n3441 = ( n3293 & ~n3439 ) | ( n3293 & n3440 ) | ( ~n3439 & n3440 ) ;
  assign n3442 = ( ~n3288 & n3306 ) | ( ~n3288 & n3441 ) | ( n3306 & n3441 ) ;
  assign n3443 = ( n3288 & n3306 ) | ( n3288 & n3441 ) | ( n3306 & n3441 ) ;
  assign n3444 = ( n3288 & n3442 ) | ( n3288 & ~n3443 ) | ( n3442 & ~n3443 ) ;
  assign n3445 = ( n3299 & n3309 ) | ( n3299 & n3444 ) | ( n3309 & n3444 ) ;
  assign n3446 = ( ~n3299 & n3309 ) | ( ~n3299 & n3444 ) | ( n3309 & n3444 ) ;
  assign n3447 = ( n3299 & ~n3445 ) | ( n3299 & n3446 ) | ( ~n3445 & n3446 ) ;
  assign n3448 = ( n3303 & n3315 ) | ( n3303 & n3447 ) | ( n3315 & n3447 ) ;
  assign n3449 = ( n3303 & ~n3315 ) | ( n3303 & n3447 ) | ( ~n3315 & n3447 ) ;
  assign n3450 = ( n3315 & ~n3448 ) | ( n3315 & n3449 ) | ( ~n3448 & n3449 ) ;
  assign n3451 = ( ~n3318 & n3433 ) | ( ~n3318 & n3450 ) | ( n3433 & n3450 ) ;
  assign n3452 = ( n3318 & n3433 ) | ( n3318 & n3450 ) | ( n3433 & n3450 ) ;
  assign n3453 = ( n3318 & n3451 ) | ( n3318 & ~n3452 ) | ( n3451 & ~n3452 ) ;
  assign n3454 = ( n3336 & n3339 ) | ( n3336 & n3453 ) | ( n3339 & n3453 ) ;
  assign n3455 = ( ~n3336 & n3339 ) | ( ~n3336 & n3453 ) | ( n3339 & n3453 ) ;
  assign n3456 = ( n3336 & ~n3454 ) | ( n3336 & n3455 ) | ( ~n3454 & n3455 ) ;
  assign n3457 = ( n3345 & n3348 ) | ( n3345 & n3402 ) | ( n3348 & n3402 ) ;
  assign n3458 = ( ~n3345 & n3348 ) | ( ~n3345 & n3402 ) | ( n3348 & n3402 ) ;
  assign n3459 = ( n3345 & ~n3457 ) | ( n3345 & n3458 ) | ( ~n3457 & n3458 ) ;
  assign n3460 = ( ~n3350 & n3426 ) | ( ~n3350 & n3459 ) | ( n3426 & n3459 ) ;
  assign n3461 = ( n3350 & n3426 ) | ( n3350 & n3459 ) | ( n3426 & n3459 ) ;
  assign n3462 = ( n3350 & n3460 ) | ( n3350 & ~n3461 ) | ( n3460 & ~n3461 ) ;
  assign n3463 = ( n3354 & n3429 ) | ( n3354 & n3462 ) | ( n3429 & n3462 ) ;
  assign n3464 = ( ~n3354 & n3429 ) | ( ~n3354 & n3462 ) | ( n3429 & n3462 ) ;
  assign n3465 = ( n3354 & ~n3463 ) | ( n3354 & n3464 ) | ( ~n3463 & n3464 ) ;
  assign n3466 = ( n3366 & n3372 ) | ( n3366 & n3393 ) | ( n3372 & n3393 ) ;
  assign n3467 = ( n3366 & ~n3372 ) | ( n3366 & n3393 ) | ( ~n3372 & n3393 ) ;
  assign n3468 = ( n3372 & ~n3466 ) | ( n3372 & n3467 ) | ( ~n3466 & n3467 ) ;
  assign n3469 = ( n3360 & ~n3408 ) | ( n3360 & n3414 ) | ( ~n3408 & n3414 ) ;
  assign n3470 = ( n3360 & n3408 ) | ( n3360 & n3414 ) | ( n3408 & n3414 ) ;
  assign n3471 = ( n3408 & n3469 ) | ( n3408 & ~n3470 ) | ( n3469 & ~n3470 ) ;
  assign n3472 = ( n3423 & n3468 ) | ( n3423 & n3471 ) | ( n3468 & n3471 ) ;
  assign n3473 = ( n3423 & ~n3468 ) | ( n3423 & n3471 ) | ( ~n3468 & n3471 ) ;
  assign n3474 = ( n3468 & ~n3472 ) | ( n3468 & n3473 ) | ( ~n3472 & n3473 ) ;
  assign n3475 = x28 & x30 ;
  assign n3476 = x1 & x57 ;
  assign n3477 = n3475 & n3476 ;
  assign n3478 = n3475 | n3476 ;
  assign n3479 = ~n3477 & n3478 ;
  assign n3480 = ( ~n3381 & n3436 ) | ( ~n3381 & n3479 ) | ( n3436 & n3479 ) ;
  assign n3481 = ( n3381 & n3436 ) | ( n3381 & n3479 ) | ( n3436 & n3479 ) ;
  assign n3482 = ( n3381 & n3480 ) | ( n3381 & ~n3481 ) | ( n3480 & ~n3481 ) ;
  assign n3483 = ( ~n3375 & n3396 ) | ( ~n3375 & n3482 ) | ( n3396 & n3482 ) ;
  assign n3484 = ( n3375 & n3396 ) | ( n3375 & n3482 ) | ( n3396 & n3482 ) ;
  assign n3485 = ( n3375 & n3483 ) | ( n3375 & ~n3484 ) | ( n3483 & ~n3484 ) ;
  assign n3486 = ( ~n3398 & n3474 ) | ( ~n3398 & n3485 ) | ( n3474 & n3485 ) ;
  assign n3487 = ( n3398 & n3474 ) | ( n3398 & n3485 ) | ( n3474 & n3485 ) ;
  assign n3488 = ( n3398 & n3486 ) | ( n3398 & ~n3487 ) | ( n3486 & ~n3487 ) ;
  assign n3489 = x17 & x41 ;
  assign n3490 = x9 & x49 ;
  assign n3491 = x16 & x42 ;
  assign n3492 = ( ~n3489 & n3490 ) | ( ~n3489 & n3491 ) | ( n3490 & n3491 ) ;
  assign n3493 = ( n3489 & n3490 ) | ( n3489 & n3491 ) | ( n3490 & n3491 ) ;
  assign n3494 = ( n3489 & n3492 ) | ( n3489 & ~n3493 ) | ( n3492 & ~n3493 ) ;
  assign n3495 = x0 & x58 ;
  assign n3496 = x4 & x54 ;
  assign n3497 = ( ~n3271 & n3495 ) | ( ~n3271 & n3496 ) | ( n3495 & n3496 ) ;
  assign n3498 = ( n3271 & n3495 ) | ( n3271 & n3496 ) | ( n3495 & n3496 ) ;
  assign n3499 = ( n3271 & n3497 ) | ( n3271 & ~n3498 ) | ( n3497 & ~n3498 ) ;
  assign n3500 = x5 & x53 ;
  assign n3501 = x21 & x37 ;
  assign n3502 = ( ~n1602 & n3500 ) | ( ~n1602 & n3501 ) | ( n3500 & n3501 ) ;
  assign n3503 = ( n1602 & n3500 ) | ( n1602 & n3501 ) | ( n3500 & n3501 ) ;
  assign n3504 = ( n1602 & n3502 ) | ( n1602 & ~n3503 ) | ( n3502 & ~n3503 ) ;
  assign n3505 = ( ~n3494 & n3499 ) | ( ~n3494 & n3504 ) | ( n3499 & n3504 ) ;
  assign n3506 = ( n3494 & n3499 ) | ( n3494 & n3504 ) | ( n3499 & n3504 ) ;
  assign n3507 = ( n3494 & n3505 ) | ( n3494 & ~n3506 ) | ( n3505 & ~n3506 ) ;
  assign n3508 = x22 & x36 ;
  assign n3509 = x23 & x35 ;
  assign n3510 = x24 & x34 ;
  assign n3511 = ( ~n3508 & n3509 ) | ( ~n3508 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3512 = ( n3508 & n3509 ) | ( n3508 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3513 = ( n3508 & n3511 ) | ( n3508 & ~n3512 ) | ( n3511 & ~n3512 ) ;
  assign n3514 = x25 & x33 ;
  assign n3515 = x26 & x32 ;
  assign n3516 = x27 & x31 ;
  assign n3517 = ( ~n3514 & n3515 ) | ( ~n3514 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3518 = ( n3514 & n3515 ) | ( n3514 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3519 = ( n3514 & n3517 ) | ( n3514 & ~n3518 ) | ( n3517 & ~n3518 ) ;
  assign n3520 = x18 & x40 ;
  assign n3521 = x7 & x51 ;
  assign n3522 = x8 & x50 ;
  assign n3523 = ( ~n3520 & n3521 ) | ( ~n3520 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3524 = ( n3520 & n3521 ) | ( n3520 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3525 = ( n3520 & n3523 ) | ( n3520 & ~n3524 ) | ( n3523 & ~n3524 ) ;
  assign n3526 = ( ~n3513 & n3519 ) | ( ~n3513 & n3525 ) | ( n3519 & n3525 ) ;
  assign n3527 = ( n3513 & n3519 ) | ( n3513 & n3525 ) | ( n3519 & n3525 ) ;
  assign n3528 = ( n3513 & n3526 ) | ( n3513 & ~n3527 ) | ( n3526 & ~n3527 ) ;
  assign n3529 = ( ~n3342 & n3507 ) | ( ~n3342 & n3528 ) | ( n3507 & n3528 ) ;
  assign n3530 = ( n3342 & n3507 ) | ( n3342 & n3528 ) | ( n3507 & n3528 ) ;
  assign n3531 = ( n3342 & n3529 ) | ( n3342 & ~n3530 ) | ( n3529 & ~n3530 ) ;
  assign n3532 = ( n3387 & n3420 ) | ( n3387 & ~n3439 ) | ( n3420 & ~n3439 ) ;
  assign n3533 = ( n3387 & n3420 ) | ( n3387 & n3439 ) | ( n3420 & n3439 ) ;
  assign n3534 = ( n3439 & n3532 ) | ( n3439 & ~n3533 ) | ( n3532 & ~n3533 ) ;
  assign n3535 = x14 & x44 ;
  assign n3536 = x13 & x45 ;
  assign n3537 = x12 & x46 ;
  assign n3538 = ( ~n3535 & n3536 ) | ( ~n3535 & n3537 ) | ( n3536 & n3537 ) ;
  assign n3539 = ( n3535 & n3536 ) | ( n3535 & n3537 ) | ( n3536 & n3537 ) ;
  assign n3540 = ( n3535 & n3538 ) | ( n3535 & ~n3539 ) | ( n3538 & ~n3539 ) ;
  assign n3541 = x10 & x48 ;
  assign n3542 = x15 & x43 ;
  assign n3543 = x11 & x47 ;
  assign n3544 = ( ~n3541 & n3542 ) | ( ~n3541 & n3543 ) | ( n3542 & n3543 ) ;
  assign n3545 = ( n3541 & n3542 ) | ( n3541 & n3543 ) | ( n3542 & n3543 ) ;
  assign n3546 = ( n3541 & n3544 ) | ( n3541 & ~n3545 ) | ( n3544 & ~n3545 ) ;
  assign n3547 = x3 & x55 ;
  assign n3548 = x19 & x39 ;
  assign n3549 = x6 & x52 ;
  assign n3550 = ( ~n3547 & n3548 ) | ( ~n3547 & n3549 ) | ( n3548 & n3549 ) ;
  assign n3551 = ( n3547 & n3548 ) | ( n3547 & n3549 ) | ( n3548 & n3549 ) ;
  assign n3552 = ( n3547 & n3550 ) | ( n3547 & ~n3551 ) | ( n3550 & ~n3551 ) ;
  assign n3553 = ( ~n3540 & n3546 ) | ( ~n3540 & n3552 ) | ( n3546 & n3552 ) ;
  assign n3554 = ( n3540 & n3546 ) | ( n3540 & n3552 ) | ( n3546 & n3552 ) ;
  assign n3555 = ( n3540 & n3553 ) | ( n3540 & ~n3554 ) | ( n3553 & ~n3554 ) ;
  assign n3556 = ( ~n3443 & n3534 ) | ( ~n3443 & n3555 ) | ( n3534 & n3555 ) ;
  assign n3557 = ( n3443 & n3534 ) | ( n3443 & n3555 ) | ( n3534 & n3555 ) ;
  assign n3558 = ( n3443 & n3556 ) | ( n3443 & ~n3557 ) | ( n3556 & ~n3557 ) ;
  assign n3559 = ( n3445 & n3531 ) | ( n3445 & n3558 ) | ( n3531 & n3558 ) ;
  assign n3560 = ( ~n3445 & n3531 ) | ( ~n3445 & n3558 ) | ( n3531 & n3558 ) ;
  assign n3561 = ( n3445 & ~n3559 ) | ( n3445 & n3560 ) | ( ~n3559 & n3560 ) ;
  assign n3562 = ( ~n3448 & n3488 ) | ( ~n3448 & n3561 ) | ( n3488 & n3561 ) ;
  assign n3563 = ( n3448 & n3488 ) | ( n3448 & n3561 ) | ( n3488 & n3561 ) ;
  assign n3564 = ( n3448 & n3562 ) | ( n3448 & ~n3563 ) | ( n3562 & ~n3563 ) ;
  assign n3565 = ( ~n3431 & n3465 ) | ( ~n3431 & n3564 ) | ( n3465 & n3564 ) ;
  assign n3566 = ( n3431 & n3465 ) | ( n3431 & n3564 ) | ( n3465 & n3564 ) ;
  assign n3567 = ( n3431 & n3565 ) | ( n3431 & ~n3566 ) | ( n3565 & ~n3566 ) ;
  assign n3568 = ( n3452 & n3454 ) | ( n3452 & n3567 ) | ( n3454 & n3567 ) ;
  assign n3569 = ( ~n3452 & n3454 ) | ( ~n3452 & n3567 ) | ( n3454 & n3567 ) ;
  assign n3570 = ( n3452 & ~n3568 ) | ( n3452 & n3569 ) | ( ~n3568 & n3569 ) ;
  assign n3571 = ( n3466 & n3470 ) | ( n3466 & n3533 ) | ( n3470 & n3533 ) ;
  assign n3572 = ( ~n3466 & n3470 ) | ( ~n3466 & n3533 ) | ( n3470 & n3533 ) ;
  assign n3573 = ( n3466 & ~n3571 ) | ( n3466 & n3572 ) | ( ~n3571 & n3572 ) ;
  assign n3574 = ( ~n3472 & n3557 ) | ( ~n3472 & n3573 ) | ( n3557 & n3573 ) ;
  assign n3575 = ( n3472 & n3557 ) | ( n3472 & n3573 ) | ( n3557 & n3573 ) ;
  assign n3576 = ( n3472 & n3574 ) | ( n3472 & ~n3575 ) | ( n3574 & ~n3575 ) ;
  assign n3577 = ( ~n3487 & n3559 ) | ( ~n3487 & n3576 ) | ( n3559 & n3576 ) ;
  assign n3578 = ( n3487 & n3559 ) | ( n3487 & n3576 ) | ( n3559 & n3576 ) ;
  assign n3579 = ( n3487 & n3577 ) | ( n3487 & ~n3578 ) | ( n3577 & ~n3578 ) ;
  assign n3580 = ( n3506 & n3527 ) | ( n3506 & n3554 ) | ( n3527 & n3554 ) ;
  assign n3581 = ( n3506 & ~n3527 ) | ( n3506 & n3554 ) | ( ~n3527 & n3554 ) ;
  assign n3582 = ( n3527 & ~n3580 ) | ( n3527 & n3581 ) | ( ~n3580 & n3581 ) ;
  assign n3583 = ( n3503 & n3512 ) | ( n3503 & n3524 ) | ( n3512 & n3524 ) ;
  assign n3584 = ( n3503 & ~n3512 ) | ( n3503 & n3524 ) | ( ~n3512 & n3524 ) ;
  assign n3585 = ( n3512 & ~n3583 ) | ( n3512 & n3584 ) | ( ~n3583 & n3584 ) ;
  assign n3586 = ( ~n3493 & n3498 ) | ( ~n3493 & n3551 ) | ( n3498 & n3551 ) ;
  assign n3587 = ( n3493 & n3498 ) | ( n3493 & n3551 ) | ( n3498 & n3551 ) ;
  assign n3588 = ( n3493 & n3586 ) | ( n3493 & ~n3587 ) | ( n3586 & ~n3587 ) ;
  assign n3589 = ( x1 & x30 ) | ( x1 & x58 ) | ( x30 & x58 ) ;
  assign n3590 = ~x1 & x30 ;
  assign n3591 = x30 & x58 ;
  assign n3592 = ( n3589 & n3590 ) | ( n3589 & ~n3591 ) | ( n3590 & ~n3591 ) ;
  assign n3593 = ( ~n3539 & n3545 ) | ( ~n3539 & n3592 ) | ( n3545 & n3592 ) ;
  assign n3594 = ( n3539 & n3545 ) | ( n3539 & n3592 ) | ( n3545 & n3592 ) ;
  assign n3595 = ( n3539 & n3593 ) | ( n3539 & ~n3594 ) | ( n3593 & ~n3594 ) ;
  assign n3596 = ( ~n3585 & n3588 ) | ( ~n3585 & n3595 ) | ( n3588 & n3595 ) ;
  assign n3597 = ( n3585 & n3588 ) | ( n3585 & n3595 ) | ( n3588 & n3595 ) ;
  assign n3598 = ( n3585 & n3596 ) | ( n3585 & ~n3597 ) | ( n3596 & ~n3597 ) ;
  assign n3599 = ( ~n3530 & n3582 ) | ( ~n3530 & n3598 ) | ( n3582 & n3598 ) ;
  assign n3600 = ( n3530 & n3582 ) | ( n3530 & n3598 ) | ( n3582 & n3598 ) ;
  assign n3601 = ( n3530 & n3599 ) | ( n3530 & ~n3600 ) | ( n3599 & ~n3600 ) ;
  assign n3602 = x3 & x57 ;
  assign n3603 = n3271 & n3602 ;
  assign n3604 = x2 & x57 ;
  assign n3605 = x3 & x56 ;
  assign n3606 = n3604 | n3605 ;
  assign n3607 = ( n3477 & n3603 ) | ( n3477 & n3606 ) | ( n3603 & n3606 ) ;
  assign n3608 = ( ~n3477 & n3603 ) | ( ~n3477 & n3606 ) | ( n3603 & n3606 ) ;
  assign n3609 = ( n3477 & ~n3607 ) | ( n3477 & n3608 ) | ( ~n3607 & n3608 ) ;
  assign n3610 = x4 & x55 ;
  assign n3611 = x5 & x54 ;
  assign n3612 = x19 & x40 ;
  assign n3613 = ( ~n3610 & n3611 ) | ( ~n3610 & n3612 ) | ( n3611 & n3612 ) ;
  assign n3614 = ( n3610 & n3611 ) | ( n3610 & n3612 ) | ( n3611 & n3612 ) ;
  assign n3615 = ( n3610 & n3613 ) | ( n3610 & ~n3614 ) | ( n3613 & ~n3614 ) ;
  assign n3616 = ( ~n3518 & n3609 ) | ( ~n3518 & n3615 ) | ( n3609 & n3615 ) ;
  assign n3617 = ( n3518 & n3609 ) | ( n3518 & n3615 ) | ( n3609 & n3615 ) ;
  assign n3618 = ( n3518 & n3616 ) | ( n3518 & ~n3617 ) | ( n3616 & ~n3617 ) ;
  assign n3619 = x8 & x51 ;
  assign n3620 = x16 & x43 ;
  assign n3621 = x17 & x42 ;
  assign n3622 = ( ~n3619 & n3620 ) | ( ~n3619 & n3621 ) | ( n3620 & n3621 ) ;
  assign n3623 = ( n3619 & n3620 ) | ( n3619 & n3621 ) | ( n3620 & n3621 ) ;
  assign n3624 = ( n3619 & n3622 ) | ( n3619 & ~n3623 ) | ( n3622 & ~n3623 ) ;
  assign n3625 = x13 & x46 ;
  assign n3626 = x29 & x30 ;
  assign n3627 = x28 & x31 ;
  assign n3628 = ( ~n3625 & n3626 ) | ( ~n3625 & n3627 ) | ( n3626 & n3627 ) ;
  assign n3629 = ( n3625 & n3626 ) | ( n3625 & n3627 ) | ( n3626 & n3627 ) ;
  assign n3630 = ( n3625 & n3628 ) | ( n3625 & ~n3629 ) | ( n3628 & ~n3629 ) ;
  assign n3631 = x11 & x48 ;
  assign n3632 = x14 & x45 ;
  assign n3633 = x12 & x47 ;
  assign n3634 = ( ~n3631 & n3632 ) | ( ~n3631 & n3633 ) | ( n3632 & n3633 ) ;
  assign n3635 = ( n3631 & n3632 ) | ( n3631 & n3633 ) | ( n3632 & n3633 ) ;
  assign n3636 = ( n3631 & n3634 ) | ( n3631 & ~n3635 ) | ( n3634 & ~n3635 ) ;
  assign n3637 = ( ~n3624 & n3630 ) | ( ~n3624 & n3636 ) | ( n3630 & n3636 ) ;
  assign n3638 = ( n3624 & n3630 ) | ( n3624 & n3636 ) | ( n3630 & n3636 ) ;
  assign n3639 = ( n3624 & n3637 ) | ( n3624 & ~n3638 ) | ( n3637 & ~n3638 ) ;
  assign n3640 = ( n3484 & n3618 ) | ( n3484 & n3639 ) | ( n3618 & n3639 ) ;
  assign n3641 = ( ~n3484 & n3618 ) | ( ~n3484 & n3639 ) | ( n3618 & n3639 ) ;
  assign n3642 = ( n3484 & ~n3640 ) | ( n3484 & n3641 ) | ( ~n3640 & n3641 ) ;
  assign n3643 = x9 & x50 ;
  assign n3644 = x15 & x44 ;
  assign n3645 = x10 & x49 ;
  assign n3646 = ( ~n3643 & n3644 ) | ( ~n3643 & n3645 ) | ( n3644 & n3645 ) ;
  assign n3647 = ( n3643 & n3644 ) | ( n3643 & n3645 ) | ( n3644 & n3645 ) ;
  assign n3648 = ( n3643 & n3646 ) | ( n3643 & ~n3647 ) | ( n3646 & ~n3647 ) ;
  assign n3649 = x6 & x53 ;
  assign n3650 = x7 & x52 ;
  assign n3651 = x18 & x41 ;
  assign n3652 = ( ~n3649 & n3650 ) | ( ~n3649 & n3651 ) | ( n3650 & n3651 ) ;
  assign n3653 = ( n3649 & n3650 ) | ( n3649 & n3651 ) | ( n3650 & n3651 ) ;
  assign n3654 = ( n3649 & n3652 ) | ( n3649 & ~n3653 ) | ( n3652 & ~n3653 ) ;
  assign n3655 = ( n3481 & n3648 ) | ( n3481 & n3654 ) | ( n3648 & n3654 ) ;
  assign n3656 = ( ~n3481 & n3648 ) | ( ~n3481 & n3654 ) | ( n3648 & n3654 ) ;
  assign n3657 = ( n3481 & ~n3655 ) | ( n3481 & n3656 ) | ( ~n3655 & n3656 ) ;
  assign n3658 = x23 & x36 ;
  assign n3659 = x24 & x35 ;
  assign n3660 = x25 & x34 ;
  assign n3661 = ( ~n3658 & n3659 ) | ( ~n3658 & n3660 ) | ( n3659 & n3660 ) ;
  assign n3662 = ( n3658 & n3659 ) | ( n3658 & n3660 ) | ( n3659 & n3660 ) ;
  assign n3663 = ( n3658 & n3661 ) | ( n3658 & ~n3662 ) | ( n3661 & ~n3662 ) ;
  assign n3664 = x26 & x33 ;
  assign n3665 = x27 & x32 ;
  assign n3666 = x0 & x59 ;
  assign n3667 = ( ~n3664 & n3665 ) | ( ~n3664 & n3666 ) | ( n3665 & n3666 ) ;
  assign n3668 = ( n3664 & n3665 ) | ( n3664 & n3666 ) | ( n3665 & n3666 ) ;
  assign n3669 = ( n3664 & n3667 ) | ( n3664 & ~n3668 ) | ( n3667 & ~n3668 ) ;
  assign n3670 = x20 & x39 ;
  assign n3671 = x21 & x38 ;
  assign n3672 = x22 & x37 ;
  assign n3673 = ( ~n3670 & n3671 ) | ( ~n3670 & n3672 ) | ( n3671 & n3672 ) ;
  assign n3674 = ( n3670 & n3671 ) | ( n3670 & n3672 ) | ( n3671 & n3672 ) ;
  assign n3675 = ( n3670 & n3673 ) | ( n3670 & ~n3674 ) | ( n3673 & ~n3674 ) ;
  assign n3676 = ( ~n3663 & n3669 ) | ( ~n3663 & n3675 ) | ( n3669 & n3675 ) ;
  assign n3677 = ( n3663 & n3669 ) | ( n3663 & n3675 ) | ( n3669 & n3675 ) ;
  assign n3678 = ( n3663 & n3676 ) | ( n3663 & ~n3677 ) | ( n3676 & ~n3677 ) ;
  assign n3679 = ( ~n3457 & n3657 ) | ( ~n3457 & n3678 ) | ( n3657 & n3678 ) ;
  assign n3680 = ( n3457 & n3657 ) | ( n3457 & n3678 ) | ( n3657 & n3678 ) ;
  assign n3681 = ( n3457 & n3679 ) | ( n3457 & ~n3680 ) | ( n3679 & ~n3680 ) ;
  assign n3682 = ( ~n3461 & n3642 ) | ( ~n3461 & n3681 ) | ( n3642 & n3681 ) ;
  assign n3683 = ( n3461 & n3642 ) | ( n3461 & n3681 ) | ( n3642 & n3681 ) ;
  assign n3684 = ( n3461 & n3682 ) | ( n3461 & ~n3683 ) | ( n3682 & ~n3683 ) ;
  assign n3685 = ( ~n3463 & n3601 ) | ( ~n3463 & n3684 ) | ( n3601 & n3684 ) ;
  assign n3686 = ( n3463 & n3601 ) | ( n3463 & n3684 ) | ( n3601 & n3684 ) ;
  assign n3687 = ( n3463 & n3685 ) | ( n3463 & ~n3686 ) | ( n3685 & ~n3686 ) ;
  assign n3688 = ( ~n3563 & n3579 ) | ( ~n3563 & n3687 ) | ( n3579 & n3687 ) ;
  assign n3689 = ( n3563 & n3579 ) | ( n3563 & n3687 ) | ( n3579 & n3687 ) ;
  assign n3690 = ( n3563 & n3688 ) | ( n3563 & ~n3689 ) | ( n3688 & ~n3689 ) ;
  assign n3691 = ( ~n3566 & n3568 ) | ( ~n3566 & n3690 ) | ( n3568 & n3690 ) ;
  assign n3692 = ( n3566 & n3568 ) | ( n3566 & n3690 ) | ( n3568 & n3690 ) ;
  assign n3693 = ( n3566 & n3691 ) | ( n3566 & ~n3692 ) | ( n3691 & ~n3692 ) ;
  assign n3694 = x58 & n1036 ;
  assign n3695 = x0 & x60 ;
  assign n3696 = x29 & x31 ;
  assign n3697 = x1 & x59 ;
  assign n3698 = n3696 & n3697 ;
  assign n3699 = n3696 | n3697 ;
  assign n3700 = ~n3698 & n3699 ;
  assign n3701 = ( n3694 & n3695 ) | ( n3694 & n3700 ) | ( n3695 & n3700 ) ;
  assign n3702 = ( ~n3694 & n3695 ) | ( ~n3694 & n3700 ) | ( n3695 & n3700 ) ;
  assign n3703 = ( n3694 & ~n3701 ) | ( n3694 & n3702 ) | ( ~n3701 & n3702 ) ;
  assign n3704 = x27 & x33 ;
  assign n3705 = x28 & x32 ;
  assign n3706 = x23 & x37 ;
  assign n3707 = ( ~n3704 & n3705 ) | ( ~n3704 & n3706 ) | ( n3705 & n3706 ) ;
  assign n3708 = ( n3704 & n3705 ) | ( n3704 & n3706 ) | ( n3705 & n3706 ) ;
  assign n3709 = ( n3704 & n3707 ) | ( n3704 & ~n3708 ) | ( n3707 & ~n3708 ) ;
  assign n3710 = ( n3594 & n3703 ) | ( n3594 & n3709 ) | ( n3703 & n3709 ) ;
  assign n3711 = ( ~n3594 & n3703 ) | ( ~n3594 & n3709 ) | ( n3703 & n3709 ) ;
  assign n3712 = ( n3594 & ~n3710 ) | ( n3594 & n3711 ) | ( ~n3710 & n3711 ) ;
  assign n3713 = x14 & x46 ;
  assign n3714 = x12 & x48 ;
  assign n3715 = x13 & x47 ;
  assign n3716 = ( ~n3713 & n3714 ) | ( ~n3713 & n3715 ) | ( n3714 & n3715 ) ;
  assign n3717 = ( n3713 & n3714 ) | ( n3713 & n3715 ) | ( n3714 & n3715 ) ;
  assign n3718 = ( n3713 & n3716 ) | ( n3713 & ~n3717 ) | ( n3716 & ~n3717 ) ;
  assign n3719 = x7 & x53 ;
  assign n3720 = x8 & x52 ;
  assign n3721 = x18 & x42 ;
  assign n3722 = ( ~n3719 & n3720 ) | ( ~n3719 & n3721 ) | ( n3720 & n3721 ) ;
  assign n3723 = ( n3719 & n3720 ) | ( n3719 & n3721 ) | ( n3720 & n3721 ) ;
  assign n3724 = ( n3719 & n3722 ) | ( n3719 & ~n3723 ) | ( n3722 & ~n3723 ) ;
  assign n3725 = x5 & x55 ;
  assign n3726 = x6 & x54 ;
  assign n3727 = x19 & x41 ;
  assign n3728 = ( ~n3725 & n3726 ) | ( ~n3725 & n3727 ) | ( n3726 & n3727 ) ;
  assign n3729 = ( n3725 & n3726 ) | ( n3725 & n3727 ) | ( n3726 & n3727 ) ;
  assign n3730 = ( n3725 & n3728 ) | ( n3725 & ~n3729 ) | ( n3728 & ~n3729 ) ;
  assign n3731 = ( ~n3718 & n3724 ) | ( ~n3718 & n3730 ) | ( n3724 & n3730 ) ;
  assign n3732 = ( n3718 & n3724 ) | ( n3718 & n3730 ) | ( n3724 & n3730 ) ;
  assign n3733 = ( n3718 & n3731 ) | ( n3718 & ~n3732 ) | ( n3731 & ~n3732 ) ;
  assign n3734 = ( ~n3597 & n3712 ) | ( ~n3597 & n3733 ) | ( n3712 & n3733 ) ;
  assign n3735 = ( n3597 & n3712 ) | ( n3597 & n3733 ) | ( n3712 & n3733 ) ;
  assign n3736 = ( n3597 & n3734 ) | ( n3597 & ~n3735 ) | ( n3734 & ~n3735 ) ;
  assign n3737 = x10 & x50 ;
  assign n3738 = x15 & x45 ;
  assign n3739 = x11 & x49 ;
  assign n3740 = ( ~n3737 & n3738 ) | ( ~n3737 & n3739 ) | ( n3738 & n3739 ) ;
  assign n3741 = ( n3737 & n3738 ) | ( n3737 & n3739 ) | ( n3738 & n3739 ) ;
  assign n3742 = ( n3737 & n3740 ) | ( n3737 & ~n3741 ) | ( n3740 & ~n3741 ) ;
  assign n3743 = x17 & x43 ;
  assign n3744 = x9 & x51 ;
  assign n3745 = x16 & x44 ;
  assign n3746 = ( ~n3743 & n3744 ) | ( ~n3743 & n3745 ) | ( n3744 & n3745 ) ;
  assign n3747 = ( n3743 & n3744 ) | ( n3743 & n3745 ) | ( n3744 & n3745 ) ;
  assign n3748 = ( n3743 & n3746 ) | ( n3743 & ~n3747 ) | ( n3746 & ~n3747 ) ;
  assign n3749 = ( n3635 & n3742 ) | ( n3635 & n3748 ) | ( n3742 & n3748 ) ;
  assign n3750 = ( ~n3635 & n3742 ) | ( ~n3635 & n3748 ) | ( n3742 & n3748 ) ;
  assign n3751 = ( n3635 & ~n3749 ) | ( n3635 & n3750 ) | ( ~n3749 & n3750 ) ;
  assign n3752 = x20 & x40 ;
  assign n3753 = x22 & x38 ;
  assign n3754 = x21 & x39 ;
  assign n3755 = ( ~n3752 & n3753 ) | ( ~n3752 & n3754 ) | ( n3753 & n3754 ) ;
  assign n3756 = ( n3752 & n3753 ) | ( n3752 & n3754 ) | ( n3753 & n3754 ) ;
  assign n3757 = ( n3752 & n3755 ) | ( n3752 & ~n3756 ) | ( n3755 & ~n3756 ) ;
  assign n3758 = x24 & x36 ;
  assign n3759 = x25 & x35 ;
  assign n3760 = x26 & x34 ;
  assign n3761 = ( ~n3758 & n3759 ) | ( ~n3758 & n3760 ) | ( n3759 & n3760 ) ;
  assign n3762 = ( n3758 & n3759 ) | ( n3758 & n3760 ) | ( n3759 & n3760 ) ;
  assign n3763 = ( n3758 & n3761 ) | ( n3758 & ~n3762 ) | ( n3761 & ~n3762 ) ;
  assign n3764 = x2 & x58 ;
  assign n3765 = x4 & x56 ;
  assign n3766 = ( ~n3602 & n3764 ) | ( ~n3602 & n3765 ) | ( n3764 & n3765 ) ;
  assign n3767 = ( n3602 & n3764 ) | ( n3602 & n3765 ) | ( n3764 & n3765 ) ;
  assign n3768 = ( n3602 & n3766 ) | ( n3602 & ~n3767 ) | ( n3766 & ~n3767 ) ;
  assign n3769 = ( ~n3757 & n3763 ) | ( ~n3757 & n3768 ) | ( n3763 & n3768 ) ;
  assign n3770 = ( n3757 & n3763 ) | ( n3757 & n3768 ) | ( n3763 & n3768 ) ;
  assign n3771 = ( n3757 & n3769 ) | ( n3757 & ~n3770 ) | ( n3769 & ~n3770 ) ;
  assign n3772 = ( ~n3571 & n3751 ) | ( ~n3571 & n3771 ) | ( n3751 & n3771 ) ;
  assign n3773 = ( n3571 & n3751 ) | ( n3571 & n3771 ) | ( n3751 & n3771 ) ;
  assign n3774 = ( n3571 & n3772 ) | ( n3571 & ~n3773 ) | ( n3772 & ~n3773 ) ;
  assign n3775 = ( n3575 & n3736 ) | ( n3575 & n3774 ) | ( n3736 & n3774 ) ;
  assign n3776 = ( ~n3575 & n3736 ) | ( ~n3575 & n3774 ) | ( n3736 & n3774 ) ;
  assign n3777 = ( n3575 & ~n3775 ) | ( n3575 & n3776 ) | ( ~n3775 & n3776 ) ;
  assign n3778 = ( n3623 & n3629 ) | ( n3623 & n3653 ) | ( n3629 & n3653 ) ;
  assign n3779 = ( ~n3623 & n3629 ) | ( ~n3623 & n3653 ) | ( n3629 & n3653 ) ;
  assign n3780 = ( n3623 & ~n3778 ) | ( n3623 & n3779 ) | ( ~n3778 & n3779 ) ;
  assign n3781 = ( n3638 & n3677 ) | ( n3638 & n3780 ) | ( n3677 & n3780 ) ;
  assign n3782 = ( n3638 & n3677 ) | ( n3638 & ~n3780 ) | ( n3677 & ~n3780 ) ;
  assign n3783 = ( n3780 & ~n3781 ) | ( n3780 & n3782 ) | ( ~n3781 & n3782 ) ;
  assign n3784 = ( n3614 & ~n3662 ) | ( n3614 & n3674 ) | ( ~n3662 & n3674 ) ;
  assign n3785 = ( n3614 & n3662 ) | ( n3614 & n3674 ) | ( n3662 & n3674 ) ;
  assign n3786 = ( n3662 & n3784 ) | ( n3662 & ~n3785 ) | ( n3784 & ~n3785 ) ;
  assign n3787 = ( n3607 & ~n3647 ) | ( n3607 & n3668 ) | ( ~n3647 & n3668 ) ;
  assign n3788 = ( n3607 & n3647 ) | ( n3607 & n3668 ) | ( n3647 & n3668 ) ;
  assign n3789 = ( n3647 & n3787 ) | ( n3647 & ~n3788 ) | ( n3787 & ~n3788 ) ;
  assign n3790 = ( ~n3655 & n3786 ) | ( ~n3655 & n3789 ) | ( n3786 & n3789 ) ;
  assign n3791 = ( n3655 & n3786 ) | ( n3655 & n3789 ) | ( n3786 & n3789 ) ;
  assign n3792 = ( n3655 & n3790 ) | ( n3655 & ~n3791 ) | ( n3790 & ~n3791 ) ;
  assign n3793 = ( n3640 & n3783 ) | ( n3640 & n3792 ) | ( n3783 & n3792 ) ;
  assign n3794 = ( ~n3640 & n3783 ) | ( ~n3640 & n3792 ) | ( n3783 & n3792 ) ;
  assign n3795 = ( n3640 & ~n3793 ) | ( n3640 & n3794 ) | ( ~n3793 & n3794 ) ;
  assign n3796 = ( ~n3578 & n3777 ) | ( ~n3578 & n3795 ) | ( n3777 & n3795 ) ;
  assign n3797 = ( n3578 & n3777 ) | ( n3578 & n3795 ) | ( n3777 & n3795 ) ;
  assign n3798 = ( n3578 & n3796 ) | ( n3578 & ~n3797 ) | ( n3796 & ~n3797 ) ;
  assign n3799 = ( ~n3583 & n3587 ) | ( ~n3583 & n3617 ) | ( n3587 & n3617 ) ;
  assign n3800 = ( n3583 & n3587 ) | ( n3583 & n3617 ) | ( n3587 & n3617 ) ;
  assign n3801 = ( n3583 & n3799 ) | ( n3583 & ~n3800 ) | ( n3799 & ~n3800 ) ;
  assign n3802 = ( ~n3580 & n3680 ) | ( ~n3580 & n3801 ) | ( n3680 & n3801 ) ;
  assign n3803 = ( n3580 & n3680 ) | ( n3580 & n3801 ) | ( n3680 & n3801 ) ;
  assign n3804 = ( n3580 & n3802 ) | ( n3580 & ~n3803 ) | ( n3802 & ~n3803 ) ;
  assign n3805 = ( ~n3600 & n3683 ) | ( ~n3600 & n3804 ) | ( n3683 & n3804 ) ;
  assign n3806 = ( n3600 & n3683 ) | ( n3600 & n3804 ) | ( n3683 & n3804 ) ;
  assign n3807 = ( n3600 & n3805 ) | ( n3600 & ~n3806 ) | ( n3805 & ~n3806 ) ;
  assign n3808 = ( ~n3686 & n3798 ) | ( ~n3686 & n3807 ) | ( n3798 & n3807 ) ;
  assign n3809 = ( n3686 & n3798 ) | ( n3686 & n3807 ) | ( n3798 & n3807 ) ;
  assign n3810 = ( n3686 & n3808 ) | ( n3686 & ~n3809 ) | ( n3808 & ~n3809 ) ;
  assign n3811 = ( n3689 & n3692 ) | ( n3689 & n3810 ) | ( n3692 & n3810 ) ;
  assign n3812 = ( ~n3689 & n3692 ) | ( ~n3689 & n3810 ) | ( n3692 & n3810 ) ;
  assign n3813 = ( n3689 & ~n3811 ) | ( n3689 & n3812 ) | ( ~n3811 & n3812 ) ;
  assign n3814 = ( ~n3701 & n3723 ) | ( ~n3701 & n3747 ) | ( n3723 & n3747 ) ;
  assign n3815 = ( n3701 & n3723 ) | ( n3701 & n3747 ) | ( n3723 & n3747 ) ;
  assign n3816 = ( n3701 & n3814 ) | ( n3701 & ~n3815 ) | ( n3814 & ~n3815 ) ;
  assign n3817 = ( ~n3710 & n3732 ) | ( ~n3710 & n3816 ) | ( n3732 & n3816 ) ;
  assign n3818 = ( n3710 & n3732 ) | ( n3710 & n3816 ) | ( n3732 & n3816 ) ;
  assign n3819 = ( n3710 & n3817 ) | ( n3710 & ~n3818 ) | ( n3817 & ~n3818 ) ;
  assign n3820 = ( n3729 & n3741 ) | ( n3729 & ~n3767 ) | ( n3741 & ~n3767 ) ;
  assign n3821 = ( n3729 & n3741 ) | ( n3729 & n3767 ) | ( n3741 & n3767 ) ;
  assign n3822 = ( n3767 & n3820 ) | ( n3767 & ~n3821 ) | ( n3820 & ~n3821 ) ;
  assign n3823 = ( n3708 & n3756 ) | ( n3708 & ~n3762 ) | ( n3756 & ~n3762 ) ;
  assign n3824 = ( n3708 & n3756 ) | ( n3708 & n3762 ) | ( n3756 & n3762 ) ;
  assign n3825 = ( n3762 & n3823 ) | ( n3762 & ~n3824 ) | ( n3823 & ~n3824 ) ;
  assign n3826 = ( n3770 & n3822 ) | ( n3770 & n3825 ) | ( n3822 & n3825 ) ;
  assign n3827 = ( n3770 & ~n3822 ) | ( n3770 & n3825 ) | ( ~n3822 & n3825 ) ;
  assign n3828 = ( n3822 & ~n3826 ) | ( n3822 & n3827 ) | ( ~n3826 & n3827 ) ;
  assign n3829 = ( ~n3735 & n3819 ) | ( ~n3735 & n3828 ) | ( n3819 & n3828 ) ;
  assign n3830 = ( n3735 & n3819 ) | ( n3735 & n3828 ) | ( n3819 & n3828 ) ;
  assign n3831 = ( n3735 & n3829 ) | ( n3735 & ~n3830 ) | ( n3829 & ~n3830 ) ;
  assign n3832 = x0 & x61 ;
  assign n3833 = x2 & x59 ;
  assign n3834 = x5 & x56 ;
  assign n3835 = ( ~n3832 & n3833 ) | ( ~n3832 & n3834 ) | ( n3833 & n3834 ) ;
  assign n3836 = ( n3832 & n3833 ) | ( n3832 & n3834 ) | ( n3833 & n3834 ) ;
  assign n3837 = ( n3832 & n3835 ) | ( n3832 & ~n3836 ) | ( n3835 & ~n3836 ) ;
  assign n3838 = x22 & x39 ;
  assign n3839 = x24 & x37 ;
  assign n3840 = x25 & x36 ;
  assign n3841 = ( ~n3838 & n3839 ) | ( ~n3838 & n3840 ) | ( n3839 & n3840 ) ;
  assign n3842 = ( n3838 & n3839 ) | ( n3838 & n3840 ) | ( n3839 & n3840 ) ;
  assign n3843 = ( n3838 & n3841 ) | ( n3838 & ~n3842 ) | ( n3841 & ~n3842 ) ;
  assign n3844 = x6 & x55 ;
  assign n3845 = x20 & x41 ;
  assign n3846 = ( ~n1761 & n3844 ) | ( ~n1761 & n3845 ) | ( n3844 & n3845 ) ;
  assign n3847 = ( n1761 & n3844 ) | ( n1761 & n3845 ) | ( n3844 & n3845 ) ;
  assign n3848 = ( n1761 & n3846 ) | ( n1761 & ~n3847 ) | ( n3846 & ~n3847 ) ;
  assign n3849 = ( ~n3837 & n3843 ) | ( ~n3837 & n3848 ) | ( n3843 & n3848 ) ;
  assign n3850 = ( n3837 & n3843 ) | ( n3837 & n3848 ) | ( n3843 & n3848 ) ;
  assign n3851 = ( n3837 & n3849 ) | ( n3837 & ~n3850 ) | ( n3849 & ~n3850 ) ;
  assign n3852 = x11 & x50 ;
  assign n3853 = x14 & x47 ;
  assign n3854 = x12 & x49 ;
  assign n3855 = ( ~n3852 & n3853 ) | ( ~n3852 & n3854 ) | ( n3853 & n3854 ) ;
  assign n3856 = ( n3852 & n3853 ) | ( n3852 & n3854 ) | ( n3853 & n3854 ) ;
  assign n3857 = ( n3852 & n3855 ) | ( n3852 & ~n3856 ) | ( n3855 & ~n3856 ) ;
  assign n3858 = x13 & x48 ;
  assign n3859 = x30 & x31 ;
  assign n3860 = x29 & x32 ;
  assign n3861 = ( ~n3858 & n3859 ) | ( ~n3858 & n3860 ) | ( n3859 & n3860 ) ;
  assign n3862 = ( n3858 & n3859 ) | ( n3858 & n3860 ) | ( n3859 & n3860 ) ;
  assign n3863 = ( n3858 & n3861 ) | ( n3858 & ~n3862 ) | ( n3861 & ~n3862 ) ;
  assign n3864 = x16 & x45 ;
  assign n3865 = x15 & x46 ;
  assign n3866 = x10 & x51 ;
  assign n3867 = ( ~n3864 & n3865 ) | ( ~n3864 & n3866 ) | ( n3865 & n3866 ) ;
  assign n3868 = ( n3864 & n3865 ) | ( n3864 & n3866 ) | ( n3865 & n3866 ) ;
  assign n3869 = ( n3864 & n3867 ) | ( n3864 & ~n3868 ) | ( n3867 & ~n3868 ) ;
  assign n3870 = ( ~n3857 & n3863 ) | ( ~n3857 & n3869 ) | ( n3863 & n3869 ) ;
  assign n3871 = ( n3857 & n3863 ) | ( n3857 & n3869 ) | ( n3863 & n3869 ) ;
  assign n3872 = ( n3857 & n3870 ) | ( n3857 & ~n3871 ) | ( n3870 & ~n3871 ) ;
  assign n3873 = ( ~n3800 & n3851 ) | ( ~n3800 & n3872 ) | ( n3851 & n3872 ) ;
  assign n3874 = ( n3800 & n3851 ) | ( n3800 & n3872 ) | ( n3851 & n3872 ) ;
  assign n3875 = ( n3800 & n3873 ) | ( n3800 & ~n3874 ) | ( n3873 & ~n3874 ) ;
  assign n3876 = ( n3793 & n3803 ) | ( n3793 & n3875 ) | ( n3803 & n3875 ) ;
  assign n3877 = ( ~n3793 & n3803 ) | ( ~n3793 & n3875 ) | ( n3803 & n3875 ) ;
  assign n3878 = ( n3793 & ~n3876 ) | ( n3793 & n3877 ) | ( ~n3876 & n3877 ) ;
  assign n3879 = ( ~n3806 & n3831 ) | ( ~n3806 & n3878 ) | ( n3831 & n3878 ) ;
  assign n3880 = ( n3806 & n3831 ) | ( n3806 & n3878 ) | ( n3831 & n3878 ) ;
  assign n3881 = ( n3806 & n3879 ) | ( n3806 & ~n3880 ) | ( n3879 & ~n3880 ) ;
  assign n3882 = x19 & x42 ;
  assign n3883 = x7 & x54 ;
  assign n3884 = x8 & x53 ;
  assign n3885 = ( ~n3882 & n3883 ) | ( ~n3882 & n3884 ) | ( n3883 & n3884 ) ;
  assign n3886 = ( n3882 & n3883 ) | ( n3882 & n3884 ) | ( n3883 & n3884 ) ;
  assign n3887 = ( n3882 & n3885 ) | ( n3882 & ~n3886 ) | ( n3885 & ~n3886 ) ;
  assign n3888 = x18 & x43 ;
  assign n3889 = x9 & x52 ;
  assign n3890 = x17 & x44 ;
  assign n3891 = ( ~n3888 & n3889 ) | ( ~n3888 & n3890 ) | ( n3889 & n3890 ) ;
  assign n3892 = ( n3888 & n3889 ) | ( n3888 & n3890 ) | ( n3889 & n3890 ) ;
  assign n3893 = ( n3888 & n3891 ) | ( n3888 & ~n3892 ) | ( n3891 & ~n3892 ) ;
  assign n3894 = x26 & x35 ;
  assign n3895 = x27 & x34 ;
  assign n3896 = x28 & x33 ;
  assign n3897 = ( ~n3894 & n3895 ) | ( ~n3894 & n3896 ) | ( n3895 & n3896 ) ;
  assign n3898 = ( n3894 & n3895 ) | ( n3894 & n3896 ) | ( n3895 & n3896 ) ;
  assign n3899 = ( n3894 & n3897 ) | ( n3894 & ~n3898 ) | ( n3897 & ~n3898 ) ;
  assign n3900 = ( n3887 & n3893 ) | ( n3887 & n3899 ) | ( n3893 & n3899 ) ;
  assign n3901 = ( ~n3887 & n3893 ) | ( ~n3887 & n3899 ) | ( n3893 & n3899 ) ;
  assign n3902 = ( n3887 & ~n3900 ) | ( n3887 & n3901 ) | ( ~n3900 & n3901 ) ;
  assign n3903 = ( n3781 & n3791 ) | ( n3781 & n3902 ) | ( n3791 & n3902 ) ;
  assign n3904 = ( ~n3781 & n3791 ) | ( ~n3781 & n3902 ) | ( n3791 & n3902 ) ;
  assign n3905 = ( n3781 & ~n3903 ) | ( n3781 & n3904 ) | ( ~n3903 & n3904 ) ;
  assign n3906 = x1 & x60 ;
  assign n3907 = x31 & ~n3698 ;
  assign n3908 = ( ~n3717 & n3906 ) | ( ~n3717 & n3907 ) | ( n3906 & n3907 ) ;
  assign n3909 = ( n3717 & n3906 ) | ( n3717 & n3907 ) | ( n3906 & n3907 ) ;
  assign n3910 = ( n3717 & n3908 ) | ( n3717 & ~n3909 ) | ( n3908 & ~n3909 ) ;
  assign n3911 = ( ~n3749 & n3785 ) | ( ~n3749 & n3910 ) | ( n3785 & n3910 ) ;
  assign n3912 = ( n3749 & n3785 ) | ( n3749 & n3910 ) | ( n3785 & n3910 ) ;
  assign n3913 = ( n3749 & n3911 ) | ( n3749 & ~n3912 ) | ( n3911 & ~n3912 ) ;
  assign n3914 = x23 & x38 ;
  assign n3915 = x4 & x57 ;
  assign n3916 = x3 & x58 ;
  assign n3917 = ( ~n3914 & n3915 ) | ( ~n3914 & n3916 ) | ( n3915 & n3916 ) ;
  assign n3918 = ( n3914 & n3915 ) | ( n3914 & n3916 ) | ( n3915 & n3916 ) ;
  assign n3919 = ( n3914 & n3917 ) | ( n3914 & ~n3918 ) | ( n3917 & ~n3918 ) ;
  assign n3920 = ( ~n3778 & n3788 ) | ( ~n3778 & n3919 ) | ( n3788 & n3919 ) ;
  assign n3921 = ( n3778 & n3788 ) | ( n3778 & n3919 ) | ( n3788 & n3919 ) ;
  assign n3922 = ( n3778 & n3920 ) | ( n3778 & ~n3921 ) | ( n3920 & ~n3921 ) ;
  assign n3923 = ( n3773 & n3913 ) | ( n3773 & n3922 ) | ( n3913 & n3922 ) ;
  assign n3924 = ( ~n3773 & n3913 ) | ( ~n3773 & n3922 ) | ( n3913 & n3922 ) ;
  assign n3925 = ( n3773 & ~n3923 ) | ( n3773 & n3924 ) | ( ~n3923 & n3924 ) ;
  assign n3926 = ( ~n3775 & n3905 ) | ( ~n3775 & n3925 ) | ( n3905 & n3925 ) ;
  assign n3927 = ( n3775 & n3905 ) | ( n3775 & n3925 ) | ( n3905 & n3925 ) ;
  assign n3928 = ( n3775 & n3926 ) | ( n3775 & ~n3927 ) | ( n3926 & ~n3927 ) ;
  assign n3929 = ( ~n3797 & n3881 ) | ( ~n3797 & n3928 ) | ( n3881 & n3928 ) ;
  assign n3930 = ( n3797 & n3881 ) | ( n3797 & n3928 ) | ( n3881 & n3928 ) ;
  assign n3931 = ( n3797 & n3929 ) | ( n3797 & ~n3930 ) | ( n3929 & ~n3930 ) ;
  assign n3932 = ( n3809 & n3811 ) | ( n3809 & n3931 ) | ( n3811 & n3931 ) ;
  assign n3933 = ( ~n3809 & n3811 ) | ( ~n3809 & n3931 ) | ( n3811 & n3931 ) ;
  assign n3934 = ( n3809 & ~n3932 ) | ( n3809 & n3933 ) | ( ~n3932 & n3933 ) ;
  assign n3935 = x3 & x59 ;
  assign n3936 = x4 & x58 ;
  assign n3937 = x5 & x57 ;
  assign n3938 = ( ~n3935 & n3936 ) | ( ~n3935 & n3937 ) | ( n3936 & n3937 ) ;
  assign n3939 = ( n3935 & n3936 ) | ( n3935 & n3937 ) | ( n3936 & n3937 ) ;
  assign n3940 = ( n3935 & n3938 ) | ( n3935 & ~n3939 ) | ( n3938 & ~n3939 ) ;
  assign n3941 = ( ~n3868 & n3892 ) | ( ~n3868 & n3940 ) | ( n3892 & n3940 ) ;
  assign n3942 = ( n3868 & n3892 ) | ( n3868 & n3940 ) | ( n3892 & n3940 ) ;
  assign n3943 = ( n3868 & n3941 ) | ( n3868 & ~n3942 ) | ( n3941 & ~n3942 ) ;
  assign n3944 = ( ~n3900 & n3921 ) | ( ~n3900 & n3943 ) | ( n3921 & n3943 ) ;
  assign n3945 = ( n3900 & n3921 ) | ( n3900 & n3943 ) | ( n3921 & n3943 ) ;
  assign n3946 = ( n3900 & n3944 ) | ( n3900 & ~n3945 ) | ( n3944 & ~n3945 ) ;
  assign n3947 = ( n3698 & ~n3908 ) | ( n3698 & n3909 ) | ( ~n3908 & n3909 ) ;
  assign n3948 = ( n3815 & n3824 ) | ( n3815 & n3947 ) | ( n3824 & n3947 ) ;
  assign n3949 = ( ~n3815 & n3824 ) | ( ~n3815 & n3947 ) | ( n3824 & n3947 ) ;
  assign n3950 = ( n3815 & ~n3948 ) | ( n3815 & n3949 ) | ( ~n3948 & n3949 ) ;
  assign n3951 = ( ~n3874 & n3946 ) | ( ~n3874 & n3950 ) | ( n3946 & n3950 ) ;
  assign n3952 = ( n3874 & n3946 ) | ( n3874 & n3950 ) | ( n3946 & n3950 ) ;
  assign n3953 = ( n3874 & n3951 ) | ( n3874 & ~n3952 ) | ( n3951 & ~n3952 ) ;
  assign n3954 = x22 & x40 ;
  assign n3955 = x23 & x39 ;
  assign n3956 = x24 & x38 ;
  assign n3957 = ( ~n3954 & n3955 ) | ( ~n3954 & n3956 ) | ( n3955 & n3956 ) ;
  assign n3958 = ( n3954 & n3955 ) | ( n3954 & n3956 ) | ( n3955 & n3956 ) ;
  assign n3959 = ( n3954 & n3957 ) | ( n3954 & ~n3958 ) | ( n3957 & ~n3958 ) ;
  assign n3960 = x27 & x35 ;
  assign n3961 = x28 & x34 ;
  assign n3962 = x29 & x33 ;
  assign n3963 = ( ~n3960 & n3961 ) | ( ~n3960 & n3962 ) | ( n3961 & n3962 ) ;
  assign n3964 = ( n3960 & n3961 ) | ( n3960 & n3962 ) | ( n3961 & n3962 ) ;
  assign n3965 = ( n3960 & n3963 ) | ( n3960 & ~n3964 ) | ( n3963 & ~n3964 ) ;
  assign n3966 = x19 & x43 ;
  assign n3967 = x8 & x54 ;
  assign n3968 = x18 & x44 ;
  assign n3969 = ( ~n3966 & n3967 ) | ( ~n3966 & n3968 ) | ( n3967 & n3968 ) ;
  assign n3970 = ( n3966 & n3967 ) | ( n3966 & n3968 ) | ( n3967 & n3968 ) ;
  assign n3971 = ( n3966 & n3969 ) | ( n3966 & ~n3970 ) | ( n3969 & ~n3970 ) ;
  assign n3972 = ( ~n3959 & n3965 ) | ( ~n3959 & n3971 ) | ( n3965 & n3971 ) ;
  assign n3973 = ( n3959 & n3965 ) | ( n3959 & n3971 ) | ( n3965 & n3971 ) ;
  assign n3974 = ( n3959 & n3972 ) | ( n3959 & ~n3973 ) | ( n3972 & ~n3973 ) ;
  assign n3975 = x31 & n3906 ;
  assign n3976 = x0 & x62 ;
  assign n3977 = x2 & x60 ;
  assign n3978 = ( ~n3975 & n3976 ) | ( ~n3975 & n3977 ) | ( n3976 & n3977 ) ;
  assign n3979 = ( n3975 & n3976 ) | ( n3975 & n3977 ) | ( n3976 & n3977 ) ;
  assign n3980 = ( n3975 & n3978 ) | ( n3975 & ~n3979 ) | ( n3978 & ~n3979 ) ;
  assign n3981 = x9 & x53 ;
  assign n3982 = x10 & x52 ;
  assign n3983 = x17 & x45 ;
  assign n3984 = ( ~n3981 & n3982 ) | ( ~n3981 & n3983 ) | ( n3982 & n3983 ) ;
  assign n3985 = ( n3981 & n3982 ) | ( n3981 & n3983 ) | ( n3982 & n3983 ) ;
  assign n3986 = ( n3981 & n3984 ) | ( n3981 & ~n3985 ) | ( n3984 & ~n3985 ) ;
  assign n3987 = x21 & x41 ;
  assign n3988 = x25 & x37 ;
  assign n3989 = x26 & x36 ;
  assign n3990 = ( ~n3987 & n3988 ) | ( ~n3987 & n3989 ) | ( n3988 & n3989 ) ;
  assign n3991 = ( n3987 & n3988 ) | ( n3987 & n3989 ) | ( n3988 & n3989 ) ;
  assign n3992 = ( n3987 & n3990 ) | ( n3987 & ~n3991 ) | ( n3990 & ~n3991 ) ;
  assign n3993 = ( ~n3980 & n3986 ) | ( ~n3980 & n3992 ) | ( n3986 & n3992 ) ;
  assign n3994 = ( n3980 & n3986 ) | ( n3980 & n3992 ) | ( n3986 & n3992 ) ;
  assign n3995 = ( n3980 & n3993 ) | ( n3980 & ~n3994 ) | ( n3993 & ~n3994 ) ;
  assign n3996 = x12 & x50 ;
  assign n3997 = x13 & x49 ;
  assign n3998 = x14 & x48 ;
  assign n3999 = ( ~n3996 & n3997 ) | ( ~n3996 & n3998 ) | ( n3997 & n3998 ) ;
  assign n4000 = ( n3996 & n3997 ) | ( n3996 & n3998 ) | ( n3997 & n3998 ) ;
  assign n4001 = ( n3996 & n3999 ) | ( n3996 & ~n4000 ) | ( n3999 & ~n4000 ) ;
  assign n4002 = x20 & x42 ;
  assign n4003 = x6 & x56 ;
  assign n4004 = x7 & x55 ;
  assign n4005 = ( ~n4002 & n4003 ) | ( ~n4002 & n4004 ) | ( n4003 & n4004 ) ;
  assign n4006 = ( n4002 & n4003 ) | ( n4002 & n4004 ) | ( n4003 & n4004 ) ;
  assign n4007 = ( n4002 & n4005 ) | ( n4002 & ~n4006 ) | ( n4005 & ~n4006 ) ;
  assign n4008 = x16 & x46 ;
  assign n4009 = x15 & x47 ;
  assign n4010 = x11 & x51 ;
  assign n4011 = ( ~n4008 & n4009 ) | ( ~n4008 & n4010 ) | ( n4009 & n4010 ) ;
  assign n4012 = ( n4008 & n4009 ) | ( n4008 & n4010 ) | ( n4009 & n4010 ) ;
  assign n4013 = ( n4008 & n4011 ) | ( n4008 & ~n4012 ) | ( n4011 & ~n4012 ) ;
  assign n4014 = ( ~n4001 & n4007 ) | ( ~n4001 & n4013 ) | ( n4007 & n4013 ) ;
  assign n4015 = ( n4001 & n4007 ) | ( n4001 & n4013 ) | ( n4007 & n4013 ) ;
  assign n4016 = ( n4001 & n4014 ) | ( n4001 & ~n4015 ) | ( n4014 & ~n4015 ) ;
  assign n4017 = ( ~n3974 & n3995 ) | ( ~n3974 & n4016 ) | ( n3995 & n4016 ) ;
  assign n4018 = ( n3974 & n3995 ) | ( n3974 & n4016 ) | ( n3995 & n4016 ) ;
  assign n4019 = ( n3974 & n4017 ) | ( n3974 & ~n4018 ) | ( n4017 & ~n4018 ) ;
  assign n4020 = ( n3830 & n3923 ) | ( n3830 & n4019 ) | ( n3923 & n4019 ) ;
  assign n4021 = ( ~n3830 & n3923 ) | ( ~n3830 & n4019 ) | ( n3923 & n4019 ) ;
  assign n4022 = ( n3830 & ~n4020 ) | ( n3830 & n4021 ) | ( ~n4020 & n4021 ) ;
  assign n4023 = ( ~n3927 & n3953 ) | ( ~n3927 & n4022 ) | ( n3953 & n4022 ) ;
  assign n4024 = ( n3927 & n3953 ) | ( n3927 & n4022 ) | ( n3953 & n4022 ) ;
  assign n4025 = ( n3927 & n4023 ) | ( n3927 & ~n4024 ) | ( n4023 & ~n4024 ) ;
  assign n4026 = ( ~n3821 & n3850 ) | ( ~n3821 & n3871 ) | ( n3850 & n3871 ) ;
  assign n4027 = ( n3821 & n3850 ) | ( n3821 & n3871 ) | ( n3850 & n3871 ) ;
  assign n4028 = ( n3821 & n4026 ) | ( n3821 & ~n4027 ) | ( n4026 & ~n4027 ) ;
  assign n4029 = ( n3836 & ~n3847 ) | ( n3836 & n3886 ) | ( ~n3847 & n3886 ) ;
  assign n4030 = ( n3836 & n3847 ) | ( n3836 & n3886 ) | ( n3847 & n3886 ) ;
  assign n4031 = ( n3847 & n4029 ) | ( n3847 & ~n4030 ) | ( n4029 & ~n4030 ) ;
  assign n4032 = ( n3842 & ~n3898 ) | ( n3842 & n3918 ) | ( ~n3898 & n3918 ) ;
  assign n4033 = ( n3842 & n3898 ) | ( n3842 & n3918 ) | ( n3898 & n3918 ) ;
  assign n4034 = ( n3898 & n4032 ) | ( n3898 & ~n4033 ) | ( n4032 & ~n4033 ) ;
  assign n4035 = x30 & x32 ;
  assign n4036 = x1 & x61 ;
  assign n4037 = n4035 & n4036 ;
  assign n4038 = n4035 | n4036 ;
  assign n4039 = ~n4037 & n4038 ;
  assign n4040 = ( ~n3856 & n3862 ) | ( ~n3856 & n4039 ) | ( n3862 & n4039 ) ;
  assign n4041 = ( n3856 & n3862 ) | ( n3856 & n4039 ) | ( n3862 & n4039 ) ;
  assign n4042 = ( n3856 & n4040 ) | ( n3856 & ~n4041 ) | ( n4040 & ~n4041 ) ;
  assign n4043 = ( n4031 & n4034 ) | ( n4031 & n4042 ) | ( n4034 & n4042 ) ;
  assign n4044 = ( ~n4031 & n4034 ) | ( ~n4031 & n4042 ) | ( n4034 & n4042 ) ;
  assign n4045 = ( n4031 & ~n4043 ) | ( n4031 & n4044 ) | ( ~n4043 & n4044 ) ;
  assign n4046 = ( ~n3903 & n4028 ) | ( ~n3903 & n4045 ) | ( n4028 & n4045 ) ;
  assign n4047 = ( n3903 & n4028 ) | ( n3903 & n4045 ) | ( n4028 & n4045 ) ;
  assign n4048 = ( n3903 & n4046 ) | ( n3903 & ~n4047 ) | ( n4046 & ~n4047 ) ;
  assign n4049 = ( n3818 & n3826 ) | ( n3818 & n3912 ) | ( n3826 & n3912 ) ;
  assign n4050 = ( n3818 & ~n3826 ) | ( n3818 & n3912 ) | ( ~n3826 & n3912 ) ;
  assign n4051 = ( n3826 & ~n4049 ) | ( n3826 & n4050 ) | ( ~n4049 & n4050 ) ;
  assign n4052 = ( ~n3876 & n4048 ) | ( ~n3876 & n4051 ) | ( n4048 & n4051 ) ;
  assign n4053 = ( n3876 & n4048 ) | ( n3876 & n4051 ) | ( n4048 & n4051 ) ;
  assign n4054 = ( n3876 & n4052 ) | ( n3876 & ~n4053 ) | ( n4052 & ~n4053 ) ;
  assign n4055 = ( ~n3880 & n4025 ) | ( ~n3880 & n4054 ) | ( n4025 & n4054 ) ;
  assign n4056 = ( n3880 & n4025 ) | ( n3880 & n4054 ) | ( n4025 & n4054 ) ;
  assign n4057 = ( n3880 & n4055 ) | ( n3880 & ~n4056 ) | ( n4055 & ~n4056 ) ;
  assign n4058 = ( n3930 & n3932 ) | ( n3930 & n4057 ) | ( n3932 & n4057 ) ;
  assign n4059 = ( ~n3930 & n3932 ) | ( ~n3930 & n4057 ) | ( n3932 & n4057 ) ;
  assign n4060 = ( n3930 & ~n4058 ) | ( n3930 & n4059 ) | ( ~n4058 & n4059 ) ;
  assign n4061 = ( n3964 & ~n3970 ) | ( n3964 & n3985 ) | ( ~n3970 & n3985 ) ;
  assign n4062 = ( n3964 & n3970 ) | ( n3964 & n3985 ) | ( n3970 & n3985 ) ;
  assign n4063 = ( n3970 & n4061 ) | ( n3970 & ~n4062 ) | ( n4061 & ~n4062 ) ;
  assign n4064 = ( n3973 & n4015 ) | ( n3973 & n4063 ) | ( n4015 & n4063 ) ;
  assign n4065 = ( ~n3973 & n4015 ) | ( ~n3973 & n4063 ) | ( n4015 & n4063 ) ;
  assign n4066 = ( n3973 & ~n4064 ) | ( n3973 & n4065 ) | ( ~n4064 & n4065 ) ;
  assign n4067 = ~x1 & x32 ;
  assign n4068 = ( x1 & x32 ) | ( x1 & x62 ) | ( x32 & x62 ) ;
  assign n4069 = x32 & x62 ;
  assign n4070 = ( n4067 & n4068 ) | ( n4067 & ~n4069 ) | ( n4068 & ~n4069 ) ;
  assign n4071 = x0 & x63 ;
  assign n4072 = ( n4037 & n4070 ) | ( n4037 & n4071 ) | ( n4070 & n4071 ) ;
  assign n4073 = ( ~n4037 & n4070 ) | ( ~n4037 & n4071 ) | ( n4070 & n4071 ) ;
  assign n4074 = ( n4037 & ~n4072 ) | ( n4037 & n4073 ) | ( ~n4072 & n4073 ) ;
  assign n4075 = x27 & x36 ;
  assign n4076 = x29 & x34 ;
  assign n4077 = x28 & x35 ;
  assign n4078 = ( ~n4075 & n4076 ) | ( ~n4075 & n4077 ) | ( n4076 & n4077 ) ;
  assign n4079 = ( n4075 & n4076 ) | ( n4075 & n4077 ) | ( n4076 & n4077 ) ;
  assign n4080 = ( n4075 & n4078 ) | ( n4075 & ~n4079 ) | ( n4078 & ~n4079 ) ;
  assign n4081 = x24 & x39 ;
  assign n4082 = x26 & x37 ;
  assign n4083 = x25 & x38 ;
  assign n4084 = ( ~n4081 & n4082 ) | ( ~n4081 & n4083 ) | ( n4082 & n4083 ) ;
  assign n4085 = ( n4081 & n4082 ) | ( n4081 & n4083 ) | ( n4082 & n4083 ) ;
  assign n4086 = ( n4081 & n4084 ) | ( n4081 & ~n4085 ) | ( n4084 & ~n4085 ) ;
  assign n4087 = ( ~n4074 & n4080 ) | ( ~n4074 & n4086 ) | ( n4080 & n4086 ) ;
  assign n4088 = ( n4074 & n4080 ) | ( n4074 & n4086 ) | ( n4080 & n4086 ) ;
  assign n4089 = ( n4074 & n4087 ) | ( n4074 & ~n4088 ) | ( n4087 & ~n4088 ) ;
  assign n4090 = ( ~n3948 & n3994 ) | ( ~n3948 & n4089 ) | ( n3994 & n4089 ) ;
  assign n4091 = ( n3948 & n3994 ) | ( n3948 & n4089 ) | ( n3994 & n4089 ) ;
  assign n4092 = ( n3948 & n4090 ) | ( n3948 & ~n4091 ) | ( n4090 & ~n4091 ) ;
  assign n4093 = ( ~n4049 & n4066 ) | ( ~n4049 & n4092 ) | ( n4066 & n4092 ) ;
  assign n4094 = ( n4049 & n4066 ) | ( n4049 & n4092 ) | ( n4066 & n4092 ) ;
  assign n4095 = ( n4049 & n4093 ) | ( n4049 & ~n4094 ) | ( n4093 & ~n4094 ) ;
  assign n4096 = x5 & x58 ;
  assign n4097 = x21 & x42 ;
  assign n4098 = x22 & x41 ;
  assign n4099 = ( ~n4096 & n4097 ) | ( ~n4096 & n4098 ) | ( n4097 & n4098 ) ;
  assign n4100 = ( n4096 & n4097 ) | ( n4096 & n4098 ) | ( n4097 & n4098 ) ;
  assign n4101 = ( n4096 & n4099 ) | ( n4096 & ~n4100 ) | ( n4099 & ~n4100 ) ;
  assign n4102 = x2 & x61 ;
  assign n4103 = x3 & x60 ;
  assign n4104 = x4 & x59 ;
  assign n4105 = ( ~n4102 & n4103 ) | ( ~n4102 & n4104 ) | ( n4103 & n4104 ) ;
  assign n4106 = ( n4102 & n4103 ) | ( n4102 & n4104 ) | ( n4103 & n4104 ) ;
  assign n4107 = ( n4102 & n4105 ) | ( n4102 & ~n4106 ) | ( n4105 & ~n4106 ) ;
  assign n4108 = ( n4012 & n4101 ) | ( n4012 & n4107 ) | ( n4101 & n4107 ) ;
  assign n4109 = ( ~n4012 & n4101 ) | ( ~n4012 & n4107 ) | ( n4101 & n4107 ) ;
  assign n4110 = ( n4012 & ~n4108 ) | ( n4012 & n4109 ) | ( ~n4108 & n4109 ) ;
  assign n4111 = x15 & x48 ;
  assign n4112 = x12 & x51 ;
  assign n4113 = x13 & x50 ;
  assign n4114 = ( ~n4111 & n4112 ) | ( ~n4111 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4115 = ( n4111 & n4112 ) | ( n4111 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4116 = ( n4111 & n4114 ) | ( n4111 & ~n4115 ) | ( n4114 & ~n4115 ) ;
  assign n4117 = x10 & x53 ;
  assign n4118 = x11 & x52 ;
  assign n4119 = x16 & x47 ;
  assign n4120 = ( ~n4117 & n4118 ) | ( ~n4117 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4121 = ( n4117 & n4118 ) | ( n4117 & n4119 ) | ( n4118 & n4119 ) ;
  assign n4122 = ( n4117 & n4120 ) | ( n4117 & ~n4121 ) | ( n4120 & ~n4121 ) ;
  assign n4123 = x18 & x45 ;
  assign n4124 = x17 & x46 ;
  assign n4125 = x9 & x54 ;
  assign n4126 = ( ~n4123 & n4124 ) | ( ~n4123 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4127 = ( n4123 & n4124 ) | ( n4123 & n4125 ) | ( n4124 & n4125 ) ;
  assign n4128 = ( n4123 & n4126 ) | ( n4123 & ~n4127 ) | ( n4126 & ~n4127 ) ;
  assign n4129 = ( ~n4116 & n4122 ) | ( ~n4116 & n4128 ) | ( n4122 & n4128 ) ;
  assign n4130 = ( n4116 & n4122 ) | ( n4116 & n4128 ) | ( n4122 & n4128 ) ;
  assign n4131 = ( n4116 & n4129 ) | ( n4116 & ~n4130 ) | ( n4129 & ~n4130 ) ;
  assign n4132 = x23 & x40 ;
  assign n4133 = x6 & x57 ;
  assign n4134 = x20 & x43 ;
  assign n4135 = ( ~n4132 & n4133 ) | ( ~n4132 & n4134 ) | ( n4133 & n4134 ) ;
  assign n4136 = ( n4132 & n4133 ) | ( n4132 & n4134 ) | ( n4133 & n4134 ) ;
  assign n4137 = ( n4132 & n4135 ) | ( n4132 & ~n4136 ) | ( n4135 & ~n4136 ) ;
  assign n4138 = x7 & x56 ;
  assign n4139 = x8 & x55 ;
  assign n4140 = x19 & x44 ;
  assign n4141 = ( ~n4138 & n4139 ) | ( ~n4138 & n4140 ) | ( n4139 & n4140 ) ;
  assign n4142 = ( n4138 & n4139 ) | ( n4138 & n4140 ) | ( n4139 & n4140 ) ;
  assign n4143 = ( n4138 & n4141 ) | ( n4138 & ~n4142 ) | ( n4141 & ~n4142 ) ;
  assign n4144 = x14 & x49 ;
  assign n4145 = x31 & x32 ;
  assign n4146 = x30 & x33 ;
  assign n4147 = ( ~n4144 & n4145 ) | ( ~n4144 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4148 = ( n4144 & n4145 ) | ( n4144 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4149 = ( n4144 & n4147 ) | ( n4144 & ~n4148 ) | ( n4147 & ~n4148 ) ;
  assign n4150 = ( ~n4137 & n4143 ) | ( ~n4137 & n4149 ) | ( n4143 & n4149 ) ;
  assign n4151 = ( n4137 & n4143 ) | ( n4137 & n4149 ) | ( n4143 & n4149 ) ;
  assign n4152 = ( n4137 & n4150 ) | ( n4137 & ~n4151 ) | ( n4150 & ~n4151 ) ;
  assign n4153 = ( n4110 & n4131 ) | ( n4110 & n4152 ) | ( n4131 & n4152 ) ;
  assign n4154 = ( ~n4110 & n4131 ) | ( ~n4110 & n4152 ) | ( n4131 & n4152 ) ;
  assign n4155 = ( n4110 & ~n4153 ) | ( n4110 & n4154 ) | ( ~n4153 & n4154 ) ;
  assign n4156 = ( ~n3952 & n4047 ) | ( ~n3952 & n4155 ) | ( n4047 & n4155 ) ;
  assign n4157 = ( n3952 & n4047 ) | ( n3952 & n4155 ) | ( n4047 & n4155 ) ;
  assign n4158 = ( n3952 & n4156 ) | ( n3952 & ~n4157 ) | ( n4156 & ~n4157 ) ;
  assign n4159 = ( ~n4053 & n4095 ) | ( ~n4053 & n4158 ) | ( n4095 & n4158 ) ;
  assign n4160 = ( n4053 & n4095 ) | ( n4053 & n4158 ) | ( n4095 & n4158 ) ;
  assign n4161 = ( n4053 & n4159 ) | ( n4053 & ~n4160 ) | ( n4159 & ~n4160 ) ;
  assign n4162 = ( n3945 & n4027 ) | ( n3945 & ~n4043 ) | ( n4027 & ~n4043 ) ;
  assign n4163 = ( n3945 & n4027 ) | ( n3945 & n4043 ) | ( n4027 & n4043 ) ;
  assign n4164 = ( n4043 & n4162 ) | ( n4043 & ~n4163 ) | ( n4162 & ~n4163 ) ;
  assign n4165 = ( n3942 & ~n4033 ) | ( n3942 & n4041 ) | ( ~n4033 & n4041 ) ;
  assign n4166 = ( n3942 & n4033 ) | ( n3942 & n4041 ) | ( n4033 & n4041 ) ;
  assign n4167 = ( n4033 & n4165 ) | ( n4033 & ~n4166 ) | ( n4165 & ~n4166 ) ;
  assign n4168 = ( n3939 & ~n3979 ) | ( n3939 & n3991 ) | ( ~n3979 & n3991 ) ;
  assign n4169 = ( n3939 & n3979 ) | ( n3939 & n3991 ) | ( n3979 & n3991 ) ;
  assign n4170 = ( n3979 & n4168 ) | ( n3979 & ~n4169 ) | ( n4168 & ~n4169 ) ;
  assign n4171 = ( n3958 & n4000 ) | ( n3958 & ~n4006 ) | ( n4000 & ~n4006 ) ;
  assign n4172 = ( n3958 & n4000 ) | ( n3958 & n4006 ) | ( n4000 & n4006 ) ;
  assign n4173 = ( n4006 & n4171 ) | ( n4006 & ~n4172 ) | ( n4171 & ~n4172 ) ;
  assign n4174 = ( ~n4030 & n4170 ) | ( ~n4030 & n4173 ) | ( n4170 & n4173 ) ;
  assign n4175 = ( n4030 & n4170 ) | ( n4030 & n4173 ) | ( n4170 & n4173 ) ;
  assign n4176 = ( n4030 & n4174 ) | ( n4030 & ~n4175 ) | ( n4174 & ~n4175 ) ;
  assign n4177 = ( ~n4018 & n4167 ) | ( ~n4018 & n4176 ) | ( n4167 & n4176 ) ;
  assign n4178 = ( n4018 & n4167 ) | ( n4018 & n4176 ) | ( n4167 & n4176 ) ;
  assign n4179 = ( n4018 & n4177 ) | ( n4018 & ~n4178 ) | ( n4177 & ~n4178 ) ;
  assign n4180 = ( ~n4020 & n4164 ) | ( ~n4020 & n4179 ) | ( n4164 & n4179 ) ;
  assign n4181 = ( n4020 & n4164 ) | ( n4020 & n4179 ) | ( n4164 & n4179 ) ;
  assign n4182 = ( n4020 & n4180 ) | ( n4020 & ~n4181 ) | ( n4180 & ~n4181 ) ;
  assign n4183 = ( n4024 & n4161 ) | ( n4024 & n4182 ) | ( n4161 & n4182 ) ;
  assign n4184 = ( ~n4024 & n4161 ) | ( ~n4024 & n4182 ) | ( n4161 & n4182 ) ;
  assign n4185 = ( n4024 & ~n4183 ) | ( n4024 & n4184 ) | ( ~n4183 & n4184 ) ;
  assign n4186 = ( n4056 & n4058 ) | ( n4056 & n4185 ) | ( n4058 & n4185 ) ;
  assign n4187 = ( ~n4056 & n4058 ) | ( ~n4056 & n4185 ) | ( n4058 & n4185 ) ;
  assign n4188 = ( n4056 & ~n4186 ) | ( n4056 & n4187 ) | ( ~n4186 & n4187 ) ;
  assign n4189 = ( ~n4085 & n4115 ) | ( ~n4085 & n4121 ) | ( n4115 & n4121 ) ;
  assign n4190 = ( n4085 & n4115 ) | ( n4085 & n4121 ) | ( n4115 & n4121 ) ;
  assign n4191 = ( n4085 & n4189 ) | ( n4085 & ~n4190 ) | ( n4189 & ~n4190 ) ;
  assign n4192 = ( n4130 & n4151 ) | ( n4130 & n4191 ) | ( n4151 & n4191 ) ;
  assign n4193 = ( ~n4130 & n4151 ) | ( ~n4130 & n4191 ) | ( n4151 & n4191 ) ;
  assign n4194 = ( n4130 & ~n4192 ) | ( n4130 & n4193 ) | ( ~n4192 & n4193 ) ;
  assign n4195 = x62 & n1206 ;
  assign n4196 = x1 & x63 ;
  assign n4197 = ( n4148 & n4195 ) | ( n4148 & n4196 ) | ( n4195 & n4196 ) ;
  assign n4198 = ( n4148 & ~n4195 ) | ( n4148 & n4196 ) | ( ~n4195 & n4196 ) ;
  assign n4199 = ( n4195 & ~n4197 ) | ( n4195 & n4198 ) | ( ~n4197 & n4198 ) ;
  assign n4200 = x13 & x51 ;
  assign n4201 = x11 & x53 ;
  assign n4202 = x12 & x52 ;
  assign n4203 = ( ~n4200 & n4201 ) | ( ~n4200 & n4202 ) | ( n4201 & n4202 ) ;
  assign n4204 = ( n4200 & n4201 ) | ( n4200 & n4202 ) | ( n4201 & n4202 ) ;
  assign n4205 = ( n4200 & n4203 ) | ( n4200 & ~n4204 ) | ( n4203 & ~n4204 ) ;
  assign n4206 = x15 & x49 ;
  assign n4207 = x9 & x55 ;
  assign n4208 = x10 & x54 ;
  assign n4209 = ( ~n4206 & n4207 ) | ( ~n4206 & n4208 ) | ( n4207 & n4208 ) ;
  assign n4210 = ( n4206 & n4207 ) | ( n4206 & n4208 ) | ( n4207 & n4208 ) ;
  assign n4211 = ( n4206 & n4209 ) | ( n4206 & ~n4210 ) | ( n4209 & ~n4210 ) ;
  assign n4212 = ( n4199 & n4205 ) | ( n4199 & n4211 ) | ( n4205 & n4211 ) ;
  assign n4213 = ( ~n4199 & n4205 ) | ( ~n4199 & n4211 ) | ( n4205 & n4211 ) ;
  assign n4214 = ( n4199 & ~n4212 ) | ( n4199 & n4213 ) | ( ~n4212 & n4213 ) ;
  assign n4215 = ( n4108 & n4166 ) | ( n4108 & n4214 ) | ( n4166 & n4214 ) ;
  assign n4216 = ( ~n4108 & n4166 ) | ( ~n4108 & n4214 ) | ( n4166 & n4214 ) ;
  assign n4217 = ( n4108 & ~n4215 ) | ( n4108 & n4216 ) | ( ~n4215 & n4216 ) ;
  assign n4218 = ( n4163 & n4194 ) | ( n4163 & n4217 ) | ( n4194 & n4217 ) ;
  assign n4219 = ( ~n4163 & n4194 ) | ( ~n4163 & n4217 ) | ( n4194 & n4217 ) ;
  assign n4220 = ( n4163 & ~n4218 ) | ( n4163 & n4219 ) | ( ~n4218 & n4219 ) ;
  assign n4221 = x2 & x62 ;
  assign n4222 = x4 & x60 ;
  assign n4223 = x3 & x61 ;
  assign n4224 = ( ~n4221 & n4222 ) | ( ~n4221 & n4223 ) | ( n4222 & n4223 ) ;
  assign n4225 = ( n4221 & n4222 ) | ( n4221 & n4223 ) | ( n4222 & n4223 ) ;
  assign n4226 = ( n4221 & n4224 ) | ( n4221 & ~n4225 ) | ( n4224 & ~n4225 ) ;
  assign n4227 = x5 & x59 ;
  assign n4228 = x18 & x46 ;
  assign n4229 = x19 & x45 ;
  assign n4230 = ( ~n4227 & n4228 ) | ( ~n4227 & n4229 ) | ( n4228 & n4229 ) ;
  assign n4231 = ( n4227 & n4228 ) | ( n4227 & n4229 ) | ( n4228 & n4229 ) ;
  assign n4232 = ( n4227 & n4230 ) | ( n4227 & ~n4231 ) | ( n4230 & ~n4231 ) ;
  assign n4233 = ( n4072 & n4226 ) | ( n4072 & n4232 ) | ( n4226 & n4232 ) ;
  assign n4234 = ( ~n4072 & n4226 ) | ( ~n4072 & n4232 ) | ( n4226 & n4232 ) ;
  assign n4235 = ( n4072 & ~n4233 ) | ( n4072 & n4234 ) | ( ~n4233 & n4234 ) ;
  assign n4236 = x23 & x41 ;
  assign n4237 = x24 & x40 ;
  assign n4238 = x25 & x39 ;
  assign n4239 = ( ~n4236 & n4237 ) | ( ~n4236 & n4238 ) | ( n4237 & n4238 ) ;
  assign n4240 = ( n4236 & n4237 ) | ( n4236 & n4238 ) | ( n4237 & n4238 ) ;
  assign n4241 = ( n4236 & n4239 ) | ( n4236 & ~n4240 ) | ( n4239 & ~n4240 ) ;
  assign n4242 = x20 & x44 ;
  assign n4243 = x22 & x42 ;
  assign n4244 = x21 & x43 ;
  assign n4245 = ( ~n4242 & n4243 ) | ( ~n4242 & n4244 ) | ( n4243 & n4244 ) ;
  assign n4246 = ( n4242 & n4243 ) | ( n4242 & n4244 ) | ( n4243 & n4244 ) ;
  assign n4247 = ( n4242 & n4245 ) | ( n4242 & ~n4246 ) | ( n4245 & ~n4246 ) ;
  assign n4248 = x6 & x58 ;
  assign n4249 = x17 & x47 ;
  assign n4250 = x7 & x57 ;
  assign n4251 = ( ~n4248 & n4249 ) | ( ~n4248 & n4250 ) | ( n4249 & n4250 ) ;
  assign n4252 = ( n4248 & n4249 ) | ( n4248 & n4250 ) | ( n4249 & n4250 ) ;
  assign n4253 = ( n4248 & n4251 ) | ( n4248 & ~n4252 ) | ( n4251 & ~n4252 ) ;
  assign n4254 = ( ~n4241 & n4247 ) | ( ~n4241 & n4253 ) | ( n4247 & n4253 ) ;
  assign n4255 = ( n4241 & n4247 ) | ( n4241 & n4253 ) | ( n4247 & n4253 ) ;
  assign n4256 = ( n4241 & n4254 ) | ( n4241 & ~n4255 ) | ( n4254 & ~n4255 ) ;
  assign n4257 = x14 & x50 ;
  assign n4258 = x31 & x33 ;
  assign n4259 = x30 & x34 ;
  assign n4260 = ( ~n4257 & n4258 ) | ( ~n4257 & n4259 ) | ( n4258 & n4259 ) ;
  assign n4261 = ( n4257 & n4258 ) | ( n4257 & n4259 ) | ( n4258 & n4259 ) ;
  assign n4262 = ( n4257 & n4260 ) | ( n4257 & ~n4261 ) | ( n4260 & ~n4261 ) ;
  assign n4263 = x27 & x37 ;
  assign n4264 = x29 & x35 ;
  assign n4265 = x28 & x36 ;
  assign n4266 = ( ~n4263 & n4264 ) | ( ~n4263 & n4265 ) | ( n4264 & n4265 ) ;
  assign n4267 = ( n4263 & n4264 ) | ( n4263 & n4265 ) | ( n4264 & n4265 ) ;
  assign n4268 = ( n4263 & n4266 ) | ( n4263 & ~n4267 ) | ( n4266 & ~n4267 ) ;
  assign n4269 = x26 & x38 ;
  assign n4270 = x16 & x48 ;
  assign n4271 = x8 & x56 ;
  assign n4272 = ( ~n4269 & n4270 ) | ( ~n4269 & n4271 ) | ( n4270 & n4271 ) ;
  assign n4273 = ( n4269 & n4270 ) | ( n4269 & n4271 ) | ( n4270 & n4271 ) ;
  assign n4274 = ( n4269 & n4272 ) | ( n4269 & ~n4273 ) | ( n4272 & ~n4273 ) ;
  assign n4275 = ( ~n4262 & n4268 ) | ( ~n4262 & n4274 ) | ( n4268 & n4274 ) ;
  assign n4276 = ( n4262 & n4268 ) | ( n4262 & n4274 ) | ( n4268 & n4274 ) ;
  assign n4277 = ( n4262 & n4275 ) | ( n4262 & ~n4276 ) | ( n4275 & ~n4276 ) ;
  assign n4278 = ( n4235 & n4256 ) | ( n4235 & n4277 ) | ( n4256 & n4277 ) ;
  assign n4279 = ( ~n4235 & n4256 ) | ( ~n4235 & n4277 ) | ( n4256 & n4277 ) ;
  assign n4280 = ( n4235 & ~n4278 ) | ( n4235 & n4279 ) | ( ~n4278 & n4279 ) ;
  assign n4281 = ( n4062 & n4169 ) | ( n4062 & n4172 ) | ( n4169 & n4172 ) ;
  assign n4282 = ( n4062 & ~n4169 ) | ( n4062 & n4172 ) | ( ~n4169 & n4172 ) ;
  assign n4283 = ( n4169 & ~n4281 ) | ( n4169 & n4282 ) | ( ~n4281 & n4282 ) ;
  assign n4284 = ( ~n4064 & n4175 ) | ( ~n4064 & n4283 ) | ( n4175 & n4283 ) ;
  assign n4285 = ( n4064 & n4175 ) | ( n4064 & n4283 ) | ( n4175 & n4283 ) ;
  assign n4286 = ( n4064 & n4284 ) | ( n4064 & ~n4285 ) | ( n4284 & ~n4285 ) ;
  assign n4287 = ( ~n4178 & n4280 ) | ( ~n4178 & n4286 ) | ( n4280 & n4286 ) ;
  assign n4288 = ( n4178 & n4280 ) | ( n4178 & n4286 ) | ( n4280 & n4286 ) ;
  assign n4289 = ( n4178 & n4287 ) | ( n4178 & ~n4288 ) | ( n4287 & ~n4288 ) ;
  assign n4290 = ( ~n4181 & n4220 ) | ( ~n4181 & n4289 ) | ( n4220 & n4289 ) ;
  assign n4291 = ( n4181 & n4220 ) | ( n4181 & n4289 ) | ( n4220 & n4289 ) ;
  assign n4292 = ( n4181 & n4290 ) | ( n4181 & ~n4291 ) | ( n4290 & ~n4291 ) ;
  assign n4293 = ( n4079 & n4127 ) | ( n4079 & n4136 ) | ( n4127 & n4136 ) ;
  assign n4294 = ( ~n4079 & n4127 ) | ( ~n4079 & n4136 ) | ( n4127 & n4136 ) ;
  assign n4295 = ( n4079 & ~n4293 ) | ( n4079 & n4294 ) | ( ~n4293 & n4294 ) ;
  assign n4296 = ( n4100 & ~n4106 ) | ( n4100 & n4142 ) | ( ~n4106 & n4142 ) ;
  assign n4297 = ( n4100 & n4106 ) | ( n4100 & n4142 ) | ( n4106 & n4142 ) ;
  assign n4298 = ( n4106 & n4296 ) | ( n4106 & ~n4297 ) | ( n4296 & ~n4297 ) ;
  assign n4299 = ( n4088 & n4295 ) | ( n4088 & n4298 ) | ( n4295 & n4298 ) ;
  assign n4300 = ( n4088 & ~n4295 ) | ( n4088 & n4298 ) | ( ~n4295 & n4298 ) ;
  assign n4301 = ( n4295 & ~n4299 ) | ( n4295 & n4300 ) | ( ~n4299 & n4300 ) ;
  assign n4302 = ( n4091 & n4153 ) | ( n4091 & n4301 ) | ( n4153 & n4301 ) ;
  assign n4303 = ( ~n4091 & n4153 ) | ( ~n4091 & n4301 ) | ( n4153 & n4301 ) ;
  assign n4304 = ( n4091 & ~n4302 ) | ( n4091 & n4303 ) | ( ~n4302 & n4303 ) ;
  assign n4305 = ( n4094 & n4157 ) | ( n4094 & n4304 ) | ( n4157 & n4304 ) ;
  assign n4306 = ( ~n4094 & n4157 ) | ( ~n4094 & n4304 ) | ( n4157 & n4304 ) ;
  assign n4307 = ( n4094 & ~n4305 ) | ( n4094 & n4306 ) | ( ~n4305 & n4306 ) ;
  assign n4308 = ( ~n4160 & n4292 ) | ( ~n4160 & n4307 ) | ( n4292 & n4307 ) ;
  assign n4309 = ( n4160 & n4292 ) | ( n4160 & n4307 ) | ( n4292 & n4307 ) ;
  assign n4310 = ( n4160 & n4308 ) | ( n4160 & ~n4309 ) | ( n4308 & ~n4309 ) ;
  assign n4311 = ( ~n4183 & n4186 ) | ( ~n4183 & n4310 ) | ( n4186 & n4310 ) ;
  assign n4312 = ( n4183 & n4186 ) | ( n4183 & n4310 ) | ( n4186 & n4310 ) ;
  assign n4313 = ( n4183 & n4311 ) | ( n4183 & ~n4312 ) | ( n4311 & ~n4312 ) ;
  assign n4314 = ( n4210 & n4240 ) | ( n4210 & n4252 ) | ( n4240 & n4252 ) ;
  assign n4315 = ( n4210 & ~n4240 ) | ( n4210 & n4252 ) | ( ~n4240 & n4252 ) ;
  assign n4316 = ( n4240 & ~n4314 ) | ( n4240 & n4315 ) | ( ~n4314 & n4315 ) ;
  assign n4317 = ( n4225 & ~n4231 ) | ( n4225 & n4273 ) | ( ~n4231 & n4273 ) ;
  assign n4318 = ( n4225 & n4231 ) | ( n4225 & n4273 ) | ( n4231 & n4273 ) ;
  assign n4319 = ( n4231 & n4317 ) | ( n4231 & ~n4318 ) | ( n4317 & ~n4318 ) ;
  assign n4320 = ( ~n4212 & n4316 ) | ( ~n4212 & n4319 ) | ( n4316 & n4319 ) ;
  assign n4321 = ( n4212 & n4316 ) | ( n4212 & n4319 ) | ( n4316 & n4319 ) ;
  assign n4322 = ( n4212 & n4320 ) | ( n4212 & ~n4321 ) | ( n4320 & ~n4321 ) ;
  assign n4323 = ( ~n4215 & n4278 ) | ( ~n4215 & n4322 ) | ( n4278 & n4322 ) ;
  assign n4324 = ( n4215 & n4278 ) | ( n4215 & n4322 ) | ( n4278 & n4322 ) ;
  assign n4325 = ( n4215 & n4323 ) | ( n4215 & ~n4324 ) | ( n4323 & ~n4324 ) ;
  assign n4326 = ( ~n4218 & n4288 ) | ( ~n4218 & n4325 ) | ( n4288 & n4325 ) ;
  assign n4327 = ( n4218 & n4288 ) | ( n4218 & n4325 ) | ( n4288 & n4325 ) ;
  assign n4328 = ( n4218 & n4326 ) | ( n4218 & ~n4327 ) | ( n4326 & ~n4327 ) ;
  assign n4329 = ( n4204 & ~n4246 ) | ( n4204 & n4267 ) | ( ~n4246 & n4267 ) ;
  assign n4330 = ( n4204 & n4246 ) | ( n4204 & n4267 ) | ( n4246 & n4267 ) ;
  assign n4331 = ( n4246 & n4329 ) | ( n4246 & ~n4330 ) | ( n4329 & ~n4330 ) ;
  assign n4332 = ( n4255 & n4276 ) | ( n4255 & n4331 ) | ( n4276 & n4331 ) ;
  assign n4333 = ( ~n4255 & n4276 ) | ( ~n4255 & n4331 ) | ( n4276 & n4331 ) ;
  assign n4334 = ( n4255 & ~n4332 ) | ( n4255 & n4333 ) | ( ~n4332 & n4333 ) ;
  assign n4335 = x4 & x61 ;
  assign n4336 = x2 & x63 ;
  assign n4337 = ( n4261 & n4335 ) | ( n4261 & n4336 ) | ( n4335 & n4336 ) ;
  assign n4338 = ( ~n4261 & n4335 ) | ( ~n4261 & n4336 ) | ( n4335 & n4336 ) ;
  assign n4339 = ( n4261 & ~n4337 ) | ( n4261 & n4338 ) | ( ~n4337 & n4338 ) ;
  assign n4340 = x12 & x53 ;
  assign n4341 = x13 & x52 ;
  assign n4342 = x18 & x47 ;
  assign n4343 = ( ~n4340 & n4341 ) | ( ~n4340 & n4342 ) | ( n4341 & n4342 ) ;
  assign n4344 = ( n4340 & n4341 ) | ( n4340 & n4342 ) | ( n4341 & n4342 ) ;
  assign n4345 = ( n4340 & n4343 ) | ( n4340 & ~n4344 ) | ( n4343 & ~n4344 ) ;
  assign n4346 = x16 & x49 ;
  assign n4347 = x14 & x51 ;
  assign n4348 = x15 & x50 ;
  assign n4349 = ( ~n4346 & n4347 ) | ( ~n4346 & n4348 ) | ( n4347 & n4348 ) ;
  assign n4350 = ( n4346 & n4347 ) | ( n4346 & n4348 ) | ( n4347 & n4348 ) ;
  assign n4351 = ( n4346 & n4349 ) | ( n4346 & ~n4350 ) | ( n4349 & ~n4350 ) ;
  assign n4352 = ( n4339 & n4345 ) | ( n4339 & n4351 ) | ( n4345 & n4351 ) ;
  assign n4353 = ( ~n4339 & n4345 ) | ( ~n4339 & n4351 ) | ( n4345 & n4351 ) ;
  assign n4354 = ( n4339 & ~n4352 ) | ( n4339 & n4353 ) | ( ~n4352 & n4353 ) ;
  assign n4355 = ( n4233 & n4281 ) | ( n4233 & n4354 ) | ( n4281 & n4354 ) ;
  assign n4356 = ( ~n4233 & n4281 ) | ( ~n4233 & n4354 ) | ( n4281 & n4354 ) ;
  assign n4357 = ( n4233 & ~n4355 ) | ( n4233 & n4356 ) | ( ~n4355 & n4356 ) ;
  assign n4358 = ( ~n4285 & n4334 ) | ( ~n4285 & n4357 ) | ( n4334 & n4357 ) ;
  assign n4359 = ( n4285 & n4334 ) | ( n4285 & n4357 ) | ( n4334 & n4357 ) ;
  assign n4360 = ( n4285 & n4358 ) | ( n4285 & ~n4359 ) | ( n4358 & ~n4359 ) ;
  assign n4361 = ( n4190 & ~n4293 ) | ( n4190 & n4297 ) | ( ~n4293 & n4297 ) ;
  assign n4362 = ( n4190 & n4293 ) | ( n4190 & n4297 ) | ( n4293 & n4297 ) ;
  assign n4363 = ( n4293 & n4361 ) | ( n4293 & ~n4362 ) | ( n4361 & ~n4362 ) ;
  assign n4364 = ( n4192 & n4299 ) | ( n4192 & n4363 ) | ( n4299 & n4363 ) ;
  assign n4365 = ( ~n4192 & n4299 ) | ( ~n4192 & n4363 ) | ( n4299 & n4363 ) ;
  assign n4366 = ( n4192 & ~n4364 ) | ( n4192 & n4365 ) | ( ~n4364 & n4365 ) ;
  assign n4367 = x5 & x60 ;
  assign n4368 = x6 & x59 ;
  assign n4369 = x7 & x58 ;
  assign n4370 = ( ~n4367 & n4368 ) | ( ~n4367 & n4369 ) | ( n4368 & n4369 ) ;
  assign n4371 = ( n4367 & n4368 ) | ( n4367 & n4369 ) | ( n4368 & n4369 ) ;
  assign n4372 = ( n4367 & n4370 ) | ( n4367 & ~n4371 ) | ( n4370 & ~n4371 ) ;
  assign n4373 = x8 & x57 ;
  assign n4374 = x22 & x43 ;
  assign n4375 = x21 & x44 ;
  assign n4376 = ( ~n4373 & n4374 ) | ( ~n4373 & n4375 ) | ( n4374 & n4375 ) ;
  assign n4377 = ( n4373 & n4374 ) | ( n4373 & n4375 ) | ( n4374 & n4375 ) ;
  assign n4378 = ( n4373 & n4376 ) | ( n4373 & ~n4377 ) | ( n4376 & ~n4377 ) ;
  assign n4379 = ( n4197 & n4372 ) | ( n4197 & n4378 ) | ( n4372 & n4378 ) ;
  assign n4380 = ( ~n4197 & n4372 ) | ( ~n4197 & n4378 ) | ( n4372 & n4378 ) ;
  assign n4381 = ( n4197 & ~n4379 ) | ( n4197 & n4380 ) | ( ~n4379 & n4380 ) ;
  assign n4382 = x26 & x39 ;
  assign n4383 = x28 & x37 ;
  assign n4384 = x27 & x38 ;
  assign n4385 = ( ~n4382 & n4383 ) | ( ~n4382 & n4384 ) | ( n4383 & n4384 ) ;
  assign n4386 = ( n4382 & n4383 ) | ( n4382 & n4384 ) | ( n4383 & n4384 ) ;
  assign n4387 = ( n4382 & n4385 ) | ( n4382 & ~n4386 ) | ( n4385 & ~n4386 ) ;
  assign n4388 = x9 & x56 ;
  assign n4389 = x10 & x55 ;
  assign n4390 = x20 & x45 ;
  assign n4391 = ( ~n4388 & n4389 ) | ( ~n4388 & n4390 ) | ( n4389 & n4390 ) ;
  assign n4392 = ( n4388 & n4389 ) | ( n4388 & n4390 ) | ( n4389 & n4390 ) ;
  assign n4393 = ( n4388 & n4391 ) | ( n4388 & ~n4392 ) | ( n4391 & ~n4392 ) ;
  assign n4394 = x23 & x42 ;
  assign n4395 = x25 & x40 ;
  assign n4396 = x24 & x41 ;
  assign n4397 = ( ~n4394 & n4395 ) | ( ~n4394 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4398 = ( n4394 & n4395 ) | ( n4394 & n4396 ) | ( n4395 & n4396 ) ;
  assign n4399 = ( n4394 & n4397 ) | ( n4394 & ~n4398 ) | ( n4397 & ~n4398 ) ;
  assign n4400 = ( ~n4387 & n4393 ) | ( ~n4387 & n4399 ) | ( n4393 & n4399 ) ;
  assign n4401 = ( n4387 & n4393 ) | ( n4387 & n4399 ) | ( n4393 & n4399 ) ;
  assign n4402 = ( n4387 & n4400 ) | ( n4387 & ~n4401 ) | ( n4400 & ~n4401 ) ;
  assign n4403 = x30 & x35 ;
  assign n4404 = x31 & x34 ;
  assign n4405 = x32 & x33 ;
  assign n4406 = ( ~n4403 & n4404 ) | ( ~n4403 & n4405 ) | ( n4404 & n4405 ) ;
  assign n4407 = ( n4403 & n4404 ) | ( n4403 & n4405 ) | ( n4404 & n4405 ) ;
  assign n4408 = ( n4403 & n4406 ) | ( n4403 & ~n4407 ) | ( n4406 & ~n4407 ) ;
  assign n4409 = x19 & x46 ;
  assign n4410 = x29 & x36 ;
  assign n4411 = x11 & x54 ;
  assign n4412 = ( ~n4409 & n4410 ) | ( ~n4409 & n4411 ) | ( n4410 & n4411 ) ;
  assign n4413 = ( n4409 & n4410 ) | ( n4409 & n4411 ) | ( n4410 & n4411 ) ;
  assign n4414 = ( n4409 & n4412 ) | ( n4409 & ~n4413 ) | ( n4412 & ~n4413 ) ;
  assign n4415 = x17 & x48 ;
  assign n4416 = x3 & x62 ;
  assign n4417 = ( ~x33 & n4415 ) | ( ~x33 & n4416 ) | ( n4415 & n4416 ) ;
  assign n4418 = ( x33 & n4415 ) | ( x33 & n4416 ) | ( n4415 & n4416 ) ;
  assign n4419 = ( x33 & n4417 ) | ( x33 & ~n4418 ) | ( n4417 & ~n4418 ) ;
  assign n4420 = ( n4408 & n4414 ) | ( n4408 & n4419 ) | ( n4414 & n4419 ) ;
  assign n4421 = ( ~n4408 & n4414 ) | ( ~n4408 & n4419 ) | ( n4414 & n4419 ) ;
  assign n4422 = ( n4408 & ~n4420 ) | ( n4408 & n4421 ) | ( ~n4420 & n4421 ) ;
  assign n4423 = ( ~n4381 & n4402 ) | ( ~n4381 & n4422 ) | ( n4402 & n4422 ) ;
  assign n4424 = ( n4381 & n4402 ) | ( n4381 & n4422 ) | ( n4402 & n4422 ) ;
  assign n4425 = ( n4381 & n4423 ) | ( n4381 & ~n4424 ) | ( n4423 & ~n4424 ) ;
  assign n4426 = ( ~n4302 & n4366 ) | ( ~n4302 & n4425 ) | ( n4366 & n4425 ) ;
  assign n4427 = ( n4302 & n4366 ) | ( n4302 & n4425 ) | ( n4366 & n4425 ) ;
  assign n4428 = ( n4302 & n4426 ) | ( n4302 & ~n4427 ) | ( n4426 & ~n4427 ) ;
  assign n4429 = ( ~n4305 & n4360 ) | ( ~n4305 & n4428 ) | ( n4360 & n4428 ) ;
  assign n4430 = ( n4305 & n4360 ) | ( n4305 & n4428 ) | ( n4360 & n4428 ) ;
  assign n4431 = ( n4305 & n4429 ) | ( n4305 & ~n4430 ) | ( n4429 & ~n4430 ) ;
  assign n4432 = ( n4291 & n4328 ) | ( n4291 & n4431 ) | ( n4328 & n4431 ) ;
  assign n4433 = ( ~n4291 & n4328 ) | ( ~n4291 & n4431 ) | ( n4328 & n4431 ) ;
  assign n4434 = ( n4291 & ~n4432 ) | ( n4291 & n4433 ) | ( ~n4432 & n4433 ) ;
  assign n4435 = ( n4309 & n4312 ) | ( n4309 & n4434 ) | ( n4312 & n4434 ) ;
  assign n4436 = ( ~n4309 & n4312 ) | ( ~n4309 & n4434 ) | ( n4312 & n4434 ) ;
  assign n4437 = ( n4309 & ~n4435 ) | ( n4309 & n4436 ) | ( ~n4435 & n4436 ) ;
  assign n4438 = x27 & x39 ;
  assign n4439 = x28 & x38 ;
  assign n4440 = x29 & x37 ;
  assign n4441 = ( ~n4438 & n4439 ) | ( ~n4438 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4442 = ( n4438 & n4439 ) | ( n4438 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4443 = ( n4438 & n4441 ) | ( n4438 & ~n4442 ) | ( n4441 & ~n4442 ) ;
  assign n4444 = x3 & x63 ;
  assign n4445 = x5 & x61 ;
  assign n4446 = x4 & x62 ;
  assign n4447 = ( ~n4444 & n4445 ) | ( ~n4444 & n4446 ) | ( n4445 & n4446 ) ;
  assign n4448 = ( n4444 & n4445 ) | ( n4444 & n4446 ) | ( n4445 & n4446 ) ;
  assign n4449 = ( n4444 & n4447 ) | ( n4444 & ~n4448 ) | ( n4447 & ~n4448 ) ;
  assign n4450 = x11 & x55 ;
  assign n4451 = x19 & x47 ;
  assign n4452 = x12 & x54 ;
  assign n4453 = ( ~n4450 & n4451 ) | ( ~n4450 & n4452 ) | ( n4451 & n4452 ) ;
  assign n4454 = ( n4450 & n4451 ) | ( n4450 & n4452 ) | ( n4451 & n4452 ) ;
  assign n4455 = ( n4450 & n4453 ) | ( n4450 & ~n4454 ) | ( n4453 & ~n4454 ) ;
  assign n4456 = ( ~n4443 & n4449 ) | ( ~n4443 & n4455 ) | ( n4449 & n4455 ) ;
  assign n4457 = ( n4443 & n4449 ) | ( n4443 & n4455 ) | ( n4449 & n4455 ) ;
  assign n4458 = ( n4443 & n4456 ) | ( n4443 & ~n4457 ) | ( n4456 & ~n4457 ) ;
  assign n4459 = x10 & x56 ;
  assign n4460 = x25 & x41 ;
  assign n4461 = x26 & x40 ;
  assign n4462 = ( ~n4459 & n4460 ) | ( ~n4459 & n4461 ) | ( n4460 & n4461 ) ;
  assign n4463 = ( n4459 & n4460 ) | ( n4459 & n4461 ) | ( n4460 & n4461 ) ;
  assign n4464 = ( n4459 & n4462 ) | ( n4459 & ~n4463 ) | ( n4462 & ~n4463 ) ;
  assign n4465 = x20 & x46 ;
  assign n4466 = x22 & x44 ;
  assign n4467 = x21 & x45 ;
  assign n4468 = ( ~n4465 & n4466 ) | ( ~n4465 & n4467 ) | ( n4466 & n4467 ) ;
  assign n4469 = ( n4465 & n4466 ) | ( n4465 & n4467 ) | ( n4466 & n4467 ) ;
  assign n4470 = ( n4465 & n4468 ) | ( n4465 & ~n4469 ) | ( n4468 & ~n4469 ) ;
  assign n4471 = x23 & x43 ;
  assign n4472 = x9 & x57 ;
  assign n4473 = x24 & x42 ;
  assign n4474 = ( ~n4471 & n4472 ) | ( ~n4471 & n4473 ) | ( n4472 & n4473 ) ;
  assign n4475 = ( n4471 & n4472 ) | ( n4471 & n4473 ) | ( n4472 & n4473 ) ;
  assign n4476 = ( n4471 & n4474 ) | ( n4471 & ~n4475 ) | ( n4474 & ~n4475 ) ;
  assign n4477 = ( ~n4464 & n4470 ) | ( ~n4464 & n4476 ) | ( n4470 & n4476 ) ;
  assign n4478 = ( n4464 & n4470 ) | ( n4464 & n4476 ) | ( n4470 & n4476 ) ;
  assign n4479 = ( n4464 & n4477 ) | ( n4464 & ~n4478 ) | ( n4477 & ~n4478 ) ;
  assign n4480 = x32 & x34 ;
  assign n4481 = x17 & x49 ;
  assign n4482 = x16 & x50 ;
  assign n4483 = ( ~n4480 & n4481 ) | ( ~n4480 & n4482 ) | ( n4481 & n4482 ) ;
  assign n4484 = ( n4480 & n4481 ) | ( n4480 & n4482 ) | ( n4481 & n4482 ) ;
  assign n4485 = ( n4480 & n4483 ) | ( n4480 & ~n4484 ) | ( n4483 & ~n4484 ) ;
  assign n4486 = x14 & x52 ;
  assign n4487 = x30 & x36 ;
  assign n4488 = x31 & x35 ;
  assign n4489 = ( ~n4486 & n4487 ) | ( ~n4486 & n4488 ) | ( n4487 & n4488 ) ;
  assign n4490 = ( n4486 & n4487 ) | ( n4486 & n4488 ) | ( n4487 & n4488 ) ;
  assign n4491 = ( n4486 & n4489 ) | ( n4486 & ~n4490 ) | ( n4489 & ~n4490 ) ;
  assign n4492 = x18 & x48 ;
  assign n4493 = x15 & x51 ;
  assign n4494 = x13 & x53 ;
  assign n4495 = ( ~n4492 & n4493 ) | ( ~n4492 & n4494 ) | ( n4493 & n4494 ) ;
  assign n4496 = ( n4492 & n4493 ) | ( n4492 & n4494 ) | ( n4493 & n4494 ) ;
  assign n4497 = ( n4492 & n4495 ) | ( n4492 & ~n4496 ) | ( n4495 & ~n4496 ) ;
  assign n4498 = ( ~n4485 & n4491 ) | ( ~n4485 & n4497 ) | ( n4491 & n4497 ) ;
  assign n4499 = ( n4485 & n4491 ) | ( n4485 & n4497 ) | ( n4491 & n4497 ) ;
  assign n4500 = ( n4485 & n4498 ) | ( n4485 & ~n4499 ) | ( n4498 & ~n4499 ) ;
  assign n4501 = ( ~n4458 & n4479 ) | ( ~n4458 & n4500 ) | ( n4479 & n4500 ) ;
  assign n4502 = ( n4458 & n4479 ) | ( n4458 & n4500 ) | ( n4479 & n4500 ) ;
  assign n4503 = ( n4458 & n4501 ) | ( n4458 & ~n4502 ) | ( n4501 & ~n4502 ) ;
  assign n4504 = ( ~n4314 & n4318 ) | ( ~n4314 & n4330 ) | ( n4318 & n4330 ) ;
  assign n4505 = ( n4314 & n4318 ) | ( n4314 & n4330 ) | ( n4318 & n4330 ) ;
  assign n4506 = ( n4314 & n4504 ) | ( n4314 & ~n4505 ) | ( n4504 & ~n4505 ) ;
  assign n4507 = ( n4321 & n4332 ) | ( n4321 & n4506 ) | ( n4332 & n4506 ) ;
  assign n4508 = ( n4321 & ~n4332 ) | ( n4321 & n4506 ) | ( ~n4332 & n4506 ) ;
  assign n4509 = ( n4332 & ~n4507 ) | ( n4332 & n4508 ) | ( ~n4507 & n4508 ) ;
  assign n4510 = ( ~n4324 & n4503 ) | ( ~n4324 & n4509 ) | ( n4503 & n4509 ) ;
  assign n4511 = ( n4324 & n4503 ) | ( n4324 & n4509 ) | ( n4503 & n4509 ) ;
  assign n4512 = ( n4324 & n4510 ) | ( n4324 & ~n4511 ) | ( n4510 & ~n4511 ) ;
  assign n4513 = ( ~n4327 & n4427 ) | ( ~n4327 & n4512 ) | ( n4427 & n4512 ) ;
  assign n4514 = ( n4327 & n4427 ) | ( n4327 & n4512 ) | ( n4427 & n4512 ) ;
  assign n4515 = ( n4327 & n4513 ) | ( n4327 & ~n4514 ) | ( n4513 & ~n4514 ) ;
  assign n4516 = x6 & x60 ;
  assign n4517 = x7 & x59 ;
  assign n4518 = x8 & x58 ;
  assign n4519 = ( ~n4516 & n4517 ) | ( ~n4516 & n4518 ) | ( n4517 & n4518 ) ;
  assign n4520 = ( n4516 & n4517 ) | ( n4516 & n4518 ) | ( n4517 & n4518 ) ;
  assign n4521 = ( n4516 & n4519 ) | ( n4516 & ~n4520 ) | ( n4519 & ~n4520 ) ;
  assign n4522 = ( ~n4337 & n4386 ) | ( ~n4337 & n4521 ) | ( n4386 & n4521 ) ;
  assign n4523 = ( n4337 & n4386 ) | ( n4337 & n4521 ) | ( n4386 & n4521 ) ;
  assign n4524 = ( n4337 & n4522 ) | ( n4337 & ~n4523 ) | ( n4522 & ~n4523 ) ;
  assign n4525 = ( ~n4352 & n4362 ) | ( ~n4352 & n4524 ) | ( n4362 & n4524 ) ;
  assign n4526 = ( n4352 & n4362 ) | ( n4352 & n4524 ) | ( n4362 & n4524 ) ;
  assign n4527 = ( n4352 & n4525 ) | ( n4352 & ~n4526 ) | ( n4525 & ~n4526 ) ;
  assign n4528 = ( n4371 & n4377 ) | ( n4371 & n4413 ) | ( n4377 & n4413 ) ;
  assign n4529 = ( n4371 & ~n4377 ) | ( n4371 & n4413 ) | ( ~n4377 & n4413 ) ;
  assign n4530 = ( n4377 & ~n4528 ) | ( n4377 & n4529 ) | ( ~n4528 & n4529 ) ;
  assign n4531 = ( n4350 & n4407 ) | ( n4350 & ~n4418 ) | ( n4407 & ~n4418 ) ;
  assign n4532 = ( n4350 & n4407 ) | ( n4350 & n4418 ) | ( n4407 & n4418 ) ;
  assign n4533 = ( n4418 & n4531 ) | ( n4418 & ~n4532 ) | ( n4531 & ~n4532 ) ;
  assign n4534 = ( ~n4420 & n4530 ) | ( ~n4420 & n4533 ) | ( n4530 & n4533 ) ;
  assign n4535 = ( n4420 & n4530 ) | ( n4420 & n4533 ) | ( n4530 & n4533 ) ;
  assign n4536 = ( n4420 & n4534 ) | ( n4420 & ~n4535 ) | ( n4534 & ~n4535 ) ;
  assign n4537 = ( n4364 & n4527 ) | ( n4364 & n4536 ) | ( n4527 & n4536 ) ;
  assign n4538 = ( ~n4364 & n4527 ) | ( ~n4364 & n4536 ) | ( n4527 & n4536 ) ;
  assign n4539 = ( n4364 & ~n4537 ) | ( n4364 & n4538 ) | ( ~n4537 & n4538 ) ;
  assign n4540 = ( n4344 & ~n4392 ) | ( n4344 & n4398 ) | ( ~n4392 & n4398 ) ;
  assign n4541 = ( n4344 & n4392 ) | ( n4344 & n4398 ) | ( n4392 & n4398 ) ;
  assign n4542 = ( n4392 & n4540 ) | ( n4392 & ~n4541 ) | ( n4540 & ~n4541 ) ;
  assign n4543 = ( ~n4379 & n4401 ) | ( ~n4379 & n4542 ) | ( n4401 & n4542 ) ;
  assign n4544 = ( n4379 & n4401 ) | ( n4379 & n4542 ) | ( n4401 & n4542 ) ;
  assign n4545 = ( n4379 & n4543 ) | ( n4379 & ~n4544 ) | ( n4543 & ~n4544 ) ;
  assign n4546 = ( ~n4355 & n4424 ) | ( ~n4355 & n4545 ) | ( n4424 & n4545 ) ;
  assign n4547 = ( n4355 & n4424 ) | ( n4355 & n4545 ) | ( n4424 & n4545 ) ;
  assign n4548 = ( n4355 & n4546 ) | ( n4355 & ~n4547 ) | ( n4546 & ~n4547 ) ;
  assign n4549 = ( n4359 & n4539 ) | ( n4359 & n4548 ) | ( n4539 & n4548 ) ;
  assign n4550 = ( ~n4359 & n4539 ) | ( ~n4359 & n4548 ) | ( n4539 & n4548 ) ;
  assign n4551 = ( n4359 & ~n4549 ) | ( n4359 & n4550 ) | ( ~n4549 & n4550 ) ;
  assign n4552 = ( ~n4430 & n4515 ) | ( ~n4430 & n4551 ) | ( n4515 & n4551 ) ;
  assign n4553 = ( n4430 & n4515 ) | ( n4430 & n4551 ) | ( n4515 & n4551 ) ;
  assign n4554 = ( n4430 & n4552 ) | ( n4430 & ~n4553 ) | ( n4552 & ~n4553 ) ;
  assign n4555 = ( ~n4432 & n4435 ) | ( ~n4432 & n4554 ) | ( n4435 & n4554 ) ;
  assign n4556 = ( n4432 & n4435 ) | ( n4432 & n4554 ) | ( n4435 & n4554 ) ;
  assign n4557 = ( n4432 & n4555 ) | ( n4432 & ~n4556 ) | ( n4555 & ~n4556 ) ;
  assign n4558 = ( n4457 & n4478 ) | ( n4457 & ~n4523 ) | ( n4478 & ~n4523 ) ;
  assign n4559 = ( n4457 & n4478 ) | ( n4457 & n4523 ) | ( n4478 & n4523 ) ;
  assign n4560 = ( n4523 & n4558 ) | ( n4523 & ~n4559 ) | ( n4558 & ~n4559 ) ;
  assign n4561 = ( n4463 & n4469 ) | ( n4463 & n4475 ) | ( n4469 & n4475 ) ;
  assign n4562 = ( ~n4463 & n4469 ) | ( ~n4463 & n4475 ) | ( n4469 & n4475 ) ;
  assign n4563 = ( n4463 & ~n4561 ) | ( n4463 & n4562 ) | ( ~n4561 & n4562 ) ;
  assign n4564 = ( ~n4442 & n4448 ) | ( ~n4442 & n4520 ) | ( n4448 & n4520 ) ;
  assign n4565 = ( n4442 & n4448 ) | ( n4442 & n4520 ) | ( n4448 & n4520 ) ;
  assign n4566 = ( n4442 & n4564 ) | ( n4442 & ~n4565 ) | ( n4564 & ~n4565 ) ;
  assign n4567 = x6 & x61 ;
  assign n4568 = ( n4484 & n4490 ) | ( n4484 & n4567 ) | ( n4490 & n4567 ) ;
  assign n4569 = ( ~n4484 & n4490 ) | ( ~n4484 & n4567 ) | ( n4490 & n4567 ) ;
  assign n4570 = ( n4484 & ~n4568 ) | ( n4484 & n4569 ) | ( ~n4568 & n4569 ) ;
  assign n4571 = ( ~n4563 & n4566 ) | ( ~n4563 & n4570 ) | ( n4566 & n4570 ) ;
  assign n4572 = ( n4563 & n4566 ) | ( n4563 & n4570 ) | ( n4566 & n4570 ) ;
  assign n4573 = ( n4563 & n4571 ) | ( n4563 & ~n4572 ) | ( n4571 & ~n4572 ) ;
  assign n4574 = ( ~n4507 & n4560 ) | ( ~n4507 & n4573 ) | ( n4560 & n4573 ) ;
  assign n4575 = ( n4507 & n4560 ) | ( n4507 & n4573 ) | ( n4560 & n4573 ) ;
  assign n4576 = ( n4507 & n4574 ) | ( n4507 & ~n4575 ) | ( n4574 & ~n4575 ) ;
  assign n4577 = x10 & x57 ;
  assign n4578 = x11 & x56 ;
  assign n4579 = x20 & x47 ;
  assign n4580 = ( ~n4577 & n4578 ) | ( ~n4577 & n4579 ) | ( n4578 & n4579 ) ;
  assign n4581 = ( n4577 & n4578 ) | ( n4577 & n4579 ) | ( n4578 & n4579 ) ;
  assign n4582 = ( n4577 & n4580 ) | ( n4577 & ~n4581 ) | ( n4580 & ~n4581 ) ;
  assign n4583 = ( ~n4454 & n4496 ) | ( ~n4454 & n4582 ) | ( n4496 & n4582 ) ;
  assign n4584 = ( n4454 & n4496 ) | ( n4454 & n4582 ) | ( n4496 & n4582 ) ;
  assign n4585 = ( n4454 & n4583 ) | ( n4454 & ~n4584 ) | ( n4583 & ~n4584 ) ;
  assign n4586 = ( ~n4499 & n4505 ) | ( ~n4499 & n4585 ) | ( n4505 & n4585 ) ;
  assign n4587 = ( n4499 & n4505 ) | ( n4499 & n4585 ) | ( n4505 & n4585 ) ;
  assign n4588 = ( n4499 & n4586 ) | ( n4499 & ~n4587 ) | ( n4586 & ~n4587 ) ;
  assign n4589 = ( ~n4502 & n4526 ) | ( ~n4502 & n4588 ) | ( n4526 & n4588 ) ;
  assign n4590 = ( n4502 & n4526 ) | ( n4502 & n4588 ) | ( n4526 & n4588 ) ;
  assign n4591 = ( n4502 & n4589 ) | ( n4502 & ~n4590 ) | ( n4589 & ~n4590 ) ;
  assign n4592 = ( ~n4537 & n4576 ) | ( ~n4537 & n4591 ) | ( n4576 & n4591 ) ;
  assign n4593 = ( n4537 & n4576 ) | ( n4537 & n4591 ) | ( n4576 & n4591 ) ;
  assign n4594 = ( n4537 & n4592 ) | ( n4537 & ~n4593 ) | ( n4592 & ~n4593 ) ;
  assign n4595 = x4 & x63 ;
  assign n4596 = x27 & x40 ;
  assign n4597 = x28 & x39 ;
  assign n4598 = ( ~n4595 & n4596 ) | ( ~n4595 & n4597 ) | ( n4596 & n4597 ) ;
  assign n4599 = ( n4595 & n4596 ) | ( n4595 & n4597 ) | ( n4596 & n4597 ) ;
  assign n4600 = ( n4595 & n4598 ) | ( n4595 & ~n4599 ) | ( n4598 & ~n4599 ) ;
  assign n4601 = x17 & x50 ;
  assign n4602 = x19 & x48 ;
  assign n4603 = x14 & x53 ;
  assign n4604 = ( ~n4601 & n4602 ) | ( ~n4601 & n4603 ) | ( n4602 & n4603 ) ;
  assign n4605 = ( n4601 & n4602 ) | ( n4601 & n4603 ) | ( n4602 & n4603 ) ;
  assign n4606 = ( n4601 & n4604 ) | ( n4601 & ~n4605 ) | ( n4604 & ~n4605 ) ;
  assign n4607 = x26 & x41 ;
  assign n4608 = x25 & x42 ;
  assign n4609 = x21 & x46 ;
  assign n4610 = ( ~n4607 & n4608 ) | ( ~n4607 & n4609 ) | ( n4608 & n4609 ) ;
  assign n4611 = ( n4607 & n4608 ) | ( n4607 & n4609 ) | ( n4608 & n4609 ) ;
  assign n4612 = ( n4607 & n4610 ) | ( n4607 & ~n4611 ) | ( n4610 & ~n4611 ) ;
  assign n4613 = ( ~n4600 & n4606 ) | ( ~n4600 & n4612 ) | ( n4606 & n4612 ) ;
  assign n4614 = ( n4600 & n4606 ) | ( n4600 & n4612 ) | ( n4606 & n4612 ) ;
  assign n4615 = ( n4600 & n4613 ) | ( n4600 & ~n4614 ) | ( n4613 & ~n4614 ) ;
  assign n4616 = x29 & x38 ;
  assign n4617 = x12 & x55 ;
  assign n4618 = x13 & x54 ;
  assign n4619 = ( ~n4616 & n4617 ) | ( ~n4616 & n4618 ) | ( n4617 & n4618 ) ;
  assign n4620 = ( n4616 & n4617 ) | ( n4616 & n4618 ) | ( n4617 & n4618 ) ;
  assign n4621 = ( n4616 & n4619 ) | ( n4616 & ~n4620 ) | ( n4619 & ~n4620 ) ;
  assign n4622 = x31 & x36 ;
  assign n4623 = x33 & x34 ;
  assign n4624 = x32 & x35 ;
  assign n4625 = ( ~n4622 & n4623 ) | ( ~n4622 & n4624 ) | ( n4623 & n4624 ) ;
  assign n4626 = ( n4622 & n4623 ) | ( n4622 & n4624 ) | ( n4623 & n4624 ) ;
  assign n4627 = ( n4622 & n4625 ) | ( n4622 & ~n4626 ) | ( n4625 & ~n4626 ) ;
  assign n4628 = x5 & x62 ;
  assign n4629 = x18 & x49 ;
  assign n4630 = ( ~x34 & n4628 ) | ( ~x34 & n4629 ) | ( n4628 & n4629 ) ;
  assign n4631 = ( x34 & n4628 ) | ( x34 & n4629 ) | ( n4628 & n4629 ) ;
  assign n4632 = ( x34 & n4630 ) | ( x34 & ~n4631 ) | ( n4630 & ~n4631 ) ;
  assign n4633 = ( ~n4621 & n4627 ) | ( ~n4621 & n4632 ) | ( n4627 & n4632 ) ;
  assign n4634 = ( n4621 & n4627 ) | ( n4621 & n4632 ) | ( n4627 & n4632 ) ;
  assign n4635 = ( n4621 & n4633 ) | ( n4621 & ~n4634 ) | ( n4633 & ~n4634 ) ;
  assign n4636 = x22 & x45 ;
  assign n4637 = x24 & x43 ;
  assign n4638 = ( ~n2111 & n4636 ) | ( ~n2111 & n4637 ) | ( n4636 & n4637 ) ;
  assign n4639 = ( n2111 & n4636 ) | ( n2111 & n4637 ) | ( n4636 & n4637 ) ;
  assign n4640 = ( n2111 & n4638 ) | ( n2111 & ~n4639 ) | ( n4638 & ~n4639 ) ;
  assign n4641 = x7 & x60 ;
  assign n4642 = x8 & x59 ;
  assign n4643 = x9 & x58 ;
  assign n4644 = ( ~n4641 & n4642 ) | ( ~n4641 & n4643 ) | ( n4642 & n4643 ) ;
  assign n4645 = ( n4641 & n4642 ) | ( n4641 & n4643 ) | ( n4642 & n4643 ) ;
  assign n4646 = ( n4641 & n4644 ) | ( n4641 & ~n4645 ) | ( n4644 & ~n4645 ) ;
  assign n4647 = x16 & x51 ;
  assign n4648 = x15 & x52 ;
  assign n4649 = x30 & x37 ;
  assign n4650 = ( ~n4647 & n4648 ) | ( ~n4647 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4651 = ( n4647 & n4648 ) | ( n4647 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4652 = ( n4647 & n4650 ) | ( n4647 & ~n4651 ) | ( n4650 & ~n4651 ) ;
  assign n4653 = ( ~n4640 & n4646 ) | ( ~n4640 & n4652 ) | ( n4646 & n4652 ) ;
  assign n4654 = ( n4640 & n4646 ) | ( n4640 & n4652 ) | ( n4646 & n4652 ) ;
  assign n4655 = ( n4640 & n4653 ) | ( n4640 & ~n4654 ) | ( n4653 & ~n4654 ) ;
  assign n4656 = ( ~n4615 & n4635 ) | ( ~n4615 & n4655 ) | ( n4635 & n4655 ) ;
  assign n4657 = ( n4615 & n4635 ) | ( n4615 & n4655 ) | ( n4635 & n4655 ) ;
  assign n4658 = ( n4615 & n4656 ) | ( n4615 & ~n4657 ) | ( n4656 & ~n4657 ) ;
  assign n4659 = ( ~n4528 & n4532 ) | ( ~n4528 & n4541 ) | ( n4532 & n4541 ) ;
  assign n4660 = ( n4528 & n4532 ) | ( n4528 & n4541 ) | ( n4532 & n4541 ) ;
  assign n4661 = ( n4528 & n4659 ) | ( n4528 & ~n4660 ) | ( n4659 & ~n4660 ) ;
  assign n4662 = ( n4535 & n4544 ) | ( n4535 & n4661 ) | ( n4544 & n4661 ) ;
  assign n4663 = ( ~n4535 & n4544 ) | ( ~n4535 & n4661 ) | ( n4544 & n4661 ) ;
  assign n4664 = ( n4535 & ~n4662 ) | ( n4535 & n4663 ) | ( ~n4662 & n4663 ) ;
  assign n4665 = ( ~n4547 & n4658 ) | ( ~n4547 & n4664 ) | ( n4658 & n4664 ) ;
  assign n4666 = ( n4547 & n4658 ) | ( n4547 & n4664 ) | ( n4658 & n4664 ) ;
  assign n4667 = ( n4547 & n4665 ) | ( n4547 & ~n4666 ) | ( n4665 & ~n4666 ) ;
  assign n4668 = ( n4511 & n4549 ) | ( n4511 & n4667 ) | ( n4549 & n4667 ) ;
  assign n4669 = ( ~n4511 & n4549 ) | ( ~n4511 & n4667 ) | ( n4549 & n4667 ) ;
  assign n4670 = ( n4511 & ~n4668 ) | ( n4511 & n4669 ) | ( ~n4668 & n4669 ) ;
  assign n4671 = ( ~n4514 & n4594 ) | ( ~n4514 & n4670 ) | ( n4594 & n4670 ) ;
  assign n4672 = ( n4514 & n4594 ) | ( n4514 & n4670 ) | ( n4594 & n4670 ) ;
  assign n4673 = ( n4514 & n4671 ) | ( n4514 & ~n4672 ) | ( n4671 & ~n4672 ) ;
  assign n4674 = ( n4553 & n4556 ) | ( n4553 & n4673 ) | ( n4556 & n4673 ) ;
  assign n4675 = ( n4553 & ~n4556 ) | ( n4553 & n4673 ) | ( ~n4556 & n4673 ) ;
  assign n4676 = ( n4556 & ~n4674 ) | ( n4556 & n4675 ) | ( ~n4674 & n4675 ) ;
  assign n4677 = ( n4559 & n4572 ) | ( n4559 & ~n4587 ) | ( n4572 & ~n4587 ) ;
  assign n4678 = ( n4559 & n4572 ) | ( n4559 & n4587 ) | ( n4572 & n4587 ) ;
  assign n4679 = ( n4587 & n4677 ) | ( n4587 & ~n4678 ) | ( n4677 & ~n4678 ) ;
  assign n4680 = x30 & x38 ;
  assign n4681 = x31 & x37 ;
  assign n4682 = x32 & x36 ;
  assign n4683 = ( ~n4680 & n4681 ) | ( ~n4680 & n4682 ) | ( n4681 & n4682 ) ;
  assign n4684 = ( n4680 & n4681 ) | ( n4680 & n4682 ) | ( n4681 & n4682 ) ;
  assign n4685 = ( n4680 & n4683 ) | ( n4680 & ~n4684 ) | ( n4683 & ~n4684 ) ;
  assign n4686 = x33 & x35 ;
  assign n4687 = x18 & x50 ;
  assign n4688 = x19 & x49 ;
  assign n4689 = ( ~n4686 & n4687 ) | ( ~n4686 & n4688 ) | ( n4687 & n4688 ) ;
  assign n4690 = ( n4686 & n4687 ) | ( n4686 & n4688 ) | ( n4687 & n4688 ) ;
  assign n4691 = ( n4686 & n4689 ) | ( n4686 & ~n4690 ) | ( n4689 & ~n4690 ) ;
  assign n4692 = x17 & x51 ;
  assign n4693 = x13 & x55 ;
  assign n4694 = x12 & x56 ;
  assign n4695 = ( ~n4692 & n4693 ) | ( ~n4692 & n4694 ) | ( n4693 & n4694 ) ;
  assign n4696 = ( n4692 & n4693 ) | ( n4692 & n4694 ) | ( n4693 & n4694 ) ;
  assign n4697 = ( n4692 & n4695 ) | ( n4692 & ~n4696 ) | ( n4695 & ~n4696 ) ;
  assign n4698 = ( n4685 & n4691 ) | ( n4685 & n4697 ) | ( n4691 & n4697 ) ;
  assign n4699 = ( ~n4685 & n4691 ) | ( ~n4685 & n4697 ) | ( n4691 & n4697 ) ;
  assign n4700 = ( n4685 & ~n4698 ) | ( n4685 & n4699 ) | ( ~n4698 & n4699 ) ;
  assign n4701 = x27 & x41 ;
  assign n4702 = x28 & x40 ;
  assign n4703 = x29 & x39 ;
  assign n4704 = ( ~n4701 & n4702 ) | ( ~n4701 & n4703 ) | ( n4702 & n4703 ) ;
  assign n4705 = ( n4701 & n4702 ) | ( n4701 & n4703 ) | ( n4702 & n4703 ) ;
  assign n4706 = ( n4701 & n4704 ) | ( n4701 & ~n4705 ) | ( n4704 & ~n4705 ) ;
  assign n4707 = x21 & x47 ;
  assign n4708 = x5 & x63 ;
  assign n4709 = x6 & x62 ;
  assign n4710 = ( ~n4707 & n4708 ) | ( ~n4707 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4711 = ( n4707 & n4708 ) | ( n4707 & n4709 ) | ( n4708 & n4709 ) ;
  assign n4712 = ( n4707 & n4710 ) | ( n4707 & ~n4711 ) | ( n4710 & ~n4711 ) ;
  assign n4713 = x9 & x59 ;
  assign n4714 = x10 & x58 ;
  assign n4715 = x11 & x57 ;
  assign n4716 = ( ~n4713 & n4714 ) | ( ~n4713 & n4715 ) | ( n4714 & n4715 ) ;
  assign n4717 = ( n4713 & n4714 ) | ( n4713 & n4715 ) | ( n4714 & n4715 ) ;
  assign n4718 = ( n4713 & n4716 ) | ( n4713 & ~n4717 ) | ( n4716 & ~n4717 ) ;
  assign n4719 = ( ~n4706 & n4712 ) | ( ~n4706 & n4718 ) | ( n4712 & n4718 ) ;
  assign n4720 = ( n4706 & n4712 ) | ( n4706 & n4718 ) | ( n4712 & n4718 ) ;
  assign n4721 = ( n4706 & n4719 ) | ( n4706 & ~n4720 ) | ( n4719 & ~n4720 ) ;
  assign n4722 = x20 & x48 ;
  assign n4723 = x23 & x45 ;
  assign n4724 = x22 & x46 ;
  assign n4725 = ( ~n4722 & n4723 ) | ( ~n4722 & n4724 ) | ( n4723 & n4724 ) ;
  assign n4726 = ( n4722 & n4723 ) | ( n4722 & n4724 ) | ( n4723 & n4724 ) ;
  assign n4727 = ( n4722 & n4725 ) | ( n4722 & ~n4726 ) | ( n4725 & ~n4726 ) ;
  assign n4728 = x24 & x44 ;
  assign n4729 = x25 & x43 ;
  assign n4730 = x26 & x42 ;
  assign n4731 = ( ~n4728 & n4729 ) | ( ~n4728 & n4730 ) | ( n4729 & n4730 ) ;
  assign n4732 = ( n4728 & n4729 ) | ( n4728 & n4730 ) | ( n4729 & n4730 ) ;
  assign n4733 = ( n4728 & n4731 ) | ( n4728 & ~n4732 ) | ( n4731 & ~n4732 ) ;
  assign n4734 = x14 & x54 ;
  assign n4735 = x16 & x52 ;
  assign n4736 = x15 & x53 ;
  assign n4737 = ( ~n4734 & n4735 ) | ( ~n4734 & n4736 ) | ( n4735 & n4736 ) ;
  assign n4738 = ( n4734 & n4735 ) | ( n4734 & n4736 ) | ( n4735 & n4736 ) ;
  assign n4739 = ( n4734 & n4737 ) | ( n4734 & ~n4738 ) | ( n4737 & ~n4738 ) ;
  assign n4740 = ( ~n4727 & n4733 ) | ( ~n4727 & n4739 ) | ( n4733 & n4739 ) ;
  assign n4741 = ( n4727 & n4733 ) | ( n4727 & n4739 ) | ( n4733 & n4739 ) ;
  assign n4742 = ( n4727 & n4740 ) | ( n4727 & ~n4741 ) | ( n4740 & ~n4741 ) ;
  assign n4743 = ( ~n4700 & n4721 ) | ( ~n4700 & n4742 ) | ( n4721 & n4742 ) ;
  assign n4744 = ( n4700 & n4721 ) | ( n4700 & n4742 ) | ( n4721 & n4742 ) ;
  assign n4745 = ( n4700 & n4743 ) | ( n4700 & ~n4744 ) | ( n4743 & ~n4744 ) ;
  assign n4746 = ( n4590 & n4679 ) | ( n4590 & n4745 ) | ( n4679 & n4745 ) ;
  assign n4747 = ( ~n4590 & n4679 ) | ( ~n4590 & n4745 ) | ( n4679 & n4745 ) ;
  assign n4748 = ( n4590 & ~n4746 ) | ( n4590 & n4747 ) | ( ~n4746 & n4747 ) ;
  assign n4749 = ( ~n4593 & n4666 ) | ( ~n4593 & n4748 ) | ( n4666 & n4748 ) ;
  assign n4750 = ( n4593 & n4666 ) | ( n4593 & n4748 ) | ( n4666 & n4748 ) ;
  assign n4751 = ( n4593 & n4749 ) | ( n4593 & ~n4750 ) | ( n4749 & ~n4750 ) ;
  assign n4752 = ( n4561 & n4584 ) | ( n4561 & n4654 ) | ( n4584 & n4654 ) ;
  assign n4753 = ( ~n4561 & n4584 ) | ( ~n4561 & n4654 ) | ( n4584 & n4654 ) ;
  assign n4754 = ( n4561 & ~n4752 ) | ( n4561 & n4753 ) | ( ~n4752 & n4753 ) ;
  assign n4755 = x8 & x60 ;
  assign n4756 = x7 & x61 ;
  assign n4757 = ( n4631 & n4755 ) | ( n4631 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4758 = ( ~n4631 & n4755 ) | ( ~n4631 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4759 = ( n4631 & ~n4757 ) | ( n4631 & n4758 ) | ( ~n4757 & n4758 ) ;
  assign n4760 = ( n4565 & n4568 ) | ( n4565 & n4759 ) | ( n4568 & n4759 ) ;
  assign n4761 = ( ~n4565 & n4568 ) | ( ~n4565 & n4759 ) | ( n4568 & n4759 ) ;
  assign n4762 = ( n4565 & ~n4760 ) | ( n4565 & n4761 ) | ( ~n4760 & n4761 ) ;
  assign n4763 = ( n4657 & n4754 ) | ( n4657 & n4762 ) | ( n4754 & n4762 ) ;
  assign n4764 = ( n4657 & ~n4754 ) | ( n4657 & n4762 ) | ( ~n4754 & n4762 ) ;
  assign n4765 = ( n4754 & ~n4763 ) | ( n4754 & n4764 ) | ( ~n4763 & n4764 ) ;
  assign n4766 = ( n4605 & ~n4611 ) | ( n4605 & n4620 ) | ( ~n4611 & n4620 ) ;
  assign n4767 = ( n4605 & n4611 ) | ( n4605 & n4620 ) | ( n4611 & n4620 ) ;
  assign n4768 = ( n4611 & n4766 ) | ( n4611 & ~n4767 ) | ( n4766 & ~n4767 ) ;
  assign n4769 = ( ~n4614 & n4634 ) | ( ~n4614 & n4768 ) | ( n4634 & n4768 ) ;
  assign n4770 = ( n4614 & n4634 ) | ( n4614 & n4768 ) | ( n4634 & n4768 ) ;
  assign n4771 = ( n4614 & n4769 ) | ( n4614 & ~n4770 ) | ( n4769 & ~n4770 ) ;
  assign n4772 = ( n4581 & ~n4639 ) | ( n4581 & n4645 ) | ( ~n4639 & n4645 ) ;
  assign n4773 = ( n4581 & n4639 ) | ( n4581 & n4645 ) | ( n4639 & n4645 ) ;
  assign n4774 = ( n4639 & n4772 ) | ( n4639 & ~n4773 ) | ( n4772 & ~n4773 ) ;
  assign n4775 = ( ~n4599 & n4626 ) | ( ~n4599 & n4651 ) | ( n4626 & n4651 ) ;
  assign n4776 = ( n4599 & n4626 ) | ( n4599 & n4651 ) | ( n4626 & n4651 ) ;
  assign n4777 = ( n4599 & n4775 ) | ( n4599 & ~n4776 ) | ( n4775 & ~n4776 ) ;
  assign n4778 = ( ~n4660 & n4774 ) | ( ~n4660 & n4777 ) | ( n4774 & n4777 ) ;
  assign n4779 = ( n4660 & n4774 ) | ( n4660 & n4777 ) | ( n4774 & n4777 ) ;
  assign n4780 = ( n4660 & n4778 ) | ( n4660 & ~n4779 ) | ( n4778 & ~n4779 ) ;
  assign n4781 = ( ~n4662 & n4771 ) | ( ~n4662 & n4780 ) | ( n4771 & n4780 ) ;
  assign n4782 = ( n4662 & n4771 ) | ( n4662 & n4780 ) | ( n4771 & n4780 ) ;
  assign n4783 = ( n4662 & n4781 ) | ( n4662 & ~n4782 ) | ( n4781 & ~n4782 ) ;
  assign n4784 = ( ~n4575 & n4765 ) | ( ~n4575 & n4783 ) | ( n4765 & n4783 ) ;
  assign n4785 = ( n4575 & n4765 ) | ( n4575 & n4783 ) | ( n4765 & n4783 ) ;
  assign n4786 = ( n4575 & n4784 ) | ( n4575 & ~n4785 ) | ( n4784 & ~n4785 ) ;
  assign n4787 = ( ~n4668 & n4751 ) | ( ~n4668 & n4786 ) | ( n4751 & n4786 ) ;
  assign n4788 = ( n4668 & n4751 ) | ( n4668 & n4786 ) | ( n4751 & n4786 ) ;
  assign n4789 = ( n4668 & n4787 ) | ( n4668 & ~n4788 ) | ( n4787 & ~n4788 ) ;
  assign n4790 = ( n4672 & n4674 ) | ( n4672 & n4789 ) | ( n4674 & n4789 ) ;
  assign n4791 = ( ~n4672 & n4674 ) | ( ~n4672 & n4789 ) | ( n4674 & n4789 ) ;
  assign n4792 = ( n4672 & ~n4790 ) | ( n4672 & n4791 ) | ( ~n4790 & n4791 ) ;
  assign n4793 = ( n4696 & ~n4705 ) | ( n4696 & n4732 ) | ( ~n4705 & n4732 ) ;
  assign n4794 = ( n4696 & n4705 ) | ( n4696 & n4732 ) | ( n4705 & n4732 ) ;
  assign n4795 = ( n4705 & n4793 ) | ( n4705 & ~n4794 ) | ( n4793 & ~n4794 ) ;
  assign n4796 = ( n4767 & n4776 ) | ( n4767 & n4795 ) | ( n4776 & n4795 ) ;
  assign n4797 = ( ~n4767 & n4776 ) | ( ~n4767 & n4795 ) | ( n4776 & n4795 ) ;
  assign n4798 = ( n4767 & ~n4796 ) | ( n4767 & n4797 ) | ( ~n4796 & n4797 ) ;
  assign n4799 = ( n4744 & n4779 ) | ( n4744 & n4798 ) | ( n4779 & n4798 ) ;
  assign n4800 = ( ~n4744 & n4779 ) | ( ~n4744 & n4798 ) | ( n4779 & n4798 ) ;
  assign n4801 = ( n4744 & ~n4799 ) | ( n4744 & n4800 ) | ( ~n4799 & n4800 ) ;
  assign n4802 = ( ~n4698 & n4741 ) | ( ~n4698 & n4760 ) | ( n4741 & n4760 ) ;
  assign n4803 = ( n4698 & n4741 ) | ( n4698 & n4760 ) | ( n4741 & n4760 ) ;
  assign n4804 = ( n4698 & n4802 ) | ( n4698 & ~n4803 ) | ( n4802 & ~n4803 ) ;
  assign n4805 = ( ~n4684 & n4690 ) | ( ~n4684 & n4738 ) | ( n4690 & n4738 ) ;
  assign n4806 = ( n4684 & n4690 ) | ( n4684 & n4738 ) | ( n4690 & n4738 ) ;
  assign n4807 = ( n4684 & n4805 ) | ( n4684 & ~n4806 ) | ( n4805 & ~n4806 ) ;
  assign n4808 = ( n4711 & ~n4717 ) | ( n4711 & n4726 ) | ( ~n4717 & n4726 ) ;
  assign n4809 = ( n4711 & n4717 ) | ( n4711 & n4726 ) | ( n4717 & n4726 ) ;
  assign n4810 = ( n4717 & n4808 ) | ( n4717 & ~n4809 ) | ( n4808 & ~n4809 ) ;
  assign n4811 = ( n4720 & n4807 ) | ( n4720 & n4810 ) | ( n4807 & n4810 ) ;
  assign n4812 = ( ~n4720 & n4807 ) | ( ~n4720 & n4810 ) | ( n4807 & n4810 ) ;
  assign n4813 = ( n4720 & ~n4811 ) | ( n4720 & n4812 ) | ( ~n4811 & n4812 ) ;
  assign n4814 = ( ~n4678 & n4804 ) | ( ~n4678 & n4813 ) | ( n4804 & n4813 ) ;
  assign n4815 = ( n4678 & n4804 ) | ( n4678 & n4813 ) | ( n4804 & n4813 ) ;
  assign n4816 = ( n4678 & n4814 ) | ( n4678 & ~n4815 ) | ( n4814 & ~n4815 ) ;
  assign n4817 = ( ~n4782 & n4801 ) | ( ~n4782 & n4816 ) | ( n4801 & n4816 ) ;
  assign n4818 = ( n4782 & n4801 ) | ( n4782 & n4816 ) | ( n4801 & n4816 ) ;
  assign n4819 = ( n4782 & n4817 ) | ( n4782 & ~n4818 ) | ( n4817 & ~n4818 ) ;
  assign n4820 = x6 & x63 ;
  assign n4821 = x26 & x43 ;
  assign n4822 = x27 & x42 ;
  assign n4823 = ( ~n4820 & n4821 ) | ( ~n4820 & n4822 ) | ( n4821 & n4822 ) ;
  assign n4824 = ( n4820 & n4821 ) | ( n4820 & n4822 ) | ( n4821 & n4822 ) ;
  assign n4825 = ( n4820 & n4823 ) | ( n4820 & ~n4824 ) | ( n4823 & ~n4824 ) ;
  assign n4826 = x23 & x46 ;
  assign n4827 = x24 & x45 ;
  assign n4828 = x25 & x44 ;
  assign n4829 = ( ~n4826 & n4827 ) | ( ~n4826 & n4828 ) | ( n4827 & n4828 ) ;
  assign n4830 = ( n4826 & n4827 ) | ( n4826 & n4828 ) | ( n4827 & n4828 ) ;
  assign n4831 = ( n4826 & n4829 ) | ( n4826 & ~n4830 ) | ( n4829 & ~n4830 ) ;
  assign n4832 = x8 & x61 ;
  assign n4833 = x9 & x60 ;
  assign n4834 = x10 & x59 ;
  assign n4835 = ( ~n4832 & n4833 ) | ( ~n4832 & n4834 ) | ( n4833 & n4834 ) ;
  assign n4836 = ( n4832 & n4833 ) | ( n4832 & n4834 ) | ( n4833 & n4834 ) ;
  assign n4837 = ( n4832 & n4835 ) | ( n4832 & ~n4836 ) | ( n4835 & ~n4836 ) ;
  assign n4838 = ( ~n4825 & n4831 ) | ( ~n4825 & n4837 ) | ( n4831 & n4837 ) ;
  assign n4839 = ( n4825 & n4831 ) | ( n4825 & n4837 ) | ( n4831 & n4837 ) ;
  assign n4840 = ( n4825 & n4838 ) | ( n4825 & ~n4839 ) | ( n4838 & ~n4839 ) ;
  assign n4841 = x14 & x55 ;
  assign n4842 = x21 & x48 ;
  assign n4843 = x22 & x47 ;
  assign n4844 = ( ~n4841 & n4842 ) | ( ~n4841 & n4843 ) | ( n4842 & n4843 ) ;
  assign n4845 = ( n4841 & n4842 ) | ( n4841 & n4843 ) | ( n4842 & n4843 ) ;
  assign n4846 = ( n4841 & n4844 ) | ( n4841 & ~n4845 ) | ( n4844 & ~n4845 ) ;
  assign n4847 = x11 & x58 ;
  assign n4848 = x12 & x57 ;
  assign n4849 = x13 & x56 ;
  assign n4850 = ( ~n4847 & n4848 ) | ( ~n4847 & n4849 ) | ( n4848 & n4849 ) ;
  assign n4851 = ( n4847 & n4848 ) | ( n4847 & n4849 ) | ( n4848 & n4849 ) ;
  assign n4852 = ( n4847 & n4850 ) | ( n4847 & ~n4851 ) | ( n4850 & ~n4851 ) ;
  assign n4853 = ( n4757 & n4846 ) | ( n4757 & n4852 ) | ( n4846 & n4852 ) ;
  assign n4854 = ( ~n4757 & n4846 ) | ( ~n4757 & n4852 ) | ( n4846 & n4852 ) ;
  assign n4855 = ( n4757 & ~n4853 ) | ( n4757 & n4854 ) | ( ~n4853 & n4854 ) ;
  assign n4856 = ( ~n4752 & n4840 ) | ( ~n4752 & n4855 ) | ( n4840 & n4855 ) ;
  assign n4857 = ( n4752 & n4840 ) | ( n4752 & n4855 ) | ( n4840 & n4855 ) ;
  assign n4858 = ( n4752 & n4856 ) | ( n4752 & ~n4857 ) | ( n4856 & ~n4857 ) ;
  assign n4859 = x28 & x41 ;
  assign n4860 = x29 & x40 ;
  assign n4861 = x30 & x39 ;
  assign n4862 = ( ~n4859 & n4860 ) | ( ~n4859 & n4861 ) | ( n4860 & n4861 ) ;
  assign n4863 = ( n4859 & n4860 ) | ( n4859 & n4861 ) | ( n4860 & n4861 ) ;
  assign n4864 = ( n4859 & n4862 ) | ( n4859 & ~n4863 ) | ( n4862 & ~n4863 ) ;
  assign n4865 = x19 & x50 ;
  assign n4866 = x18 & x51 ;
  assign n4867 = x17 & x52 ;
  assign n4868 = ( ~n4865 & n4866 ) | ( ~n4865 & n4867 ) | ( n4866 & n4867 ) ;
  assign n4869 = ( n4865 & n4866 ) | ( n4865 & n4867 ) | ( n4866 & n4867 ) ;
  assign n4870 = ( n4865 & n4868 ) | ( n4865 & ~n4869 ) | ( n4868 & ~n4869 ) ;
  assign n4871 = ( n4773 & n4864 ) | ( n4773 & n4870 ) | ( n4864 & n4870 ) ;
  assign n4872 = ( ~n4773 & n4864 ) | ( ~n4773 & n4870 ) | ( n4864 & n4870 ) ;
  assign n4873 = ( n4773 & ~n4871 ) | ( n4773 & n4872 ) | ( ~n4871 & n4872 ) ;
  assign n4874 = x34 & x35 ;
  assign n4875 = x7 & x62 ;
  assign n4876 = ( x35 & n4874 ) | ( x35 & n4875 ) | ( n4874 & n4875 ) ;
  assign n4877 = ( x35 & ~n4874 ) | ( x35 & n4875 ) | ( ~n4874 & n4875 ) ;
  assign n4878 = ( n4874 & ~n4876 ) | ( n4874 & n4877 ) | ( ~n4876 & n4877 ) ;
  assign n4879 = x31 & x38 ;
  assign n4880 = x32 & x37 ;
  assign n4881 = x33 & x36 ;
  assign n4882 = ( ~n4879 & n4880 ) | ( ~n4879 & n4881 ) | ( n4880 & n4881 ) ;
  assign n4883 = ( n4879 & n4880 ) | ( n4879 & n4881 ) | ( n4880 & n4881 ) ;
  assign n4884 = ( n4879 & n4882 ) | ( n4879 & ~n4883 ) | ( n4882 & ~n4883 ) ;
  assign n4885 = x16 & x53 ;
  assign n4886 = x15 & x54 ;
  assign n4887 = x20 & x49 ;
  assign n4888 = ( ~n4885 & n4886 ) | ( ~n4885 & n4887 ) | ( n4886 & n4887 ) ;
  assign n4889 = ( n4885 & n4886 ) | ( n4885 & n4887 ) | ( n4886 & n4887 ) ;
  assign n4890 = ( n4885 & n4888 ) | ( n4885 & ~n4889 ) | ( n4888 & ~n4889 ) ;
  assign n4891 = ( n4878 & n4884 ) | ( n4878 & n4890 ) | ( n4884 & n4890 ) ;
  assign n4892 = ( ~n4878 & n4884 ) | ( ~n4878 & n4890 ) | ( n4884 & n4890 ) ;
  assign n4893 = ( n4878 & ~n4891 ) | ( n4878 & n4892 ) | ( ~n4891 & n4892 ) ;
  assign n4894 = ( ~n4770 & n4873 ) | ( ~n4770 & n4893 ) | ( n4873 & n4893 ) ;
  assign n4895 = ( n4770 & n4873 ) | ( n4770 & n4893 ) | ( n4873 & n4893 ) ;
  assign n4896 = ( n4770 & n4894 ) | ( n4770 & ~n4895 ) | ( n4894 & ~n4895 ) ;
  assign n4897 = ( ~n4763 & n4858 ) | ( ~n4763 & n4896 ) | ( n4858 & n4896 ) ;
  assign n4898 = ( n4763 & n4858 ) | ( n4763 & n4896 ) | ( n4858 & n4896 ) ;
  assign n4899 = ( n4763 & n4897 ) | ( n4763 & ~n4898 ) | ( n4897 & ~n4898 ) ;
  assign n4900 = ( ~n4746 & n4785 ) | ( ~n4746 & n4899 ) | ( n4785 & n4899 ) ;
  assign n4901 = ( n4746 & n4785 ) | ( n4746 & n4899 ) | ( n4785 & n4899 ) ;
  assign n4902 = ( n4746 & n4900 ) | ( n4746 & ~n4901 ) | ( n4900 & ~n4901 ) ;
  assign n4903 = ( ~n4750 & n4819 ) | ( ~n4750 & n4902 ) | ( n4819 & n4902 ) ;
  assign n4904 = ( n4750 & n4819 ) | ( n4750 & n4902 ) | ( n4819 & n4902 ) ;
  assign n4905 = ( n4750 & n4903 ) | ( n4750 & ~n4904 ) | ( n4903 & ~n4904 ) ;
  assign n4906 = ( n4788 & n4790 ) | ( n4788 & n4905 ) | ( n4790 & n4905 ) ;
  assign n4907 = ( ~n4788 & n4790 ) | ( ~n4788 & n4905 ) | ( n4790 & n4905 ) ;
  assign n4908 = ( n4788 & ~n4906 ) | ( n4788 & n4907 ) | ( ~n4906 & n4907 ) ;
  assign n4909 = ( n4836 & ~n4845 ) | ( n4836 & n4851 ) | ( ~n4845 & n4851 ) ;
  assign n4910 = ( n4836 & n4845 ) | ( n4836 & n4851 ) | ( n4845 & n4851 ) ;
  assign n4911 = ( n4845 & n4909 ) | ( n4845 & ~n4910 ) | ( n4909 & ~n4910 ) ;
  assign n4912 = ( n4794 & n4809 ) | ( n4794 & n4911 ) | ( n4809 & n4911 ) ;
  assign n4913 = ( ~n4794 & n4809 ) | ( ~n4794 & n4911 ) | ( n4809 & n4911 ) ;
  assign n4914 = ( n4794 & ~n4912 ) | ( n4794 & n4913 ) | ( ~n4912 & n4913 ) ;
  assign n4915 = ( n4803 & n4857 ) | ( n4803 & n4914 ) | ( n4857 & n4914 ) ;
  assign n4916 = ( ~n4803 & n4857 ) | ( ~n4803 & n4914 ) | ( n4857 & n4914 ) ;
  assign n4917 = ( n4803 & ~n4915 ) | ( n4803 & n4916 ) | ( ~n4915 & n4916 ) ;
  assign n4918 = ( n4815 & n4898 ) | ( n4815 & n4917 ) | ( n4898 & n4917 ) ;
  assign n4919 = ( n4815 & n4898 ) | ( n4815 & ~n4917 ) | ( n4898 & ~n4917 ) ;
  assign n4920 = ( n4917 & ~n4918 ) | ( n4917 & n4919 ) | ( ~n4918 & n4919 ) ;
  assign n4921 = ( ~n4824 & n4830 ) | ( ~n4824 & n4863 ) | ( n4830 & n4863 ) ;
  assign n4922 = ( n4824 & n4830 ) | ( n4824 & n4863 ) | ( n4830 & n4863 ) ;
  assign n4923 = ( n4824 & n4921 ) | ( n4824 & ~n4922 ) | ( n4921 & ~n4922 ) ;
  assign n4924 = x8 & x62 ;
  assign n4925 = ( n4876 & n4883 ) | ( n4876 & n4924 ) | ( n4883 & n4924 ) ;
  assign n4926 = ( n4876 & ~n4883 ) | ( n4876 & n4924 ) | ( ~n4883 & n4924 ) ;
  assign n4927 = ( n4883 & ~n4925 ) | ( n4883 & n4926 ) | ( ~n4925 & n4926 ) ;
  assign n4928 = ( ~n4871 & n4923 ) | ( ~n4871 & n4927 ) | ( n4923 & n4927 ) ;
  assign n4929 = ( n4871 & n4923 ) | ( n4871 & n4927 ) | ( n4923 & n4927 ) ;
  assign n4930 = ( n4871 & n4928 ) | ( n4871 & ~n4929 ) | ( n4928 & ~n4929 ) ;
  assign n4931 = ( n4839 & ~n4853 ) | ( n4839 & n4891 ) | ( ~n4853 & n4891 ) ;
  assign n4932 = ( n4839 & n4853 ) | ( n4839 & n4891 ) | ( n4853 & n4891 ) ;
  assign n4933 = ( n4853 & n4931 ) | ( n4853 & ~n4932 ) | ( n4931 & ~n4932 ) ;
  assign n4934 = ( ~n4895 & n4930 ) | ( ~n4895 & n4933 ) | ( n4930 & n4933 ) ;
  assign n4935 = ( n4895 & n4930 ) | ( n4895 & n4933 ) | ( n4930 & n4933 ) ;
  assign n4936 = ( n4895 & n4934 ) | ( n4895 & ~n4935 ) | ( n4934 & ~n4935 ) ;
  assign n4937 = x32 & x38 ;
  assign n4938 = x33 & x37 ;
  assign n4939 = x34 & x36 ;
  assign n4940 = ( ~n4937 & n4938 ) | ( ~n4937 & n4939 ) | ( n4938 & n4939 ) ;
  assign n4941 = ( n4937 & n4938 ) | ( n4937 & n4939 ) | ( n4938 & n4939 ) ;
  assign n4942 = ( n4937 & n4940 ) | ( n4937 & ~n4941 ) | ( n4940 & ~n4941 ) ;
  assign n4943 = ( ~n4869 & n4889 ) | ( ~n4869 & n4942 ) | ( n4889 & n4942 ) ;
  assign n4944 = ( n4869 & n4889 ) | ( n4869 & n4942 ) | ( n4889 & n4942 ) ;
  assign n4945 = ( n4869 & n4943 ) | ( n4869 & ~n4944 ) | ( n4943 & ~n4944 ) ;
  assign n4946 = x12 & x58 ;
  assign n4947 = x13 & x57 ;
  assign n4948 = ( ~n2370 & n4946 ) | ( ~n2370 & n4947 ) | ( n4946 & n4947 ) ;
  assign n4949 = ( n2370 & n4946 ) | ( n2370 & n4947 ) | ( n4946 & n4947 ) ;
  assign n4950 = ( n2370 & n4948 ) | ( n2370 & ~n4949 ) | ( n4948 & ~n4949 ) ;
  assign n4951 = x18 & x52 ;
  assign n4952 = x17 & x53 ;
  assign n4953 = x16 & x54 ;
  assign n4954 = ( ~n4951 & n4952 ) | ( ~n4951 & n4953 ) | ( n4952 & n4953 ) ;
  assign n4955 = ( n4951 & n4952 ) | ( n4951 & n4953 ) | ( n4952 & n4953 ) ;
  assign n4956 = ( n4951 & n4954 ) | ( n4951 & ~n4955 ) | ( n4954 & ~n4955 ) ;
  assign n4957 = x9 & x61 ;
  assign n4958 = x10 & x60 ;
  assign n4959 = x11 & x59 ;
  assign n4960 = ( ~n4957 & n4958 ) | ( ~n4957 & n4959 ) | ( n4958 & n4959 ) ;
  assign n4961 = ( n4957 & n4958 ) | ( n4957 & n4959 ) | ( n4958 & n4959 ) ;
  assign n4962 = ( n4957 & n4960 ) | ( n4957 & ~n4961 ) | ( n4960 & ~n4961 ) ;
  assign n4963 = ( ~n4950 & n4956 ) | ( ~n4950 & n4962 ) | ( n4956 & n4962 ) ;
  assign n4964 = ( n4950 & n4956 ) | ( n4950 & n4962 ) | ( n4956 & n4962 ) ;
  assign n4965 = ( n4950 & n4963 ) | ( n4950 & ~n4964 ) | ( n4963 & ~n4964 ) ;
  assign n4966 = ( n4796 & n4945 ) | ( n4796 & n4965 ) | ( n4945 & n4965 ) ;
  assign n4967 = ( ~n4796 & n4945 ) | ( ~n4796 & n4965 ) | ( n4945 & n4965 ) ;
  assign n4968 = ( n4796 & ~n4966 ) | ( n4796 & n4967 ) | ( ~n4966 & n4967 ) ;
  assign n4969 = x28 & x42 ;
  assign n4970 = x23 & x47 ;
  assign n4971 = x7 & x63 ;
  assign n4972 = ( ~n4969 & n4970 ) | ( ~n4969 & n4971 ) | ( n4970 & n4971 ) ;
  assign n4973 = ( n4969 & n4970 ) | ( n4969 & n4971 ) | ( n4970 & n4971 ) ;
  assign n4974 = ( n4969 & n4972 ) | ( n4969 & ~n4973 ) | ( n4972 & ~n4973 ) ;
  assign n4975 = x29 & x41 ;
  assign n4976 = x30 & x40 ;
  assign n4977 = x31 & x39 ;
  assign n4978 = ( ~n4975 & n4976 ) | ( ~n4975 & n4977 ) | ( n4976 & n4977 ) ;
  assign n4979 = ( n4975 & n4976 ) | ( n4975 & n4977 ) | ( n4976 & n4977 ) ;
  assign n4980 = ( n4975 & n4978 ) | ( n4975 & ~n4979 ) | ( n4978 & ~n4979 ) ;
  assign n4981 = ( ~n4806 & n4974 ) | ( ~n4806 & n4980 ) | ( n4974 & n4980 ) ;
  assign n4982 = ( n4806 & n4974 ) | ( n4806 & n4980 ) | ( n4974 & n4980 ) ;
  assign n4983 = ( n4806 & n4981 ) | ( n4806 & ~n4982 ) | ( n4981 & ~n4982 ) ;
  assign n4984 = x21 & x49 ;
  assign n4985 = x19 & x51 ;
  assign n4986 = x20 & x50 ;
  assign n4987 = ( ~n4984 & n4985 ) | ( ~n4984 & n4986 ) | ( n4985 & n4986 ) ;
  assign n4988 = ( n4984 & n4985 ) | ( n4984 & n4986 ) | ( n4985 & n4986 ) ;
  assign n4989 = ( n4984 & n4987 ) | ( n4984 & ~n4988 ) | ( n4987 & ~n4988 ) ;
  assign n4990 = x25 & x45 ;
  assign n4991 = x27 & x43 ;
  assign n4992 = x26 & x44 ;
  assign n4993 = ( ~n4990 & n4991 ) | ( ~n4990 & n4992 ) | ( n4991 & n4992 ) ;
  assign n4994 = ( n4990 & n4991 ) | ( n4990 & n4992 ) | ( n4991 & n4992 ) ;
  assign n4995 = ( n4990 & n4993 ) | ( n4990 & ~n4994 ) | ( n4993 & ~n4994 ) ;
  assign n4996 = x22 & x48 ;
  assign n4997 = x14 & x56 ;
  assign n4998 = x15 & x55 ;
  assign n4999 = ( ~n4996 & n4997 ) | ( ~n4996 & n4998 ) | ( n4997 & n4998 ) ;
  assign n5000 = ( n4996 & n4997 ) | ( n4996 & n4998 ) | ( n4997 & n4998 ) ;
  assign n5001 = ( n4996 & n4999 ) | ( n4996 & ~n5000 ) | ( n4999 & ~n5000 ) ;
  assign n5002 = ( ~n4989 & n4995 ) | ( ~n4989 & n5001 ) | ( n4995 & n5001 ) ;
  assign n5003 = ( n4989 & n4995 ) | ( n4989 & n5001 ) | ( n4995 & n5001 ) ;
  assign n5004 = ( n4989 & n5002 ) | ( n4989 & ~n5003 ) | ( n5002 & ~n5003 ) ;
  assign n5005 = ( n4811 & n4983 ) | ( n4811 & n5004 ) | ( n4983 & n5004 ) ;
  assign n5006 = ( ~n4811 & n4983 ) | ( ~n4811 & n5004 ) | ( n4983 & n5004 ) ;
  assign n5007 = ( n4811 & ~n5005 ) | ( n4811 & n5006 ) | ( ~n5005 & n5006 ) ;
  assign n5008 = ( n4799 & n4968 ) | ( n4799 & n5007 ) | ( n4968 & n5007 ) ;
  assign n5009 = ( ~n4799 & n4968 ) | ( ~n4799 & n5007 ) | ( n4968 & n5007 ) ;
  assign n5010 = ( n4799 & ~n5008 ) | ( n4799 & n5009 ) | ( ~n5008 & n5009 ) ;
  assign n5011 = ( ~n4818 & n4936 ) | ( ~n4818 & n5010 ) | ( n4936 & n5010 ) ;
  assign n5012 = ( n4818 & n4936 ) | ( n4818 & n5010 ) | ( n4936 & n5010 ) ;
  assign n5013 = ( n4818 & n5011 ) | ( n4818 & ~n5012 ) | ( n5011 & ~n5012 ) ;
  assign n5014 = ( n4901 & n4920 ) | ( n4901 & n5013 ) | ( n4920 & n5013 ) ;
  assign n5015 = ( ~n4901 & n4920 ) | ( ~n4901 & n5013 ) | ( n4920 & n5013 ) ;
  assign n5016 = ( n4901 & ~n5014 ) | ( n4901 & n5015 ) | ( ~n5014 & n5015 ) ;
  assign n5017 = ( n4904 & n4906 ) | ( n4904 & n5016 ) | ( n4906 & n5016 ) ;
  assign n5018 = ( ~n4904 & n4906 ) | ( ~n4904 & n5016 ) | ( n4906 & n5016 ) ;
  assign n5019 = ( n4904 & ~n5017 ) | ( n4904 & n5018 ) | ( ~n5017 & n5018 ) ;
  assign n5020 = ( n4922 & n4925 ) | ( n4922 & n4944 ) | ( n4925 & n4944 ) ;
  assign n5021 = ( n4922 & ~n4925 ) | ( n4922 & n4944 ) | ( ~n4925 & n4944 ) ;
  assign n5022 = ( n4925 & ~n5020 ) | ( n4925 & n5021 ) | ( ~n5020 & n5021 ) ;
  assign n5023 = ( ~n4929 & n4966 ) | ( ~n4929 & n5022 ) | ( n4966 & n5022 ) ;
  assign n5024 = ( n4929 & n4966 ) | ( n4929 & n5022 ) | ( n4966 & n5022 ) ;
  assign n5025 = ( n4929 & n5023 ) | ( n4929 & ~n5024 ) | ( n5023 & ~n5024 ) ;
  assign n5026 = ( ~n4935 & n5008 ) | ( ~n4935 & n5025 ) | ( n5008 & n5025 ) ;
  assign n5027 = ( n4935 & n5008 ) | ( n4935 & n5025 ) | ( n5008 & n5025 ) ;
  assign n5028 = ( n4935 & n5026 ) | ( n4935 & ~n5027 ) | ( n5026 & ~n5027 ) ;
  assign n5029 = x11 & x60 ;
  assign n5030 = x8 & x63 ;
  assign n5031 = x10 & x61 ;
  assign n5032 = ( ~n5029 & n5030 ) | ( ~n5029 & n5031 ) | ( n5030 & n5031 ) ;
  assign n5033 = ( n5029 & n5030 ) | ( n5029 & n5031 ) | ( n5030 & n5031 ) ;
  assign n5034 = ( n5029 & n5032 ) | ( n5029 & ~n5033 ) | ( n5032 & ~n5033 ) ;
  assign n5035 = ( ~n4941 & n4955 ) | ( ~n4941 & n5034 ) | ( n4955 & n5034 ) ;
  assign n5036 = ( n4941 & n4955 ) | ( n4941 & n5034 ) | ( n4955 & n5034 ) ;
  assign n5037 = ( n4941 & n5035 ) | ( n4941 & ~n5036 ) | ( n5035 & ~n5036 ) ;
  assign n5038 = x21 & x50 ;
  assign n5039 = x20 & x51 ;
  assign n5040 = x19 & x52 ;
  assign n5041 = ( ~n5038 & n5039 ) | ( ~n5038 & n5040 ) | ( n5039 & n5040 ) ;
  assign n5042 = ( n5038 & n5039 ) | ( n5038 & n5040 ) | ( n5039 & n5040 ) ;
  assign n5043 = ( n5038 & n5041 ) | ( n5038 & ~n5042 ) | ( n5041 & ~n5042 ) ;
  assign n5044 = x22 & x49 ;
  assign n5045 = x9 & x62 ;
  assign n5046 = ( ~x36 & n5044 ) | ( ~x36 & n5045 ) | ( n5044 & n5045 ) ;
  assign n5047 = ( x36 & n5044 ) | ( x36 & n5045 ) | ( n5044 & n5045 ) ;
  assign n5048 = ( x36 & n5046 ) | ( x36 & ~n5047 ) | ( n5046 & ~n5047 ) ;
  assign n5049 = x34 & x37 ;
  assign n5050 = x33 & x38 ;
  assign n5051 = x35 & x36 ;
  assign n5052 = ( ~n5049 & n5050 ) | ( ~n5049 & n5051 ) | ( n5050 & n5051 ) ;
  assign n5053 = ( n5049 & n5050 ) | ( n5049 & n5051 ) | ( n5050 & n5051 ) ;
  assign n5054 = ( n5049 & n5052 ) | ( n5049 & ~n5053 ) | ( n5052 & ~n5053 ) ;
  assign n5055 = ( ~n5043 & n5048 ) | ( ~n5043 & n5054 ) | ( n5048 & n5054 ) ;
  assign n5056 = ( n5043 & n5048 ) | ( n5043 & n5054 ) | ( n5048 & n5054 ) ;
  assign n5057 = ( n5043 & n5055 ) | ( n5043 & ~n5056 ) | ( n5055 & ~n5056 ) ;
  assign n5058 = ( n4912 & n5037 ) | ( n4912 & n5057 ) | ( n5037 & n5057 ) ;
  assign n5059 = ( ~n4912 & n5037 ) | ( ~n4912 & n5057 ) | ( n5037 & n5057 ) ;
  assign n5060 = ( n4912 & ~n5058 ) | ( n4912 & n5059 ) | ( ~n5058 & n5059 ) ;
  assign n5061 = x30 & x41 ;
  assign n5062 = x31 & x40 ;
  assign n5063 = x32 & x39 ;
  assign n5064 = ( ~n5061 & n5062 ) | ( ~n5061 & n5063 ) | ( n5062 & n5063 ) ;
  assign n5065 = ( n5061 & n5062 ) | ( n5061 & n5063 ) | ( n5062 & n5063 ) ;
  assign n5066 = ( n5061 & n5064 ) | ( n5061 & ~n5065 ) | ( n5064 & ~n5065 ) ;
  assign n5067 = x23 & x48 ;
  assign n5068 = x17 & x54 ;
  assign n5069 = x18 & x53 ;
  assign n5070 = ( ~n5067 & n5068 ) | ( ~n5067 & n5069 ) | ( n5068 & n5069 ) ;
  assign n5071 = ( n5067 & n5068 ) | ( n5067 & n5069 ) | ( n5068 & n5069 ) ;
  assign n5072 = ( n5067 & n5070 ) | ( n5067 & ~n5071 ) | ( n5070 & ~n5071 ) ;
  assign n5073 = x27 & x44 ;
  assign n5074 = x28 & x43 ;
  assign n5075 = x29 & x42 ;
  assign n5076 = ( ~n5073 & n5074 ) | ( ~n5073 & n5075 ) | ( n5074 & n5075 ) ;
  assign n5077 = ( n5073 & n5074 ) | ( n5073 & n5075 ) | ( n5074 & n5075 ) ;
  assign n5078 = ( n5073 & n5076 ) | ( n5073 & ~n5077 ) | ( n5076 & ~n5077 ) ;
  assign n5079 = ( ~n5066 & n5072 ) | ( ~n5066 & n5078 ) | ( n5072 & n5078 ) ;
  assign n5080 = ( n5066 & n5072 ) | ( n5066 & n5078 ) | ( n5072 & n5078 ) ;
  assign n5081 = ( n5066 & n5079 ) | ( n5066 & ~n5080 ) | ( n5079 & ~n5080 ) ;
  assign n5082 = x14 & x57 ;
  assign n5083 = x15 & x56 ;
  assign n5084 = x16 & x55 ;
  assign n5085 = ( ~n5082 & n5083 ) | ( ~n5082 & n5084 ) | ( n5083 & n5084 ) ;
  assign n5086 = ( n5082 & n5083 ) | ( n5082 & n5084 ) | ( n5083 & n5084 ) ;
  assign n5087 = ( n5082 & n5085 ) | ( n5082 & ~n5086 ) | ( n5085 & ~n5086 ) ;
  assign n5088 = x24 & x47 ;
  assign n5089 = x25 & x46 ;
  assign n5090 = x26 & x45 ;
  assign n5091 = ( ~n5088 & n5089 ) | ( ~n5088 & n5090 ) | ( n5089 & n5090 ) ;
  assign n5092 = ( n5088 & n5089 ) | ( n5088 & n5090 ) | ( n5089 & n5090 ) ;
  assign n5093 = ( n5088 & n5091 ) | ( n5088 & ~n5092 ) | ( n5091 & ~n5092 ) ;
  assign n5094 = x13 & x58 ;
  assign n5095 = x12 & x59 ;
  assign n5096 = ( n4988 & n5094 ) | ( n4988 & n5095 ) | ( n5094 & n5095 ) ;
  assign n5097 = ( ~n4988 & n5094 ) | ( ~n4988 & n5095 ) | ( n5094 & n5095 ) ;
  assign n5098 = ( n4988 & ~n5096 ) | ( n4988 & n5097 ) | ( ~n5096 & n5097 ) ;
  assign n5099 = ( ~n5087 & n5093 ) | ( ~n5087 & n5098 ) | ( n5093 & n5098 ) ;
  assign n5100 = ( n5087 & n5093 ) | ( n5087 & n5098 ) | ( n5093 & n5098 ) ;
  assign n5101 = ( n5087 & n5099 ) | ( n5087 & ~n5100 ) | ( n5099 & ~n5100 ) ;
  assign n5102 = ( ~n4932 & n5081 ) | ( ~n4932 & n5101 ) | ( n5081 & n5101 ) ;
  assign n5103 = ( n4932 & n5081 ) | ( n4932 & n5101 ) | ( n5081 & n5101 ) ;
  assign n5104 = ( n4932 & n5102 ) | ( n4932 & ~n5103 ) | ( n5102 & ~n5103 ) ;
  assign n5105 = ( ~n4915 & n5060 ) | ( ~n4915 & n5104 ) | ( n5060 & n5104 ) ;
  assign n5106 = ( n4915 & n5060 ) | ( n4915 & n5104 ) | ( n5060 & n5104 ) ;
  assign n5107 = ( n4915 & n5105 ) | ( n4915 & ~n5106 ) | ( n5105 & ~n5106 ) ;
  assign n5108 = ( ~n4910 & n4964 ) | ( ~n4910 & n5003 ) | ( n4964 & n5003 ) ;
  assign n5109 = ( n4910 & n4964 ) | ( n4910 & n5003 ) | ( n4964 & n5003 ) ;
  assign n5110 = ( n4910 & n5108 ) | ( n4910 & ~n5109 ) | ( n5108 & ~n5109 ) ;
  assign n5111 = ( n4949 & ~n4961 ) | ( n4949 & n4994 ) | ( ~n4961 & n4994 ) ;
  assign n5112 = ( n4949 & n4961 ) | ( n4949 & n4994 ) | ( n4961 & n4994 ) ;
  assign n5113 = ( n4961 & n5111 ) | ( n4961 & ~n5112 ) | ( n5111 & ~n5112 ) ;
  assign n5114 = ( n4973 & ~n4979 ) | ( n4973 & n5000 ) | ( ~n4979 & n5000 ) ;
  assign n5115 = ( n4973 & n4979 ) | ( n4973 & n5000 ) | ( n4979 & n5000 ) ;
  assign n5116 = ( n4979 & n5114 ) | ( n4979 & ~n5115 ) | ( n5114 & ~n5115 ) ;
  assign n5117 = ( ~n4982 & n5113 ) | ( ~n4982 & n5116 ) | ( n5113 & n5116 ) ;
  assign n5118 = ( n4982 & n5113 ) | ( n4982 & n5116 ) | ( n5113 & n5116 ) ;
  assign n5119 = ( n4982 & n5117 ) | ( n4982 & ~n5118 ) | ( n5117 & ~n5118 ) ;
  assign n5120 = ( n5005 & n5110 ) | ( n5005 & n5119 ) | ( n5110 & n5119 ) ;
  assign n5121 = ( ~n5005 & n5110 ) | ( ~n5005 & n5119 ) | ( n5110 & n5119 ) ;
  assign n5122 = ( n5005 & ~n5120 ) | ( n5005 & n5121 ) | ( ~n5120 & n5121 ) ;
  assign n5123 = ( ~n4918 & n5107 ) | ( ~n4918 & n5122 ) | ( n5107 & n5122 ) ;
  assign n5124 = ( n4918 & n5107 ) | ( n4918 & n5122 ) | ( n5107 & n5122 ) ;
  assign n5125 = ( n4918 & n5123 ) | ( n4918 & ~n5124 ) | ( n5123 & ~n5124 ) ;
  assign n5126 = ( ~n5012 & n5028 ) | ( ~n5012 & n5125 ) | ( n5028 & n5125 ) ;
  assign n5127 = ( n5012 & n5028 ) | ( n5012 & n5125 ) | ( n5028 & n5125 ) ;
  assign n5128 = ( n5012 & n5126 ) | ( n5012 & ~n5127 ) | ( n5126 & ~n5127 ) ;
  assign n5129 = ( n5014 & n5017 ) | ( n5014 & n5128 ) | ( n5017 & n5128 ) ;
  assign n5130 = ( ~n5014 & n5017 ) | ( ~n5014 & n5128 ) | ( n5017 & n5128 ) ;
  assign n5131 = ( n5014 & ~n5129 ) | ( n5014 & n5130 ) | ( ~n5129 & n5130 ) ;
  assign n5132 = ( n5056 & n5080 ) | ( n5056 & n5112 ) | ( n5080 & n5112 ) ;
  assign n5133 = ( n5056 & n5080 ) | ( n5056 & ~n5112 ) | ( n5080 & ~n5112 ) ;
  assign n5134 = ( n5112 & ~n5132 ) | ( n5112 & n5133 ) | ( ~n5132 & n5133 ) ;
  assign n5135 = ( n5065 & n5071 ) | ( n5065 & n5077 ) | ( n5071 & n5077 ) ;
  assign n5136 = ( ~n5065 & n5071 ) | ( ~n5065 & n5077 ) | ( n5071 & n5077 ) ;
  assign n5137 = ( n5065 & ~n5135 ) | ( n5065 & n5136 ) | ( ~n5135 & n5136 ) ;
  assign n5138 = ( ~n5042 & n5047 ) | ( ~n5042 & n5053 ) | ( n5047 & n5053 ) ;
  assign n5139 = ( n5042 & n5047 ) | ( n5042 & n5053 ) | ( n5047 & n5053 ) ;
  assign n5140 = ( n5042 & n5138 ) | ( n5042 & ~n5139 ) | ( n5138 & ~n5139 ) ;
  assign n5141 = ( ~n5100 & n5137 ) | ( ~n5100 & n5140 ) | ( n5137 & n5140 ) ;
  assign n5142 = ( n5100 & n5137 ) | ( n5100 & n5140 ) | ( n5137 & n5140 ) ;
  assign n5143 = ( n5100 & n5141 ) | ( n5100 & ~n5142 ) | ( n5141 & ~n5142 ) ;
  assign n5144 = ( ~n5103 & n5134 ) | ( ~n5103 & n5143 ) | ( n5134 & n5143 ) ;
  assign n5145 = ( n5103 & n5134 ) | ( n5103 & n5143 ) | ( n5134 & n5143 ) ;
  assign n5146 = ( n5103 & n5144 ) | ( n5103 & ~n5145 ) | ( n5144 & ~n5145 ) ;
  assign n5147 = x12 & x60 ;
  assign n5148 = x24 & x48 ;
  assign n5149 = x25 & x47 ;
  assign n5150 = ( ~n5147 & n5148 ) | ( ~n5147 & n5149 ) | ( n5148 & n5149 ) ;
  assign n5151 = ( n5147 & n5148 ) | ( n5147 & n5149 ) | ( n5148 & n5149 ) ;
  assign n5152 = ( n5147 & n5150 ) | ( n5147 & ~n5151 ) | ( n5150 & ~n5151 ) ;
  assign n5153 = x9 & x63 ;
  assign n5154 = x10 & x62 ;
  assign n5155 = x11 & x61 ;
  assign n5156 = ( ~n5153 & n5154 ) | ( ~n5153 & n5155 ) | ( n5154 & n5155 ) ;
  assign n5157 = ( n5153 & n5154 ) | ( n5153 & n5155 ) | ( n5154 & n5155 ) ;
  assign n5158 = ( n5153 & n5156 ) | ( n5153 & ~n5157 ) | ( n5156 & ~n5157 ) ;
  assign n5159 = ( n5096 & n5152 ) | ( n5096 & n5158 ) | ( n5152 & n5158 ) ;
  assign n5160 = ( ~n5096 & n5152 ) | ( ~n5096 & n5158 ) | ( n5152 & n5158 ) ;
  assign n5161 = ( n5096 & ~n5159 ) | ( n5096 & n5160 ) | ( ~n5159 & n5160 ) ;
  assign n5162 = x35 & x37 ;
  assign n5163 = x21 & x51 ;
  assign n5164 = x22 & x50 ;
  assign n5165 = ( ~n5162 & n5163 ) | ( ~n5162 & n5164 ) | ( n5163 & n5164 ) ;
  assign n5166 = ( n5162 & n5163 ) | ( n5162 & n5164 ) | ( n5163 & n5164 ) ;
  assign n5167 = ( n5162 & n5165 ) | ( n5162 & ~n5166 ) | ( n5165 & ~n5166 ) ;
  assign n5168 = x17 & x55 ;
  assign n5169 = x18 & x54 ;
  assign n5170 = x20 & x52 ;
  assign n5171 = ( ~n5168 & n5169 ) | ( ~n5168 & n5170 ) | ( n5169 & n5170 ) ;
  assign n5172 = ( n5168 & n5169 ) | ( n5168 & n5170 ) | ( n5169 & n5170 ) ;
  assign n5173 = ( n5168 & n5171 ) | ( n5168 & ~n5172 ) | ( n5171 & ~n5172 ) ;
  assign n5174 = x16 & x56 ;
  assign n5175 = x32 & x40 ;
  assign n5176 = x23 & x49 ;
  assign n5177 = ( ~n5174 & n5175 ) | ( ~n5174 & n5176 ) | ( n5175 & n5176 ) ;
  assign n5178 = ( n5174 & n5175 ) | ( n5174 & n5176 ) | ( n5175 & n5176 ) ;
  assign n5179 = ( n5174 & n5177 ) | ( n5174 & ~n5178 ) | ( n5177 & ~n5178 ) ;
  assign n5180 = ( ~n5167 & n5173 ) | ( ~n5167 & n5179 ) | ( n5173 & n5179 ) ;
  assign n5181 = ( n5167 & n5173 ) | ( n5167 & n5179 ) | ( n5173 & n5179 ) ;
  assign n5182 = ( n5167 & n5180 ) | ( n5167 & ~n5181 ) | ( n5180 & ~n5181 ) ;
  assign n5183 = ( ~n5109 & n5161 ) | ( ~n5109 & n5182 ) | ( n5161 & n5182 ) ;
  assign n5184 = ( n5109 & n5161 ) | ( n5109 & n5182 ) | ( n5161 & n5182 ) ;
  assign n5185 = ( n5109 & n5183 ) | ( n5109 & ~n5184 ) | ( n5183 & ~n5184 ) ;
  assign n5186 = ( ~n5033 & n5086 ) | ( ~n5033 & n5092 ) | ( n5086 & n5092 ) ;
  assign n5187 = ( n5033 & n5086 ) | ( n5033 & n5092 ) | ( n5086 & n5092 ) ;
  assign n5188 = ( n5033 & n5186 ) | ( n5033 & ~n5187 ) | ( n5186 & ~n5187 ) ;
  assign n5189 = x26 & x46 ;
  assign n5190 = x27 & x45 ;
  assign n5191 = x28 & x44 ;
  assign n5192 = ( ~n5189 & n5190 ) | ( ~n5189 & n5191 ) | ( n5190 & n5191 ) ;
  assign n5193 = ( n5189 & n5190 ) | ( n5189 & n5191 ) | ( n5190 & n5191 ) ;
  assign n5194 = ( n5189 & n5192 ) | ( n5189 & ~n5193 ) | ( n5192 & ~n5193 ) ;
  assign n5195 = x19 & x53 ;
  assign n5196 = x34 & x38 ;
  assign n5197 = x33 & x39 ;
  assign n5198 = ( ~n5195 & n5196 ) | ( ~n5195 & n5197 ) | ( n5196 & n5197 ) ;
  assign n5199 = ( n5195 & n5196 ) | ( n5195 & n5197 ) | ( n5196 & n5197 ) ;
  assign n5200 = ( n5195 & n5198 ) | ( n5195 & ~n5199 ) | ( n5198 & ~n5199 ) ;
  assign n5201 = x13 & x59 ;
  assign n5202 = x14 & x58 ;
  assign n5203 = x15 & x57 ;
  assign n5204 = ( ~n5201 & n5202 ) | ( ~n5201 & n5203 ) | ( n5202 & n5203 ) ;
  assign n5205 = ( n5201 & n5202 ) | ( n5201 & n5203 ) | ( n5202 & n5203 ) ;
  assign n5206 = ( n5201 & n5204 ) | ( n5201 & ~n5205 ) | ( n5204 & ~n5205 ) ;
  assign n5207 = ( ~n5194 & n5200 ) | ( ~n5194 & n5206 ) | ( n5200 & n5206 ) ;
  assign n5208 = ( n5194 & n5200 ) | ( n5194 & n5206 ) | ( n5200 & n5206 ) ;
  assign n5209 = ( n5194 & n5207 ) | ( n5194 & ~n5208 ) | ( n5207 & ~n5208 ) ;
  assign n5210 = ( ~n5020 & n5188 ) | ( ~n5020 & n5209 ) | ( n5188 & n5209 ) ;
  assign n5211 = ( n5020 & n5188 ) | ( n5020 & n5209 ) | ( n5188 & n5209 ) ;
  assign n5212 = ( n5020 & n5210 ) | ( n5020 & ~n5211 ) | ( n5210 & ~n5211 ) ;
  assign n5213 = ( n5024 & n5185 ) | ( n5024 & n5212 ) | ( n5185 & n5212 ) ;
  assign n5214 = ( ~n5024 & n5185 ) | ( ~n5024 & n5212 ) | ( n5185 & n5212 ) ;
  assign n5215 = ( n5024 & ~n5213 ) | ( n5024 & n5214 ) | ( ~n5213 & n5214 ) ;
  assign n5216 = ( ~n5027 & n5146 ) | ( ~n5027 & n5215 ) | ( n5146 & n5215 ) ;
  assign n5217 = ( n5027 & n5146 ) | ( n5027 & n5215 ) | ( n5146 & n5215 ) ;
  assign n5218 = ( n5027 & n5216 ) | ( n5027 & ~n5217 ) | ( n5216 & ~n5217 ) ;
  assign n5219 = x29 & x43 ;
  assign n5220 = x31 & x41 ;
  assign n5221 = x30 & x42 ;
  assign n5222 = ( ~n5219 & n5220 ) | ( ~n5219 & n5221 ) | ( n5220 & n5221 ) ;
  assign n5223 = ( n5219 & n5220 ) | ( n5219 & n5221 ) | ( n5220 & n5221 ) ;
  assign n5224 = ( n5219 & n5222 ) | ( n5219 & ~n5223 ) | ( n5222 & ~n5223 ) ;
  assign n5225 = ( n5036 & n5115 ) | ( n5036 & n5224 ) | ( n5115 & n5224 ) ;
  assign n5226 = ( ~n5036 & n5115 ) | ( ~n5036 & n5224 ) | ( n5115 & n5224 ) ;
  assign n5227 = ( n5036 & ~n5225 ) | ( n5036 & n5226 ) | ( ~n5225 & n5226 ) ;
  assign n5228 = ( ~n5058 & n5118 ) | ( ~n5058 & n5227 ) | ( n5118 & n5227 ) ;
  assign n5229 = ( n5058 & n5118 ) | ( n5058 & n5227 ) | ( n5118 & n5227 ) ;
  assign n5230 = ( n5058 & n5228 ) | ( n5058 & ~n5229 ) | ( n5228 & ~n5229 ) ;
  assign n5231 = ( ~n5106 & n5120 ) | ( ~n5106 & n5230 ) | ( n5120 & n5230 ) ;
  assign n5232 = ( n5106 & n5120 ) | ( n5106 & n5230 ) | ( n5120 & n5230 ) ;
  assign n5233 = ( n5106 & n5231 ) | ( n5106 & ~n5232 ) | ( n5231 & ~n5232 ) ;
  assign n5234 = ( ~n5124 & n5218 ) | ( ~n5124 & n5233 ) | ( n5218 & n5233 ) ;
  assign n5235 = ( n5124 & n5218 ) | ( n5124 & n5233 ) | ( n5218 & n5233 ) ;
  assign n5236 = ( n5124 & n5234 ) | ( n5124 & ~n5235 ) | ( n5234 & ~n5235 ) ;
  assign n5237 = ( n5127 & n5129 ) | ( n5127 & n5236 ) | ( n5129 & n5236 ) ;
  assign n5238 = ( n5127 & ~n5129 ) | ( n5127 & n5236 ) | ( ~n5129 & n5236 ) ;
  assign n5239 = ( n5129 & ~n5237 ) | ( n5129 & n5238 ) | ( ~n5237 & n5238 ) ;
  assign n5240 = x31 & x42 ;
  assign n5241 = x32 & x41 ;
  assign n5242 = x33 & x40 ;
  assign n5243 = ( ~n5240 & n5241 ) | ( ~n5240 & n5242 ) | ( n5241 & n5242 ) ;
  assign n5244 = ( n5240 & n5241 ) | ( n5240 & n5242 ) | ( n5241 & n5242 ) ;
  assign n5245 = ( n5240 & n5243 ) | ( n5240 & ~n5244 ) | ( n5243 & ~n5244 ) ;
  assign n5246 = ( n5135 & n5187 ) | ( n5135 & n5245 ) | ( n5187 & n5245 ) ;
  assign n5247 = ( ~n5135 & n5187 ) | ( ~n5135 & n5245 ) | ( n5187 & n5245 ) ;
  assign n5248 = ( n5135 & ~n5246 ) | ( n5135 & n5247 ) | ( ~n5246 & n5247 ) ;
  assign n5249 = ( n5142 & n5211 ) | ( n5142 & n5248 ) | ( n5211 & n5248 ) ;
  assign n5250 = ( n5142 & n5211 ) | ( n5142 & ~n5248 ) | ( n5211 & ~n5248 ) ;
  assign n5251 = ( n5248 & ~n5249 ) | ( n5248 & n5250 ) | ( ~n5249 & n5250 ) ;
  assign n5252 = ( n5145 & n5213 ) | ( n5145 & n5251 ) | ( n5213 & n5251 ) ;
  assign n5253 = ( ~n5145 & n5213 ) | ( ~n5145 & n5251 ) | ( n5213 & n5251 ) ;
  assign n5254 = ( n5145 & ~n5252 ) | ( n5145 & n5253 ) | ( ~n5252 & n5253 ) ;
  assign n5255 = ( n5139 & ~n5159 ) | ( n5139 & n5208 ) | ( ~n5159 & n5208 ) ;
  assign n5256 = ( n5139 & n5159 ) | ( n5139 & n5208 ) | ( n5159 & n5208 ) ;
  assign n5257 = ( n5159 & n5255 ) | ( n5159 & ~n5256 ) | ( n5255 & ~n5256 ) ;
  assign n5258 = ( n5151 & ~n5157 ) | ( n5151 & n5172 ) | ( ~n5157 & n5172 ) ;
  assign n5259 = ( n5151 & n5157 ) | ( n5151 & n5172 ) | ( n5157 & n5172 ) ;
  assign n5260 = ( n5157 & n5258 ) | ( n5157 & ~n5259 ) | ( n5258 & ~n5259 ) ;
  assign n5261 = x13 & x60 ;
  assign n5262 = ( ~n5166 & n5199 ) | ( ~n5166 & n5261 ) | ( n5199 & n5261 ) ;
  assign n5263 = ( n5166 & n5199 ) | ( n5166 & n5261 ) | ( n5199 & n5261 ) ;
  assign n5264 = ( n5166 & n5262 ) | ( n5166 & ~n5263 ) | ( n5262 & ~n5263 ) ;
  assign n5265 = ( ~n5181 & n5260 ) | ( ~n5181 & n5264 ) | ( n5260 & n5264 ) ;
  assign n5266 = ( n5181 & n5260 ) | ( n5181 & n5264 ) | ( n5260 & n5264 ) ;
  assign n5267 = ( n5181 & n5265 ) | ( n5181 & ~n5266 ) | ( n5265 & ~n5266 ) ;
  assign n5268 = ( ~n5184 & n5257 ) | ( ~n5184 & n5267 ) | ( n5257 & n5267 ) ;
  assign n5269 = ( n5184 & n5257 ) | ( n5184 & n5267 ) | ( n5257 & n5267 ) ;
  assign n5270 = ( n5184 & n5268 ) | ( n5184 & ~n5269 ) | ( n5268 & ~n5269 ) ;
  assign n5271 = x18 & x55 ;
  assign n5272 = x19 & x54 ;
  assign n5273 = x24 & x49 ;
  assign n5274 = ( ~n5271 & n5272 ) | ( ~n5271 & n5273 ) | ( n5272 & n5273 ) ;
  assign n5275 = ( n5271 & n5272 ) | ( n5271 & n5273 ) | ( n5272 & n5273 ) ;
  assign n5276 = ( n5271 & n5274 ) | ( n5271 & ~n5275 ) | ( n5274 & ~n5275 ) ;
  assign n5277 = x22 & x51 ;
  assign n5278 = x20 & x53 ;
  assign n5279 = x21 & x52 ;
  assign n5280 = ( ~n5277 & n5278 ) | ( ~n5277 & n5279 ) | ( n5278 & n5279 ) ;
  assign n5281 = ( n5277 & n5278 ) | ( n5277 & n5279 ) | ( n5278 & n5279 ) ;
  assign n5282 = ( n5277 & n5280 ) | ( n5277 & ~n5281 ) | ( n5280 & ~n5281 ) ;
  assign n5283 = x23 & x50 ;
  assign n5284 = x11 & x62 ;
  assign n5285 = ( ~x37 & n5283 ) | ( ~x37 & n5284 ) | ( n5283 & n5284 ) ;
  assign n5286 = ( x37 & n5283 ) | ( x37 & n5284 ) | ( n5283 & n5284 ) ;
  assign n5287 = ( x37 & n5285 ) | ( x37 & ~n5286 ) | ( n5285 & ~n5286 ) ;
  assign n5288 = ( ~n5276 & n5282 ) | ( ~n5276 & n5287 ) | ( n5282 & n5287 ) ;
  assign n5289 = ( n5276 & n5282 ) | ( n5276 & n5287 ) | ( n5282 & n5287 ) ;
  assign n5290 = ( n5276 & n5288 ) | ( n5276 & ~n5289 ) | ( n5288 & ~n5289 ) ;
  assign n5291 = x17 & x56 ;
  assign n5292 = x26 & x47 ;
  assign n5293 = x27 & x46 ;
  assign n5294 = ( ~n5291 & n5292 ) | ( ~n5291 & n5293 ) | ( n5292 & n5293 ) ;
  assign n5295 = ( n5291 & n5292 ) | ( n5291 & n5293 ) | ( n5292 & n5293 ) ;
  assign n5296 = ( n5291 & n5294 ) | ( n5291 & ~n5295 ) | ( n5294 & ~n5295 ) ;
  assign n5297 = x14 & x59 ;
  assign n5298 = x15 & x58 ;
  assign n5299 = x16 & x57 ;
  assign n5300 = ( ~n5297 & n5298 ) | ( ~n5297 & n5299 ) | ( n5298 & n5299 ) ;
  assign n5301 = ( n5297 & n5298 ) | ( n5297 & n5299 ) | ( n5298 & n5299 ) ;
  assign n5302 = ( n5297 & n5300 ) | ( n5297 & ~n5301 ) | ( n5300 & ~n5301 ) ;
  assign n5303 = ( n5178 & n5296 ) | ( n5178 & n5302 ) | ( n5296 & n5302 ) ;
  assign n5304 = ( ~n5178 & n5296 ) | ( ~n5178 & n5302 ) | ( n5296 & n5302 ) ;
  assign n5305 = ( n5178 & ~n5303 ) | ( n5178 & n5304 ) | ( ~n5303 & n5304 ) ;
  assign n5306 = ( ~n5132 & n5290 ) | ( ~n5132 & n5305 ) | ( n5290 & n5305 ) ;
  assign n5307 = ( n5132 & n5290 ) | ( n5132 & n5305 ) | ( n5290 & n5305 ) ;
  assign n5308 = ( n5132 & n5306 ) | ( n5132 & ~n5307 ) | ( n5306 & ~n5307 ) ;
  assign n5309 = ( ~n5193 & n5205 ) | ( ~n5193 & n5223 ) | ( n5205 & n5223 ) ;
  assign n5310 = ( n5193 & n5205 ) | ( n5193 & n5223 ) | ( n5205 & n5223 ) ;
  assign n5311 = ( n5193 & n5309 ) | ( n5193 & ~n5310 ) | ( n5309 & ~n5310 ) ;
  assign n5312 = x28 & x45 ;
  assign n5313 = x29 & x44 ;
  assign n5314 = x30 & x43 ;
  assign n5315 = ( ~n5312 & n5313 ) | ( ~n5312 & n5314 ) | ( n5313 & n5314 ) ;
  assign n5316 = ( n5312 & n5313 ) | ( n5312 & n5314 ) | ( n5313 & n5314 ) ;
  assign n5317 = ( n5312 & n5315 ) | ( n5312 & ~n5316 ) | ( n5315 & ~n5316 ) ;
  assign n5318 = x34 & x39 ;
  assign n5319 = x36 & x37 ;
  assign n5320 = x35 & x38 ;
  assign n5321 = ( ~n5318 & n5319 ) | ( ~n5318 & n5320 ) | ( n5319 & n5320 ) ;
  assign n5322 = ( n5318 & n5319 ) | ( n5318 & n5320 ) | ( n5319 & n5320 ) ;
  assign n5323 = ( n5318 & n5321 ) | ( n5318 & ~n5322 ) | ( n5321 & ~n5322 ) ;
  assign n5324 = x25 & x48 ;
  assign n5325 = x10 & x63 ;
  assign n5326 = x12 & x61 ;
  assign n5327 = ( ~n5324 & n5325 ) | ( ~n5324 & n5326 ) | ( n5325 & n5326 ) ;
  assign n5328 = ( n5324 & n5325 ) | ( n5324 & n5326 ) | ( n5325 & n5326 ) ;
  assign n5329 = ( n5324 & n5327 ) | ( n5324 & ~n5328 ) | ( n5327 & ~n5328 ) ;
  assign n5330 = ( ~n5317 & n5323 ) | ( ~n5317 & n5329 ) | ( n5323 & n5329 ) ;
  assign n5331 = ( n5317 & n5323 ) | ( n5317 & n5329 ) | ( n5323 & n5329 ) ;
  assign n5332 = ( n5317 & n5330 ) | ( n5317 & ~n5331 ) | ( n5330 & ~n5331 ) ;
  assign n5333 = ( ~n5225 & n5311 ) | ( ~n5225 & n5332 ) | ( n5311 & n5332 ) ;
  assign n5334 = ( n5225 & n5311 ) | ( n5225 & n5332 ) | ( n5311 & n5332 ) ;
  assign n5335 = ( n5225 & n5333 ) | ( n5225 & ~n5334 ) | ( n5333 & ~n5334 ) ;
  assign n5336 = ( n5229 & n5308 ) | ( n5229 & n5335 ) | ( n5308 & n5335 ) ;
  assign n5337 = ( ~n5229 & n5308 ) | ( ~n5229 & n5335 ) | ( n5308 & n5335 ) ;
  assign n5338 = ( n5229 & ~n5336 ) | ( n5229 & n5337 ) | ( ~n5336 & n5337 ) ;
  assign n5339 = ( ~n5232 & n5270 ) | ( ~n5232 & n5338 ) | ( n5270 & n5338 ) ;
  assign n5340 = ( n5232 & n5270 ) | ( n5232 & n5338 ) | ( n5270 & n5338 ) ;
  assign n5341 = ( n5232 & n5339 ) | ( n5232 & ~n5340 ) | ( n5339 & ~n5340 ) ;
  assign n5342 = ( ~n5217 & n5254 ) | ( ~n5217 & n5341 ) | ( n5254 & n5341 ) ;
  assign n5343 = ( n5217 & n5254 ) | ( n5217 & n5341 ) | ( n5254 & n5341 ) ;
  assign n5344 = ( n5217 & n5342 ) | ( n5217 & ~n5343 ) | ( n5342 & ~n5343 ) ;
  assign n5345 = ( ~n5235 & n5237 ) | ( ~n5235 & n5344 ) | ( n5237 & n5344 ) ;
  assign n5346 = ( n5235 & n5237 ) | ( n5235 & n5344 ) | ( n5237 & n5344 ) ;
  assign n5347 = ( n5235 & n5345 ) | ( n5235 & ~n5346 ) | ( n5345 & ~n5346 ) ;
  assign n5348 = x14 & x60 ;
  assign n5349 = x16 & x58 ;
  assign n5350 = x15 & x59 ;
  assign n5351 = ( ~n5348 & n5349 ) | ( ~n5348 & n5350 ) | ( n5349 & n5350 ) ;
  assign n5352 = ( n5348 & n5349 ) | ( n5348 & n5350 ) | ( n5349 & n5350 ) ;
  assign n5353 = ( n5348 & n5351 ) | ( n5348 & ~n5352 ) | ( n5351 & ~n5352 ) ;
  assign n5354 = ( ~n5244 & n5322 ) | ( ~n5244 & n5353 ) | ( n5322 & n5353 ) ;
  assign n5355 = ( n5244 & n5322 ) | ( n5244 & n5353 ) | ( n5322 & n5353 ) ;
  assign n5356 = ( n5244 & n5354 ) | ( n5244 & ~n5355 ) | ( n5354 & ~n5355 ) ;
  assign n5357 = ( ~n5246 & n5289 ) | ( ~n5246 & n5356 ) | ( n5289 & n5356 ) ;
  assign n5358 = ( n5246 & n5289 ) | ( n5246 & n5356 ) | ( n5289 & n5356 ) ;
  assign n5359 = ( n5246 & n5357 ) | ( n5246 & ~n5358 ) | ( n5357 & ~n5358 ) ;
  assign n5360 = ( n5307 & n5334 ) | ( n5307 & n5359 ) | ( n5334 & n5359 ) ;
  assign n5361 = ( ~n5307 & n5334 ) | ( ~n5307 & n5359 ) | ( n5334 & n5359 ) ;
  assign n5362 = ( n5307 & ~n5360 ) | ( n5307 & n5361 ) | ( ~n5360 & n5361 ) ;
  assign n5363 = ( n5275 & n5281 ) | ( n5275 & n5328 ) | ( n5281 & n5328 ) ;
  assign n5364 = ( ~n5275 & n5281 ) | ( ~n5275 & n5328 ) | ( n5281 & n5328 ) ;
  assign n5365 = ( n5275 & ~n5363 ) | ( n5275 & n5364 ) | ( ~n5363 & n5364 ) ;
  assign n5366 = ( n5295 & ~n5301 ) | ( n5295 & n5316 ) | ( ~n5301 & n5316 ) ;
  assign n5367 = ( n5295 & n5301 ) | ( n5295 & n5316 ) | ( n5301 & n5316 ) ;
  assign n5368 = ( n5301 & n5366 ) | ( n5301 & ~n5367 ) | ( n5366 & ~n5367 ) ;
  assign n5369 = ( n5331 & n5365 ) | ( n5331 & n5368 ) | ( n5365 & n5368 ) ;
  assign n5370 = ( n5331 & ~n5365 ) | ( n5331 & n5368 ) | ( ~n5365 & n5368 ) ;
  assign n5371 = ( n5365 & ~n5369 ) | ( n5365 & n5370 ) | ( ~n5369 & n5370 ) ;
  assign n5372 = x13 & x61 ;
  assign n5373 = x12 & x62 ;
  assign n5374 = ( n5286 & n5372 ) | ( n5286 & n5373 ) | ( n5372 & n5373 ) ;
  assign n5375 = ( ~n5286 & n5372 ) | ( ~n5286 & n5373 ) | ( n5372 & n5373 ) ;
  assign n5376 = ( n5286 & ~n5374 ) | ( n5286 & n5375 ) | ( ~n5374 & n5375 ) ;
  assign n5377 = x17 & x57 ;
  assign n5378 = x30 & x44 ;
  assign n5379 = x29 & x45 ;
  assign n5380 = ( ~n5377 & n5378 ) | ( ~n5377 & n5379 ) | ( n5378 & n5379 ) ;
  assign n5381 = ( n5377 & n5378 ) | ( n5377 & n5379 ) | ( n5378 & n5379 ) ;
  assign n5382 = ( n5377 & n5380 ) | ( n5377 & ~n5381 ) | ( n5380 & ~n5381 ) ;
  assign n5383 = ( ~n5310 & n5376 ) | ( ~n5310 & n5382 ) | ( n5376 & n5382 ) ;
  assign n5384 = ( n5310 & n5376 ) | ( n5310 & n5382 ) | ( n5376 & n5382 ) ;
  assign n5385 = ( n5310 & n5383 ) | ( n5310 & ~n5384 ) | ( n5383 & ~n5384 ) ;
  assign n5386 = x11 & x63 ;
  assign n5387 = x31 & x43 ;
  assign n5388 = x32 & x42 ;
  assign n5389 = ( ~n5386 & n5387 ) | ( ~n5386 & n5388 ) | ( n5387 & n5388 ) ;
  assign n5390 = ( n5386 & n5387 ) | ( n5386 & n5388 ) | ( n5387 & n5388 ) ;
  assign n5391 = ( n5386 & n5389 ) | ( n5386 & ~n5390 ) | ( n5389 & ~n5390 ) ;
  assign n5392 = x26 & x48 ;
  assign n5393 = x27 & x47 ;
  assign n5394 = x28 & x46 ;
  assign n5395 = ( ~n5392 & n5393 ) | ( ~n5392 & n5394 ) | ( n5393 & n5394 ) ;
  assign n5396 = ( n5392 & n5393 ) | ( n5392 & n5394 ) | ( n5393 & n5394 ) ;
  assign n5397 = ( n5392 & n5395 ) | ( n5392 & ~n5396 ) | ( n5395 & ~n5396 ) ;
  assign n5398 = x33 & x41 ;
  assign n5399 = x18 & x56 ;
  assign n5400 = x25 & x49 ;
  assign n5401 = ( ~n5398 & n5399 ) | ( ~n5398 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5402 = ( n5398 & n5399 ) | ( n5398 & n5400 ) | ( n5399 & n5400 ) ;
  assign n5403 = ( n5398 & n5401 ) | ( n5398 & ~n5402 ) | ( n5401 & ~n5402 ) ;
  assign n5404 = ( ~n5391 & n5397 ) | ( ~n5391 & n5403 ) | ( n5397 & n5403 ) ;
  assign n5405 = ( n5391 & n5397 ) | ( n5391 & n5403 ) | ( n5397 & n5403 ) ;
  assign n5406 = ( n5391 & n5404 ) | ( n5391 & ~n5405 ) | ( n5404 & ~n5405 ) ;
  assign n5407 = x20 & x54 ;
  assign n5408 = x34 & x40 ;
  assign n5409 = x35 & x39 ;
  assign n5410 = ( ~n5407 & n5408 ) | ( ~n5407 & n5409 ) | ( n5408 & n5409 ) ;
  assign n5411 = ( n5407 & n5408 ) | ( n5407 & n5409 ) | ( n5408 & n5409 ) ;
  assign n5412 = ( n5407 & n5410 ) | ( n5407 & ~n5411 ) | ( n5410 & ~n5411 ) ;
  assign n5413 = x36 & x38 ;
  assign n5414 = x23 & x51 ;
  assign n5415 = x24 & x50 ;
  assign n5416 = ( ~n5413 & n5414 ) | ( ~n5413 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5417 = ( n5413 & n5414 ) | ( n5413 & n5415 ) | ( n5414 & n5415 ) ;
  assign n5418 = ( n5413 & n5416 ) | ( n5413 & ~n5417 ) | ( n5416 & ~n5417 ) ;
  assign n5419 = x22 & x52 ;
  assign n5420 = x19 & x55 ;
  assign n5421 = x21 & x53 ;
  assign n5422 = ( ~n5419 & n5420 ) | ( ~n5419 & n5421 ) | ( n5420 & n5421 ) ;
  assign n5423 = ( n5419 & n5420 ) | ( n5419 & n5421 ) | ( n5420 & n5421 ) ;
  assign n5424 = ( n5419 & n5422 ) | ( n5419 & ~n5423 ) | ( n5422 & ~n5423 ) ;
  assign n5425 = ( ~n5412 & n5418 ) | ( ~n5412 & n5424 ) | ( n5418 & n5424 ) ;
  assign n5426 = ( n5412 & n5418 ) | ( n5412 & n5424 ) | ( n5418 & n5424 ) ;
  assign n5427 = ( n5412 & n5425 ) | ( n5412 & ~n5426 ) | ( n5425 & ~n5426 ) ;
  assign n5428 = ( n5385 & n5406 ) | ( n5385 & n5427 ) | ( n5406 & n5427 ) ;
  assign n5429 = ( ~n5385 & n5406 ) | ( ~n5385 & n5427 ) | ( n5406 & n5427 ) ;
  assign n5430 = ( n5385 & ~n5428 ) | ( n5385 & n5429 ) | ( ~n5428 & n5429 ) ;
  assign n5431 = ( ~n5249 & n5371 ) | ( ~n5249 & n5430 ) | ( n5371 & n5430 ) ;
  assign n5432 = ( n5249 & n5371 ) | ( n5249 & n5430 ) | ( n5371 & n5430 ) ;
  assign n5433 = ( n5249 & n5431 ) | ( n5249 & ~n5432 ) | ( n5431 & ~n5432 ) ;
  assign n5434 = ( n5252 & n5362 ) | ( n5252 & n5433 ) | ( n5362 & n5433 ) ;
  assign n5435 = ( ~n5252 & n5362 ) | ( ~n5252 & n5433 ) | ( n5362 & n5433 ) ;
  assign n5436 = ( n5252 & ~n5434 ) | ( n5252 & n5435 ) | ( ~n5434 & n5435 ) ;
  assign n5437 = ( ~n5259 & n5263 ) | ( ~n5259 & n5303 ) | ( n5263 & n5303 ) ;
  assign n5438 = ( n5259 & n5263 ) | ( n5259 & n5303 ) | ( n5263 & n5303 ) ;
  assign n5439 = ( n5259 & n5437 ) | ( n5259 & ~n5438 ) | ( n5437 & ~n5438 ) ;
  assign n5440 = ( n5256 & n5266 ) | ( n5256 & n5439 ) | ( n5266 & n5439 ) ;
  assign n5441 = ( n5256 & ~n5266 ) | ( n5256 & n5439 ) | ( ~n5266 & n5439 ) ;
  assign n5442 = ( n5266 & ~n5440 ) | ( n5266 & n5441 ) | ( ~n5440 & n5441 ) ;
  assign n5443 = ( n5269 & n5336 ) | ( n5269 & n5442 ) | ( n5336 & n5442 ) ;
  assign n5444 = ( ~n5269 & n5336 ) | ( ~n5269 & n5442 ) | ( n5336 & n5442 ) ;
  assign n5445 = ( n5269 & ~n5443 ) | ( n5269 & n5444 ) | ( ~n5443 & n5444 ) ;
  assign n5446 = ( ~n5340 & n5436 ) | ( ~n5340 & n5445 ) | ( n5436 & n5445 ) ;
  assign n5447 = ( n5340 & n5436 ) | ( n5340 & n5445 ) | ( n5436 & n5445 ) ;
  assign n5448 = ( n5340 & n5446 ) | ( n5340 & ~n5447 ) | ( n5446 & ~n5447 ) ;
  assign n5449 = ( n5343 & n5346 ) | ( n5343 & n5448 ) | ( n5346 & n5448 ) ;
  assign n5450 = ( ~n5343 & n5346 ) | ( ~n5343 & n5448 ) | ( n5346 & n5448 ) ;
  assign n5451 = ( n5343 & ~n5449 ) | ( n5343 & n5450 ) | ( ~n5449 & n5450 ) ;
  assign n5452 = ( n5411 & n5417 ) | ( n5411 & n5423 ) | ( n5417 & n5423 ) ;
  assign n5453 = ( ~n5411 & n5417 ) | ( ~n5411 & n5423 ) | ( n5417 & n5423 ) ;
  assign n5454 = ( n5411 & ~n5452 ) | ( n5411 & n5453 ) | ( ~n5452 & n5453 ) ;
  assign n5455 = ( ~n5374 & n5390 ) | ( ~n5374 & n5402 ) | ( n5390 & n5402 ) ;
  assign n5456 = ( n5374 & n5390 ) | ( n5374 & n5402 ) | ( n5390 & n5402 ) ;
  assign n5457 = ( n5374 & n5455 ) | ( n5374 & ~n5456 ) | ( n5455 & ~n5456 ) ;
  assign n5458 = ( ~n5384 & n5454 ) | ( ~n5384 & n5457 ) | ( n5454 & n5457 ) ;
  assign n5459 = ( n5384 & n5454 ) | ( n5384 & n5457 ) | ( n5454 & n5457 ) ;
  assign n5460 = ( n5384 & n5458 ) | ( n5384 & ~n5459 ) | ( n5458 & ~n5459 ) ;
  assign n5461 = ( n5355 & n5363 ) | ( n5355 & n5367 ) | ( n5363 & n5367 ) ;
  assign n5462 = ( n5355 & ~n5363 ) | ( n5355 & n5367 ) | ( ~n5363 & n5367 ) ;
  assign n5463 = ( n5363 & ~n5461 ) | ( n5363 & n5462 ) | ( ~n5461 & n5462 ) ;
  assign n5464 = ( ~n5428 & n5460 ) | ( ~n5428 & n5463 ) | ( n5460 & n5463 ) ;
  assign n5465 = ( n5428 & n5460 ) | ( n5428 & n5463 ) | ( n5460 & n5463 ) ;
  assign n5466 = ( n5428 & n5464 ) | ( n5428 & ~n5465 ) | ( n5464 & ~n5465 ) ;
  assign n5467 = ( n5352 & ~n5381 ) | ( n5352 & n5396 ) | ( ~n5381 & n5396 ) ;
  assign n5468 = ( n5352 & n5381 ) | ( n5352 & n5396 ) | ( n5381 & n5396 ) ;
  assign n5469 = ( n5381 & n5467 ) | ( n5381 & ~n5468 ) | ( n5467 & ~n5468 ) ;
  assign n5470 = ( n5405 & n5426 ) | ( n5405 & n5469 ) | ( n5426 & n5469 ) ;
  assign n5471 = ( ~n5405 & n5426 ) | ( ~n5405 & n5469 ) | ( n5426 & n5469 ) ;
  assign n5472 = ( n5405 & ~n5470 ) | ( n5405 & n5471 ) | ( ~n5470 & n5471 ) ;
  assign n5473 = x37 & x38 ;
  assign n5474 = x13 & x62 ;
  assign n5475 = ( x38 & n5473 ) | ( x38 & n5474 ) | ( n5473 & n5474 ) ;
  assign n5476 = ( x38 & ~n5473 ) | ( x38 & n5474 ) | ( ~n5473 & n5474 ) ;
  assign n5477 = ( n5473 & ~n5475 ) | ( n5473 & n5476 ) | ( ~n5475 & n5476 ) ;
  assign n5478 = x23 & x52 ;
  assign n5479 = x35 & x40 ;
  assign n5480 = x36 & x39 ;
  assign n5481 = ( ~n5478 & n5479 ) | ( ~n5478 & n5480 ) | ( n5479 & n5480 ) ;
  assign n5482 = ( n5478 & n5479 ) | ( n5478 & n5480 ) | ( n5479 & n5480 ) ;
  assign n5483 = ( n5478 & n5481 ) | ( n5478 & ~n5482 ) | ( n5481 & ~n5482 ) ;
  assign n5484 = x30 & x45 ;
  assign n5485 = x12 & x63 ;
  assign n5486 = x19 & x56 ;
  assign n5487 = ( ~n5484 & n5485 ) | ( ~n5484 & n5486 ) | ( n5485 & n5486 ) ;
  assign n5488 = ( n5484 & n5485 ) | ( n5484 & n5486 ) | ( n5485 & n5486 ) ;
  assign n5489 = ( n5484 & n5487 ) | ( n5484 & ~n5488 ) | ( n5487 & ~n5488 ) ;
  assign n5490 = ( n5477 & n5483 ) | ( n5477 & n5489 ) | ( n5483 & n5489 ) ;
  assign n5491 = ( ~n5477 & n5483 ) | ( ~n5477 & n5489 ) | ( n5483 & n5489 ) ;
  assign n5492 = ( n5477 & ~n5490 ) | ( n5477 & n5491 ) | ( ~n5490 & n5491 ) ;
  assign n5493 = x17 & x58 ;
  assign n5494 = x26 & x49 ;
  assign n5495 = x18 & x57 ;
  assign n5496 = ( ~n5493 & n5494 ) | ( ~n5493 & n5495 ) | ( n5494 & n5495 ) ;
  assign n5497 = ( n5493 & n5494 ) | ( n5493 & n5495 ) | ( n5494 & n5495 ) ;
  assign n5498 = ( n5493 & n5496 ) | ( n5493 & ~n5497 ) | ( n5496 & ~n5497 ) ;
  assign n5499 = x27 & x48 ;
  assign n5500 = x28 & x47 ;
  assign n5501 = x29 & x46 ;
  assign n5502 = ( ~n5499 & n5500 ) | ( ~n5499 & n5501 ) | ( n5500 & n5501 ) ;
  assign n5503 = ( n5499 & n5500 ) | ( n5499 & n5501 ) | ( n5500 & n5501 ) ;
  assign n5504 = ( n5499 & n5502 ) | ( n5499 & ~n5503 ) | ( n5502 & ~n5503 ) ;
  assign n5505 = x14 & x61 ;
  assign n5506 = x16 & x59 ;
  assign n5507 = x15 & x60 ;
  assign n5508 = ( ~n5505 & n5506 ) | ( ~n5505 & n5507 ) | ( n5506 & n5507 ) ;
  assign n5509 = ( n5505 & n5506 ) | ( n5505 & n5507 ) | ( n5506 & n5507 ) ;
  assign n5510 = ( n5505 & n5508 ) | ( n5505 & ~n5509 ) | ( n5508 & ~n5509 ) ;
  assign n5511 = ( ~n5498 & n5504 ) | ( ~n5498 & n5510 ) | ( n5504 & n5510 ) ;
  assign n5512 = ( n5498 & n5504 ) | ( n5498 & n5510 ) | ( n5504 & n5510 ) ;
  assign n5513 = ( n5498 & n5511 ) | ( n5498 & ~n5512 ) | ( n5511 & ~n5512 ) ;
  assign n5514 = ( n5438 & n5492 ) | ( n5438 & n5513 ) | ( n5492 & n5513 ) ;
  assign n5515 = ( ~n5438 & n5492 ) | ( ~n5438 & n5513 ) | ( n5492 & n5513 ) ;
  assign n5516 = ( n5438 & ~n5514 ) | ( n5438 & n5515 ) | ( ~n5514 & n5515 ) ;
  assign n5517 = ( ~n5440 & n5472 ) | ( ~n5440 & n5516 ) | ( n5472 & n5516 ) ;
  assign n5518 = ( n5440 & n5472 ) | ( n5440 & n5516 ) | ( n5472 & n5516 ) ;
  assign n5519 = ( n5440 & n5517 ) | ( n5440 & ~n5518 ) | ( n5517 & ~n5518 ) ;
  assign n5520 = ( ~n5443 & n5466 ) | ( ~n5443 & n5519 ) | ( n5466 & n5519 ) ;
  assign n5521 = ( n5443 & n5466 ) | ( n5443 & n5519 ) | ( n5466 & n5519 ) ;
  assign n5522 = ( n5443 & n5520 ) | ( n5443 & ~n5521 ) | ( n5520 & ~n5521 ) ;
  assign n5523 = x34 & x41 ;
  assign n5524 = x20 & x55 ;
  assign n5525 = x25 & x50 ;
  assign n5526 = ( ~n5523 & n5524 ) | ( ~n5523 & n5525 ) | ( n5524 & n5525 ) ;
  assign n5527 = ( n5523 & n5524 ) | ( n5523 & n5525 ) | ( n5524 & n5525 ) ;
  assign n5528 = ( n5523 & n5526 ) | ( n5523 & ~n5527 ) | ( n5526 & ~n5527 ) ;
  assign n5529 = x21 & x54 ;
  assign n5530 = x24 & x51 ;
  assign n5531 = x22 & x53 ;
  assign n5532 = ( ~n5529 & n5530 ) | ( ~n5529 & n5531 ) | ( n5530 & n5531 ) ;
  assign n5533 = ( n5529 & n5530 ) | ( n5529 & n5531 ) | ( n5530 & n5531 ) ;
  assign n5534 = ( n5529 & n5532 ) | ( n5529 & ~n5533 ) | ( n5532 & ~n5533 ) ;
  assign n5535 = x31 & x44 ;
  assign n5536 = x32 & x43 ;
  assign n5537 = x33 & x42 ;
  assign n5538 = ( ~n5535 & n5536 ) | ( ~n5535 & n5537 ) | ( n5536 & n5537 ) ;
  assign n5539 = ( n5535 & n5536 ) | ( n5535 & n5537 ) | ( n5536 & n5537 ) ;
  assign n5540 = ( n5535 & n5538 ) | ( n5535 & ~n5539 ) | ( n5538 & ~n5539 ) ;
  assign n5541 = ( ~n5528 & n5534 ) | ( ~n5528 & n5540 ) | ( n5534 & n5540 ) ;
  assign n5542 = ( n5528 & n5534 ) | ( n5528 & n5540 ) | ( n5534 & n5540 ) ;
  assign n5543 = ( n5528 & n5541 ) | ( n5528 & ~n5542 ) | ( n5541 & ~n5542 ) ;
  assign n5544 = ( n5358 & n5369 ) | ( n5358 & n5543 ) | ( n5369 & n5543 ) ;
  assign n5545 = ( ~n5358 & n5369 ) | ( ~n5358 & n5543 ) | ( n5369 & n5543 ) ;
  assign n5546 = ( n5358 & ~n5544 ) | ( n5358 & n5545 ) | ( ~n5544 & n5545 ) ;
  assign n5547 = ( n5360 & n5432 ) | ( n5360 & n5546 ) | ( n5432 & n5546 ) ;
  assign n5548 = ( ~n5360 & n5432 ) | ( ~n5360 & n5546 ) | ( n5432 & n5546 ) ;
  assign n5549 = ( n5360 & ~n5547 ) | ( n5360 & n5548 ) | ( ~n5547 & n5548 ) ;
  assign n5550 = ( ~n5434 & n5522 ) | ( ~n5434 & n5549 ) | ( n5522 & n5549 ) ;
  assign n5551 = ( n5434 & n5522 ) | ( n5434 & n5549 ) | ( n5522 & n5549 ) ;
  assign n5552 = ( n5434 & n5550 ) | ( n5434 & ~n5551 ) | ( n5550 & ~n5551 ) ;
  assign n5553 = ( ~n5447 & n5449 ) | ( ~n5447 & n5552 ) | ( n5449 & n5552 ) ;
  assign n5554 = ( n5447 & n5449 ) | ( n5447 & n5552 ) | ( n5449 & n5552 ) ;
  assign n5555 = ( n5447 & n5553 ) | ( n5447 & ~n5554 ) | ( n5553 & ~n5554 ) ;
  assign n5556 = x20 & x56 ;
  assign n5557 = x21 & x55 ;
  assign n5558 = x22 & x54 ;
  assign n5559 = ( ~n5556 & n5557 ) | ( ~n5556 & n5558 ) | ( n5557 & n5558 ) ;
  assign n5560 = ( n5556 & n5557 ) | ( n5556 & n5558 ) | ( n5557 & n5558 ) ;
  assign n5561 = ( n5556 & n5559 ) | ( n5556 & ~n5560 ) | ( n5559 & ~n5560 ) ;
  assign n5562 = x33 & x43 ;
  assign n5563 = x19 & x57 ;
  assign n5564 = x23 & x53 ;
  assign n5565 = ( ~n5562 & n5563 ) | ( ~n5562 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5566 = ( n5562 & n5563 ) | ( n5562 & n5564 ) | ( n5563 & n5564 ) ;
  assign n5567 = ( n5562 & n5565 ) | ( n5562 & ~n5566 ) | ( n5565 & ~n5566 ) ;
  assign n5568 = x13 & x63 ;
  assign n5569 = x31 & x45 ;
  assign n5570 = x32 & x44 ;
  assign n5571 = ( ~n5568 & n5569 ) | ( ~n5568 & n5570 ) | ( n5569 & n5570 ) ;
  assign n5572 = ( n5568 & n5569 ) | ( n5568 & n5570 ) | ( n5569 & n5570 ) ;
  assign n5573 = ( n5568 & n5571 ) | ( n5568 & ~n5572 ) | ( n5571 & ~n5572 ) ;
  assign n5574 = ( ~n5561 & n5567 ) | ( ~n5561 & n5573 ) | ( n5567 & n5573 ) ;
  assign n5575 = ( n5561 & n5567 ) | ( n5561 & n5573 ) | ( n5567 & n5573 ) ;
  assign n5576 = ( n5561 & n5574 ) | ( n5561 & ~n5575 ) | ( n5574 & ~n5575 ) ;
  assign n5577 = ( n5459 & n5470 ) | ( n5459 & n5576 ) | ( n5470 & n5576 ) ;
  assign n5578 = ( ~n5459 & n5470 ) | ( ~n5459 & n5576 ) | ( n5470 & n5576 ) ;
  assign n5579 = ( n5459 & ~n5577 ) | ( n5459 & n5578 ) | ( ~n5577 & n5578 ) ;
  assign n5580 = ( ~n5465 & n5518 ) | ( ~n5465 & n5579 ) | ( n5518 & n5579 ) ;
  assign n5581 = ( n5465 & n5518 ) | ( n5465 & n5579 ) | ( n5518 & n5579 ) ;
  assign n5582 = ( n5465 & n5580 ) | ( n5465 & ~n5581 ) | ( n5580 & ~n5581 ) ;
  assign n5583 = ( n5452 & n5456 ) | ( n5452 & n5468 ) | ( n5456 & n5468 ) ;
  assign n5584 = ( ~n5452 & n5456 ) | ( ~n5452 & n5468 ) | ( n5456 & n5468 ) ;
  assign n5585 = ( n5452 & ~n5583 ) | ( n5452 & n5584 ) | ( ~n5583 & n5584 ) ;
  assign n5586 = ( n5488 & ~n5503 ) | ( n5488 & n5527 ) | ( ~n5503 & n5527 ) ;
  assign n5587 = ( n5488 & n5503 ) | ( n5488 & n5527 ) | ( n5503 & n5527 ) ;
  assign n5588 = ( n5503 & n5586 ) | ( n5503 & ~n5587 ) | ( n5586 & ~n5587 ) ;
  assign n5589 = x14 & x62 ;
  assign n5590 = ( n5475 & n5482 ) | ( n5475 & n5589 ) | ( n5482 & n5589 ) ;
  assign n5591 = ( n5475 & ~n5482 ) | ( n5475 & n5589 ) | ( ~n5482 & n5589 ) ;
  assign n5592 = ( n5482 & ~n5590 ) | ( n5482 & n5591 ) | ( ~n5590 & n5591 ) ;
  assign n5593 = ( n5542 & n5588 ) | ( n5542 & n5592 ) | ( n5588 & n5592 ) ;
  assign n5594 = ( ~n5542 & n5588 ) | ( ~n5542 & n5592 ) | ( n5588 & n5592 ) ;
  assign n5595 = ( n5542 & ~n5593 ) | ( n5542 & n5594 ) | ( ~n5593 & n5594 ) ;
  assign n5596 = ( ~n5514 & n5585 ) | ( ~n5514 & n5595 ) | ( n5585 & n5595 ) ;
  assign n5597 = ( n5514 & n5585 ) | ( n5514 & n5595 ) | ( n5585 & n5595 ) ;
  assign n5598 = ( n5514 & n5596 ) | ( n5514 & ~n5597 ) | ( n5596 & ~n5597 ) ;
  assign n5599 = ( n5497 & ~n5509 ) | ( n5497 & n5539 ) | ( ~n5509 & n5539 ) ;
  assign n5600 = ( n5497 & n5509 ) | ( n5497 & n5539 ) | ( n5509 & n5539 ) ;
  assign n5601 = ( n5509 & n5599 ) | ( n5509 & ~n5600 ) | ( n5599 & ~n5600 ) ;
  assign n5602 = ( ~n5490 & n5512 ) | ( ~n5490 & n5601 ) | ( n5512 & n5601 ) ;
  assign n5603 = ( n5490 & n5512 ) | ( n5490 & n5601 ) | ( n5512 & n5601 ) ;
  assign n5604 = ( n5490 & n5602 ) | ( n5490 & ~n5603 ) | ( n5602 & ~n5603 ) ;
  assign n5605 = x34 & x42 ;
  assign n5606 = x36 & x40 ;
  assign n5607 = x35 & x41 ;
  assign n5608 = ( ~n5605 & n5606 ) | ( ~n5605 & n5607 ) | ( n5606 & n5607 ) ;
  assign n5609 = ( n5605 & n5606 ) | ( n5605 & n5607 ) | ( n5606 & n5607 ) ;
  assign n5610 = ( n5605 & n5608 ) | ( n5605 & ~n5609 ) | ( n5608 & ~n5609 ) ;
  assign n5611 = x37 & x39 ;
  assign n5612 = x25 & x51 ;
  assign n5613 = x24 & x52 ;
  assign n5614 = ( ~n5611 & n5612 ) | ( ~n5611 & n5613 ) | ( n5612 & n5613 ) ;
  assign n5615 = ( n5611 & n5612 ) | ( n5611 & n5613 ) | ( n5612 & n5613 ) ;
  assign n5616 = ( n5611 & n5614 ) | ( n5611 & ~n5615 ) | ( n5614 & ~n5615 ) ;
  assign n5617 = x28 & x48 ;
  assign n5618 = x29 & x47 ;
  assign n5619 = x30 & x46 ;
  assign n5620 = ( ~n5617 & n5618 ) | ( ~n5617 & n5619 ) | ( n5618 & n5619 ) ;
  assign n5621 = ( n5617 & n5618 ) | ( n5617 & n5619 ) | ( n5618 & n5619 ) ;
  assign n5622 = ( n5617 & n5620 ) | ( n5617 & ~n5621 ) | ( n5620 & ~n5621 ) ;
  assign n5623 = ( ~n5610 & n5616 ) | ( ~n5610 & n5622 ) | ( n5616 & n5622 ) ;
  assign n5624 = ( n5610 & n5616 ) | ( n5610 & n5622 ) | ( n5616 & n5622 ) ;
  assign n5625 = ( n5610 & n5623 ) | ( n5610 & ~n5624 ) | ( n5623 & ~n5624 ) ;
  assign n5626 = x18 & x58 ;
  assign n5627 = x26 & x50 ;
  assign n5628 = x27 & x49 ;
  assign n5629 = ( ~n5626 & n5627 ) | ( ~n5626 & n5628 ) | ( n5627 & n5628 ) ;
  assign n5630 = ( n5626 & n5627 ) | ( n5626 & n5628 ) | ( n5627 & n5628 ) ;
  assign n5631 = ( n5626 & n5629 ) | ( n5626 & ~n5630 ) | ( n5629 & ~n5630 ) ;
  assign n5632 = x15 & x61 ;
  assign n5633 = x16 & x60 ;
  assign n5634 = x17 & x59 ;
  assign n5635 = ( ~n5632 & n5633 ) | ( ~n5632 & n5634 ) | ( n5633 & n5634 ) ;
  assign n5636 = ( n5632 & n5633 ) | ( n5632 & n5634 ) | ( n5633 & n5634 ) ;
  assign n5637 = ( n5632 & n5635 ) | ( n5632 & ~n5636 ) | ( n5635 & ~n5636 ) ;
  assign n5638 = ( n5533 & n5631 ) | ( n5533 & n5637 ) | ( n5631 & n5637 ) ;
  assign n5639 = ( ~n5533 & n5631 ) | ( ~n5533 & n5637 ) | ( n5631 & n5637 ) ;
  assign n5640 = ( n5533 & ~n5638 ) | ( n5533 & n5639 ) | ( ~n5638 & n5639 ) ;
  assign n5641 = ( ~n5461 & n5625 ) | ( ~n5461 & n5640 ) | ( n5625 & n5640 ) ;
  assign n5642 = ( n5461 & n5625 ) | ( n5461 & n5640 ) | ( n5625 & n5640 ) ;
  assign n5643 = ( n5461 & n5641 ) | ( n5461 & ~n5642 ) | ( n5641 & ~n5642 ) ;
  assign n5644 = ( ~n5544 & n5604 ) | ( ~n5544 & n5643 ) | ( n5604 & n5643 ) ;
  assign n5645 = ( n5544 & n5604 ) | ( n5544 & n5643 ) | ( n5604 & n5643 ) ;
  assign n5646 = ( n5544 & n5644 ) | ( n5544 & ~n5645 ) | ( n5644 & ~n5645 ) ;
  assign n5647 = ( n5547 & n5598 ) | ( n5547 & n5646 ) | ( n5598 & n5646 ) ;
  assign n5648 = ( ~n5547 & n5598 ) | ( ~n5547 & n5646 ) | ( n5598 & n5646 ) ;
  assign n5649 = ( n5547 & ~n5647 ) | ( n5547 & n5648 ) | ( ~n5647 & n5648 ) ;
  assign n5650 = ( ~n5521 & n5582 ) | ( ~n5521 & n5649 ) | ( n5582 & n5649 ) ;
  assign n5651 = ( n5521 & n5582 ) | ( n5521 & n5649 ) | ( n5582 & n5649 ) ;
  assign n5652 = ( n5521 & n5650 ) | ( n5521 & ~n5651 ) | ( n5650 & ~n5651 ) ;
  assign n5653 = ( n5551 & n5554 ) | ( n5551 & n5652 ) | ( n5554 & n5652 ) ;
  assign n5654 = ( ~n5551 & n5554 ) | ( ~n5551 & n5652 ) | ( n5554 & n5652 ) ;
  assign n5655 = ( n5551 & ~n5653 ) | ( n5551 & n5654 ) | ( ~n5653 & n5654 ) ;
  assign n5656 = x22 & x55 ;
  assign n5657 = x34 & x43 ;
  assign n5658 = x26 & x51 ;
  assign n5659 = ( ~n5656 & n5657 ) | ( ~n5656 & n5658 ) | ( n5657 & n5658 ) ;
  assign n5660 = ( n5656 & n5657 ) | ( n5656 & n5658 ) | ( n5657 & n5658 ) ;
  assign n5661 = ( n5656 & n5659 ) | ( n5656 & ~n5660 ) | ( n5659 & ~n5660 ) ;
  assign n5662 = x16 & x61 ;
  assign n5663 = x32 & x45 ;
  assign n5664 = x33 & x44 ;
  assign n5665 = ( ~n5662 & n5663 ) | ( ~n5662 & n5664 ) | ( n5663 & n5664 ) ;
  assign n5666 = ( n5662 & n5663 ) | ( n5662 & n5664 ) | ( n5663 & n5664 ) ;
  assign n5667 = ( n5662 & n5665 ) | ( n5662 & ~n5666 ) | ( n5665 & ~n5666 ) ;
  assign n5668 = x25 & x52 ;
  assign n5669 = x24 & x53 ;
  assign n5670 = x23 & x54 ;
  assign n5671 = ( ~n5668 & n5669 ) | ( ~n5668 & n5670 ) | ( n5669 & n5670 ) ;
  assign n5672 = ( n5668 & n5669 ) | ( n5668 & n5670 ) | ( n5669 & n5670 ) ;
  assign n5673 = ( n5668 & n5671 ) | ( n5668 & ~n5672 ) | ( n5671 & ~n5672 ) ;
  assign n5674 = ( ~n5661 & n5667 ) | ( ~n5661 & n5673 ) | ( n5667 & n5673 ) ;
  assign n5675 = ( n5661 & n5667 ) | ( n5661 & n5673 ) | ( n5667 & n5673 ) ;
  assign n5676 = ( n5661 & n5674 ) | ( n5661 & ~n5675 ) | ( n5674 & ~n5675 ) ;
  assign n5677 = ( ~n5593 & n5603 ) | ( ~n5593 & n5676 ) | ( n5603 & n5676 ) ;
  assign n5678 = ( n5593 & n5603 ) | ( n5593 & n5676 ) | ( n5603 & n5676 ) ;
  assign n5679 = ( n5593 & n5677 ) | ( n5593 & ~n5678 ) | ( n5677 & ~n5678 ) ;
  assign n5680 = ( n5597 & n5645 ) | ( n5597 & n5679 ) | ( n5645 & n5679 ) ;
  assign n5681 = ( ~n5597 & n5645 ) | ( ~n5597 & n5679 ) | ( n5645 & n5679 ) ;
  assign n5682 = ( n5597 & ~n5680 ) | ( n5597 & n5681 ) | ( ~n5680 & n5681 ) ;
  assign n5683 = x17 & x60 ;
  assign n5684 = x18 & x59 ;
  assign n5685 = ( n5615 & n5683 ) | ( n5615 & n5684 ) | ( n5683 & n5684 ) ;
  assign n5686 = ( ~n5615 & n5683 ) | ( ~n5615 & n5684 ) | ( n5683 & n5684 ) ;
  assign n5687 = ( n5615 & ~n5685 ) | ( n5615 & n5686 ) | ( ~n5685 & n5686 ) ;
  assign n5688 = ( n5587 & n5600 ) | ( n5587 & n5687 ) | ( n5600 & n5687 ) ;
  assign n5689 = ( ~n5587 & n5600 ) | ( ~n5587 & n5687 ) | ( n5600 & n5687 ) ;
  assign n5690 = ( n5587 & ~n5688 ) | ( n5587 & n5689 ) | ( ~n5688 & n5689 ) ;
  assign n5691 = ( n5560 & ~n5572 ) | ( n5560 & n5621 ) | ( ~n5572 & n5621 ) ;
  assign n5692 = ( n5560 & n5572 ) | ( n5560 & n5621 ) | ( n5572 & n5621 ) ;
  assign n5693 = ( n5572 & n5691 ) | ( n5572 & ~n5692 ) | ( n5691 & ~n5692 ) ;
  assign n5694 = ( n5566 & ~n5630 ) | ( n5566 & n5636 ) | ( ~n5630 & n5636 ) ;
  assign n5695 = ( n5566 & n5630 ) | ( n5566 & n5636 ) | ( n5630 & n5636 ) ;
  assign n5696 = ( n5630 & n5694 ) | ( n5630 & ~n5695 ) | ( n5694 & ~n5695 ) ;
  assign n5697 = ( ~n5575 & n5693 ) | ( ~n5575 & n5696 ) | ( n5693 & n5696 ) ;
  assign n5698 = ( n5575 & n5693 ) | ( n5575 & n5696 ) | ( n5693 & n5696 ) ;
  assign n5699 = ( n5575 & n5697 ) | ( n5575 & ~n5698 ) | ( n5697 & ~n5698 ) ;
  assign n5700 = ( ~n5642 & n5690 ) | ( ~n5642 & n5699 ) | ( n5690 & n5699 ) ;
  assign n5701 = ( n5642 & n5690 ) | ( n5642 & n5699 ) | ( n5690 & n5699 ) ;
  assign n5702 = ( n5642 & n5700 ) | ( n5642 & ~n5701 ) | ( n5700 & ~n5701 ) ;
  assign n5703 = ( ~n5590 & n5624 ) | ( ~n5590 & n5638 ) | ( n5624 & n5638 ) ;
  assign n5704 = ( n5590 & n5624 ) | ( n5590 & n5638 ) | ( n5624 & n5638 ) ;
  assign n5705 = ( n5590 & n5703 ) | ( n5590 & ~n5704 ) | ( n5703 & ~n5704 ) ;
  assign n5706 = x38 & x39 ;
  assign n5707 = x15 & x62 ;
  assign n5708 = ( x39 & n5706 ) | ( x39 & n5707 ) | ( n5706 & n5707 ) ;
  assign n5709 = ( x39 & ~n5706 ) | ( x39 & n5707 ) | ( ~n5706 & n5707 ) ;
  assign n5710 = ( n5706 & ~n5708 ) | ( n5706 & n5709 ) | ( ~n5708 & n5709 ) ;
  assign n5711 = x35 & x42 ;
  assign n5712 = x36 & x41 ;
  assign n5713 = x37 & x40 ;
  assign n5714 = ( ~n5711 & n5712 ) | ( ~n5711 & n5713 ) | ( n5712 & n5713 ) ;
  assign n5715 = ( n5711 & n5712 ) | ( n5711 & n5713 ) | ( n5712 & n5713 ) ;
  assign n5716 = ( n5711 & n5714 ) | ( n5711 & ~n5715 ) | ( n5714 & ~n5715 ) ;
  assign n5717 = x30 & x47 ;
  assign n5718 = x14 & x63 ;
  assign n5719 = x31 & x46 ;
  assign n5720 = ( ~n5717 & n5718 ) | ( ~n5717 & n5719 ) | ( n5718 & n5719 ) ;
  assign n5721 = ( n5717 & n5718 ) | ( n5717 & n5719 ) | ( n5718 & n5719 ) ;
  assign n5722 = ( n5717 & n5720 ) | ( n5717 & ~n5721 ) | ( n5720 & ~n5721 ) ;
  assign n5723 = ( n5710 & n5716 ) | ( n5710 & n5722 ) | ( n5716 & n5722 ) ;
  assign n5724 = ( ~n5710 & n5716 ) | ( ~n5710 & n5722 ) | ( n5716 & n5722 ) ;
  assign n5725 = ( n5710 & ~n5723 ) | ( n5710 & n5724 ) | ( ~n5723 & n5724 ) ;
  assign n5726 = x27 & x50 ;
  assign n5727 = x28 & x49 ;
  assign n5728 = x29 & x48 ;
  assign n5729 = ( ~n5726 & n5727 ) | ( ~n5726 & n5728 ) | ( n5727 & n5728 ) ;
  assign n5730 = ( n5726 & n5727 ) | ( n5726 & n5728 ) | ( n5727 & n5728 ) ;
  assign n5731 = ( n5726 & n5729 ) | ( n5726 & ~n5730 ) | ( n5729 & ~n5730 ) ;
  assign n5732 = x19 & x58 ;
  assign n5733 = x20 & x57 ;
  assign n5734 = x21 & x56 ;
  assign n5735 = ( ~n5732 & n5733 ) | ( ~n5732 & n5734 ) | ( n5733 & n5734 ) ;
  assign n5736 = ( n5732 & n5733 ) | ( n5732 & n5734 ) | ( n5733 & n5734 ) ;
  assign n5737 = ( n5732 & n5735 ) | ( n5732 & ~n5736 ) | ( n5735 & ~n5736 ) ;
  assign n5738 = ( n5609 & n5731 ) | ( n5609 & n5737 ) | ( n5731 & n5737 ) ;
  assign n5739 = ( ~n5609 & n5731 ) | ( ~n5609 & n5737 ) | ( n5731 & n5737 ) ;
  assign n5740 = ( n5609 & ~n5738 ) | ( n5609 & n5739 ) | ( ~n5738 & n5739 ) ;
  assign n5741 = ( ~n5583 & n5725 ) | ( ~n5583 & n5740 ) | ( n5725 & n5740 ) ;
  assign n5742 = ( n5583 & n5725 ) | ( n5583 & n5740 ) | ( n5725 & n5740 ) ;
  assign n5743 = ( n5583 & n5741 ) | ( n5583 & ~n5742 ) | ( n5741 & ~n5742 ) ;
  assign n5744 = ( ~n5577 & n5705 ) | ( ~n5577 & n5743 ) | ( n5705 & n5743 ) ;
  assign n5745 = ( n5577 & n5705 ) | ( n5577 & n5743 ) | ( n5705 & n5743 ) ;
  assign n5746 = ( n5577 & n5744 ) | ( n5577 & ~n5745 ) | ( n5744 & ~n5745 ) ;
  assign n5747 = ( ~n5581 & n5702 ) | ( ~n5581 & n5746 ) | ( n5702 & n5746 ) ;
  assign n5748 = ( n5581 & n5702 ) | ( n5581 & n5746 ) | ( n5702 & n5746 ) ;
  assign n5749 = ( n5581 & n5747 ) | ( n5581 & ~n5748 ) | ( n5747 & ~n5748 ) ;
  assign n5750 = ( ~n5647 & n5682 ) | ( ~n5647 & n5749 ) | ( n5682 & n5749 ) ;
  assign n5751 = ( n5647 & n5682 ) | ( n5647 & n5749 ) | ( n5682 & n5749 ) ;
  assign n5752 = ( n5647 & n5750 ) | ( n5647 & ~n5751 ) | ( n5750 & ~n5751 ) ;
  assign n5753 = ( n5651 & n5653 ) | ( n5651 & n5752 ) | ( n5653 & n5752 ) ;
  assign n5754 = ( ~n5651 & n5653 ) | ( ~n5651 & n5752 ) | ( n5653 & n5752 ) ;
  assign n5755 = ( n5651 & ~n5753 ) | ( n5651 & n5754 ) | ( ~n5753 & n5754 ) ;
  assign n5756 = ( n5675 & n5723 ) | ( n5675 & ~n5738 ) | ( n5723 & ~n5738 ) ;
  assign n5757 = ( n5675 & n5723 ) | ( n5675 & n5738 ) | ( n5723 & n5738 ) ;
  assign n5758 = ( n5738 & n5756 ) | ( n5738 & ~n5757 ) | ( n5756 & ~n5757 ) ;
  assign n5759 = ( ~n5672 & n5708 ) | ( ~n5672 & n5715 ) | ( n5708 & n5715 ) ;
  assign n5760 = ( n5672 & n5708 ) | ( n5672 & n5715 ) | ( n5708 & n5715 ) ;
  assign n5761 = ( n5672 & n5759 ) | ( n5672 & ~n5760 ) | ( n5759 & ~n5760 ) ;
  assign n5762 = ( n5666 & ~n5721 ) | ( n5666 & n5730 ) | ( ~n5721 & n5730 ) ;
  assign n5763 = ( n5666 & n5721 ) | ( n5666 & n5730 ) | ( n5721 & n5730 ) ;
  assign n5764 = ( n5721 & n5762 ) | ( n5721 & ~n5763 ) | ( n5762 & ~n5763 ) ;
  assign n5765 = ( ~n5695 & n5761 ) | ( ~n5695 & n5764 ) | ( n5761 & n5764 ) ;
  assign n5766 = ( n5695 & n5761 ) | ( n5695 & n5764 ) | ( n5761 & n5764 ) ;
  assign n5767 = ( n5695 & n5765 ) | ( n5695 & ~n5766 ) | ( n5765 & ~n5766 ) ;
  assign n5768 = ( ~n5698 & n5758 ) | ( ~n5698 & n5767 ) | ( n5758 & n5767 ) ;
  assign n5769 = ( n5698 & n5758 ) | ( n5698 & n5767 ) | ( n5758 & n5767 ) ;
  assign n5770 = ( n5698 & n5768 ) | ( n5698 & ~n5769 ) | ( n5768 & ~n5769 ) ;
  assign n5771 = x37 & x41 ;
  assign n5772 = x38 & x40 ;
  assign n5773 = x26 & x52 ;
  assign n5774 = ( ~n5771 & n5772 ) | ( ~n5771 & n5773 ) | ( n5772 & n5773 ) ;
  assign n5775 = ( n5771 & n5772 ) | ( n5771 & n5773 ) | ( n5772 & n5773 ) ;
  assign n5776 = ( n5771 & n5774 ) | ( n5771 & ~n5775 ) | ( n5774 & ~n5775 ) ;
  assign n5777 = x23 & x55 ;
  assign n5778 = x35 & x43 ;
  assign n5779 = x36 & x42 ;
  assign n5780 = ( ~n5777 & n5778 ) | ( ~n5777 & n5779 ) | ( n5778 & n5779 ) ;
  assign n5781 = ( n5777 & n5778 ) | ( n5777 & n5779 ) | ( n5778 & n5779 ) ;
  assign n5782 = ( n5777 & n5780 ) | ( n5777 & ~n5781 ) | ( n5780 & ~n5781 ) ;
  assign n5783 = ( n5692 & n5776 ) | ( n5692 & n5782 ) | ( n5776 & n5782 ) ;
  assign n5784 = ( ~n5692 & n5776 ) | ( ~n5692 & n5782 ) | ( n5776 & n5782 ) ;
  assign n5785 = ( n5692 & ~n5783 ) | ( n5692 & n5784 ) | ( ~n5783 & n5784 ) ;
  assign n5786 = ( n5660 & ~n5685 ) | ( n5660 & n5736 ) | ( ~n5685 & n5736 ) ;
  assign n5787 = ( n5660 & n5685 ) | ( n5660 & n5736 ) | ( n5685 & n5736 ) ;
  assign n5788 = ( n5685 & n5786 ) | ( n5685 & ~n5787 ) | ( n5786 & ~n5787 ) ;
  assign n5789 = ( ~n5688 & n5785 ) | ( ~n5688 & n5788 ) | ( n5785 & n5788 ) ;
  assign n5790 = ( n5688 & n5785 ) | ( n5688 & n5788 ) | ( n5785 & n5788 ) ;
  assign n5791 = ( n5688 & n5789 ) | ( n5688 & ~n5790 ) | ( n5789 & ~n5790 ) ;
  assign n5792 = ( n5678 & n5742 ) | ( n5678 & n5791 ) | ( n5742 & n5791 ) ;
  assign n5793 = ( ~n5678 & n5742 ) | ( ~n5678 & n5791 ) | ( n5742 & n5791 ) ;
  assign n5794 = ( n5678 & ~n5792 ) | ( n5678 & n5793 ) | ( ~n5792 & n5793 ) ;
  assign n5795 = ( ~n5680 & n5770 ) | ( ~n5680 & n5794 ) | ( n5770 & n5794 ) ;
  assign n5796 = ( n5680 & n5770 ) | ( n5680 & n5794 ) | ( n5770 & n5794 ) ;
  assign n5797 = ( n5680 & n5795 ) | ( n5680 & ~n5796 ) | ( n5795 & ~n5796 ) ;
  assign n5798 = x15 & x63 ;
  assign n5799 = x16 & x62 ;
  assign n5800 = x17 & x61 ;
  assign n5801 = ( ~n5798 & n5799 ) | ( ~n5798 & n5800 ) | ( n5799 & n5800 ) ;
  assign n5802 = ( n5798 & n5799 ) | ( n5798 & n5800 ) | ( n5799 & n5800 ) ;
  assign n5803 = ( n5798 & n5801 ) | ( n5798 & ~n5802 ) | ( n5801 & ~n5802 ) ;
  assign n5804 = x27 & x51 ;
  assign n5805 = x29 & x49 ;
  assign n5806 = x28 & x50 ;
  assign n5807 = ( ~n5804 & n5805 ) | ( ~n5804 & n5806 ) | ( n5805 & n5806 ) ;
  assign n5808 = ( n5804 & n5805 ) | ( n5804 & n5806 ) | ( n5805 & n5806 ) ;
  assign n5809 = ( n5804 & n5807 ) | ( n5804 & ~n5808 ) | ( n5807 & ~n5808 ) ;
  assign n5810 = x18 & x60 ;
  assign n5811 = x21 & x57 ;
  assign n5812 = x19 & x59 ;
  assign n5813 = ( ~n5810 & n5811 ) | ( ~n5810 & n5812 ) | ( n5811 & n5812 ) ;
  assign n5814 = ( n5810 & n5811 ) | ( n5810 & n5812 ) | ( n5811 & n5812 ) ;
  assign n5815 = ( n5810 & n5813 ) | ( n5810 & ~n5814 ) | ( n5813 & ~n5814 ) ;
  assign n5816 = ( ~n5803 & n5809 ) | ( ~n5803 & n5815 ) | ( n5809 & n5815 ) ;
  assign n5817 = ( n5803 & n5809 ) | ( n5803 & n5815 ) | ( n5809 & n5815 ) ;
  assign n5818 = ( n5803 & n5816 ) | ( n5803 & ~n5817 ) | ( n5816 & ~n5817 ) ;
  assign n5819 = x20 & x58 ;
  assign n5820 = x30 & x48 ;
  assign n5821 = x31 & x47 ;
  assign n5822 = ( ~n5819 & n5820 ) | ( ~n5819 & n5821 ) | ( n5820 & n5821 ) ;
  assign n5823 = ( n5819 & n5820 ) | ( n5819 & n5821 ) | ( n5820 & n5821 ) ;
  assign n5824 = ( n5819 & n5822 ) | ( n5819 & ~n5823 ) | ( n5822 & ~n5823 ) ;
  assign n5825 = x25 & x53 ;
  assign n5826 = x24 & x54 ;
  assign n5827 = x22 & x56 ;
  assign n5828 = ( ~n5825 & n5826 ) | ( ~n5825 & n5827 ) | ( n5826 & n5827 ) ;
  assign n5829 = ( n5825 & n5826 ) | ( n5825 & n5827 ) | ( n5826 & n5827 ) ;
  assign n5830 = ( n5825 & n5828 ) | ( n5825 & ~n5829 ) | ( n5828 & ~n5829 ) ;
  assign n5831 = x32 & x46 ;
  assign n5832 = x33 & x45 ;
  assign n5833 = x34 & x44 ;
  assign n5834 = ( ~n5831 & n5832 ) | ( ~n5831 & n5833 ) | ( n5832 & n5833 ) ;
  assign n5835 = ( n5831 & n5832 ) | ( n5831 & n5833 ) | ( n5832 & n5833 ) ;
  assign n5836 = ( n5831 & n5834 ) | ( n5831 & ~n5835 ) | ( n5834 & ~n5835 ) ;
  assign n5837 = ( ~n5824 & n5830 ) | ( ~n5824 & n5836 ) | ( n5830 & n5836 ) ;
  assign n5838 = ( n5824 & n5830 ) | ( n5824 & n5836 ) | ( n5830 & n5836 ) ;
  assign n5839 = ( n5824 & n5837 ) | ( n5824 & ~n5838 ) | ( n5837 & ~n5838 ) ;
  assign n5840 = ( n5704 & n5818 ) | ( n5704 & n5839 ) | ( n5818 & n5839 ) ;
  assign n5841 = ( ~n5704 & n5818 ) | ( ~n5704 & n5839 ) | ( n5818 & n5839 ) ;
  assign n5842 = ( n5704 & ~n5840 ) | ( n5704 & n5841 ) | ( ~n5840 & n5841 ) ;
  assign n5843 = ( n5701 & n5745 ) | ( n5701 & n5842 ) | ( n5745 & n5842 ) ;
  assign n5844 = ( ~n5701 & n5745 ) | ( ~n5701 & n5842 ) | ( n5745 & n5842 ) ;
  assign n5845 = ( n5701 & ~n5843 ) | ( n5701 & n5844 ) | ( ~n5843 & n5844 ) ;
  assign n5846 = ( n5748 & n5797 ) | ( n5748 & n5845 ) | ( n5797 & n5845 ) ;
  assign n5847 = ( ~n5748 & n5797 ) | ( ~n5748 & n5845 ) | ( n5797 & n5845 ) ;
  assign n5848 = ( n5748 & ~n5846 ) | ( n5748 & n5847 ) | ( ~n5846 & n5847 ) ;
  assign n5849 = ( n5751 & n5753 ) | ( n5751 & n5848 ) | ( n5753 & n5848 ) ;
  assign n5850 = ( n5751 & ~n5753 ) | ( n5751 & n5848 ) | ( ~n5753 & n5848 ) ;
  assign n5851 = ( n5753 & ~n5849 ) | ( n5753 & n5850 ) | ( ~n5849 & n5850 ) ;
  assign n5852 = x36 & x43 ;
  assign n5853 = x23 & x56 ;
  assign n5854 = ( ~n2905 & n5852 ) | ( ~n2905 & n5853 ) | ( n5852 & n5853 ) ;
  assign n5855 = ( n2905 & n5852 ) | ( n2905 & n5853 ) | ( n5852 & n5853 ) ;
  assign n5856 = ( n2905 & n5854 ) | ( n2905 & ~n5855 ) | ( n5854 & ~n5855 ) ;
  assign n5857 = x16 & x63 ;
  assign n5858 = x34 & x45 ;
  assign n5859 = x35 & x44 ;
  assign n5860 = ( ~n5857 & n5858 ) | ( ~n5857 & n5859 ) | ( n5858 & n5859 ) ;
  assign n5861 = ( n5857 & n5858 ) | ( n5857 & n5859 ) | ( n5858 & n5859 ) ;
  assign n5862 = ( n5857 & n5860 ) | ( n5857 & ~n5861 ) | ( n5860 & ~n5861 ) ;
  assign n5863 = ( n5787 & n5856 ) | ( n5787 & n5862 ) | ( n5856 & n5862 ) ;
  assign n5864 = ( ~n5787 & n5856 ) | ( ~n5787 & n5862 ) | ( n5856 & n5862 ) ;
  assign n5865 = ( n5787 & ~n5863 ) | ( n5787 & n5864 ) | ( ~n5863 & n5864 ) ;
  assign n5866 = ( n5808 & ~n5814 ) | ( n5808 & n5829 ) | ( ~n5814 & n5829 ) ;
  assign n5867 = ( n5808 & n5814 ) | ( n5808 & n5829 ) | ( n5814 & n5829 ) ;
  assign n5868 = ( n5814 & n5866 ) | ( n5814 & ~n5867 ) | ( n5866 & ~n5867 ) ;
  assign n5869 = ( n5783 & n5865 ) | ( n5783 & n5868 ) | ( n5865 & n5868 ) ;
  assign n5870 = ( n5783 & ~n5865 ) | ( n5783 & n5868 ) | ( ~n5865 & n5868 ) ;
  assign n5871 = ( n5865 & ~n5869 ) | ( n5865 & n5870 ) | ( ~n5869 & n5870 ) ;
  assign n5872 = ( n5802 & n5823 ) | ( n5802 & n5835 ) | ( n5823 & n5835 ) ;
  assign n5873 = ( n5802 & ~n5823 ) | ( n5802 & n5835 ) | ( ~n5823 & n5835 ) ;
  assign n5874 = ( n5823 & ~n5872 ) | ( n5823 & n5873 ) | ( ~n5872 & n5873 ) ;
  assign n5875 = x18 & x61 ;
  assign n5876 = ( ~n5775 & n5781 ) | ( ~n5775 & n5875 ) | ( n5781 & n5875 ) ;
  assign n5877 = ( n5775 & n5781 ) | ( n5775 & n5875 ) | ( n5781 & n5875 ) ;
  assign n5878 = ( n5775 & n5876 ) | ( n5775 & ~n5877 ) | ( n5876 & ~n5877 ) ;
  assign n5879 = ( ~n5838 & n5874 ) | ( ~n5838 & n5878 ) | ( n5874 & n5878 ) ;
  assign n5880 = ( n5838 & n5874 ) | ( n5838 & n5878 ) | ( n5874 & n5878 ) ;
  assign n5881 = ( n5838 & n5879 ) | ( n5838 & ~n5880 ) | ( n5879 & ~n5880 ) ;
  assign n5882 = ( n5840 & n5871 ) | ( n5840 & n5881 ) | ( n5871 & n5881 ) ;
  assign n5883 = ( ~n5840 & n5871 ) | ( ~n5840 & n5881 ) | ( n5871 & n5881 ) ;
  assign n5884 = ( n5840 & ~n5882 ) | ( n5840 & n5883 ) | ( ~n5882 & n5883 ) ;
  assign n5885 = ( n5792 & n5843 ) | ( n5792 & n5884 ) | ( n5843 & n5884 ) ;
  assign n5886 = ( ~n5792 & n5843 ) | ( ~n5792 & n5884 ) | ( n5843 & n5884 ) ;
  assign n5887 = ( n5792 & ~n5885 ) | ( n5792 & n5886 ) | ( ~n5885 & n5886 ) ;
  assign n5888 = ( n5760 & n5763 ) | ( n5760 & n5817 ) | ( n5763 & n5817 ) ;
  assign n5889 = ( ~n5760 & n5763 ) | ( ~n5760 & n5817 ) | ( n5763 & n5817 ) ;
  assign n5890 = ( n5760 & ~n5888 ) | ( n5760 & n5889 ) | ( ~n5888 & n5889 ) ;
  assign n5891 = ( n5757 & n5790 ) | ( n5757 & n5890 ) | ( n5790 & n5890 ) ;
  assign n5892 = ( n5757 & ~n5790 ) | ( n5757 & n5890 ) | ( ~n5790 & n5890 ) ;
  assign n5893 = ( n5790 & ~n5891 ) | ( n5790 & n5892 ) | ( ~n5891 & n5892 ) ;
  assign n5894 = x31 & x48 ;
  assign n5895 = x33 & x46 ;
  assign n5896 = x32 & x47 ;
  assign n5897 = ( ~n5894 & n5895 ) | ( ~n5894 & n5896 ) | ( n5895 & n5896 ) ;
  assign n5898 = ( n5894 & n5895 ) | ( n5894 & n5896 ) | ( n5895 & n5896 ) ;
  assign n5899 = ( n5894 & n5897 ) | ( n5894 & ~n5898 ) | ( n5897 & ~n5898 ) ;
  assign n5900 = x22 & x57 ;
  assign n5901 = x29 & x50 ;
  assign n5902 = x30 & x49 ;
  assign n5903 = ( ~n5900 & n5901 ) | ( ~n5900 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5904 = ( n5900 & n5901 ) | ( n5900 & n5902 ) | ( n5901 & n5902 ) ;
  assign n5905 = ( n5900 & n5903 ) | ( n5900 & ~n5904 ) | ( n5903 & ~n5904 ) ;
  assign n5906 = x19 & x60 ;
  assign n5907 = x20 & x59 ;
  assign n5908 = x21 & x58 ;
  assign n5909 = ( ~n5906 & n5907 ) | ( ~n5906 & n5908 ) | ( n5907 & n5908 ) ;
  assign n5910 = ( n5906 & n5907 ) | ( n5906 & n5908 ) | ( n5907 & n5908 ) ;
  assign n5911 = ( n5906 & n5909 ) | ( n5906 & ~n5910 ) | ( n5909 & ~n5910 ) ;
  assign n5912 = ( ~n5899 & n5905 ) | ( ~n5899 & n5911 ) | ( n5905 & n5911 ) ;
  assign n5913 = ( n5899 & n5905 ) | ( n5899 & n5911 ) | ( n5905 & n5911 ) ;
  assign n5914 = ( n5899 & n5912 ) | ( n5899 & ~n5913 ) | ( n5912 & ~n5913 ) ;
  assign n5915 = x24 & x55 ;
  assign n5916 = x26 & x53 ;
  assign n5917 = x25 & x54 ;
  assign n5918 = ( ~n5915 & n5916 ) | ( ~n5915 & n5917 ) | ( n5916 & n5917 ) ;
  assign n5919 = ( n5915 & n5916 ) | ( n5915 & n5917 ) | ( n5916 & n5917 ) ;
  assign n5920 = ( n5915 & n5918 ) | ( n5915 & ~n5919 ) | ( n5918 & ~n5919 ) ;
  assign n5921 = x37 & x42 ;
  assign n5922 = x39 & x40 ;
  assign n5923 = x38 & x41 ;
  assign n5924 = ( ~n5921 & n5922 ) | ( ~n5921 & n5923 ) | ( n5922 & n5923 ) ;
  assign n5925 = ( n5921 & n5922 ) | ( n5921 & n5923 ) | ( n5922 & n5923 ) ;
  assign n5926 = ( n5921 & n5924 ) | ( n5921 & ~n5925 ) | ( n5924 & ~n5925 ) ;
  assign n5927 = x28 & x51 ;
  assign n5928 = x17 & x62 ;
  assign n5929 = ( ~x40 & n5927 ) | ( ~x40 & n5928 ) | ( n5927 & n5928 ) ;
  assign n5930 = ( x40 & n5927 ) | ( x40 & n5928 ) | ( n5927 & n5928 ) ;
  assign n5931 = ( x40 & n5929 ) | ( x40 & ~n5930 ) | ( n5929 & ~n5930 ) ;
  assign n5932 = ( ~n5920 & n5926 ) | ( ~n5920 & n5931 ) | ( n5926 & n5931 ) ;
  assign n5933 = ( n5920 & n5926 ) | ( n5920 & n5931 ) | ( n5926 & n5931 ) ;
  assign n5934 = ( n5920 & n5932 ) | ( n5920 & ~n5933 ) | ( n5932 & ~n5933 ) ;
  assign n5935 = ( n5766 & n5914 ) | ( n5766 & n5934 ) | ( n5914 & n5934 ) ;
  assign n5936 = ( ~n5766 & n5914 ) | ( ~n5766 & n5934 ) | ( n5914 & n5934 ) ;
  assign n5937 = ( n5766 & ~n5935 ) | ( n5766 & n5936 ) | ( ~n5935 & n5936 ) ;
  assign n5938 = ( n5769 & n5893 ) | ( n5769 & n5937 ) | ( n5893 & n5937 ) ;
  assign n5939 = ( ~n5769 & n5893 ) | ( ~n5769 & n5937 ) | ( n5893 & n5937 ) ;
  assign n5940 = ( n5769 & ~n5938 ) | ( n5769 & n5939 ) | ( ~n5938 & n5939 ) ;
  assign n5941 = ( ~n5796 & n5887 ) | ( ~n5796 & n5940 ) | ( n5887 & n5940 ) ;
  assign n5942 = ( n5796 & n5887 ) | ( n5796 & n5940 ) | ( n5887 & n5940 ) ;
  assign n5943 = ( n5796 & n5941 ) | ( n5796 & ~n5942 ) | ( n5941 & ~n5942 ) ;
  assign n5944 = ( n5846 & n5849 ) | ( n5846 & n5943 ) | ( n5849 & n5943 ) ;
  assign n5945 = ( ~n5846 & n5849 ) | ( ~n5846 & n5943 ) | ( n5849 & n5943 ) ;
  assign n5946 = ( n5846 & ~n5944 ) | ( n5846 & n5945 ) | ( ~n5944 & n5945 ) ;
  assign n5947 = x20 & x60 ;
  assign n5948 = x21 & x59 ;
  assign n5949 = x22 & x58 ;
  assign n5950 = ( ~n5947 & n5948 ) | ( ~n5947 & n5949 ) | ( n5948 & n5949 ) ;
  assign n5951 = ( n5947 & n5948 ) | ( n5947 & n5949 ) | ( n5948 & n5949 ) ;
  assign n5952 = ( n5947 & n5950 ) | ( n5947 & ~n5951 ) | ( n5950 & ~n5951 ) ;
  assign n5953 = x30 & x50 ;
  assign n5954 = x31 & x49 ;
  assign n5955 = x32 & x48 ;
  assign n5956 = ( ~n5953 & n5954 ) | ( ~n5953 & n5955 ) | ( n5954 & n5955 ) ;
  assign n5957 = ( n5953 & n5954 ) | ( n5953 & n5955 ) | ( n5954 & n5955 ) ;
  assign n5958 = ( n5953 & n5956 ) | ( n5953 & ~n5957 ) | ( n5956 & ~n5957 ) ;
  assign n5959 = ( n5925 & n5952 ) | ( n5925 & n5958 ) | ( n5952 & n5958 ) ;
  assign n5960 = ( ~n5925 & n5952 ) | ( ~n5925 & n5958 ) | ( n5952 & n5958 ) ;
  assign n5961 = ( n5925 & ~n5959 ) | ( n5925 & n5960 ) | ( ~n5959 & n5960 ) ;
  assign n5962 = x19 & x61 ;
  assign n5963 = x18 & x62 ;
  assign n5964 = ( n5930 & n5962 ) | ( n5930 & n5963 ) | ( n5962 & n5963 ) ;
  assign n5965 = ( ~n5930 & n5962 ) | ( ~n5930 & n5963 ) | ( n5962 & n5963 ) ;
  assign n5966 = ( n5930 & ~n5964 ) | ( n5930 & n5965 ) | ( ~n5964 & n5965 ) ;
  assign n5967 = x34 & x46 ;
  assign n5968 = x35 & x45 ;
  assign n5969 = x36 & x44 ;
  assign n5970 = ( ~n5967 & n5968 ) | ( ~n5967 & n5969 ) | ( n5968 & n5969 ) ;
  assign n5971 = ( n5967 & n5968 ) | ( n5967 & n5969 ) | ( n5968 & n5969 ) ;
  assign n5972 = ( n5967 & n5970 ) | ( n5967 & ~n5971 ) | ( n5970 & ~n5971 ) ;
  assign n5973 = x33 & x47 ;
  assign n5974 = x17 & x63 ;
  assign n5975 = x29 & x51 ;
  assign n5976 = ( ~n5973 & n5974 ) | ( ~n5973 & n5975 ) | ( n5974 & n5975 ) ;
  assign n5977 = ( n5973 & n5974 ) | ( n5973 & n5975 ) | ( n5974 & n5975 ) ;
  assign n5978 = ( n5973 & n5976 ) | ( n5973 & ~n5977 ) | ( n5976 & ~n5977 ) ;
  assign n5979 = ( n5966 & n5972 ) | ( n5966 & n5978 ) | ( n5972 & n5978 ) ;
  assign n5980 = ( ~n5966 & n5972 ) | ( ~n5966 & n5978 ) | ( n5972 & n5978 ) ;
  assign n5981 = ( n5966 & ~n5979 ) | ( n5966 & n5980 ) | ( ~n5979 & n5980 ) ;
  assign n5982 = x23 & x57 ;
  assign n5983 = x24 & x56 ;
  assign n5984 = x26 & x54 ;
  assign n5985 = ( ~n5982 & n5983 ) | ( ~n5982 & n5984 ) | ( n5983 & n5984 ) ;
  assign n5986 = ( n5982 & n5983 ) | ( n5982 & n5984 ) | ( n5983 & n5984 ) ;
  assign n5987 = ( n5982 & n5985 ) | ( n5982 & ~n5986 ) | ( n5985 & ~n5986 ) ;
  assign n5988 = x39 & x41 ;
  assign n5989 = x27 & x53 ;
  assign n5990 = x28 & x52 ;
  assign n5991 = ( ~n5988 & n5989 ) | ( ~n5988 & n5990 ) | ( n5989 & n5990 ) ;
  assign n5992 = ( n5988 & n5989 ) | ( n5988 & n5990 ) | ( n5989 & n5990 ) ;
  assign n5993 = ( n5988 & n5991 ) | ( n5988 & ~n5992 ) | ( n5991 & ~n5992 ) ;
  assign n5994 = x25 & x55 ;
  assign n5995 = x37 & x43 ;
  assign n5996 = x38 & x42 ;
  assign n5997 = ( ~n5994 & n5995 ) | ( ~n5994 & n5996 ) | ( n5995 & n5996 ) ;
  assign n5998 = ( n5994 & n5995 ) | ( n5994 & n5996 ) | ( n5995 & n5996 ) ;
  assign n5999 = ( n5994 & n5997 ) | ( n5994 & ~n5998 ) | ( n5997 & ~n5998 ) ;
  assign n6000 = ( ~n5987 & n5993 ) | ( ~n5987 & n5999 ) | ( n5993 & n5999 ) ;
  assign n6001 = ( n5987 & n5993 ) | ( n5987 & n5999 ) | ( n5993 & n5999 ) ;
  assign n6002 = ( n5987 & n6000 ) | ( n5987 & ~n6001 ) | ( n6000 & ~n6001 ) ;
  assign n6003 = ( ~n5961 & n5981 ) | ( ~n5961 & n6002 ) | ( n5981 & n6002 ) ;
  assign n6004 = ( n5961 & n5981 ) | ( n5961 & n6002 ) | ( n5981 & n6002 ) ;
  assign n6005 = ( n5961 & n6003 ) | ( n5961 & ~n6004 ) | ( n6003 & ~n6004 ) ;
  assign n6006 = ( ~n5882 & n5891 ) | ( ~n5882 & n6005 ) | ( n5891 & n6005 ) ;
  assign n6007 = ( n5882 & n5891 ) | ( n5882 & n6005 ) | ( n5891 & n6005 ) ;
  assign n6008 = ( n5882 & n6006 ) | ( n5882 & ~n6007 ) | ( n6006 & ~n6007 ) ;
  assign n6009 = ( n5855 & ~n5861 ) | ( n5855 & n5919 ) | ( ~n5861 & n5919 ) ;
  assign n6010 = ( n5855 & n5861 ) | ( n5855 & n5919 ) | ( n5861 & n5919 ) ;
  assign n6011 = ( n5861 & n6009 ) | ( n5861 & ~n6010 ) | ( n6009 & ~n6010 ) ;
  assign n6012 = ( n5863 & n5888 ) | ( n5863 & n6011 ) | ( n5888 & n6011 ) ;
  assign n6013 = ( n5863 & ~n5888 ) | ( n5863 & n6011 ) | ( ~n5888 & n6011 ) ;
  assign n6014 = ( n5888 & ~n6012 ) | ( n5888 & n6013 ) | ( ~n6012 & n6013 ) ;
  assign n6015 = ( ~n5898 & n5904 ) | ( ~n5898 & n5910 ) | ( n5904 & n5910 ) ;
  assign n6016 = ( n5898 & n5904 ) | ( n5898 & n5910 ) | ( n5904 & n5910 ) ;
  assign n6017 = ( n5898 & n6015 ) | ( n5898 & ~n6016 ) | ( n6015 & ~n6016 ) ;
  assign n6018 = ( n5913 & n5933 ) | ( n5913 & n6017 ) | ( n5933 & n6017 ) ;
  assign n6019 = ( ~n5913 & n5933 ) | ( ~n5913 & n6017 ) | ( n5933 & n6017 ) ;
  assign n6020 = ( n5913 & ~n6018 ) | ( n5913 & n6019 ) | ( ~n6018 & n6019 ) ;
  assign n6021 = ( ~n5935 & n6014 ) | ( ~n5935 & n6020 ) | ( n6014 & n6020 ) ;
  assign n6022 = ( n5935 & n6014 ) | ( n5935 & n6020 ) | ( n6014 & n6020 ) ;
  assign n6023 = ( n5935 & n6021 ) | ( n5935 & ~n6022 ) | ( n6021 & ~n6022 ) ;
  assign n6024 = ( n5867 & n5872 ) | ( n5867 & n5877 ) | ( n5872 & n5877 ) ;
  assign n6025 = ( n5867 & ~n5872 ) | ( n5867 & n5877 ) | ( ~n5872 & n5877 ) ;
  assign n6026 = ( n5872 & ~n6024 ) | ( n5872 & n6025 ) | ( ~n6024 & n6025 ) ;
  assign n6027 = ( ~n5869 & n5880 ) | ( ~n5869 & n6026 ) | ( n5880 & n6026 ) ;
  assign n6028 = ( n5869 & n5880 ) | ( n5869 & n6026 ) | ( n5880 & n6026 ) ;
  assign n6029 = ( n5869 & n6027 ) | ( n5869 & ~n6028 ) | ( n6027 & ~n6028 ) ;
  assign n6030 = ( n5938 & n6023 ) | ( n5938 & n6029 ) | ( n6023 & n6029 ) ;
  assign n6031 = ( ~n5938 & n6023 ) | ( ~n5938 & n6029 ) | ( n6023 & n6029 ) ;
  assign n6032 = ( n5938 & ~n6030 ) | ( n5938 & n6031 ) | ( ~n6030 & n6031 ) ;
  assign n6033 = ( n5885 & n6008 ) | ( n5885 & n6032 ) | ( n6008 & n6032 ) ;
  assign n6034 = ( ~n5885 & n6008 ) | ( ~n5885 & n6032 ) | ( n6008 & n6032 ) ;
  assign n6035 = ( n5885 & ~n6033 ) | ( n5885 & n6034 ) | ( ~n6033 & n6034 ) ;
  assign n6036 = ( n5942 & n5944 ) | ( n5942 & n6035 ) | ( n5944 & n6035 ) ;
  assign n6037 = ( ~n5942 & n5944 ) | ( ~n5942 & n6035 ) | ( n5944 & n6035 ) ;
  assign n6038 = ( n5942 & ~n6036 ) | ( n5942 & n6037 ) | ( ~n6036 & n6037 ) ;
  assign n6039 = ( n5951 & n5957 ) | ( n5951 & ~n5977 ) | ( n5957 & ~n5977 ) ;
  assign n6040 = ( n5951 & n5957 ) | ( n5951 & n5977 ) | ( n5957 & n5977 ) ;
  assign n6041 = ( n5977 & n6039 ) | ( n5977 & ~n6040 ) | ( n6039 & ~n6040 ) ;
  assign n6042 = x30 & x51 ;
  assign n6043 = x32 & x49 ;
  assign n6044 = x31 & x50 ;
  assign n6045 = ( ~n6042 & n6043 ) | ( ~n6042 & n6044 ) | ( n6043 & n6044 ) ;
  assign n6046 = ( n6042 & n6043 ) | ( n6042 & n6044 ) | ( n6043 & n6044 ) ;
  assign n6047 = ( n6042 & n6045 ) | ( n6042 & ~n6046 ) | ( n6045 & ~n6046 ) ;
  assign n6048 = ( ~n5964 & n5971 ) | ( ~n5964 & n6047 ) | ( n5971 & n6047 ) ;
  assign n6049 = ( n5964 & n5971 ) | ( n5964 & n6047 ) | ( n5971 & n6047 ) ;
  assign n6050 = ( n5964 & n6048 ) | ( n5964 & ~n6049 ) | ( n6048 & ~n6049 ) ;
  assign n6051 = ( ~n5979 & n6041 ) | ( ~n5979 & n6050 ) | ( n6041 & n6050 ) ;
  assign n6052 = ( n5979 & n6041 ) | ( n5979 & n6050 ) | ( n6041 & n6050 ) ;
  assign n6053 = ( n5979 & n6051 ) | ( n5979 & ~n6052 ) | ( n6051 & ~n6052 ) ;
  assign n6054 = ( n5986 & n5992 ) | ( n5986 & n5998 ) | ( n5992 & n5998 ) ;
  assign n6055 = ( n5986 & n5992 ) | ( n5986 & ~n5998 ) | ( n5992 & ~n5998 ) ;
  assign n6056 = ( n5998 & ~n6054 ) | ( n5998 & n6055 ) | ( ~n6054 & n6055 ) ;
  assign n6057 = ( ~n5959 & n6001 ) | ( ~n5959 & n6056 ) | ( n6001 & n6056 ) ;
  assign n6058 = ( n5959 & n6001 ) | ( n5959 & n6056 ) | ( n6001 & n6056 ) ;
  assign n6059 = ( n5959 & n6057 ) | ( n5959 & ~n6058 ) | ( n6057 & ~n6058 ) ;
  assign n6060 = ( n6004 & n6053 ) | ( n6004 & n6059 ) | ( n6053 & n6059 ) ;
  assign n6061 = ( ~n6004 & n6053 ) | ( ~n6004 & n6059 ) | ( n6053 & n6059 ) ;
  assign n6062 = ( n6004 & ~n6060 ) | ( n6004 & n6061 ) | ( ~n6060 & n6061 ) ;
  assign n6063 = x27 & x54 ;
  assign n6064 = x38 & x43 ;
  assign n6065 = x39 & x42 ;
  assign n6066 = ( ~n6063 & n6064 ) | ( ~n6063 & n6065 ) | ( n6064 & n6065 ) ;
  assign n6067 = ( n6063 & n6064 ) | ( n6063 & n6065 ) | ( n6064 & n6065 ) ;
  assign n6068 = ( n6063 & n6066 ) | ( n6063 & ~n6067 ) | ( n6066 & ~n6067 ) ;
  assign n6069 = ( ~n6010 & n6016 ) | ( ~n6010 & n6068 ) | ( n6016 & n6068 ) ;
  assign n6070 = ( n6010 & n6016 ) | ( n6010 & n6068 ) | ( n6016 & n6068 ) ;
  assign n6071 = ( n6010 & n6069 ) | ( n6010 & ~n6070 ) | ( n6069 & ~n6070 ) ;
  assign n6072 = ( ~n6012 & n6018 ) | ( ~n6012 & n6071 ) | ( n6018 & n6071 ) ;
  assign n6073 = ( n6012 & n6018 ) | ( n6012 & n6071 ) | ( n6018 & n6071 ) ;
  assign n6074 = ( n6012 & n6072 ) | ( n6012 & ~n6073 ) | ( n6072 & ~n6073 ) ;
  assign n6075 = ( n6007 & n6062 ) | ( n6007 & n6074 ) | ( n6062 & n6074 ) ;
  assign n6076 = ( ~n6007 & n6062 ) | ( ~n6007 & n6074 ) | ( n6062 & n6074 ) ;
  assign n6077 = ( n6007 & ~n6075 ) | ( n6007 & n6076 ) | ( ~n6075 & n6076 ) ;
  assign n6078 = x40 & x41 ;
  assign n6079 = x19 & x62 ;
  assign n6080 = ( x41 & n6078 ) | ( x41 & n6079 ) | ( n6078 & n6079 ) ;
  assign n6081 = ( x41 & ~n6078 ) | ( x41 & n6079 ) | ( ~n6078 & n6079 ) ;
  assign n6082 = ( n6078 & ~n6080 ) | ( n6078 & n6081 ) | ( ~n6080 & n6081 ) ;
  assign n6083 = x24 & x57 ;
  assign n6084 = x33 & x48 ;
  assign n6085 = x34 & x47 ;
  assign n6086 = ( ~n6083 & n6084 ) | ( ~n6083 & n6085 ) | ( n6084 & n6085 ) ;
  assign n6087 = ( n6083 & n6084 ) | ( n6083 & n6085 ) | ( n6084 & n6085 ) ;
  assign n6088 = ( n6083 & n6086 ) | ( n6083 & ~n6087 ) | ( n6086 & ~n6087 ) ;
  assign n6089 = x22 & x59 ;
  assign n6090 = x25 & x56 ;
  assign n6091 = x23 & x58 ;
  assign n6092 = ( ~n6089 & n6090 ) | ( ~n6089 & n6091 ) | ( n6090 & n6091 ) ;
  assign n6093 = ( n6089 & n6090 ) | ( n6089 & n6091 ) | ( n6090 & n6091 ) ;
  assign n6094 = ( n6089 & n6092 ) | ( n6089 & ~n6093 ) | ( n6092 & ~n6093 ) ;
  assign n6095 = ( n6082 & n6088 ) | ( n6082 & n6094 ) | ( n6088 & n6094 ) ;
  assign n6096 = ( ~n6082 & n6088 ) | ( ~n6082 & n6094 ) | ( n6088 & n6094 ) ;
  assign n6097 = ( n6082 & ~n6095 ) | ( n6082 & n6096 ) | ( ~n6095 & n6096 ) ;
  assign n6098 = x35 & x46 ;
  assign n6099 = x36 & x45 ;
  assign n6100 = x37 & x44 ;
  assign n6101 = ( ~n6098 & n6099 ) | ( ~n6098 & n6100 ) | ( n6099 & n6100 ) ;
  assign n6102 = ( n6098 & n6099 ) | ( n6098 & n6100 ) | ( n6099 & n6100 ) ;
  assign n6103 = ( n6098 & n6101 ) | ( n6098 & ~n6102 ) | ( n6101 & ~n6102 ) ;
  assign n6104 = x18 & x63 ;
  assign n6105 = x20 & x61 ;
  assign n6106 = x21 & x60 ;
  assign n6107 = ( ~n6104 & n6105 ) | ( ~n6104 & n6106 ) | ( n6105 & n6106 ) ;
  assign n6108 = ( n6104 & n6105 ) | ( n6104 & n6106 ) | ( n6105 & n6106 ) ;
  assign n6109 = ( n6104 & n6107 ) | ( n6104 & ~n6108 ) | ( n6107 & ~n6108 ) ;
  assign n6110 = x26 & x55 ;
  assign n6111 = x28 & x53 ;
  assign n6112 = x29 & x52 ;
  assign n6113 = ( ~n6110 & n6111 ) | ( ~n6110 & n6112 ) | ( n6111 & n6112 ) ;
  assign n6114 = ( n6110 & n6111 ) | ( n6110 & n6112 ) | ( n6111 & n6112 ) ;
  assign n6115 = ( n6110 & n6113 ) | ( n6110 & ~n6114 ) | ( n6113 & ~n6114 ) ;
  assign n6116 = ( n6103 & n6109 ) | ( n6103 & n6115 ) | ( n6109 & n6115 ) ;
  assign n6117 = ( ~n6103 & n6109 ) | ( ~n6103 & n6115 ) | ( n6109 & n6115 ) ;
  assign n6118 = ( n6103 & ~n6116 ) | ( n6103 & n6117 ) | ( ~n6116 & n6117 ) ;
  assign n6119 = ( ~n6024 & n6097 ) | ( ~n6024 & n6118 ) | ( n6097 & n6118 ) ;
  assign n6120 = ( n6024 & n6097 ) | ( n6024 & n6118 ) | ( n6097 & n6118 ) ;
  assign n6121 = ( n6024 & n6119 ) | ( n6024 & ~n6120 ) | ( n6119 & ~n6120 ) ;
  assign n6122 = ( ~n6022 & n6028 ) | ( ~n6022 & n6121 ) | ( n6028 & n6121 ) ;
  assign n6123 = ( n6022 & n6028 ) | ( n6022 & n6121 ) | ( n6028 & n6121 ) ;
  assign n6124 = ( n6022 & n6122 ) | ( n6022 & ~n6123 ) | ( n6122 & ~n6123 ) ;
  assign n6125 = ( ~n6030 & n6077 ) | ( ~n6030 & n6124 ) | ( n6077 & n6124 ) ;
  assign n6126 = ( n6030 & n6077 ) | ( n6030 & n6124 ) | ( n6077 & n6124 ) ;
  assign n6127 = ( n6030 & n6125 ) | ( n6030 & ~n6126 ) | ( n6125 & ~n6126 ) ;
  assign n6128 = ( ~n6033 & n6036 ) | ( ~n6033 & n6127 ) | ( n6036 & n6127 ) ;
  assign n6129 = ( n6033 & n6036 ) | ( n6033 & n6127 ) | ( n6036 & n6127 ) ;
  assign n6130 = ( n6033 & n6128 ) | ( n6033 & ~n6129 ) | ( n6128 & ~n6129 ) ;
  assign n6131 = x19 & x63 ;
  assign n6132 = ( n6067 & n6080 ) | ( n6067 & n6131 ) | ( n6080 & n6131 ) ;
  assign n6133 = ( ~n6067 & n6080 ) | ( ~n6067 & n6131 ) | ( n6080 & n6131 ) ;
  assign n6134 = ( n6067 & ~n6132 ) | ( n6067 & n6133 ) | ( ~n6132 & n6133 ) ;
  assign n6135 = ( n6049 & n6095 ) | ( n6049 & n6134 ) | ( n6095 & n6134 ) ;
  assign n6136 = ( n6049 & ~n6095 ) | ( n6049 & n6134 ) | ( ~n6095 & n6134 ) ;
  assign n6137 = ( n6095 & ~n6135 ) | ( n6095 & n6136 ) | ( ~n6135 & n6136 ) ;
  assign n6138 = ( n6046 & n6087 ) | ( n6046 & ~n6114 ) | ( n6087 & ~n6114 ) ;
  assign n6139 = ( n6046 & n6087 ) | ( n6046 & n6114 ) | ( n6087 & n6114 ) ;
  assign n6140 = ( n6114 & n6138 ) | ( n6114 & ~n6139 ) | ( n6138 & ~n6139 ) ;
  assign n6141 = ( n6093 & ~n6102 ) | ( n6093 & n6108 ) | ( ~n6102 & n6108 ) ;
  assign n6142 = ( n6093 & n6102 ) | ( n6093 & n6108 ) | ( n6102 & n6108 ) ;
  assign n6143 = ( n6102 & n6141 ) | ( n6102 & ~n6142 ) | ( n6141 & ~n6142 ) ;
  assign n6144 = ( ~n6116 & n6140 ) | ( ~n6116 & n6143 ) | ( n6140 & n6143 ) ;
  assign n6145 = ( n6116 & n6140 ) | ( n6116 & n6143 ) | ( n6140 & n6143 ) ;
  assign n6146 = ( n6116 & n6144 ) | ( n6116 & ~n6145 ) | ( n6144 & ~n6145 ) ;
  assign n6147 = ( ~n6120 & n6137 ) | ( ~n6120 & n6146 ) | ( n6137 & n6146 ) ;
  assign n6148 = ( n6120 & n6137 ) | ( n6120 & n6146 ) | ( n6137 & n6146 ) ;
  assign n6149 = ( n6120 & n6147 ) | ( n6120 & ~n6148 ) | ( n6147 & ~n6148 ) ;
  assign n6150 = x27 & x55 ;
  assign n6151 = x25 & x57 ;
  assign n6152 = ( ~n3115 & n6150 ) | ( ~n3115 & n6151 ) | ( n6150 & n6151 ) ;
  assign n6153 = ( n3115 & n6150 ) | ( n3115 & n6151 ) | ( n6150 & n6151 ) ;
  assign n6154 = ( n3115 & n6152 ) | ( n3115 & ~n6153 ) | ( n6152 & ~n6153 ) ;
  assign n6155 = ( ~n6040 & n6054 ) | ( ~n6040 & n6154 ) | ( n6054 & n6154 ) ;
  assign n6156 = ( n6040 & n6054 ) | ( n6040 & n6154 ) | ( n6054 & n6154 ) ;
  assign n6157 = ( n6040 & n6155 ) | ( n6040 & ~n6156 ) | ( n6155 & ~n6156 ) ;
  assign n6158 = ( ~n6052 & n6058 ) | ( ~n6052 & n6157 ) | ( n6058 & n6157 ) ;
  assign n6159 = ( n6052 & n6058 ) | ( n6052 & n6157 ) | ( n6058 & n6157 ) ;
  assign n6160 = ( n6052 & n6158 ) | ( n6052 & ~n6159 ) | ( n6158 & ~n6159 ) ;
  assign n6161 = ( ~n6123 & n6149 ) | ( ~n6123 & n6160 ) | ( n6149 & n6160 ) ;
  assign n6162 = ( n6123 & n6149 ) | ( n6123 & n6160 ) | ( n6149 & n6160 ) ;
  assign n6163 = ( n6123 & n6161 ) | ( n6123 & ~n6162 ) | ( n6161 & ~n6162 ) ;
  assign n6164 = x21 & x61 ;
  assign n6165 = x20 & x62 ;
  assign n6166 = x31 & x51 ;
  assign n6167 = ( ~n6164 & n6165 ) | ( ~n6164 & n6166 ) | ( n6165 & n6166 ) ;
  assign n6168 = ( n6164 & n6165 ) | ( n6164 & n6166 ) | ( n6165 & n6166 ) ;
  assign n6169 = ( n6164 & n6167 ) | ( n6164 & ~n6168 ) | ( n6167 & ~n6168 ) ;
  assign n6170 = x22 & x60 ;
  assign n6171 = x24 & x58 ;
  assign n6172 = x23 & x59 ;
  assign n6173 = ( ~n6170 & n6171 ) | ( ~n6170 & n6172 ) | ( n6171 & n6172 ) ;
  assign n6174 = ( n6170 & n6171 ) | ( n6170 & n6172 ) | ( n6171 & n6172 ) ;
  assign n6175 = ( n6170 & n6173 ) | ( n6170 & ~n6174 ) | ( n6173 & ~n6174 ) ;
  assign n6176 = x32 & x50 ;
  assign n6177 = x34 & x48 ;
  assign n6178 = x33 & x49 ;
  assign n6179 = ( ~n6176 & n6177 ) | ( ~n6176 & n6178 ) | ( n6177 & n6178 ) ;
  assign n6180 = ( n6176 & n6177 ) | ( n6176 & n6178 ) | ( n6177 & n6178 ) ;
  assign n6181 = ( n6176 & n6179 ) | ( n6176 & ~n6180 ) | ( n6179 & ~n6180 ) ;
  assign n6182 = ( ~n6169 & n6175 ) | ( ~n6169 & n6181 ) | ( n6175 & n6181 ) ;
  assign n6183 = ( n6169 & n6175 ) | ( n6169 & n6181 ) | ( n6175 & n6181 ) ;
  assign n6184 = ( n6169 & n6182 ) | ( n6169 & ~n6183 ) | ( n6182 & ~n6183 ) ;
  assign n6185 = x35 & x47 ;
  assign n6186 = x37 & x45 ;
  assign n6187 = x36 & x46 ;
  assign n6188 = ( ~n6185 & n6186 ) | ( ~n6185 & n6187 ) | ( n6186 & n6187 ) ;
  assign n6189 = ( n6185 & n6186 ) | ( n6185 & n6187 ) | ( n6186 & n6187 ) ;
  assign n6190 = ( n6185 & n6188 ) | ( n6185 & ~n6189 ) | ( n6188 & ~n6189 ) ;
  assign n6191 = x40 & x42 ;
  assign n6192 = x29 & x53 ;
  assign n6193 = x30 & x52 ;
  assign n6194 = ( ~n6191 & n6192 ) | ( ~n6191 & n6193 ) | ( n6192 & n6193 ) ;
  assign n6195 = ( n6191 & n6192 ) | ( n6191 & n6193 ) | ( n6192 & n6193 ) ;
  assign n6196 = ( n6191 & n6194 ) | ( n6191 & ~n6195 ) | ( n6194 & ~n6195 ) ;
  assign n6197 = x26 & x56 ;
  assign n6198 = x39 & x43 ;
  assign n6199 = x38 & x44 ;
  assign n6200 = ( ~n6197 & n6198 ) | ( ~n6197 & n6199 ) | ( n6198 & n6199 ) ;
  assign n6201 = ( n6197 & n6198 ) | ( n6197 & n6199 ) | ( n6198 & n6199 ) ;
  assign n6202 = ( n6197 & n6200 ) | ( n6197 & ~n6201 ) | ( n6200 & ~n6201 ) ;
  assign n6203 = ( ~n6190 & n6196 ) | ( ~n6190 & n6202 ) | ( n6196 & n6202 ) ;
  assign n6204 = ( n6190 & n6196 ) | ( n6190 & n6202 ) | ( n6196 & n6202 ) ;
  assign n6205 = ( n6190 & n6203 ) | ( n6190 & ~n6204 ) | ( n6203 & ~n6204 ) ;
  assign n6206 = ( n6070 & n6184 ) | ( n6070 & n6205 ) | ( n6184 & n6205 ) ;
  assign n6207 = ( ~n6070 & n6184 ) | ( ~n6070 & n6205 ) | ( n6184 & n6205 ) ;
  assign n6208 = ( n6070 & ~n6206 ) | ( n6070 & n6207 ) | ( ~n6206 & n6207 ) ;
  assign n6209 = ( n6060 & n6073 ) | ( n6060 & n6208 ) | ( n6073 & n6208 ) ;
  assign n6210 = ( ~n6060 & n6073 ) | ( ~n6060 & n6208 ) | ( n6073 & n6208 ) ;
  assign n6211 = ( n6060 & ~n6209 ) | ( n6060 & n6210 ) | ( ~n6209 & n6210 ) ;
  assign n6212 = ( ~n6075 & n6163 ) | ( ~n6075 & n6211 ) | ( n6163 & n6211 ) ;
  assign n6213 = ( n6075 & n6163 ) | ( n6075 & n6211 ) | ( n6163 & n6211 ) ;
  assign n6214 = ( n6075 & n6212 ) | ( n6075 & ~n6213 ) | ( n6212 & ~n6213 ) ;
  assign n6215 = ( n6126 & n6129 ) | ( n6126 & n6214 ) | ( n6129 & n6214 ) ;
  assign n6216 = ( ~n6126 & n6129 ) | ( ~n6126 & n6214 ) | ( n6129 & n6214 ) ;
  assign n6217 = ( n6126 & ~n6215 ) | ( n6126 & n6216 ) | ( ~n6215 & n6216 ) ;
  assign n6218 = x41 & x42 ;
  assign n6219 = x21 & x62 ;
  assign n6220 = ( x42 & n6218 ) | ( x42 & n6219 ) | ( n6218 & n6219 ) ;
  assign n6221 = ( x42 & ~n6218 ) | ( x42 & n6219 ) | ( ~n6218 & n6219 ) ;
  assign n6222 = ( n6218 & ~n6220 ) | ( n6218 & n6221 ) | ( ~n6220 & n6221 ) ;
  assign n6223 = x33 & x50 ;
  assign n6224 = x34 & x49 ;
  assign n6225 = x35 & x48 ;
  assign n6226 = ( ~n6223 & n6224 ) | ( ~n6223 & n6225 ) | ( n6224 & n6225 ) ;
  assign n6227 = ( n6223 & n6224 ) | ( n6223 & n6225 ) | ( n6224 & n6225 ) ;
  assign n6228 = ( n6223 & n6226 ) | ( n6223 & ~n6227 ) | ( n6226 & ~n6227 ) ;
  assign n6229 = x29 & x54 ;
  assign n6230 = x39 & x44 ;
  assign n6231 = x40 & x43 ;
  assign n6232 = ( ~n6229 & n6230 ) | ( ~n6229 & n6231 ) | ( n6230 & n6231 ) ;
  assign n6233 = ( n6229 & n6230 ) | ( n6229 & n6231 ) | ( n6230 & n6231 ) ;
  assign n6234 = ( n6229 & n6232 ) | ( n6229 & ~n6233 ) | ( n6232 & ~n6233 ) ;
  assign n6235 = ( n6222 & n6228 ) | ( n6222 & n6234 ) | ( n6228 & n6234 ) ;
  assign n6236 = ( ~n6222 & n6228 ) | ( ~n6222 & n6234 ) | ( n6228 & n6234 ) ;
  assign n6237 = ( n6222 & ~n6235 ) | ( n6222 & n6236 ) | ( ~n6235 & n6236 ) ;
  assign n6238 = x27 & x56 ;
  assign n6239 = x20 & x63 ;
  assign n6240 = x22 & x61 ;
  assign n6241 = ( ~n6238 & n6239 ) | ( ~n6238 & n6240 ) | ( n6239 & n6240 ) ;
  assign n6242 = ( n6238 & n6239 ) | ( n6238 & n6240 ) | ( n6239 & n6240 ) ;
  assign n6243 = ( n6238 & n6241 ) | ( n6238 & ~n6242 ) | ( n6241 & ~n6242 ) ;
  assign n6244 = x36 & x47 ;
  assign n6245 = x37 & x46 ;
  assign n6246 = x38 & x45 ;
  assign n6247 = ( ~n6244 & n6245 ) | ( ~n6244 & n6246 ) | ( n6245 & n6246 ) ;
  assign n6248 = ( n6244 & n6245 ) | ( n6244 & n6246 ) | ( n6245 & n6246 ) ;
  assign n6249 = ( n6244 & n6247 ) | ( n6244 & ~n6248 ) | ( n6247 & ~n6248 ) ;
  assign n6250 = x25 & x58 ;
  assign n6251 = x26 & x57 ;
  assign n6252 = x32 & x51 ;
  assign n6253 = ( ~n6250 & n6251 ) | ( ~n6250 & n6252 ) | ( n6251 & n6252 ) ;
  assign n6254 = ( n6250 & n6251 ) | ( n6250 & n6252 ) | ( n6251 & n6252 ) ;
  assign n6255 = ( n6250 & n6253 ) | ( n6250 & ~n6254 ) | ( n6253 & ~n6254 ) ;
  assign n6256 = ( ~n6243 & n6249 ) | ( ~n6243 & n6255 ) | ( n6249 & n6255 ) ;
  assign n6257 = ( n6243 & n6249 ) | ( n6243 & n6255 ) | ( n6249 & n6255 ) ;
  assign n6258 = ( n6243 & n6256 ) | ( n6243 & ~n6257 ) | ( n6256 & ~n6257 ) ;
  assign n6259 = ( ~n6156 & n6237 ) | ( ~n6156 & n6258 ) | ( n6237 & n6258 ) ;
  assign n6260 = ( n6156 & n6237 ) | ( n6156 & n6258 ) | ( n6237 & n6258 ) ;
  assign n6261 = ( n6156 & n6259 ) | ( n6156 & ~n6260 ) | ( n6259 & ~n6260 ) ;
  assign n6262 = ( ~n6148 & n6159 ) | ( ~n6148 & n6261 ) | ( n6159 & n6261 ) ;
  assign n6263 = ( n6148 & n6159 ) | ( n6148 & n6261 ) | ( n6159 & n6261 ) ;
  assign n6264 = ( n6148 & n6262 ) | ( n6148 & ~n6263 ) | ( n6262 & ~n6263 ) ;
  assign n6265 = ( ~n6139 & n6142 ) | ( ~n6139 & n6183 ) | ( n6142 & n6183 ) ;
  assign n6266 = ( n6139 & n6142 ) | ( n6139 & n6183 ) | ( n6142 & n6183 ) ;
  assign n6267 = ( n6139 & n6265 ) | ( n6139 & ~n6266 ) | ( n6265 & ~n6266 ) ;
  assign n6268 = x31 & x52 ;
  assign n6269 = x30 & x53 ;
  assign n6270 = x28 & x55 ;
  assign n6271 = ( ~n6268 & n6269 ) | ( ~n6268 & n6270 ) | ( n6269 & n6270 ) ;
  assign n6272 = ( n6268 & n6269 ) | ( n6268 & n6270 ) | ( n6269 & n6270 ) ;
  assign n6273 = ( n6268 & n6271 ) | ( n6268 & ~n6272 ) | ( n6271 & ~n6272 ) ;
  assign n6274 = x24 & x59 ;
  assign n6275 = x23 & x60 ;
  assign n6276 = ( n6195 & n6274 ) | ( n6195 & n6275 ) | ( n6274 & n6275 ) ;
  assign n6277 = ( ~n6195 & n6274 ) | ( ~n6195 & n6275 ) | ( n6274 & n6275 ) ;
  assign n6278 = ( n6195 & ~n6276 ) | ( n6195 & n6277 ) | ( ~n6276 & n6277 ) ;
  assign n6279 = ( ~n6132 & n6273 ) | ( ~n6132 & n6278 ) | ( n6273 & n6278 ) ;
  assign n6280 = ( n6132 & n6273 ) | ( n6132 & n6278 ) | ( n6273 & n6278 ) ;
  assign n6281 = ( n6132 & n6279 ) | ( n6132 & ~n6280 ) | ( n6279 & ~n6280 ) ;
  assign n6282 = ( ~n6135 & n6267 ) | ( ~n6135 & n6281 ) | ( n6267 & n6281 ) ;
  assign n6283 = ( n6135 & n6267 ) | ( n6135 & n6281 ) | ( n6267 & n6281 ) ;
  assign n6284 = ( n6135 & n6282 ) | ( n6135 & ~n6283 ) | ( n6282 & ~n6283 ) ;
  assign n6285 = ( n6174 & ~n6189 ) | ( n6174 & n6201 ) | ( ~n6189 & n6201 ) ;
  assign n6286 = ( n6174 & n6189 ) | ( n6174 & n6201 ) | ( n6189 & n6201 ) ;
  assign n6287 = ( n6189 & n6285 ) | ( n6189 & ~n6286 ) | ( n6285 & ~n6286 ) ;
  assign n6288 = ( n6153 & n6168 ) | ( n6153 & ~n6180 ) | ( n6168 & ~n6180 ) ;
  assign n6289 = ( n6153 & n6168 ) | ( n6153 & n6180 ) | ( n6168 & n6180 ) ;
  assign n6290 = ( n6180 & n6288 ) | ( n6180 & ~n6289 ) | ( n6288 & ~n6289 ) ;
  assign n6291 = ( n6204 & n6287 ) | ( n6204 & n6290 ) | ( n6287 & n6290 ) ;
  assign n6292 = ( ~n6204 & n6287 ) | ( ~n6204 & n6290 ) | ( n6287 & n6290 ) ;
  assign n6293 = ( n6204 & ~n6291 ) | ( n6204 & n6292 ) | ( ~n6291 & n6292 ) ;
  assign n6294 = ( n6145 & n6206 ) | ( n6145 & n6293 ) | ( n6206 & n6293 ) ;
  assign n6295 = ( ~n6145 & n6206 ) | ( ~n6145 & n6293 ) | ( n6206 & n6293 ) ;
  assign n6296 = ( n6145 & ~n6294 ) | ( n6145 & n6295 ) | ( ~n6294 & n6295 ) ;
  assign n6297 = ( ~n6209 & n6284 ) | ( ~n6209 & n6296 ) | ( n6284 & n6296 ) ;
  assign n6298 = ( n6209 & n6284 ) | ( n6209 & n6296 ) | ( n6284 & n6296 ) ;
  assign n6299 = ( n6209 & n6297 ) | ( n6209 & ~n6298 ) | ( n6297 & ~n6298 ) ;
  assign n6300 = ( ~n6162 & n6264 ) | ( ~n6162 & n6299 ) | ( n6264 & n6299 ) ;
  assign n6301 = ( n6162 & n6264 ) | ( n6162 & n6299 ) | ( n6264 & n6299 ) ;
  assign n6302 = ( n6162 & n6300 ) | ( n6162 & ~n6301 ) | ( n6300 & ~n6301 ) ;
  assign n6303 = ( ~n6213 & n6215 ) | ( ~n6213 & n6302 ) | ( n6215 & n6302 ) ;
  assign n6304 = ( n6213 & n6215 ) | ( n6213 & n6302 ) | ( n6215 & n6302 ) ;
  assign n6305 = ( n6213 & n6303 ) | ( n6213 & ~n6304 ) | ( n6303 & ~n6304 ) ;
  assign n6306 = x26 & x58 ;
  assign n6307 = x31 & x53 ;
  assign n6308 = x32 & x52 ;
  assign n6309 = ( ~n6306 & n6307 ) | ( ~n6306 & n6308 ) | ( n6307 & n6308 ) ;
  assign n6310 = ( n6306 & n6307 ) | ( n6306 & n6308 ) | ( n6307 & n6308 ) ;
  assign n6311 = ( n6306 & n6309 ) | ( n6306 & ~n6310 ) | ( n6309 & ~n6310 ) ;
  assign n6312 = ( ~n6242 & n6276 ) | ( ~n6242 & n6311 ) | ( n6276 & n6311 ) ;
  assign n6313 = ( n6242 & n6276 ) | ( n6242 & n6311 ) | ( n6276 & n6311 ) ;
  assign n6314 = ( n6242 & n6312 ) | ( n6242 & ~n6313 ) | ( n6312 & ~n6313 ) ;
  assign n6315 = ( ~n6266 & n6280 ) | ( ~n6266 & n6314 ) | ( n6280 & n6314 ) ;
  assign n6316 = ( n6266 & n6280 ) | ( n6266 & n6314 ) | ( n6280 & n6314 ) ;
  assign n6317 = ( n6266 & n6315 ) | ( n6266 & ~n6316 ) | ( n6315 & ~n6316 ) ;
  assign n6318 = ( n6227 & ~n6248 ) | ( n6227 & n6254 ) | ( ~n6248 & n6254 ) ;
  assign n6319 = ( n6227 & n6248 ) | ( n6227 & n6254 ) | ( n6248 & n6254 ) ;
  assign n6320 = ( n6248 & n6318 ) | ( n6248 & ~n6319 ) | ( n6318 & ~n6319 ) ;
  assign n6321 = ( ~n6286 & n6289 ) | ( ~n6286 & n6320 ) | ( n6289 & n6320 ) ;
  assign n6322 = ( n6286 & n6289 ) | ( n6286 & n6320 ) | ( n6289 & n6320 ) ;
  assign n6323 = ( n6286 & n6321 ) | ( n6286 & ~n6322 ) | ( n6321 & ~n6322 ) ;
  assign n6324 = x34 & x50 ;
  assign n6325 = x35 & x49 ;
  assign n6326 = x36 & x48 ;
  assign n6327 = ( ~n6324 & n6325 ) | ( ~n6324 & n6326 ) | ( n6325 & n6326 ) ;
  assign n6328 = ( n6324 & n6325 ) | ( n6324 & n6326 ) | ( n6325 & n6326 ) ;
  assign n6329 = ( n6324 & n6327 ) | ( n6324 & ~n6328 ) | ( n6327 & ~n6328 ) ;
  assign n6330 = x33 & x51 ;
  assign n6331 = x24 & x60 ;
  assign n6332 = x25 & x59 ;
  assign n6333 = ( ~n6330 & n6331 ) | ( ~n6330 & n6332 ) | ( n6331 & n6332 ) ;
  assign n6334 = ( n6330 & n6331 ) | ( n6330 & n6332 ) | ( n6331 & n6332 ) ;
  assign n6335 = ( n6330 & n6333 ) | ( n6330 & ~n6334 ) | ( n6333 & ~n6334 ) ;
  assign n6336 = x21 & x63 ;
  assign n6337 = x22 & x62 ;
  assign n6338 = x23 & x61 ;
  assign n6339 = ( ~n6336 & n6337 ) | ( ~n6336 & n6338 ) | ( n6337 & n6338 ) ;
  assign n6340 = ( n6336 & n6337 ) | ( n6336 & n6338 ) | ( n6337 & n6338 ) ;
  assign n6341 = ( n6336 & n6339 ) | ( n6336 & ~n6340 ) | ( n6339 & ~n6340 ) ;
  assign n6342 = ( ~n6329 & n6335 ) | ( ~n6329 & n6341 ) | ( n6335 & n6341 ) ;
  assign n6343 = ( n6329 & n6335 ) | ( n6329 & n6341 ) | ( n6335 & n6341 ) ;
  assign n6344 = ( n6329 & n6342 ) | ( n6329 & ~n6343 ) | ( n6342 & ~n6343 ) ;
  assign n6345 = x37 & x47 ;
  assign n6346 = x27 & x57 ;
  assign n6347 = x30 & x54 ;
  assign n6348 = ( ~n6345 & n6346 ) | ( ~n6345 & n6347 ) | ( n6346 & n6347 ) ;
  assign n6349 = ( n6345 & n6346 ) | ( n6345 & n6347 ) | ( n6346 & n6347 ) ;
  assign n6350 = ( n6345 & n6348 ) | ( n6345 & ~n6349 ) | ( n6348 & ~n6349 ) ;
  assign n6351 = x38 & x46 ;
  assign n6352 = x28 & x56 ;
  assign n6353 = x29 & x55 ;
  assign n6354 = ( ~n6351 & n6352 ) | ( ~n6351 & n6353 ) | ( n6352 & n6353 ) ;
  assign n6355 = ( n6351 & n6352 ) | ( n6351 & n6353 ) | ( n6352 & n6353 ) ;
  assign n6356 = ( n6351 & n6354 ) | ( n6351 & ~n6355 ) | ( n6354 & ~n6355 ) ;
  assign n6357 = x39 & x45 ;
  assign n6358 = x40 & x44 ;
  assign n6359 = x41 & x43 ;
  assign n6360 = ( ~n6357 & n6358 ) | ( ~n6357 & n6359 ) | ( n6358 & n6359 ) ;
  assign n6361 = ( n6357 & n6358 ) | ( n6357 & n6359 ) | ( n6358 & n6359 ) ;
  assign n6362 = ( n6357 & n6360 ) | ( n6357 & ~n6361 ) | ( n6360 & ~n6361 ) ;
  assign n6363 = ( ~n6350 & n6356 ) | ( ~n6350 & n6362 ) | ( n6356 & n6362 ) ;
  assign n6364 = ( n6350 & n6356 ) | ( n6350 & n6362 ) | ( n6356 & n6362 ) ;
  assign n6365 = ( n6350 & n6363 ) | ( n6350 & ~n6364 ) | ( n6363 & ~n6364 ) ;
  assign n6366 = ( ~n6323 & n6344 ) | ( ~n6323 & n6365 ) | ( n6344 & n6365 ) ;
  assign n6367 = ( n6323 & n6344 ) | ( n6323 & n6365 ) | ( n6344 & n6365 ) ;
  assign n6368 = ( n6323 & n6366 ) | ( n6323 & ~n6367 ) | ( n6366 & ~n6367 ) ;
  assign n6369 = ( n6283 & n6317 ) | ( n6283 & n6368 ) | ( n6317 & n6368 ) ;
  assign n6370 = ( ~n6283 & n6317 ) | ( ~n6283 & n6368 ) | ( n6317 & n6368 ) ;
  assign n6371 = ( n6283 & ~n6369 ) | ( n6283 & n6370 ) | ( ~n6369 & n6370 ) ;
  assign n6372 = ( n6220 & ~n6233 ) | ( n6220 & n6272 ) | ( ~n6233 & n6272 ) ;
  assign n6373 = ( n6220 & n6233 ) | ( n6220 & n6272 ) | ( n6233 & n6272 ) ;
  assign n6374 = ( n6233 & n6372 ) | ( n6233 & ~n6373 ) | ( n6372 & ~n6373 ) ;
  assign n6375 = ( ~n6235 & n6257 ) | ( ~n6235 & n6374 ) | ( n6257 & n6374 ) ;
  assign n6376 = ( n6235 & n6257 ) | ( n6235 & n6374 ) | ( n6257 & n6374 ) ;
  assign n6377 = ( n6235 & n6375 ) | ( n6235 & ~n6376 ) | ( n6375 & ~n6376 ) ;
  assign n6378 = ( n6260 & n6291 ) | ( n6260 & n6377 ) | ( n6291 & n6377 ) ;
  assign n6379 = ( ~n6260 & n6291 ) | ( ~n6260 & n6377 ) | ( n6291 & n6377 ) ;
  assign n6380 = ( n6260 & ~n6378 ) | ( n6260 & n6379 ) | ( ~n6378 & n6379 ) ;
  assign n6381 = ( n6263 & n6294 ) | ( n6263 & n6380 ) | ( n6294 & n6380 ) ;
  assign n6382 = ( ~n6263 & n6294 ) | ( ~n6263 & n6380 ) | ( n6294 & n6380 ) ;
  assign n6383 = ( n6263 & ~n6381 ) | ( n6263 & n6382 ) | ( ~n6381 & n6382 ) ;
  assign n6384 = ( ~n6298 & n6371 ) | ( ~n6298 & n6383 ) | ( n6371 & n6383 ) ;
  assign n6385 = ( n6298 & n6371 ) | ( n6298 & n6383 ) | ( n6371 & n6383 ) ;
  assign n6386 = ( n6298 & n6384 ) | ( n6298 & ~n6385 ) | ( n6384 & ~n6385 ) ;
  assign n6387 = ( n6301 & n6304 ) | ( n6301 & n6386 ) | ( n6304 & n6386 ) ;
  assign n6388 = ( ~n6301 & n6304 ) | ( ~n6301 & n6386 ) | ( n6304 & n6386 ) ;
  assign n6389 = ( n6301 & ~n6387 ) | ( n6301 & n6388 ) | ( ~n6387 & n6388 ) ;
  assign n6390 = ( n6313 & ~n6319 ) | ( n6313 & n6373 ) | ( ~n6319 & n6373 ) ;
  assign n6391 = ( n6313 & n6319 ) | ( n6313 & n6373 ) | ( n6319 & n6373 ) ;
  assign n6392 = ( n6319 & n6390 ) | ( n6319 & ~n6391 ) | ( n6390 & ~n6391 ) ;
  assign n6393 = ( n6316 & n6367 ) | ( n6316 & n6392 ) | ( n6367 & n6392 ) ;
  assign n6394 = ( n6316 & n6367 ) | ( n6316 & ~n6392 ) | ( n6367 & ~n6392 ) ;
  assign n6395 = ( n6392 & ~n6393 ) | ( n6392 & n6394 ) | ( ~n6393 & n6394 ) ;
  assign n6396 = ( n6369 & n6378 ) | ( n6369 & n6395 ) | ( n6378 & n6395 ) ;
  assign n6397 = ( ~n6369 & n6378 ) | ( ~n6369 & n6395 ) | ( n6378 & n6395 ) ;
  assign n6398 = ( n6369 & ~n6396 ) | ( n6369 & n6397 ) | ( ~n6396 & n6397 ) ;
  assign n6399 = x42 & x43 ;
  assign n6400 = x23 & x62 ;
  assign n6401 = ( x43 & n6399 ) | ( x43 & n6400 ) | ( n6399 & n6400 ) ;
  assign n6402 = ( x43 & ~n6399 ) | ( x43 & n6400 ) | ( ~n6399 & n6400 ) ;
  assign n6403 = ( n6399 & ~n6401 ) | ( n6399 & n6402 ) | ( ~n6401 & n6402 ) ;
  assign n6404 = x29 & x56 ;
  assign n6405 = x30 & x55 ;
  assign n6406 = x31 & x54 ;
  assign n6407 = ( ~n6404 & n6405 ) | ( ~n6404 & n6406 ) | ( n6405 & n6406 ) ;
  assign n6408 = ( n6404 & n6405 ) | ( n6404 & n6406 ) | ( n6405 & n6406 ) ;
  assign n6409 = ( n6404 & n6407 ) | ( n6404 & ~n6408 ) | ( n6407 & ~n6408 ) ;
  assign n6410 = x36 & x49 ;
  assign n6411 = x37 & x48 ;
  assign n6412 = x38 & x47 ;
  assign n6413 = ( ~n6410 & n6411 ) | ( ~n6410 & n6412 ) | ( n6411 & n6412 ) ;
  assign n6414 = ( n6410 & n6411 ) | ( n6410 & n6412 ) | ( n6411 & n6412 ) ;
  assign n6415 = ( n6410 & n6413 ) | ( n6410 & ~n6414 ) | ( n6413 & ~n6414 ) ;
  assign n6416 = ( n6403 & n6409 ) | ( n6403 & n6415 ) | ( n6409 & n6415 ) ;
  assign n6417 = ( ~n6403 & n6409 ) | ( ~n6403 & n6415 ) | ( n6409 & n6415 ) ;
  assign n6418 = ( n6403 & ~n6416 ) | ( n6403 & n6417 ) | ( ~n6416 & n6417 ) ;
  assign n6419 = x39 & x46 ;
  assign n6420 = x41 & x44 ;
  assign n6421 = x40 & x45 ;
  assign n6422 = ( ~n6419 & n6420 ) | ( ~n6419 & n6421 ) | ( n6420 & n6421 ) ;
  assign n6423 = ( n6419 & n6420 ) | ( n6419 & n6421 ) | ( n6420 & n6421 ) ;
  assign n6424 = ( n6419 & n6422 ) | ( n6419 & ~n6423 ) | ( n6422 & ~n6423 ) ;
  assign n6425 = x22 & x63 ;
  assign n6426 = x35 & x50 ;
  assign n6427 = x28 & x57 ;
  assign n6428 = ( ~n6425 & n6426 ) | ( ~n6425 & n6427 ) | ( n6426 & n6427 ) ;
  assign n6429 = ( n6425 & n6426 ) | ( n6425 & n6427 ) | ( n6426 & n6427 ) ;
  assign n6430 = ( n6425 & n6428 ) | ( n6425 & ~n6429 ) | ( n6428 & ~n6429 ) ;
  assign n6431 = x32 & x53 ;
  assign n6432 = x33 & x52 ;
  assign n6433 = x34 & x51 ;
  assign n6434 = ( ~n6431 & n6432 ) | ( ~n6431 & n6433 ) | ( n6432 & n6433 ) ;
  assign n6435 = ( n6431 & n6432 ) | ( n6431 & n6433 ) | ( n6432 & n6433 ) ;
  assign n6436 = ( n6431 & n6434 ) | ( n6431 & ~n6435 ) | ( n6434 & ~n6435 ) ;
  assign n6437 = ( ~n6424 & n6430 ) | ( ~n6424 & n6436 ) | ( n6430 & n6436 ) ;
  assign n6438 = ( n6424 & n6430 ) | ( n6424 & n6436 ) | ( n6430 & n6436 ) ;
  assign n6439 = ( n6424 & n6437 ) | ( n6424 & ~n6438 ) | ( n6437 & ~n6438 ) ;
  assign n6440 = ( n6376 & n6418 ) | ( n6376 & n6439 ) | ( n6418 & n6439 ) ;
  assign n6441 = ( ~n6376 & n6418 ) | ( ~n6376 & n6439 ) | ( n6418 & n6439 ) ;
  assign n6442 = ( n6376 & ~n6440 ) | ( n6376 & n6441 ) | ( ~n6440 & n6441 ) ;
  assign n6443 = ( ~n6328 & n6334 ) | ( ~n6328 & n6340 ) | ( n6334 & n6340 ) ;
  assign n6444 = ( n6328 & n6334 ) | ( n6328 & n6340 ) | ( n6334 & n6340 ) ;
  assign n6445 = ( n6328 & n6443 ) | ( n6328 & ~n6444 ) | ( n6443 & ~n6444 ) ;
  assign n6446 = ( n6343 & n6364 ) | ( n6343 & n6445 ) | ( n6364 & n6445 ) ;
  assign n6447 = ( ~n6343 & n6364 ) | ( ~n6343 & n6445 ) | ( n6364 & n6445 ) ;
  assign n6448 = ( n6343 & ~n6446 ) | ( n6343 & n6447 ) | ( ~n6446 & n6447 ) ;
  assign n6449 = x24 & x61 ;
  assign n6450 = ( ~n6355 & n6361 ) | ( ~n6355 & n6449 ) | ( n6361 & n6449 ) ;
  assign n6451 = ( n6355 & n6361 ) | ( n6355 & n6449 ) | ( n6361 & n6449 ) ;
  assign n6452 = ( n6355 & n6450 ) | ( n6355 & ~n6451 ) | ( n6450 & ~n6451 ) ;
  assign n6453 = x25 & x60 ;
  assign n6454 = x26 & x59 ;
  assign n6455 = x27 & x58 ;
  assign n6456 = ( ~n6453 & n6454 ) | ( ~n6453 & n6455 ) | ( n6454 & n6455 ) ;
  assign n6457 = ( n6453 & n6454 ) | ( n6453 & n6455 ) | ( n6454 & n6455 ) ;
  assign n6458 = ( n6453 & n6456 ) | ( n6453 & ~n6457 ) | ( n6456 & ~n6457 ) ;
  assign n6459 = ( ~n6310 & n6349 ) | ( ~n6310 & n6458 ) | ( n6349 & n6458 ) ;
  assign n6460 = ( n6310 & n6349 ) | ( n6310 & n6458 ) | ( n6349 & n6458 ) ;
  assign n6461 = ( n6310 & n6459 ) | ( n6310 & ~n6460 ) | ( n6459 & ~n6460 ) ;
  assign n6462 = ( n6322 & n6452 ) | ( n6322 & n6461 ) | ( n6452 & n6461 ) ;
  assign n6463 = ( ~n6322 & n6452 ) | ( ~n6322 & n6461 ) | ( n6452 & n6461 ) ;
  assign n6464 = ( n6322 & ~n6462 ) | ( n6322 & n6463 ) | ( ~n6462 & n6463 ) ;
  assign n6465 = ( ~n6442 & n6448 ) | ( ~n6442 & n6464 ) | ( n6448 & n6464 ) ;
  assign n6466 = ( n6442 & n6448 ) | ( n6442 & n6464 ) | ( n6448 & n6464 ) ;
  assign n6467 = ( n6442 & n6465 ) | ( n6442 & ~n6466 ) | ( n6465 & ~n6466 ) ;
  assign n6468 = ( n6381 & n6398 ) | ( n6381 & n6467 ) | ( n6398 & n6467 ) ;
  assign n6469 = ( ~n6381 & n6398 ) | ( ~n6381 & n6467 ) | ( n6398 & n6467 ) ;
  assign n6470 = ( n6381 & ~n6468 ) | ( n6381 & n6469 ) | ( ~n6468 & n6469 ) ;
  assign n6471 = ( ~n6385 & n6387 ) | ( ~n6385 & n6470 ) | ( n6387 & n6470 ) ;
  assign n6472 = ( n6385 & n6387 ) | ( n6385 & n6470 ) | ( n6387 & n6470 ) ;
  assign n6473 = ( n6385 & n6471 ) | ( n6385 & ~n6472 ) | ( n6471 & ~n6472 ) ;
  assign n6474 = x25 & x61 ;
  assign n6475 = x24 & x62 ;
  assign n6476 = ( ~n6401 & n6474 ) | ( ~n6401 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6477 = ( n6401 & n6474 ) | ( n6401 & n6475 ) | ( n6474 & n6475 ) ;
  assign n6478 = ( n6401 & n6476 ) | ( n6401 & ~n6477 ) | ( n6476 & ~n6477 ) ;
  assign n6479 = ( n6444 & n6451 ) | ( n6444 & n6478 ) | ( n6451 & n6478 ) ;
  assign n6480 = ( n6444 & ~n6451 ) | ( n6444 & n6478 ) | ( ~n6451 & n6478 ) ;
  assign n6481 = ( n6451 & ~n6479 ) | ( n6451 & n6480 ) | ( ~n6479 & n6480 ) ;
  assign n6482 = ( ~n6440 & n6462 ) | ( ~n6440 & n6481 ) | ( n6462 & n6481 ) ;
  assign n6483 = ( n6440 & n6462 ) | ( n6440 & n6481 ) | ( n6462 & n6481 ) ;
  assign n6484 = ( n6440 & n6482 ) | ( n6440 & ~n6483 ) | ( n6482 & ~n6483 ) ;
  assign n6485 = ( ~n6393 & n6466 ) | ( ~n6393 & n6484 ) | ( n6466 & n6484 ) ;
  assign n6486 = ( n6393 & n6466 ) | ( n6393 & n6484 ) | ( n6466 & n6484 ) ;
  assign n6487 = ( n6393 & n6485 ) | ( n6393 & ~n6486 ) | ( n6485 & ~n6486 ) ;
  assign n6488 = ( ~n6408 & n6414 ) | ( ~n6408 & n6423 ) | ( n6414 & n6423 ) ;
  assign n6489 = ( n6408 & n6414 ) | ( n6408 & n6423 ) | ( n6414 & n6423 ) ;
  assign n6490 = ( n6408 & n6488 ) | ( n6408 & ~n6489 ) | ( n6488 & ~n6489 ) ;
  assign n6491 = ( n6429 & ~n6435 ) | ( n6429 & n6457 ) | ( ~n6435 & n6457 ) ;
  assign n6492 = ( n6429 & n6435 ) | ( n6429 & n6457 ) | ( n6435 & n6457 ) ;
  assign n6493 = ( n6435 & n6491 ) | ( n6435 & ~n6492 ) | ( n6491 & ~n6492 ) ;
  assign n6494 = ( n6391 & n6490 ) | ( n6391 & n6493 ) | ( n6490 & n6493 ) ;
  assign n6495 = ( ~n6391 & n6490 ) | ( ~n6391 & n6493 ) | ( n6490 & n6493 ) ;
  assign n6496 = ( n6391 & ~n6494 ) | ( n6391 & n6495 ) | ( ~n6494 & n6495 ) ;
  assign n6497 = ( n6416 & n6438 ) | ( n6416 & ~n6460 ) | ( n6438 & ~n6460 ) ;
  assign n6498 = ( n6416 & n6438 ) | ( n6416 & n6460 ) | ( n6438 & n6460 ) ;
  assign n6499 = ( n6460 & n6497 ) | ( n6460 & ~n6498 ) | ( n6497 & ~n6498 ) ;
  assign n6500 = x23 & x63 ;
  assign n6501 = x36 & x50 ;
  assign n6502 = x37 & x49 ;
  assign n6503 = ( ~n6500 & n6501 ) | ( ~n6500 & n6502 ) | ( n6501 & n6502 ) ;
  assign n6504 = ( n6500 & n6501 ) | ( n6500 & n6502 ) | ( n6501 & n6502 ) ;
  assign n6505 = ( n6500 & n6503 ) | ( n6500 & ~n6504 ) | ( n6503 & ~n6504 ) ;
  assign n6506 = x38 & x48 ;
  assign n6507 = x31 & x55 ;
  assign n6508 = x29 & x57 ;
  assign n6509 = ( ~n6506 & n6507 ) | ( ~n6506 & n6508 ) | ( n6507 & n6508 ) ;
  assign n6510 = ( n6506 & n6507 ) | ( n6506 & n6508 ) | ( n6507 & n6508 ) ;
  assign n6511 = ( n6506 & n6509 ) | ( n6506 & ~n6510 ) | ( n6509 & ~n6510 ) ;
  assign n6512 = x33 & x53 ;
  assign n6513 = x34 & x52 ;
  assign n6514 = x35 & x51 ;
  assign n6515 = ( ~n6512 & n6513 ) | ( ~n6512 & n6514 ) | ( n6513 & n6514 ) ;
  assign n6516 = ( n6512 & n6513 ) | ( n6512 & n6514 ) | ( n6513 & n6514 ) ;
  assign n6517 = ( n6512 & n6515 ) | ( n6512 & ~n6516 ) | ( n6515 & ~n6516 ) ;
  assign n6518 = ( ~n6505 & n6511 ) | ( ~n6505 & n6517 ) | ( n6511 & n6517 ) ;
  assign n6519 = ( n6505 & n6511 ) | ( n6505 & n6517 ) | ( n6511 & n6517 ) ;
  assign n6520 = ( n6505 & n6518 ) | ( n6505 & ~n6519 ) | ( n6518 & ~n6519 ) ;
  assign n6521 = x26 & x60 ;
  assign n6522 = x27 & x59 ;
  assign n6523 = x28 & x58 ;
  assign n6524 = ( ~n6521 & n6522 ) | ( ~n6521 & n6523 ) | ( n6522 & n6523 ) ;
  assign n6525 = ( n6521 & n6522 ) | ( n6521 & n6523 ) | ( n6522 & n6523 ) ;
  assign n6526 = ( n6521 & n6524 ) | ( n6521 & ~n6525 ) | ( n6524 & ~n6525 ) ;
  assign n6527 = x30 & x56 ;
  assign n6528 = x40 & x46 ;
  assign n6529 = x39 & x47 ;
  assign n6530 = ( ~n6527 & n6528 ) | ( ~n6527 & n6529 ) | ( n6528 & n6529 ) ;
  assign n6531 = ( n6527 & n6528 ) | ( n6527 & n6529 ) | ( n6528 & n6529 ) ;
  assign n6532 = ( n6527 & n6530 ) | ( n6527 & ~n6531 ) | ( n6530 & ~n6531 ) ;
  assign n6533 = x41 & x45 ;
  assign n6534 = x42 & x44 ;
  assign n6535 = x32 & x54 ;
  assign n6536 = ( ~n6533 & n6534 ) | ( ~n6533 & n6535 ) | ( n6534 & n6535 ) ;
  assign n6537 = ( n6533 & n6534 ) | ( n6533 & n6535 ) | ( n6534 & n6535 ) ;
  assign n6538 = ( n6533 & n6536 ) | ( n6533 & ~n6537 ) | ( n6536 & ~n6537 ) ;
  assign n6539 = ( ~n6526 & n6532 ) | ( ~n6526 & n6538 ) | ( n6532 & n6538 ) ;
  assign n6540 = ( n6526 & n6532 ) | ( n6526 & n6538 ) | ( n6532 & n6538 ) ;
  assign n6541 = ( n6526 & n6539 ) | ( n6526 & ~n6540 ) | ( n6539 & ~n6540 ) ;
  assign n6542 = ( n6446 & n6520 ) | ( n6446 & n6541 ) | ( n6520 & n6541 ) ;
  assign n6543 = ( ~n6446 & n6520 ) | ( ~n6446 & n6541 ) | ( n6520 & n6541 ) ;
  assign n6544 = ( n6446 & ~n6542 ) | ( n6446 & n6543 ) | ( ~n6542 & n6543 ) ;
  assign n6545 = ( n6496 & n6499 ) | ( n6496 & n6544 ) | ( n6499 & n6544 ) ;
  assign n6546 = ( ~n6496 & n6499 ) | ( ~n6496 & n6544 ) | ( n6499 & n6544 ) ;
  assign n6547 = ( n6496 & ~n6545 ) | ( n6496 & n6546 ) | ( ~n6545 & n6546 ) ;
  assign n6548 = ( ~n6396 & n6487 ) | ( ~n6396 & n6547 ) | ( n6487 & n6547 ) ;
  assign n6549 = ( n6396 & n6487 ) | ( n6396 & n6547 ) | ( n6487 & n6547 ) ;
  assign n6550 = ( n6396 & n6548 ) | ( n6396 & ~n6549 ) | ( n6548 & ~n6549 ) ;
  assign n6551 = ( ~n6468 & n6472 ) | ( ~n6468 & n6550 ) | ( n6472 & n6550 ) ;
  assign n6552 = ( n6468 & n6472 ) | ( n6468 & n6550 ) | ( n6472 & n6550 ) ;
  assign n6553 = ( n6468 & n6551 ) | ( n6468 & ~n6552 ) | ( n6551 & ~n6552 ) ;
  assign n6554 = ( ~n6489 & n6519 ) | ( ~n6489 & n6540 ) | ( n6519 & n6540 ) ;
  assign n6555 = ( n6489 & n6519 ) | ( n6489 & n6540 ) | ( n6519 & n6540 ) ;
  assign n6556 = ( n6489 & n6554 ) | ( n6489 & ~n6555 ) | ( n6554 & ~n6555 ) ;
  assign n6557 = ( ~n6483 & n6542 ) | ( ~n6483 & n6556 ) | ( n6542 & n6556 ) ;
  assign n6558 = ( n6483 & n6542 ) | ( n6483 & n6556 ) | ( n6542 & n6556 ) ;
  assign n6559 = ( n6483 & n6557 ) | ( n6483 & ~n6558 ) | ( n6557 & ~n6558 ) ;
  assign n6560 = x40 & x47 ;
  assign n6561 = x31 & x56 ;
  assign n6562 = x33 & x54 ;
  assign n6563 = ( ~n6560 & n6561 ) | ( ~n6560 & n6562 ) | ( n6561 & n6562 ) ;
  assign n6564 = ( n6560 & n6561 ) | ( n6560 & n6562 ) | ( n6561 & n6562 ) ;
  assign n6565 = ( n6560 & n6563 ) | ( n6560 & ~n6564 ) | ( n6563 & ~n6564 ) ;
  assign n6566 = x43 & x44 ;
  assign n6567 = x25 & x62 ;
  assign n6568 = ( x44 & n6566 ) | ( x44 & n6567 ) | ( n6566 & n6567 ) ;
  assign n6569 = ( x44 & ~n6566 ) | ( x44 & n6567 ) | ( ~n6566 & n6567 ) ;
  assign n6570 = ( n6566 & ~n6568 ) | ( n6566 & n6569 ) | ( ~n6568 & n6569 ) ;
  assign n6571 = ( ~n6492 & n6565 ) | ( ~n6492 & n6570 ) | ( n6565 & n6570 ) ;
  assign n6572 = ( n6492 & n6565 ) | ( n6492 & n6570 ) | ( n6565 & n6570 ) ;
  assign n6573 = ( n6492 & n6571 ) | ( n6492 & ~n6572 ) | ( n6571 & ~n6572 ) ;
  assign n6574 = x32 & x55 ;
  assign n6575 = x41 & x46 ;
  assign n6576 = x42 & x45 ;
  assign n6577 = ( ~n6574 & n6575 ) | ( ~n6574 & n6576 ) | ( n6575 & n6576 ) ;
  assign n6578 = ( n6574 & n6575 ) | ( n6574 & n6576 ) | ( n6575 & n6576 ) ;
  assign n6579 = ( n6574 & n6577 ) | ( n6574 & ~n6578 ) | ( n6577 & ~n6578 ) ;
  assign n6580 = x37 & x50 ;
  assign n6581 = x38 & x49 ;
  assign n6582 = x39 & x48 ;
  assign n6583 = ( ~n6580 & n6581 ) | ( ~n6580 & n6582 ) | ( n6581 & n6582 ) ;
  assign n6584 = ( n6580 & n6581 ) | ( n6580 & n6582 ) | ( n6581 & n6582 ) ;
  assign n6585 = ( n6580 & n6583 ) | ( n6580 & ~n6584 ) | ( n6583 & ~n6584 ) ;
  assign n6586 = x24 & x63 ;
  assign n6587 = x26 & x61 ;
  assign n6588 = x27 & x60 ;
  assign n6589 = ( ~n6586 & n6587 ) | ( ~n6586 & n6588 ) | ( n6587 & n6588 ) ;
  assign n6590 = ( n6586 & n6587 ) | ( n6586 & n6588 ) | ( n6587 & n6588 ) ;
  assign n6591 = ( n6586 & n6589 ) | ( n6586 & ~n6590 ) | ( n6589 & ~n6590 ) ;
  assign n6592 = ( ~n6579 & n6585 ) | ( ~n6579 & n6591 ) | ( n6585 & n6591 ) ;
  assign n6593 = ( n6579 & n6585 ) | ( n6579 & n6591 ) | ( n6585 & n6591 ) ;
  assign n6594 = ( n6579 & n6592 ) | ( n6579 & ~n6593 ) | ( n6592 & ~n6593 ) ;
  assign n6595 = x30 & x57 ;
  assign n6596 = x28 & x59 ;
  assign n6597 = x34 & x53 ;
  assign n6598 = ( ~n6595 & n6596 ) | ( ~n6595 & n6597 ) | ( n6596 & n6597 ) ;
  assign n6599 = ( n6595 & n6596 ) | ( n6595 & n6597 ) | ( n6596 & n6597 ) ;
  assign n6600 = ( n6595 & n6598 ) | ( n6595 & ~n6599 ) | ( n6598 & ~n6599 ) ;
  assign n6601 = x35 & x52 ;
  assign n6602 = x29 & x58 ;
  assign n6603 = x36 & x51 ;
  assign n6604 = ( ~n6601 & n6602 ) | ( ~n6601 & n6603 ) | ( n6602 & n6603 ) ;
  assign n6605 = ( n6601 & n6602 ) | ( n6601 & n6603 ) | ( n6602 & n6603 ) ;
  assign n6606 = ( n6601 & n6604 ) | ( n6601 & ~n6605 ) | ( n6604 & ~n6605 ) ;
  assign n6607 = ( n6477 & n6600 ) | ( n6477 & n6606 ) | ( n6600 & n6606 ) ;
  assign n6608 = ( ~n6477 & n6600 ) | ( ~n6477 & n6606 ) | ( n6600 & n6606 ) ;
  assign n6609 = ( n6477 & ~n6607 ) | ( n6477 & n6608 ) | ( ~n6607 & n6608 ) ;
  assign n6610 = ( ~n6573 & n6594 ) | ( ~n6573 & n6609 ) | ( n6594 & n6609 ) ;
  assign n6611 = ( n6573 & n6594 ) | ( n6573 & n6609 ) | ( n6594 & n6609 ) ;
  assign n6612 = ( n6573 & n6610 ) | ( n6573 & ~n6611 ) | ( n6610 & ~n6611 ) ;
  assign n6613 = ( n6510 & ~n6531 ) | ( n6510 & n6537 ) | ( ~n6531 & n6537 ) ;
  assign n6614 = ( n6510 & n6531 ) | ( n6510 & n6537 ) | ( n6531 & n6537 ) ;
  assign n6615 = ( n6531 & n6613 ) | ( n6531 & ~n6614 ) | ( n6613 & ~n6614 ) ;
  assign n6616 = ( n6504 & ~n6516 ) | ( n6504 & n6525 ) | ( ~n6516 & n6525 ) ;
  assign n6617 = ( n6504 & n6516 ) | ( n6504 & n6525 ) | ( n6516 & n6525 ) ;
  assign n6618 = ( n6516 & n6616 ) | ( n6516 & ~n6617 ) | ( n6616 & ~n6617 ) ;
  assign n6619 = ( ~n6479 & n6615 ) | ( ~n6479 & n6618 ) | ( n6615 & n6618 ) ;
  assign n6620 = ( n6479 & n6615 ) | ( n6479 & n6618 ) | ( n6615 & n6618 ) ;
  assign n6621 = ( n6479 & n6619 ) | ( n6479 & ~n6620 ) | ( n6619 & ~n6620 ) ;
  assign n6622 = ( ~n6494 & n6498 ) | ( ~n6494 & n6621 ) | ( n6498 & n6621 ) ;
  assign n6623 = ( n6494 & n6498 ) | ( n6494 & n6621 ) | ( n6498 & n6621 ) ;
  assign n6624 = ( n6494 & n6622 ) | ( n6494 & ~n6623 ) | ( n6622 & ~n6623 ) ;
  assign n6625 = ( ~n6545 & n6612 ) | ( ~n6545 & n6624 ) | ( n6612 & n6624 ) ;
  assign n6626 = ( n6545 & n6612 ) | ( n6545 & n6624 ) | ( n6612 & n6624 ) ;
  assign n6627 = ( n6545 & n6625 ) | ( n6545 & ~n6626 ) | ( n6625 & ~n6626 ) ;
  assign n6628 = ( ~n6486 & n6559 ) | ( ~n6486 & n6627 ) | ( n6559 & n6627 ) ;
  assign n6629 = ( n6486 & n6559 ) | ( n6486 & n6627 ) | ( n6559 & n6627 ) ;
  assign n6630 = ( n6486 & n6628 ) | ( n6486 & ~n6629 ) | ( n6628 & ~n6629 ) ;
  assign n6631 = ( ~n6549 & n6552 ) | ( ~n6549 & n6630 ) | ( n6552 & n6630 ) ;
  assign n6632 = ( n6549 & n6552 ) | ( n6549 & n6630 ) | ( n6552 & n6630 ) ;
  assign n6633 = ( n6549 & n6631 ) | ( n6549 & ~n6632 ) | ( n6631 & ~n6632 ) ;
  assign n6634 = ( n6593 & ~n6607 ) | ( n6593 & n6617 ) | ( ~n6607 & n6617 ) ;
  assign n6635 = ( n6593 & n6607 ) | ( n6593 & n6617 ) | ( n6607 & n6617 ) ;
  assign n6636 = ( n6607 & n6634 ) | ( n6607 & ~n6635 ) | ( n6634 & ~n6635 ) ;
  assign n6637 = ( ~n6611 & n6623 ) | ( ~n6611 & n6636 ) | ( n6623 & n6636 ) ;
  assign n6638 = ( n6611 & n6623 ) | ( n6611 & n6636 ) | ( n6623 & n6636 ) ;
  assign n6639 = ( n6611 & n6637 ) | ( n6611 & ~n6638 ) | ( n6637 & ~n6638 ) ;
  assign n6640 = ( n6584 & ~n6590 ) | ( n6584 & n6599 ) | ( ~n6590 & n6599 ) ;
  assign n6641 = ( n6584 & n6590 ) | ( n6584 & n6599 ) | ( n6590 & n6599 ) ;
  assign n6642 = ( n6590 & n6640 ) | ( n6590 & ~n6641 ) | ( n6640 & ~n6641 ) ;
  assign n6643 = x43 & x45 ;
  assign n6644 = x33 & x55 ;
  assign n6645 = x34 & x54 ;
  assign n6646 = ( ~n6643 & n6644 ) | ( ~n6643 & n6645 ) | ( n6644 & n6645 ) ;
  assign n6647 = ( n6643 & n6644 ) | ( n6643 & n6645 ) | ( n6644 & n6645 ) ;
  assign n6648 = ( n6643 & n6646 ) | ( n6643 & ~n6647 ) | ( n6646 & ~n6647 ) ;
  assign n6649 = ( ~n6564 & n6605 ) | ( ~n6564 & n6648 ) | ( n6605 & n6648 ) ;
  assign n6650 = ( n6564 & n6605 ) | ( n6564 & n6648 ) | ( n6605 & n6648 ) ;
  assign n6651 = ( n6564 & n6649 ) | ( n6564 & ~n6650 ) | ( n6649 & ~n6650 ) ;
  assign n6652 = ( ~n6572 & n6642 ) | ( ~n6572 & n6651 ) | ( n6642 & n6651 ) ;
  assign n6653 = ( n6572 & n6642 ) | ( n6572 & n6651 ) | ( n6642 & n6651 ) ;
  assign n6654 = ( n6572 & n6652 ) | ( n6572 & ~n6653 ) | ( n6652 & ~n6653 ) ;
  assign n6655 = ( ~n6555 & n6620 ) | ( ~n6555 & n6654 ) | ( n6620 & n6654 ) ;
  assign n6656 = ( n6555 & n6620 ) | ( n6555 & n6654 ) | ( n6620 & n6654 ) ;
  assign n6657 = ( n6555 & n6655 ) | ( n6555 & ~n6656 ) | ( n6655 & ~n6656 ) ;
  assign n6658 = x40 & x48 ;
  assign n6659 = x32 & x56 ;
  assign n6660 = ( ~n3591 & n6658 ) | ( ~n3591 & n6659 ) | ( n6658 & n6659 ) ;
  assign n6661 = ( n3591 & n6658 ) | ( n3591 & n6659 ) | ( n6658 & n6659 ) ;
  assign n6662 = ( n3591 & n6660 ) | ( n3591 & ~n6661 ) | ( n6660 & ~n6661 ) ;
  assign n6663 = x29 & x59 ;
  assign n6664 = x39 & x49 ;
  assign n6665 = x38 & x50 ;
  assign n6666 = ( ~n6663 & n6664 ) | ( ~n6663 & n6665 ) | ( n6664 & n6665 ) ;
  assign n6667 = ( n6663 & n6664 ) | ( n6663 & n6665 ) | ( n6664 & n6665 ) ;
  assign n6668 = ( n6663 & n6666 ) | ( n6663 & ~n6667 ) | ( n6666 & ~n6667 ) ;
  assign n6669 = ( n6614 & n6662 ) | ( n6614 & n6668 ) | ( n6662 & n6668 ) ;
  assign n6670 = ( ~n6614 & n6662 ) | ( ~n6614 & n6668 ) | ( n6662 & n6668 ) ;
  assign n6671 = ( n6614 & ~n6669 ) | ( n6614 & n6670 ) | ( ~n6669 & n6670 ) ;
  assign n6672 = x25 & x63 ;
  assign n6673 = ( n6568 & n6578 ) | ( n6568 & n6672 ) | ( n6578 & n6672 ) ;
  assign n6674 = ( n6568 & ~n6578 ) | ( n6568 & n6672 ) | ( ~n6578 & n6672 ) ;
  assign n6675 = ( n6578 & ~n6673 ) | ( n6578 & n6674 ) | ( ~n6673 & n6674 ) ;
  assign n6676 = x35 & x53 ;
  assign n6677 = x37 & x51 ;
  assign n6678 = x36 & x52 ;
  assign n6679 = ( ~n6676 & n6677 ) | ( ~n6676 & n6678 ) | ( n6677 & n6678 ) ;
  assign n6680 = ( n6676 & n6677 ) | ( n6676 & n6678 ) | ( n6677 & n6678 ) ;
  assign n6681 = ( n6676 & n6679 ) | ( n6676 & ~n6680 ) | ( n6679 & ~n6680 ) ;
  assign n6682 = x31 & x57 ;
  assign n6683 = x42 & x46 ;
  assign n6684 = x41 & x47 ;
  assign n6685 = ( ~n6682 & n6683 ) | ( ~n6682 & n6684 ) | ( n6683 & n6684 ) ;
  assign n6686 = ( n6682 & n6683 ) | ( n6682 & n6684 ) | ( n6683 & n6684 ) ;
  assign n6687 = ( n6682 & n6685 ) | ( n6682 & ~n6686 ) | ( n6685 & ~n6686 ) ;
  assign n6688 = x26 & x62 ;
  assign n6689 = x27 & x61 ;
  assign n6690 = x28 & x60 ;
  assign n6691 = ( ~n6688 & n6689 ) | ( ~n6688 & n6690 ) | ( n6689 & n6690 ) ;
  assign n6692 = ( n6688 & n6689 ) | ( n6688 & n6690 ) | ( n6689 & n6690 ) ;
  assign n6693 = ( n6688 & n6691 ) | ( n6688 & ~n6692 ) | ( n6691 & ~n6692 ) ;
  assign n6694 = ( ~n6681 & n6687 ) | ( ~n6681 & n6693 ) | ( n6687 & n6693 ) ;
  assign n6695 = ( n6681 & n6687 ) | ( n6681 & n6693 ) | ( n6687 & n6693 ) ;
  assign n6696 = ( n6681 & n6694 ) | ( n6681 & ~n6695 ) | ( n6694 & ~n6695 ) ;
  assign n6697 = ( ~n6671 & n6675 ) | ( ~n6671 & n6696 ) | ( n6675 & n6696 ) ;
  assign n6698 = ( n6671 & n6675 ) | ( n6671 & n6696 ) | ( n6675 & n6696 ) ;
  assign n6699 = ( n6671 & n6697 ) | ( n6671 & ~n6698 ) | ( n6697 & ~n6698 ) ;
  assign n6700 = ( ~n6558 & n6657 ) | ( ~n6558 & n6699 ) | ( n6657 & n6699 ) ;
  assign n6701 = ( n6558 & n6657 ) | ( n6558 & n6699 ) | ( n6657 & n6699 ) ;
  assign n6702 = ( n6558 & n6700 ) | ( n6558 & ~n6701 ) | ( n6700 & ~n6701 ) ;
  assign n6703 = ( ~n6626 & n6639 ) | ( ~n6626 & n6702 ) | ( n6639 & n6702 ) ;
  assign n6704 = ( n6626 & n6639 ) | ( n6626 & n6702 ) | ( n6639 & n6702 ) ;
  assign n6705 = ( n6626 & n6703 ) | ( n6626 & ~n6704 ) | ( n6703 & ~n6704 ) ;
  assign n6706 = ( ~n6629 & n6632 ) | ( ~n6629 & n6705 ) | ( n6632 & n6705 ) ;
  assign n6707 = ( n6629 & n6632 ) | ( n6629 & n6705 ) | ( n6632 & n6705 ) ;
  assign n6708 = ( n6629 & n6706 ) | ( n6629 & ~n6707 ) | ( n6706 & ~n6707 ) ;
  assign n6709 = ( n6641 & ~n6650 ) | ( n6641 & n6673 ) | ( ~n6650 & n6673 ) ;
  assign n6710 = ( n6641 & n6650 ) | ( n6641 & n6673 ) | ( n6650 & n6673 ) ;
  assign n6711 = ( n6650 & n6709 ) | ( n6650 & ~n6710 ) | ( n6709 & ~n6710 ) ;
  assign n6712 = ( ~n6635 & n6653 ) | ( ~n6635 & n6711 ) | ( n6653 & n6711 ) ;
  assign n6713 = ( n6635 & n6653 ) | ( n6635 & n6711 ) | ( n6653 & n6711 ) ;
  assign n6714 = ( n6635 & n6712 ) | ( n6635 & ~n6713 ) | ( n6712 & ~n6713 ) ;
  assign n6715 = ( n6661 & n6680 ) | ( n6661 & n6692 ) | ( n6680 & n6692 ) ;
  assign n6716 = ( ~n6661 & n6680 ) | ( ~n6661 & n6692 ) | ( n6680 & n6692 ) ;
  assign n6717 = ( n6661 & ~n6715 ) | ( n6661 & n6716 ) | ( ~n6715 & n6716 ) ;
  assign n6718 = x30 & x59 ;
  assign n6719 = x32 & x57 ;
  assign n6720 = x31 & x58 ;
  assign n6721 = ( ~n6718 & n6719 ) | ( ~n6718 & n6720 ) | ( n6719 & n6720 ) ;
  assign n6722 = ( n6718 & n6719 ) | ( n6718 & n6720 ) | ( n6719 & n6720 ) ;
  assign n6723 = ( n6718 & n6721 ) | ( n6718 & ~n6722 ) | ( n6721 & ~n6722 ) ;
  assign n6724 = x36 & x53 ;
  assign n6725 = x37 & x52 ;
  assign n6726 = x38 & x51 ;
  assign n6727 = ( ~n6724 & n6725 ) | ( ~n6724 & n6726 ) | ( n6725 & n6726 ) ;
  assign n6728 = ( n6724 & n6725 ) | ( n6724 & n6726 ) | ( n6725 & n6726 ) ;
  assign n6729 = ( n6724 & n6727 ) | ( n6724 & ~n6728 ) | ( n6727 & ~n6728 ) ;
  assign n6730 = x41 & x48 ;
  assign n6731 = x33 & x56 ;
  assign n6732 = x35 & x54 ;
  assign n6733 = ( ~n6730 & n6731 ) | ( ~n6730 & n6732 ) | ( n6731 & n6732 ) ;
  assign n6734 = ( n6730 & n6731 ) | ( n6730 & n6732 ) | ( n6731 & n6732 ) ;
  assign n6735 = ( n6730 & n6733 ) | ( n6730 & ~n6734 ) | ( n6733 & ~n6734 ) ;
  assign n6736 = ( ~n6723 & n6729 ) | ( ~n6723 & n6735 ) | ( n6729 & n6735 ) ;
  assign n6737 = ( n6723 & n6729 ) | ( n6723 & n6735 ) | ( n6729 & n6735 ) ;
  assign n6738 = ( n6723 & n6736 ) | ( n6723 & ~n6737 ) | ( n6736 & ~n6737 ) ;
  assign n6739 = x28 & x61 ;
  assign n6740 = x29 & x60 ;
  assign n6741 = ( n6647 & n6739 ) | ( n6647 & n6740 ) | ( n6739 & n6740 ) ;
  assign n6742 = ( ~n6647 & n6739 ) | ( ~n6647 & n6740 ) | ( n6739 & n6740 ) ;
  assign n6743 = ( n6647 & ~n6741 ) | ( n6647 & n6742 ) | ( ~n6741 & n6742 ) ;
  assign n6744 = x34 & x55 ;
  assign n6745 = x42 & x47 ;
  assign n6746 = x43 & x46 ;
  assign n6747 = ( ~n6744 & n6745 ) | ( ~n6744 & n6746 ) | ( n6745 & n6746 ) ;
  assign n6748 = ( n6744 & n6745 ) | ( n6744 & n6746 ) | ( n6745 & n6746 ) ;
  assign n6749 = ( n6744 & n6747 ) | ( n6744 & ~n6748 ) | ( n6747 & ~n6748 ) ;
  assign n6750 = x44 & x45 ;
  assign n6751 = x27 & x62 ;
  assign n6752 = ( x45 & n6750 ) | ( x45 & n6751 ) | ( n6750 & n6751 ) ;
  assign n6753 = ( x45 & ~n6750 ) | ( x45 & n6751 ) | ( ~n6750 & n6751 ) ;
  assign n6754 = ( n6750 & ~n6752 ) | ( n6750 & n6753 ) | ( ~n6752 & n6753 ) ;
  assign n6755 = ( ~n6743 & n6749 ) | ( ~n6743 & n6754 ) | ( n6749 & n6754 ) ;
  assign n6756 = ( n6743 & n6749 ) | ( n6743 & n6754 ) | ( n6749 & n6754 ) ;
  assign n6757 = ( n6743 & n6755 ) | ( n6743 & ~n6756 ) | ( n6755 & ~n6756 ) ;
  assign n6758 = ( ~n6717 & n6738 ) | ( ~n6717 & n6757 ) | ( n6738 & n6757 ) ;
  assign n6759 = ( n6717 & n6738 ) | ( n6717 & n6757 ) | ( n6738 & n6757 ) ;
  assign n6760 = ( n6717 & n6758 ) | ( n6717 & ~n6759 ) | ( n6758 & ~n6759 ) ;
  assign n6761 = ( ~n6638 & n6714 ) | ( ~n6638 & n6760 ) | ( n6714 & n6760 ) ;
  assign n6762 = ( n6638 & n6714 ) | ( n6638 & n6760 ) | ( n6714 & n6760 ) ;
  assign n6763 = ( n6638 & n6761 ) | ( n6638 & ~n6762 ) | ( n6761 & ~n6762 ) ;
  assign n6764 = x26 & x63 ;
  assign n6765 = x39 & x50 ;
  assign n6766 = x40 & x49 ;
  assign n6767 = ( ~n6764 & n6765 ) | ( ~n6764 & n6766 ) | ( n6765 & n6766 ) ;
  assign n6768 = ( n6764 & n6765 ) | ( n6764 & n6766 ) | ( n6765 & n6766 ) ;
  assign n6769 = ( n6764 & n6767 ) | ( n6764 & ~n6768 ) | ( n6767 & ~n6768 ) ;
  assign n6770 = ( ~n6667 & n6686 ) | ( ~n6667 & n6769 ) | ( n6686 & n6769 ) ;
  assign n6771 = ( n6667 & n6686 ) | ( n6667 & n6769 ) | ( n6686 & n6769 ) ;
  assign n6772 = ( n6667 & n6770 ) | ( n6667 & ~n6771 ) | ( n6770 & ~n6771 ) ;
  assign n6773 = ( ~n6669 & n6695 ) | ( ~n6669 & n6772 ) | ( n6695 & n6772 ) ;
  assign n6774 = ( n6669 & n6695 ) | ( n6669 & n6772 ) | ( n6695 & n6772 ) ;
  assign n6775 = ( n6669 & n6773 ) | ( n6669 & ~n6774 ) | ( n6773 & ~n6774 ) ;
  assign n6776 = ( n6656 & n6698 ) | ( n6656 & n6775 ) | ( n6698 & n6775 ) ;
  assign n6777 = ( ~n6656 & n6698 ) | ( ~n6656 & n6775 ) | ( n6698 & n6775 ) ;
  assign n6778 = ( n6656 & ~n6776 ) | ( n6656 & n6777 ) | ( ~n6776 & n6777 ) ;
  assign n6779 = ( n6701 & n6763 ) | ( n6701 & n6778 ) | ( n6763 & n6778 ) ;
  assign n6780 = ( ~n6701 & n6763 ) | ( ~n6701 & n6778 ) | ( n6763 & n6778 ) ;
  assign n6781 = ( n6701 & ~n6779 ) | ( n6701 & n6780 ) | ( ~n6779 & n6780 ) ;
  assign n6782 = ( ~n6704 & n6707 ) | ( ~n6704 & n6781 ) | ( n6707 & n6781 ) ;
  assign n6783 = ( n6704 & n6707 ) | ( n6704 & n6781 ) | ( n6707 & n6781 ) ;
  assign n6784 = ( n6704 & n6782 ) | ( n6704 & ~n6783 ) | ( n6782 & ~n6783 ) ;
  assign n6785 = ( ~n6722 & n6728 ) | ( ~n6722 & n6768 ) | ( n6728 & n6768 ) ;
  assign n6786 = ( n6722 & n6728 ) | ( n6722 & n6768 ) | ( n6728 & n6768 ) ;
  assign n6787 = ( n6722 & n6785 ) | ( n6722 & ~n6786 ) | ( n6785 & ~n6786 ) ;
  assign n6788 = x36 & x54 ;
  assign n6789 = x38 & x52 ;
  assign n6790 = x37 & x53 ;
  assign n6791 = ( ~n6788 & n6789 ) | ( ~n6788 & n6790 ) | ( n6789 & n6790 ) ;
  assign n6792 = ( n6788 & n6789 ) | ( n6788 & n6790 ) | ( n6789 & n6790 ) ;
  assign n6793 = ( n6788 & n6791 ) | ( n6788 & ~n6792 ) | ( n6791 & ~n6792 ) ;
  assign n6794 = x42 & x48 ;
  assign n6795 = x43 & x47 ;
  assign n6796 = x44 & x46 ;
  assign n6797 = ( ~n6794 & n6795 ) | ( ~n6794 & n6796 ) | ( n6795 & n6796 ) ;
  assign n6798 = ( n6794 & n6795 ) | ( n6794 & n6796 ) | ( n6795 & n6796 ) ;
  assign n6799 = ( n6794 & n6797 ) | ( n6794 & ~n6798 ) | ( n6797 & ~n6798 ) ;
  assign n6800 = x35 & x55 ;
  assign n6801 = x33 & x57 ;
  assign n6802 = x34 & x56 ;
  assign n6803 = ( ~n6800 & n6801 ) | ( ~n6800 & n6802 ) | ( n6801 & n6802 ) ;
  assign n6804 = ( n6800 & n6801 ) | ( n6800 & n6802 ) | ( n6801 & n6802 ) ;
  assign n6805 = ( n6800 & n6803 ) | ( n6800 & ~n6804 ) | ( n6803 & ~n6804 ) ;
  assign n6806 = ( ~n6793 & n6799 ) | ( ~n6793 & n6805 ) | ( n6799 & n6805 ) ;
  assign n6807 = ( n6793 & n6799 ) | ( n6793 & n6805 ) | ( n6799 & n6805 ) ;
  assign n6808 = ( n6793 & n6806 ) | ( n6793 & ~n6807 ) | ( n6806 & ~n6807 ) ;
  assign n6809 = ( ~n6710 & n6787 ) | ( ~n6710 & n6808 ) | ( n6787 & n6808 ) ;
  assign n6810 = ( n6710 & n6787 ) | ( n6710 & n6808 ) | ( n6787 & n6808 ) ;
  assign n6811 = ( n6710 & n6809 ) | ( n6710 & ~n6810 ) | ( n6809 & ~n6810 ) ;
  assign n6812 = x39 & x51 ;
  assign n6813 = x40 & x50 ;
  assign n6814 = x41 & x49 ;
  assign n6815 = ( ~n6812 & n6813 ) | ( ~n6812 & n6814 ) | ( n6813 & n6814 ) ;
  assign n6816 = ( n6812 & n6813 ) | ( n6812 & n6814 ) | ( n6813 & n6814 ) ;
  assign n6817 = ( n6812 & n6815 ) | ( n6812 & ~n6816 ) | ( n6815 & ~n6816 ) ;
  assign n6818 = ( ~n6715 & n6771 ) | ( ~n6715 & n6817 ) | ( n6771 & n6817 ) ;
  assign n6819 = ( n6715 & n6771 ) | ( n6715 & n6817 ) | ( n6771 & n6817 ) ;
  assign n6820 = ( n6715 & n6818 ) | ( n6715 & ~n6819 ) | ( n6818 & ~n6819 ) ;
  assign n6821 = x30 & x60 ;
  assign n6822 = x32 & x58 ;
  assign n6823 = x31 & x59 ;
  assign n6824 = ( ~n6821 & n6822 ) | ( ~n6821 & n6823 ) | ( n6822 & n6823 ) ;
  assign n6825 = ( n6821 & n6822 ) | ( n6821 & n6823 ) | ( n6822 & n6823 ) ;
  assign n6826 = ( n6821 & n6824 ) | ( n6821 & ~n6825 ) | ( n6824 & ~n6825 ) ;
  assign n6827 = x27 & x63 ;
  assign n6828 = x29 & x61 ;
  assign n6829 = x28 & x62 ;
  assign n6830 = ( ~n6827 & n6828 ) | ( ~n6827 & n6829 ) | ( n6828 & n6829 ) ;
  assign n6831 = ( n6827 & n6828 ) | ( n6827 & n6829 ) | ( n6828 & n6829 ) ;
  assign n6832 = ( n6827 & n6830 ) | ( n6827 & ~n6831 ) | ( n6830 & ~n6831 ) ;
  assign n6833 = ( n6741 & n6826 ) | ( n6741 & n6832 ) | ( n6826 & n6832 ) ;
  assign n6834 = ( ~n6741 & n6826 ) | ( ~n6741 & n6832 ) | ( n6826 & n6832 ) ;
  assign n6835 = ( n6741 & ~n6833 ) | ( n6741 & n6834 ) | ( ~n6833 & n6834 ) ;
  assign n6836 = ( n6774 & n6820 ) | ( n6774 & n6835 ) | ( n6820 & n6835 ) ;
  assign n6837 = ( ~n6774 & n6820 ) | ( ~n6774 & n6835 ) | ( n6820 & n6835 ) ;
  assign n6838 = ( n6774 & ~n6836 ) | ( n6774 & n6837 ) | ( ~n6836 & n6837 ) ;
  assign n6839 = ( ~n6776 & n6811 ) | ( ~n6776 & n6838 ) | ( n6811 & n6838 ) ;
  assign n6840 = ( n6776 & n6811 ) | ( n6776 & n6838 ) | ( n6811 & n6838 ) ;
  assign n6841 = ( n6776 & n6839 ) | ( n6776 & ~n6840 ) | ( n6839 & ~n6840 ) ;
  assign n6842 = ( ~n6734 & n6748 ) | ( ~n6734 & n6752 ) | ( n6748 & n6752 ) ;
  assign n6843 = ( n6734 & n6748 ) | ( n6734 & n6752 ) | ( n6748 & n6752 ) ;
  assign n6844 = ( n6734 & n6842 ) | ( n6734 & ~n6843 ) | ( n6842 & ~n6843 ) ;
  assign n6845 = ( ~n6737 & n6756 ) | ( ~n6737 & n6844 ) | ( n6756 & n6844 ) ;
  assign n6846 = ( n6737 & n6756 ) | ( n6737 & n6844 ) | ( n6756 & n6844 ) ;
  assign n6847 = ( n6737 & n6845 ) | ( n6737 & ~n6846 ) | ( n6845 & ~n6846 ) ;
  assign n6848 = ( ~n6713 & n6759 ) | ( ~n6713 & n6847 ) | ( n6759 & n6847 ) ;
  assign n6849 = ( n6713 & n6759 ) | ( n6713 & n6847 ) | ( n6759 & n6847 ) ;
  assign n6850 = ( n6713 & n6848 ) | ( n6713 & ~n6849 ) | ( n6848 & ~n6849 ) ;
  assign n6851 = ( n6762 & n6841 ) | ( n6762 & n6850 ) | ( n6841 & n6850 ) ;
  assign n6852 = ( ~n6762 & n6841 ) | ( ~n6762 & n6850 ) | ( n6841 & n6850 ) ;
  assign n6853 = ( n6762 & ~n6851 ) | ( n6762 & n6852 ) | ( ~n6851 & n6852 ) ;
  assign n6854 = ( ~n6779 & n6783 ) | ( ~n6779 & n6853 ) | ( n6783 & n6853 ) ;
  assign n6855 = ( n6779 & n6783 ) | ( n6779 & n6853 ) | ( n6783 & n6853 ) ;
  assign n6856 = ( n6779 & n6854 ) | ( n6779 & ~n6855 ) | ( n6854 & ~n6855 ) ;
  assign n6857 = ( n6792 & n6825 ) | ( n6792 & n6831 ) | ( n6825 & n6831 ) ;
  assign n6858 = ( n6792 & ~n6825 ) | ( n6792 & n6831 ) | ( ~n6825 & n6831 ) ;
  assign n6859 = ( n6825 & ~n6857 ) | ( n6825 & n6858 ) | ( ~n6857 & n6858 ) ;
  assign n6860 = x45 & x46 ;
  assign n6861 = x29 & x62 ;
  assign n6862 = ( x46 & n6860 ) | ( x46 & n6861 ) | ( n6860 & n6861 ) ;
  assign n6863 = ( x46 & ~n6860 ) | ( x46 & n6861 ) | ( ~n6860 & n6861 ) ;
  assign n6864 = ( n6860 & ~n6862 ) | ( n6860 & n6863 ) | ( ~n6862 & n6863 ) ;
  assign n6865 = x35 & x56 ;
  assign n6866 = x44 & x47 ;
  assign n6867 = x43 & x48 ;
  assign n6868 = ( ~n6865 & n6866 ) | ( ~n6865 & n6867 ) | ( n6866 & n6867 ) ;
  assign n6869 = ( n6865 & n6866 ) | ( n6865 & n6867 ) | ( n6866 & n6867 ) ;
  assign n6870 = ( n6865 & n6868 ) | ( n6865 & ~n6869 ) | ( n6868 & ~n6869 ) ;
  assign n6871 = x28 & x63 ;
  assign n6872 = x41 & x50 ;
  assign n6873 = x40 & x51 ;
  assign n6874 = ( ~n6871 & n6872 ) | ( ~n6871 & n6873 ) | ( n6872 & n6873 ) ;
  assign n6875 = ( n6871 & n6872 ) | ( n6871 & n6873 ) | ( n6872 & n6873 ) ;
  assign n6876 = ( n6871 & n6874 ) | ( n6871 & ~n6875 ) | ( n6874 & ~n6875 ) ;
  assign n6877 = ( n6864 & n6870 ) | ( n6864 & n6876 ) | ( n6870 & n6876 ) ;
  assign n6878 = ( ~n6864 & n6870 ) | ( ~n6864 & n6876 ) | ( n6870 & n6876 ) ;
  assign n6879 = ( n6864 & ~n6877 ) | ( n6864 & n6878 ) | ( ~n6877 & n6878 ) ;
  assign n6880 = ( ~n6819 & n6859 ) | ( ~n6819 & n6879 ) | ( n6859 & n6879 ) ;
  assign n6881 = ( n6819 & n6859 ) | ( n6819 & n6879 ) | ( n6859 & n6879 ) ;
  assign n6882 = ( n6819 & n6880 ) | ( n6819 & ~n6881 ) | ( n6880 & ~n6881 ) ;
  assign n6883 = x42 & x49 ;
  assign n6884 = x34 & x57 ;
  assign n6885 = x36 & x55 ;
  assign n6886 = ( ~n6883 & n6884 ) | ( ~n6883 & n6885 ) | ( n6884 & n6885 ) ;
  assign n6887 = ( n6883 & n6884 ) | ( n6883 & n6885 ) | ( n6884 & n6885 ) ;
  assign n6888 = ( n6883 & n6886 ) | ( n6883 & ~n6887 ) | ( n6886 & ~n6887 ) ;
  assign n6889 = ( ~n6786 & n6843 ) | ( ~n6786 & n6888 ) | ( n6843 & n6888 ) ;
  assign n6890 = ( n6786 & n6843 ) | ( n6786 & n6888 ) | ( n6843 & n6888 ) ;
  assign n6891 = ( n6786 & n6889 ) | ( n6786 & ~n6890 ) | ( n6889 & ~n6890 ) ;
  assign n6892 = x37 & x54 ;
  assign n6893 = x38 & x53 ;
  assign n6894 = x39 & x52 ;
  assign n6895 = ( ~n6892 & n6893 ) | ( ~n6892 & n6894 ) | ( n6893 & n6894 ) ;
  assign n6896 = ( n6892 & n6893 ) | ( n6892 & n6894 ) | ( n6893 & n6894 ) ;
  assign n6897 = ( n6892 & n6895 ) | ( n6892 & ~n6896 ) | ( n6895 & ~n6896 ) ;
  assign n6898 = x31 & x60 ;
  assign n6899 = x32 & x59 ;
  assign n6900 = x33 & x58 ;
  assign n6901 = ( ~n6898 & n6899 ) | ( ~n6898 & n6900 ) | ( n6899 & n6900 ) ;
  assign n6902 = ( n6898 & n6899 ) | ( n6898 & n6900 ) | ( n6899 & n6900 ) ;
  assign n6903 = ( n6898 & n6901 ) | ( n6898 & ~n6902 ) | ( n6901 & ~n6902 ) ;
  assign n6904 = ( n6816 & n6897 ) | ( n6816 & n6903 ) | ( n6897 & n6903 ) ;
  assign n6905 = ( ~n6816 & n6897 ) | ( ~n6816 & n6903 ) | ( n6897 & n6903 ) ;
  assign n6906 = ( n6816 & ~n6904 ) | ( n6816 & n6905 ) | ( ~n6904 & n6905 ) ;
  assign n6907 = ( ~n6846 & n6891 ) | ( ~n6846 & n6906 ) | ( n6891 & n6906 ) ;
  assign n6908 = ( n6846 & n6891 ) | ( n6846 & n6906 ) | ( n6891 & n6906 ) ;
  assign n6909 = ( n6846 & n6907 ) | ( n6846 & ~n6908 ) | ( n6907 & ~n6908 ) ;
  assign n6910 = ( ~n6849 & n6882 ) | ( ~n6849 & n6909 ) | ( n6882 & n6909 ) ;
  assign n6911 = ( n6849 & n6882 ) | ( n6849 & n6909 ) | ( n6882 & n6909 ) ;
  assign n6912 = ( n6849 & n6910 ) | ( n6849 & ~n6911 ) | ( n6910 & ~n6911 ) ;
  assign n6913 = x30 & x61 ;
  assign n6914 = ( ~n6798 & n6804 ) | ( ~n6798 & n6913 ) | ( n6804 & n6913 ) ;
  assign n6915 = ( n6798 & n6804 ) | ( n6798 & n6913 ) | ( n6804 & n6913 ) ;
  assign n6916 = ( n6798 & n6914 ) | ( n6798 & ~n6915 ) | ( n6914 & ~n6915 ) ;
  assign n6917 = ( ~n6807 & n6833 ) | ( ~n6807 & n6916 ) | ( n6833 & n6916 ) ;
  assign n6918 = ( n6807 & n6833 ) | ( n6807 & n6916 ) | ( n6833 & n6916 ) ;
  assign n6919 = ( n6807 & n6917 ) | ( n6807 & ~n6918 ) | ( n6917 & ~n6918 ) ;
  assign n6920 = ( n6810 & n6836 ) | ( n6810 & n6919 ) | ( n6836 & n6919 ) ;
  assign n6921 = ( ~n6810 & n6836 ) | ( ~n6810 & n6919 ) | ( n6836 & n6919 ) ;
  assign n6922 = ( n6810 & ~n6920 ) | ( n6810 & n6921 ) | ( ~n6920 & n6921 ) ;
  assign n6923 = ( n6840 & n6912 ) | ( n6840 & n6922 ) | ( n6912 & n6922 ) ;
  assign n6924 = ( ~n6840 & n6912 ) | ( ~n6840 & n6922 ) | ( n6912 & n6922 ) ;
  assign n6925 = ( n6840 & ~n6923 ) | ( n6840 & n6924 ) | ( ~n6923 & n6924 ) ;
  assign n6926 = ( ~n6851 & n6855 ) | ( ~n6851 & n6925 ) | ( n6855 & n6925 ) ;
  assign n6927 = ( n6851 & n6855 ) | ( n6851 & n6925 ) | ( n6855 & n6925 ) ;
  assign n6928 = ( n6851 & n6926 ) | ( n6851 & ~n6927 ) | ( n6926 & ~n6927 ) ;
  assign n6929 = x39 & x53 ;
  assign n6930 = x41 & x51 ;
  assign n6931 = x40 & x52 ;
  assign n6932 = ( ~n6929 & n6930 ) | ( ~n6929 & n6931 ) | ( n6930 & n6931 ) ;
  assign n6933 = ( n6929 & n6930 ) | ( n6929 & n6931 ) | ( n6930 & n6931 ) ;
  assign n6934 = ( n6929 & n6932 ) | ( n6929 & ~n6933 ) | ( n6932 & ~n6933 ) ;
  assign n6935 = x31 & x61 ;
  assign n6936 = x30 & x62 ;
  assign n6937 = ( ~n6862 & n6935 ) | ( ~n6862 & n6936 ) | ( n6935 & n6936 ) ;
  assign n6938 = ( n6862 & n6935 ) | ( n6862 & n6936 ) | ( n6935 & n6936 ) ;
  assign n6939 = ( n6862 & n6937 ) | ( n6862 & ~n6938 ) | ( n6937 & ~n6938 ) ;
  assign n6940 = ( n6915 & n6934 ) | ( n6915 & n6939 ) | ( n6934 & n6939 ) ;
  assign n6941 = ( ~n6915 & n6934 ) | ( ~n6915 & n6939 ) | ( n6934 & n6939 ) ;
  assign n6942 = ( n6915 & ~n6940 ) | ( n6915 & n6941 ) | ( ~n6940 & n6941 ) ;
  assign n6943 = x34 & x58 ;
  assign n6944 = x42 & x50 ;
  assign n6945 = x35 & x57 ;
  assign n6946 = ( ~n6943 & n6944 ) | ( ~n6943 & n6945 ) | ( n6944 & n6945 ) ;
  assign n6947 = ( n6943 & n6944 ) | ( n6943 & n6945 ) | ( n6944 & n6945 ) ;
  assign n6948 = ( n6943 & n6946 ) | ( n6943 & ~n6947 ) | ( n6946 & ~n6947 ) ;
  assign n6949 = x43 & x49 ;
  assign n6950 = x44 & x48 ;
  assign n6951 = x45 & x47 ;
  assign n6952 = ( ~n6949 & n6950 ) | ( ~n6949 & n6951 ) | ( n6950 & n6951 ) ;
  assign n6953 = ( n6949 & n6950 ) | ( n6949 & n6951 ) | ( n6950 & n6951 ) ;
  assign n6954 = ( n6949 & n6952 ) | ( n6949 & ~n6953 ) | ( n6952 & ~n6953 ) ;
  assign n6955 = x29 & x63 ;
  assign n6956 = x33 & x59 ;
  assign n6957 = x36 & x56 ;
  assign n6958 = ( ~n6955 & n6956 ) | ( ~n6955 & n6957 ) | ( n6956 & n6957 ) ;
  assign n6959 = ( n6955 & n6956 ) | ( n6955 & n6957 ) | ( n6956 & n6957 ) ;
  assign n6960 = ( n6955 & n6958 ) | ( n6955 & ~n6959 ) | ( n6958 & ~n6959 ) ;
  assign n6961 = ( ~n6948 & n6954 ) | ( ~n6948 & n6960 ) | ( n6954 & n6960 ) ;
  assign n6962 = ( n6948 & n6954 ) | ( n6948 & n6960 ) | ( n6954 & n6960 ) ;
  assign n6963 = ( n6948 & n6961 ) | ( n6948 & ~n6962 ) | ( n6961 & ~n6962 ) ;
  assign n6964 = ( ~n6918 & n6942 ) | ( ~n6918 & n6963 ) | ( n6942 & n6963 ) ;
  assign n6965 = ( n6918 & n6942 ) | ( n6918 & n6963 ) | ( n6942 & n6963 ) ;
  assign n6966 = ( n6918 & n6964 ) | ( n6918 & ~n6965 ) | ( n6964 & ~n6965 ) ;
  assign n6967 = ( ~n6908 & n6920 ) | ( ~n6908 & n6966 ) | ( n6920 & n6966 ) ;
  assign n6968 = ( n6908 & n6920 ) | ( n6908 & n6966 ) | ( n6920 & n6966 ) ;
  assign n6969 = ( n6908 & n6967 ) | ( n6908 & ~n6968 ) | ( n6967 & ~n6968 ) ;
  assign n6970 = ( n6857 & n6877 ) | ( n6857 & n6904 ) | ( n6877 & n6904 ) ;
  assign n6971 = ( ~n6857 & n6877 ) | ( ~n6857 & n6904 ) | ( n6877 & n6904 ) ;
  assign n6972 = ( n6857 & ~n6970 ) | ( n6857 & n6971 ) | ( ~n6970 & n6971 ) ;
  assign n6973 = ( n6875 & ~n6896 ) | ( n6875 & n6902 ) | ( ~n6896 & n6902 ) ;
  assign n6974 = ( n6875 & n6896 ) | ( n6875 & n6902 ) | ( n6896 & n6902 ) ;
  assign n6975 = ( n6896 & n6973 ) | ( n6896 & ~n6974 ) | ( n6973 & ~n6974 ) ;
  assign n6976 = x32 & x60 ;
  assign n6977 = x37 & x55 ;
  assign n6978 = x38 & x54 ;
  assign n6979 = ( ~n6976 & n6977 ) | ( ~n6976 & n6978 ) | ( n6977 & n6978 ) ;
  assign n6980 = ( n6976 & n6977 ) | ( n6976 & n6978 ) | ( n6977 & n6978 ) ;
  assign n6981 = ( n6976 & n6979 ) | ( n6976 & ~n6980 ) | ( n6979 & ~n6980 ) ;
  assign n6982 = ( ~n6869 & n6887 ) | ( ~n6869 & n6981 ) | ( n6887 & n6981 ) ;
  assign n6983 = ( n6869 & n6887 ) | ( n6869 & n6981 ) | ( n6887 & n6981 ) ;
  assign n6984 = ( n6869 & n6982 ) | ( n6869 & ~n6983 ) | ( n6982 & ~n6983 ) ;
  assign n6985 = ( ~n6890 & n6975 ) | ( ~n6890 & n6984 ) | ( n6975 & n6984 ) ;
  assign n6986 = ( n6890 & n6975 ) | ( n6890 & n6984 ) | ( n6975 & n6984 ) ;
  assign n6987 = ( n6890 & n6985 ) | ( n6890 & ~n6986 ) | ( n6985 & ~n6986 ) ;
  assign n6988 = ( ~n6881 & n6972 ) | ( ~n6881 & n6987 ) | ( n6972 & n6987 ) ;
  assign n6989 = ( n6881 & n6972 ) | ( n6881 & n6987 ) | ( n6972 & n6987 ) ;
  assign n6990 = ( n6881 & n6988 ) | ( n6881 & ~n6989 ) | ( n6988 & ~n6989 ) ;
  assign n6991 = ( n6911 & n6969 ) | ( n6911 & n6990 ) | ( n6969 & n6990 ) ;
  assign n6992 = ( ~n6911 & n6969 ) | ( ~n6911 & n6990 ) | ( n6969 & n6990 ) ;
  assign n6993 = ( n6911 & ~n6991 ) | ( n6911 & n6992 ) | ( ~n6991 & n6992 ) ;
  assign n6994 = ( n6923 & n6927 ) | ( n6923 & n6993 ) | ( n6927 & n6993 ) ;
  assign n6995 = ( n6923 & n6927 ) | ( n6923 & ~n6993 ) | ( n6927 & ~n6993 ) ;
  assign n6996 = ( n6993 & ~n6994 ) | ( n6993 & n6995 ) | ( ~n6994 & n6995 ) ;
  assign n6997 = ( n6962 & n6974 ) | ( n6962 & n6983 ) | ( n6974 & n6983 ) ;
  assign n6998 = ( n6962 & ~n6974 ) | ( n6962 & n6983 ) | ( ~n6974 & n6983 ) ;
  assign n6999 = ( n6974 & ~n6997 ) | ( n6974 & n6998 ) | ( ~n6997 & n6998 ) ;
  assign n7000 = ( n6933 & ~n6947 ) | ( n6933 & n6953 ) | ( ~n6947 & n6953 ) ;
  assign n7001 = ( n6933 & n6947 ) | ( n6933 & n6953 ) | ( n6947 & n6953 ) ;
  assign n7002 = ( n6947 & n7000 ) | ( n6947 & ~n7001 ) | ( n7000 & ~n7001 ) ;
  assign n7003 = ( ~n6938 & n6959 ) | ( ~n6938 & n6980 ) | ( n6959 & n6980 ) ;
  assign n7004 = ( n6938 & n6959 ) | ( n6938 & n6980 ) | ( n6959 & n6980 ) ;
  assign n7005 = ( n6938 & n7003 ) | ( n6938 & ~n7004 ) | ( n7003 & ~n7004 ) ;
  assign n7006 = ( ~n6940 & n7002 ) | ( ~n6940 & n7005 ) | ( n7002 & n7005 ) ;
  assign n7007 = ( n6940 & n7002 ) | ( n6940 & n7005 ) | ( n7002 & n7005 ) ;
  assign n7008 = ( n6940 & n7006 ) | ( n6940 & ~n7007 ) | ( n7006 & ~n7007 ) ;
  assign n7009 = ( ~n6986 & n6999 ) | ( ~n6986 & n7008 ) | ( n6999 & n7008 ) ;
  assign n7010 = ( n6986 & n6999 ) | ( n6986 & n7008 ) | ( n6999 & n7008 ) ;
  assign n7011 = ( n6986 & n7009 ) | ( n6986 & ~n7010 ) | ( n7009 & ~n7010 ) ;
  assign n7012 = x34 & x59 ;
  assign n7013 = x41 & x52 ;
  assign n7014 = x40 & x53 ;
  assign n7015 = ( ~n7012 & n7013 ) | ( ~n7012 & n7014 ) | ( n7013 & n7014 ) ;
  assign n7016 = ( n7012 & n7013 ) | ( n7012 & n7014 ) | ( n7013 & n7014 ) ;
  assign n7017 = ( n7012 & n7015 ) | ( n7012 & ~n7016 ) | ( n7015 & ~n7016 ) ;
  assign n7018 = x35 & x58 ;
  assign n7019 = x36 & x57 ;
  assign n7020 = x39 & x54 ;
  assign n7021 = ( ~n7018 & n7019 ) | ( ~n7018 & n7020 ) | ( n7019 & n7020 ) ;
  assign n7022 = ( n7018 & n7019 ) | ( n7018 & n7020 ) | ( n7019 & n7020 ) ;
  assign n7023 = ( n7018 & n7021 ) | ( n7018 & ~n7022 ) | ( n7021 & ~n7022 ) ;
  assign n7024 = x30 & x63 ;
  assign n7025 = x32 & x61 ;
  assign n7026 = x33 & x60 ;
  assign n7027 = ( ~n7024 & n7025 ) | ( ~n7024 & n7026 ) | ( n7025 & n7026 ) ;
  assign n7028 = ( n7024 & n7025 ) | ( n7024 & n7026 ) | ( n7025 & n7026 ) ;
  assign n7029 = ( n7024 & n7027 ) | ( n7024 & ~n7028 ) | ( n7027 & ~n7028 ) ;
  assign n7030 = ( ~n7017 & n7023 ) | ( ~n7017 & n7029 ) | ( n7023 & n7029 ) ;
  assign n7031 = ( n7017 & n7023 ) | ( n7017 & n7029 ) | ( n7023 & n7029 ) ;
  assign n7032 = ( n7017 & n7030 ) | ( n7017 & ~n7031 ) | ( n7030 & ~n7031 ) ;
  assign n7033 = x46 & x47 ;
  assign n7034 = x31 & x62 ;
  assign n7035 = ( x47 & n7033 ) | ( x47 & n7034 ) | ( n7033 & n7034 ) ;
  assign n7036 = ( x47 & ~n7033 ) | ( x47 & n7034 ) | ( ~n7033 & n7034 ) ;
  assign n7037 = ( n7033 & ~n7035 ) | ( n7033 & n7036 ) | ( ~n7035 & n7036 ) ;
  assign n7038 = x42 & x51 ;
  assign n7039 = x44 & x49 ;
  assign n7040 = x43 & x50 ;
  assign n7041 = ( ~n7038 & n7039 ) | ( ~n7038 & n7040 ) | ( n7039 & n7040 ) ;
  assign n7042 = ( n7038 & n7039 ) | ( n7038 & n7040 ) | ( n7039 & n7040 ) ;
  assign n7043 = ( n7038 & n7041 ) | ( n7038 & ~n7042 ) | ( n7041 & ~n7042 ) ;
  assign n7044 = x37 & x56 ;
  assign n7045 = x45 & x48 ;
  assign n7046 = x38 & x55 ;
  assign n7047 = ( ~n7044 & n7045 ) | ( ~n7044 & n7046 ) | ( n7045 & n7046 ) ;
  assign n7048 = ( n7044 & n7045 ) | ( n7044 & n7046 ) | ( n7045 & n7046 ) ;
  assign n7049 = ( n7044 & n7047 ) | ( n7044 & ~n7048 ) | ( n7047 & ~n7048 ) ;
  assign n7050 = ( n7037 & n7043 ) | ( n7037 & n7049 ) | ( n7043 & n7049 ) ;
  assign n7051 = ( ~n7037 & n7043 ) | ( ~n7037 & n7049 ) | ( n7043 & n7049 ) ;
  assign n7052 = ( n7037 & ~n7050 ) | ( n7037 & n7051 ) | ( ~n7050 & n7051 ) ;
  assign n7053 = ( ~n6970 & n7032 ) | ( ~n6970 & n7052 ) | ( n7032 & n7052 ) ;
  assign n7054 = ( n6970 & n7032 ) | ( n6970 & n7052 ) | ( n7032 & n7052 ) ;
  assign n7055 = ( n6970 & n7053 ) | ( n6970 & ~n7054 ) | ( n7053 & ~n7054 ) ;
  assign n7056 = ( n6965 & n6989 ) | ( n6965 & n7055 ) | ( n6989 & n7055 ) ;
  assign n7057 = ( ~n6965 & n6989 ) | ( ~n6965 & n7055 ) | ( n6989 & n7055 ) ;
  assign n7058 = ( n6965 & ~n7056 ) | ( n6965 & n7057 ) | ( ~n7056 & n7057 ) ;
  assign n7059 = ( n6968 & n7011 ) | ( n6968 & n7058 ) | ( n7011 & n7058 ) ;
  assign n7060 = ( ~n6968 & n7011 ) | ( ~n6968 & n7058 ) | ( n7011 & n7058 ) ;
  assign n7061 = ( n6968 & ~n7059 ) | ( n6968 & n7060 ) | ( ~n7059 & n7060 ) ;
  assign n7062 = ( n6991 & n6994 ) | ( n6991 & n7061 ) | ( n6994 & n7061 ) ;
  assign n7063 = ( ~n6991 & n6994 ) | ( ~n6991 & n7061 ) | ( n6994 & n7061 ) ;
  assign n7064 = ( n6991 & ~n7062 ) | ( n6991 & n7063 ) | ( ~n7062 & n7063 ) ;
  assign n7065 = ( ~n7016 & n7022 ) | ( ~n7016 & n7028 ) | ( n7022 & n7028 ) ;
  assign n7066 = ( n7016 & n7022 ) | ( n7016 & n7028 ) | ( n7022 & n7028 ) ;
  assign n7067 = ( n7016 & n7065 ) | ( n7016 & ~n7066 ) | ( n7065 & ~n7066 ) ;
  assign n7068 = x31 & x63 ;
  assign n7069 = ( n7035 & n7048 ) | ( n7035 & n7068 ) | ( n7048 & n7068 ) ;
  assign n7070 = ( n7035 & ~n7048 ) | ( n7035 & n7068 ) | ( ~n7048 & n7068 ) ;
  assign n7071 = ( n7048 & ~n7069 ) | ( n7048 & n7070 ) | ( ~n7069 & n7070 ) ;
  assign n7072 = ( n7050 & n7067 ) | ( n7050 & n7071 ) | ( n7067 & n7071 ) ;
  assign n7073 = ( ~n7050 & n7067 ) | ( ~n7050 & n7071 ) | ( n7067 & n7071 ) ;
  assign n7074 = ( n7050 & ~n7072 ) | ( n7050 & n7073 ) | ( ~n7072 & n7073 ) ;
  assign n7075 = x40 & x54 ;
  assign n7076 = x41 & x53 ;
  assign n7077 = x42 & x52 ;
  assign n7078 = ( ~n7075 & n7076 ) | ( ~n7075 & n7077 ) | ( n7076 & n7077 ) ;
  assign n7079 = ( n7075 & n7076 ) | ( n7075 & n7077 ) | ( n7076 & n7077 ) ;
  assign n7080 = ( n7075 & n7078 ) | ( n7075 & ~n7079 ) | ( n7078 & ~n7079 ) ;
  assign n7081 = x36 & x58 ;
  assign n7082 = x44 & x50 ;
  assign n7083 = x43 & x51 ;
  assign n7084 = ( ~n7081 & n7082 ) | ( ~n7081 & n7083 ) | ( n7082 & n7083 ) ;
  assign n7085 = ( n7081 & n7082 ) | ( n7081 & n7083 ) | ( n7082 & n7083 ) ;
  assign n7086 = ( n7081 & n7084 ) | ( n7081 & ~n7085 ) | ( n7084 & ~n7085 ) ;
  assign n7087 = x45 & x49 ;
  assign n7088 = x46 & x48 ;
  assign n7089 = x38 & x56 ;
  assign n7090 = ( ~n7087 & n7088 ) | ( ~n7087 & n7089 ) | ( n7088 & n7089 ) ;
  assign n7091 = ( n7087 & n7088 ) | ( n7087 & n7089 ) | ( n7088 & n7089 ) ;
  assign n7092 = ( n7087 & n7090 ) | ( n7087 & ~n7091 ) | ( n7090 & ~n7091 ) ;
  assign n7093 = ( n7080 & n7086 ) | ( n7080 & n7092 ) | ( n7086 & n7092 ) ;
  assign n7094 = ( ~n7080 & n7086 ) | ( ~n7080 & n7092 ) | ( n7086 & n7092 ) ;
  assign n7095 = ( n7080 & ~n7093 ) | ( n7080 & n7094 ) | ( ~n7093 & n7094 ) ;
  assign n7096 = x33 & x61 ;
  assign n7097 = x35 & x59 ;
  assign n7098 = ( ~n4069 & n7096 ) | ( ~n4069 & n7097 ) | ( n7096 & n7097 ) ;
  assign n7099 = ( n4069 & n7096 ) | ( n4069 & n7097 ) | ( n7096 & n7097 ) ;
  assign n7100 = ( n4069 & n7098 ) | ( n4069 & ~n7099 ) | ( n7098 & ~n7099 ) ;
  assign n7101 = x37 & x57 ;
  assign n7102 = x34 & x60 ;
  assign n7103 = x39 & x55 ;
  assign n7104 = ( ~n7101 & n7102 ) | ( ~n7101 & n7103 ) | ( n7102 & n7103 ) ;
  assign n7105 = ( n7101 & n7102 ) | ( n7101 & n7103 ) | ( n7102 & n7103 ) ;
  assign n7106 = ( n7101 & n7104 ) | ( n7101 & ~n7105 ) | ( n7104 & ~n7105 ) ;
  assign n7107 = ( n7042 & n7100 ) | ( n7042 & n7106 ) | ( n7100 & n7106 ) ;
  assign n7108 = ( ~n7042 & n7100 ) | ( ~n7042 & n7106 ) | ( n7100 & n7106 ) ;
  assign n7109 = ( n7042 & ~n7107 ) | ( n7042 & n7108 ) | ( ~n7107 & n7108 ) ;
  assign n7110 = ( ~n6997 & n7095 ) | ( ~n6997 & n7109 ) | ( n7095 & n7109 ) ;
  assign n7111 = ( n6997 & n7095 ) | ( n6997 & n7109 ) | ( n7095 & n7109 ) ;
  assign n7112 = ( n6997 & n7110 ) | ( n6997 & ~n7111 ) | ( n7110 & ~n7111 ) ;
  assign n7113 = ( ~n7010 & n7074 ) | ( ~n7010 & n7112 ) | ( n7074 & n7112 ) ;
  assign n7114 = ( n7010 & n7074 ) | ( n7010 & n7112 ) | ( n7074 & n7112 ) ;
  assign n7115 = ( n7010 & n7113 ) | ( n7010 & ~n7114 ) | ( n7113 & ~n7114 ) ;
  assign n7116 = ( n7001 & ~n7004 ) | ( n7001 & n7031 ) | ( ~n7004 & n7031 ) ;
  assign n7117 = ( n7001 & n7004 ) | ( n7001 & n7031 ) | ( n7004 & n7031 ) ;
  assign n7118 = ( n7004 & n7116 ) | ( n7004 & ~n7117 ) | ( n7116 & ~n7117 ) ;
  assign n7119 = ( n7007 & n7054 ) | ( n7007 & n7118 ) | ( n7054 & n7118 ) ;
  assign n7120 = ( n7007 & n7054 ) | ( n7007 & ~n7118 ) | ( n7054 & ~n7118 ) ;
  assign n7121 = ( n7118 & ~n7119 ) | ( n7118 & n7120 ) | ( ~n7119 & n7120 ) ;
  assign n7122 = ( n7056 & n7115 ) | ( n7056 & n7121 ) | ( n7115 & n7121 ) ;
  assign n7123 = ( ~n7056 & n7115 ) | ( ~n7056 & n7121 ) | ( n7115 & n7121 ) ;
  assign n7124 = ( n7056 & ~n7122 ) | ( n7056 & n7123 ) | ( ~n7122 & n7123 ) ;
  assign n7125 = ( ~n7059 & n7062 ) | ( ~n7059 & n7124 ) | ( n7062 & n7124 ) ;
  assign n7126 = ( n7059 & n7062 ) | ( n7059 & n7124 ) | ( n7062 & n7124 ) ;
  assign n7127 = ( n7059 & n7125 ) | ( n7059 & ~n7126 ) | ( n7125 & ~n7126 ) ;
  assign n7128 = x36 & x59 ;
  assign n7129 = x35 & x60 ;
  assign n7130 = ( n7091 & n7128 ) | ( n7091 & n7129 ) | ( n7128 & n7129 ) ;
  assign n7131 = ( ~n7091 & n7128 ) | ( ~n7091 & n7129 ) | ( n7128 & n7129 ) ;
  assign n7132 = ( n7091 & ~n7130 ) | ( n7091 & n7131 ) | ( ~n7130 & n7131 ) ;
  assign n7133 = ( n7066 & n7069 ) | ( n7066 & n7132 ) | ( n7069 & n7132 ) ;
  assign n7134 = ( ~n7066 & n7069 ) | ( ~n7066 & n7132 ) | ( n7069 & n7132 ) ;
  assign n7135 = ( n7066 & ~n7133 ) | ( n7066 & n7134 ) | ( ~n7133 & n7134 ) ;
  assign n7136 = ( ~n7072 & n7111 ) | ( ~n7072 & n7135 ) | ( n7111 & n7135 ) ;
  assign n7137 = ( n7072 & n7111 ) | ( n7072 & n7135 ) | ( n7111 & n7135 ) ;
  assign n7138 = ( n7072 & n7136 ) | ( n7072 & ~n7137 ) | ( n7136 & ~n7137 ) ;
  assign n7139 = ( n7079 & ~n7099 ) | ( n7079 & n7105 ) | ( ~n7099 & n7105 ) ;
  assign n7140 = ( n7079 & n7099 ) | ( n7079 & n7105 ) | ( n7099 & n7105 ) ;
  assign n7141 = ( n7099 & n7139 ) | ( n7099 & ~n7140 ) | ( n7139 & ~n7140 ) ;
  assign n7142 = ( ~n7093 & n7107 ) | ( ~n7093 & n7141 ) | ( n7107 & n7141 ) ;
  assign n7143 = ( n7093 & n7107 ) | ( n7093 & n7141 ) | ( n7107 & n7141 ) ;
  assign n7144 = ( n7093 & n7142 ) | ( n7093 & ~n7143 ) | ( n7142 & ~n7143 ) ;
  assign n7145 = x47 & x48 ;
  assign n7146 = x33 & x62 ;
  assign n7147 = ( x48 & n7145 ) | ( x48 & n7146 ) | ( n7145 & n7146 ) ;
  assign n7148 = ( x48 & ~n7145 ) | ( x48 & n7146 ) | ( ~n7145 & n7146 ) ;
  assign n7149 = ( n7145 & ~n7147 ) | ( n7145 & n7148 ) | ( ~n7147 & n7148 ) ;
  assign n7150 = x42 & x53 ;
  assign n7151 = x44 & x51 ;
  assign n7152 = x43 & x52 ;
  assign n7153 = ( ~n7150 & n7151 ) | ( ~n7150 & n7152 ) | ( n7151 & n7152 ) ;
  assign n7154 = ( n7150 & n7151 ) | ( n7150 & n7152 ) | ( n7151 & n7152 ) ;
  assign n7155 = ( n7150 & n7153 ) | ( n7150 & ~n7154 ) | ( n7153 & ~n7154 ) ;
  assign n7156 = x39 & x56 ;
  assign n7157 = x45 & x50 ;
  assign n7158 = x46 & x49 ;
  assign n7159 = ( ~n7156 & n7157 ) | ( ~n7156 & n7158 ) | ( n7157 & n7158 ) ;
  assign n7160 = ( n7156 & n7157 ) | ( n7156 & n7158 ) | ( n7157 & n7158 ) ;
  assign n7161 = ( n7156 & n7159 ) | ( n7156 & ~n7160 ) | ( n7159 & ~n7160 ) ;
  assign n7162 = ( n7149 & n7155 ) | ( n7149 & n7161 ) | ( n7155 & n7161 ) ;
  assign n7163 = ( ~n7149 & n7155 ) | ( ~n7149 & n7161 ) | ( n7155 & n7161 ) ;
  assign n7164 = ( n7149 & ~n7162 ) | ( n7149 & n7163 ) | ( ~n7162 & n7163 ) ;
  assign n7165 = x37 & x58 ;
  assign n7166 = x38 & x57 ;
  assign n7167 = x40 & x55 ;
  assign n7168 = ( ~n7165 & n7166 ) | ( ~n7165 & n7167 ) | ( n7166 & n7167 ) ;
  assign n7169 = ( n7165 & n7166 ) | ( n7165 & n7167 ) | ( n7166 & n7167 ) ;
  assign n7170 = ( n7165 & n7168 ) | ( n7165 & ~n7169 ) | ( n7168 & ~n7169 ) ;
  assign n7171 = x41 & x54 ;
  assign n7172 = x32 & x63 ;
  assign n7173 = x34 & x61 ;
  assign n7174 = ( ~n7171 & n7172 ) | ( ~n7171 & n7173 ) | ( n7172 & n7173 ) ;
  assign n7175 = ( n7171 & n7172 ) | ( n7171 & n7173 ) | ( n7172 & n7173 ) ;
  assign n7176 = ( n7171 & n7174 ) | ( n7171 & ~n7175 ) | ( n7174 & ~n7175 ) ;
  assign n7177 = ( n7085 & n7170 ) | ( n7085 & n7176 ) | ( n7170 & n7176 ) ;
  assign n7178 = ( ~n7085 & n7170 ) | ( ~n7085 & n7176 ) | ( n7170 & n7176 ) ;
  assign n7179 = ( n7085 & ~n7177 ) | ( n7085 & n7178 ) | ( ~n7177 & n7178 ) ;
  assign n7180 = ( ~n7117 & n7164 ) | ( ~n7117 & n7179 ) | ( n7164 & n7179 ) ;
  assign n7181 = ( n7117 & n7164 ) | ( n7117 & n7179 ) | ( n7164 & n7179 ) ;
  assign n7182 = ( n7117 & n7180 ) | ( n7117 & ~n7181 ) | ( n7180 & ~n7181 ) ;
  assign n7183 = ( ~n7119 & n7144 ) | ( ~n7119 & n7182 ) | ( n7144 & n7182 ) ;
  assign n7184 = ( n7119 & n7144 ) | ( n7119 & n7182 ) | ( n7144 & n7182 ) ;
  assign n7185 = ( n7119 & n7183 ) | ( n7119 & ~n7184 ) | ( n7183 & ~n7184 ) ;
  assign n7186 = ( ~n7114 & n7138 ) | ( ~n7114 & n7185 ) | ( n7138 & n7185 ) ;
  assign n7187 = ( n7114 & n7138 ) | ( n7114 & n7185 ) | ( n7138 & n7185 ) ;
  assign n7188 = ( n7114 & n7186 ) | ( n7114 & ~n7187 ) | ( n7186 & ~n7187 ) ;
  assign n7189 = ( ~n7122 & n7126 ) | ( ~n7122 & n7188 ) | ( n7126 & n7188 ) ;
  assign n7190 = ( n7122 & n7126 ) | ( n7122 & n7188 ) | ( n7126 & n7188 ) ;
  assign n7191 = ( n7122 & n7189 ) | ( n7122 & ~n7190 ) | ( n7189 & ~n7190 ) ;
  assign n7192 = ( n7130 & n7169 ) | ( n7130 & n7175 ) | ( n7169 & n7175 ) ;
  assign n7193 = ( ~n7130 & n7169 ) | ( ~n7130 & n7175 ) | ( n7169 & n7175 ) ;
  assign n7194 = ( n7130 & ~n7192 ) | ( n7130 & n7193 ) | ( ~n7192 & n7193 ) ;
  assign n7195 = x41 & x55 ;
  assign n7196 = x42 & x54 ;
  assign n7197 = x43 & x53 ;
  assign n7198 = ( ~n7195 & n7196 ) | ( ~n7195 & n7197 ) | ( n7196 & n7197 ) ;
  assign n7199 = ( n7195 & n7196 ) | ( n7195 & n7197 ) | ( n7196 & n7197 ) ;
  assign n7200 = ( n7195 & n7198 ) | ( n7195 & ~n7199 ) | ( n7198 & ~n7199 ) ;
  assign n7201 = x33 & x63 ;
  assign n7202 = x34 & x62 ;
  assign n7203 = x35 & x61 ;
  assign n7204 = ( ~n7201 & n7202 ) | ( ~n7201 & n7203 ) | ( n7202 & n7203 ) ;
  assign n7205 = ( n7201 & n7202 ) | ( n7201 & n7203 ) | ( n7202 & n7203 ) ;
  assign n7206 = ( n7201 & n7204 ) | ( n7201 & ~n7205 ) | ( n7204 & ~n7205 ) ;
  assign n7207 = ( ~n7140 & n7200 ) | ( ~n7140 & n7206 ) | ( n7200 & n7206 ) ;
  assign n7208 = ( n7140 & n7200 ) | ( n7140 & n7206 ) | ( n7200 & n7206 ) ;
  assign n7209 = ( n7140 & n7207 ) | ( n7140 & ~n7208 ) | ( n7207 & ~n7208 ) ;
  assign n7210 = ( ~n7133 & n7194 ) | ( ~n7133 & n7209 ) | ( n7194 & n7209 ) ;
  assign n7211 = ( n7133 & n7194 ) | ( n7133 & n7209 ) | ( n7194 & n7209 ) ;
  assign n7212 = ( n7133 & n7210 ) | ( n7133 & ~n7211 ) | ( n7210 & ~n7211 ) ;
  assign n7213 = ( n7147 & ~n7154 ) | ( n7147 & n7160 ) | ( ~n7154 & n7160 ) ;
  assign n7214 = ( n7147 & n7154 ) | ( n7147 & n7160 ) | ( n7154 & n7160 ) ;
  assign n7215 = ( n7154 & n7213 ) | ( n7154 & ~n7214 ) | ( n7213 & ~n7214 ) ;
  assign n7216 = ( ~n7162 & n7177 ) | ( ~n7162 & n7215 ) | ( n7177 & n7215 ) ;
  assign n7217 = ( n7162 & n7177 ) | ( n7162 & n7215 ) | ( n7177 & n7215 ) ;
  assign n7218 = ( n7162 & n7216 ) | ( n7162 & ~n7217 ) | ( n7216 & ~n7217 ) ;
  assign n7219 = ( ~n7137 & n7212 ) | ( ~n7137 & n7218 ) | ( n7212 & n7218 ) ;
  assign n7220 = ( n7137 & n7212 ) | ( n7137 & n7218 ) | ( n7212 & n7218 ) ;
  assign n7221 = ( n7137 & n7219 ) | ( n7137 & ~n7220 ) | ( n7219 & ~n7220 ) ;
  assign n7222 = x44 & x52 ;
  assign n7223 = x39 & x57 ;
  assign n7224 = x38 & x58 ;
  assign n7225 = ( ~n7222 & n7223 ) | ( ~n7222 & n7224 ) | ( n7223 & n7224 ) ;
  assign n7226 = ( n7222 & n7223 ) | ( n7222 & n7224 ) | ( n7223 & n7224 ) ;
  assign n7227 = ( n7222 & n7225 ) | ( n7222 & ~n7226 ) | ( n7225 & ~n7226 ) ;
  assign n7228 = x45 & x51 ;
  assign n7229 = x46 & x50 ;
  assign n7230 = x47 & x49 ;
  assign n7231 = ( ~n7228 & n7229 ) | ( ~n7228 & n7230 ) | ( n7229 & n7230 ) ;
  assign n7232 = ( n7228 & n7229 ) | ( n7228 & n7230 ) | ( n7229 & n7230 ) ;
  assign n7233 = ( n7228 & n7231 ) | ( n7228 & ~n7232 ) | ( n7231 & ~n7232 ) ;
  assign n7234 = x36 & x60 ;
  assign n7235 = x37 & x59 ;
  assign n7236 = x40 & x56 ;
  assign n7237 = ( ~n7234 & n7235 ) | ( ~n7234 & n7236 ) | ( n7235 & n7236 ) ;
  assign n7238 = ( n7234 & n7235 ) | ( n7234 & n7236 ) | ( n7235 & n7236 ) ;
  assign n7239 = ( n7234 & n7237 ) | ( n7234 & ~n7238 ) | ( n7237 & ~n7238 ) ;
  assign n7240 = ( ~n7227 & n7233 ) | ( ~n7227 & n7239 ) | ( n7233 & n7239 ) ;
  assign n7241 = ( n7227 & n7233 ) | ( n7227 & n7239 ) | ( n7233 & n7239 ) ;
  assign n7242 = ( n7227 & n7240 ) | ( n7227 & ~n7241 ) | ( n7240 & ~n7241 ) ;
  assign n7243 = ( ~n7143 & n7181 ) | ( ~n7143 & n7242 ) | ( n7181 & n7242 ) ;
  assign n7244 = ( n7143 & n7181 ) | ( n7143 & n7242 ) | ( n7181 & n7242 ) ;
  assign n7245 = ( n7143 & n7243 ) | ( n7143 & ~n7244 ) | ( n7243 & ~n7244 ) ;
  assign n7246 = ( n7184 & n7221 ) | ( n7184 & n7245 ) | ( n7221 & n7245 ) ;
  assign n7247 = ( ~n7184 & n7221 ) | ( ~n7184 & n7245 ) | ( n7221 & n7245 ) ;
  assign n7248 = ( n7184 & ~n7246 ) | ( n7184 & n7247 ) | ( ~n7246 & n7247 ) ;
  assign n7249 = ( n7187 & n7190 ) | ( n7187 & n7248 ) | ( n7190 & n7248 ) ;
  assign n7250 = ( ~n7187 & n7190 ) | ( ~n7187 & n7248 ) | ( n7190 & n7248 ) ;
  assign n7251 = ( n7187 & ~n7249 ) | ( n7187 & n7250 ) | ( ~n7249 & n7250 ) ;
  assign n7252 = x36 & x61 ;
  assign n7253 = ( n7226 & n7232 ) | ( n7226 & n7252 ) | ( n7232 & n7252 ) ;
  assign n7254 = ( ~n7226 & n7232 ) | ( ~n7226 & n7252 ) | ( n7232 & n7252 ) ;
  assign n7255 = ( n7226 & ~n7253 ) | ( n7226 & n7254 ) | ( ~n7253 & n7254 ) ;
  assign n7256 = ( ~n7192 & n7241 ) | ( ~n7192 & n7255 ) | ( n7241 & n7255 ) ;
  assign n7257 = ( n7192 & n7241 ) | ( n7192 & n7255 ) | ( n7241 & n7255 ) ;
  assign n7258 = ( n7192 & n7256 ) | ( n7192 & ~n7257 ) | ( n7256 & ~n7257 ) ;
  assign n7259 = x40 & x57 ;
  assign n7260 = x47 & x50 ;
  assign n7261 = x46 & x51 ;
  assign n7262 = ( ~n7259 & n7260 ) | ( ~n7259 & n7261 ) | ( n7260 & n7261 ) ;
  assign n7263 = ( n7259 & n7260 ) | ( n7259 & n7261 ) | ( n7260 & n7261 ) ;
  assign n7264 = ( n7259 & n7262 ) | ( n7259 & ~n7263 ) | ( n7262 & ~n7263 ) ;
  assign n7265 = x48 & x49 ;
  assign n7266 = x35 & x62 ;
  assign n7267 = ( x49 & n7265 ) | ( x49 & n7266 ) | ( n7265 & n7266 ) ;
  assign n7268 = ( x49 & ~n7265 ) | ( x49 & n7266 ) | ( ~n7265 & n7266 ) ;
  assign n7269 = ( n7265 & ~n7267 ) | ( n7265 & n7268 ) | ( ~n7267 & n7268 ) ;
  assign n7270 = ( ~n7214 & n7264 ) | ( ~n7214 & n7269 ) | ( n7264 & n7269 ) ;
  assign n7271 = ( n7214 & n7264 ) | ( n7214 & n7269 ) | ( n7264 & n7269 ) ;
  assign n7272 = ( n7214 & n7270 ) | ( n7214 & ~n7271 ) | ( n7270 & ~n7271 ) ;
  assign n7273 = ( n7199 & ~n7205 ) | ( n7199 & n7238 ) | ( ~n7205 & n7238 ) ;
  assign n7274 = ( n7199 & n7205 ) | ( n7199 & n7238 ) | ( n7205 & n7238 ) ;
  assign n7275 = ( n7205 & n7273 ) | ( n7205 & ~n7274 ) | ( n7273 & ~n7274 ) ;
  assign n7276 = ( ~n7208 & n7272 ) | ( ~n7208 & n7275 ) | ( n7272 & n7275 ) ;
  assign n7277 = ( n7208 & n7272 ) | ( n7208 & n7275 ) | ( n7272 & n7275 ) ;
  assign n7278 = ( n7208 & n7276 ) | ( n7208 & ~n7277 ) | ( n7276 & ~n7277 ) ;
  assign n7279 = ( n7244 & n7258 ) | ( n7244 & n7278 ) | ( n7258 & n7278 ) ;
  assign n7280 = ( ~n7244 & n7258 ) | ( ~n7244 & n7278 ) | ( n7258 & n7278 ) ;
  assign n7281 = ( n7244 & ~n7279 ) | ( n7244 & n7280 ) | ( ~n7279 & n7280 ) ;
  assign n7282 = x43 & x54 ;
  assign n7283 = x45 & x52 ;
  assign n7284 = x44 & x53 ;
  assign n7285 = ( ~n7282 & n7283 ) | ( ~n7282 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7286 = ( n7282 & n7283 ) | ( n7282 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7287 = ( n7282 & n7285 ) | ( n7282 & ~n7286 ) | ( n7285 & ~n7286 ) ;
  assign n7288 = x34 & x63 ;
  assign n7289 = x41 & x56 ;
  assign n7290 = x42 & x55 ;
  assign n7291 = ( ~n7288 & n7289 ) | ( ~n7288 & n7290 ) | ( n7289 & n7290 ) ;
  assign n7292 = ( n7288 & n7289 ) | ( n7288 & n7290 ) | ( n7289 & n7290 ) ;
  assign n7293 = ( n7288 & n7291 ) | ( n7288 & ~n7292 ) | ( n7291 & ~n7292 ) ;
  assign n7294 = x37 & x60 ;
  assign n7295 = x39 & x58 ;
  assign n7296 = x38 & x59 ;
  assign n7297 = ( ~n7294 & n7295 ) | ( ~n7294 & n7296 ) | ( n7295 & n7296 ) ;
  assign n7298 = ( n7294 & n7295 ) | ( n7294 & n7296 ) | ( n7295 & n7296 ) ;
  assign n7299 = ( n7294 & n7297 ) | ( n7294 & ~n7298 ) | ( n7297 & ~n7298 ) ;
  assign n7300 = ( ~n7287 & n7293 ) | ( ~n7287 & n7299 ) | ( n7293 & n7299 ) ;
  assign n7301 = ( n7287 & n7293 ) | ( n7287 & n7299 ) | ( n7293 & n7299 ) ;
  assign n7302 = ( n7287 & n7300 ) | ( n7287 & ~n7301 ) | ( n7300 & ~n7301 ) ;
  assign n7303 = ( ~n7211 & n7217 ) | ( ~n7211 & n7302 ) | ( n7217 & n7302 ) ;
  assign n7304 = ( n7211 & n7217 ) | ( n7211 & n7302 ) | ( n7217 & n7302 ) ;
  assign n7305 = ( n7211 & n7303 ) | ( n7211 & ~n7304 ) | ( n7303 & ~n7304 ) ;
  assign n7306 = ( n7220 & n7281 ) | ( n7220 & n7305 ) | ( n7281 & n7305 ) ;
  assign n7307 = ( n7220 & ~n7281 ) | ( n7220 & n7305 ) | ( ~n7281 & n7305 ) ;
  assign n7308 = ( n7281 & ~n7306 ) | ( n7281 & n7307 ) | ( ~n7306 & n7307 ) ;
  assign n7309 = ( n7246 & n7249 ) | ( n7246 & n7308 ) | ( n7249 & n7308 ) ;
  assign n7310 = ( ~n7246 & n7249 ) | ( ~n7246 & n7308 ) | ( n7249 & n7308 ) ;
  assign n7311 = ( n7246 & ~n7309 ) | ( n7246 & n7310 ) | ( ~n7309 & n7310 ) ;
  assign n7312 = ( ~n7286 & n7292 ) | ( ~n7286 & n7298 ) | ( n7292 & n7298 ) ;
  assign n7313 = ( n7286 & n7292 ) | ( n7286 & n7298 ) | ( n7292 & n7298 ) ;
  assign n7314 = ( n7286 & n7312 ) | ( n7286 & ~n7313 ) | ( n7312 & ~n7313 ) ;
  assign n7315 = x36 & x62 ;
  assign n7316 = x37 & x61 ;
  assign n7317 = ( ~n7267 & n7315 ) | ( ~n7267 & n7316 ) | ( n7315 & n7316 ) ;
  assign n7318 = ( n7267 & n7315 ) | ( n7267 & n7316 ) | ( n7315 & n7316 ) ;
  assign n7319 = ( n7267 & n7317 ) | ( n7267 & ~n7318 ) | ( n7317 & ~n7318 ) ;
  assign n7320 = x46 & x52 ;
  assign n7321 = x47 & x51 ;
  assign n7322 = x48 & x50 ;
  assign n7323 = ( ~n7320 & n7321 ) | ( ~n7320 & n7322 ) | ( n7321 & n7322 ) ;
  assign n7324 = ( n7320 & n7321 ) | ( n7320 & n7322 ) | ( n7321 & n7322 ) ;
  assign n7325 = ( n7320 & n7323 ) | ( n7320 & ~n7324 ) | ( n7323 & ~n7324 ) ;
  assign n7326 = x45 & x53 ;
  assign n7327 = x39 & x59 ;
  assign n7328 = x40 & x58 ;
  assign n7329 = ( ~n7326 & n7327 ) | ( ~n7326 & n7328 ) | ( n7327 & n7328 ) ;
  assign n7330 = ( n7326 & n7327 ) | ( n7326 & n7328 ) | ( n7327 & n7328 ) ;
  assign n7331 = ( n7326 & n7329 ) | ( n7326 & ~n7330 ) | ( n7329 & ~n7330 ) ;
  assign n7332 = ( ~n7319 & n7325 ) | ( ~n7319 & n7331 ) | ( n7325 & n7331 ) ;
  assign n7333 = ( n7319 & n7325 ) | ( n7319 & n7331 ) | ( n7325 & n7331 ) ;
  assign n7334 = ( n7319 & n7332 ) | ( n7319 & ~n7333 ) | ( n7332 & ~n7333 ) ;
  assign n7335 = ( ~n7271 & n7314 ) | ( ~n7271 & n7334 ) | ( n7314 & n7334 ) ;
  assign n7336 = ( n7271 & n7314 ) | ( n7271 & n7334 ) | ( n7314 & n7334 ) ;
  assign n7337 = ( n7271 & n7335 ) | ( n7271 & ~n7336 ) | ( n7335 & ~n7336 ) ;
  assign n7338 = ( n7253 & ~n7274 ) | ( n7253 & n7301 ) | ( ~n7274 & n7301 ) ;
  assign n7339 = ( n7253 & n7274 ) | ( n7253 & n7301 ) | ( n7274 & n7301 ) ;
  assign n7340 = ( n7274 & n7338 ) | ( n7274 & ~n7339 ) | ( n7338 & ~n7339 ) ;
  assign n7341 = ( ~n7304 & n7337 ) | ( ~n7304 & n7340 ) | ( n7337 & n7340 ) ;
  assign n7342 = ( n7304 & n7337 ) | ( n7304 & n7340 ) | ( n7337 & n7340 ) ;
  assign n7343 = ( n7304 & n7341 ) | ( n7304 & ~n7342 ) | ( n7341 & ~n7342 ) ;
  assign n7344 = x35 & x63 ;
  assign n7345 = x43 & x55 ;
  assign n7346 = x44 & x54 ;
  assign n7347 = ( ~n7344 & n7345 ) | ( ~n7344 & n7346 ) | ( n7345 & n7346 ) ;
  assign n7348 = ( n7344 & n7345 ) | ( n7344 & n7346 ) | ( n7345 & n7346 ) ;
  assign n7349 = ( n7344 & n7347 ) | ( n7344 & ~n7348 ) | ( n7347 & ~n7348 ) ;
  assign n7350 = x38 & x60 ;
  assign n7351 = x41 & x57 ;
  assign n7352 = x42 & x56 ;
  assign n7353 = ( ~n7350 & n7351 ) | ( ~n7350 & n7352 ) | ( n7351 & n7352 ) ;
  assign n7354 = ( n7350 & n7351 ) | ( n7350 & n7352 ) | ( n7351 & n7352 ) ;
  assign n7355 = ( n7350 & n7353 ) | ( n7350 & ~n7354 ) | ( n7353 & ~n7354 ) ;
  assign n7356 = ( n7263 & n7349 ) | ( n7263 & n7355 ) | ( n7349 & n7355 ) ;
  assign n7357 = ( ~n7263 & n7349 ) | ( ~n7263 & n7355 ) | ( n7349 & n7355 ) ;
  assign n7358 = ( n7263 & ~n7356 ) | ( n7263 & n7357 ) | ( ~n7356 & n7357 ) ;
  assign n7359 = ( n7257 & n7277 ) | ( n7257 & n7358 ) | ( n7277 & n7358 ) ;
  assign n7360 = ( ~n7257 & n7277 ) | ( ~n7257 & n7358 ) | ( n7277 & n7358 ) ;
  assign n7361 = ( n7257 & ~n7359 ) | ( n7257 & n7360 ) | ( ~n7359 & n7360 ) ;
  assign n7362 = ( ~n7279 & n7343 ) | ( ~n7279 & n7361 ) | ( n7343 & n7361 ) ;
  assign n7363 = ( n7279 & n7343 ) | ( n7279 & n7361 ) | ( n7343 & n7361 ) ;
  assign n7364 = ( n7279 & n7362 ) | ( n7279 & ~n7363 ) | ( n7362 & ~n7363 ) ;
  assign n7365 = ( ~n7306 & n7309 ) | ( ~n7306 & n7364 ) | ( n7309 & n7364 ) ;
  assign n7366 = ( n7306 & n7309 ) | ( n7306 & n7364 ) | ( n7309 & n7364 ) ;
  assign n7367 = ( n7306 & n7365 ) | ( n7306 & ~n7366 ) | ( n7365 & ~n7366 ) ;
  assign n7368 = x49 & x50 ;
  assign n7369 = x37 & x62 ;
  assign n7370 = ( x50 & n7368 ) | ( x50 & n7369 ) | ( n7368 & n7369 ) ;
  assign n7371 = ( x50 & ~n7368 ) | ( x50 & n7369 ) | ( ~n7368 & n7369 ) ;
  assign n7372 = ( n7368 & ~n7370 ) | ( n7368 & n7371 ) | ( ~n7370 & n7371 ) ;
  assign n7373 = ( ~n7313 & n7356 ) | ( ~n7313 & n7372 ) | ( n7356 & n7372 ) ;
  assign n7374 = ( n7313 & n7356 ) | ( n7313 & n7372 ) | ( n7356 & n7372 ) ;
  assign n7375 = ( n7313 & n7373 ) | ( n7313 & ~n7374 ) | ( n7373 & ~n7374 ) ;
  assign n7376 = ( n7324 & ~n7330 ) | ( n7324 & n7348 ) | ( ~n7330 & n7348 ) ;
  assign n7377 = ( n7324 & n7330 ) | ( n7324 & n7348 ) | ( n7330 & n7348 ) ;
  assign n7378 = ( n7330 & n7376 ) | ( n7330 & ~n7377 ) | ( n7376 & ~n7377 ) ;
  assign n7379 = x36 & x63 ;
  assign n7380 = x39 & x60 ;
  assign n7381 = x38 & x61 ;
  assign n7382 = ( ~n7379 & n7380 ) | ( ~n7379 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7383 = ( n7379 & n7380 ) | ( n7379 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7384 = ( n7379 & n7382 ) | ( n7379 & ~n7383 ) | ( n7382 & ~n7383 ) ;
  assign n7385 = ( ~n7318 & n7354 ) | ( ~n7318 & n7384 ) | ( n7354 & n7384 ) ;
  assign n7386 = ( n7318 & n7354 ) | ( n7318 & n7384 ) | ( n7354 & n7384 ) ;
  assign n7387 = ( n7318 & n7385 ) | ( n7318 & ~n7386 ) | ( n7385 & ~n7386 ) ;
  assign n7388 = ( ~n7333 & n7378 ) | ( ~n7333 & n7387 ) | ( n7378 & n7387 ) ;
  assign n7389 = ( n7333 & n7378 ) | ( n7333 & n7387 ) | ( n7378 & n7387 ) ;
  assign n7390 = ( n7333 & n7388 ) | ( n7333 & ~n7389 ) | ( n7388 & ~n7389 ) ;
  assign n7391 = ( ~n7359 & n7375 ) | ( ~n7359 & n7390 ) | ( n7375 & n7390 ) ;
  assign n7392 = ( n7359 & n7375 ) | ( n7359 & n7390 ) | ( n7375 & n7390 ) ;
  assign n7393 = ( n7359 & n7391 ) | ( n7359 & ~n7392 ) | ( n7391 & ~n7392 ) ;
  assign n7394 = x48 & x51 ;
  assign n7395 = x42 & x57 ;
  assign n7396 = x43 & x56 ;
  assign n7397 = ( ~n7394 & n7395 ) | ( ~n7394 & n7396 ) | ( n7395 & n7396 ) ;
  assign n7398 = ( n7394 & n7395 ) | ( n7394 & n7396 ) | ( n7395 & n7396 ) ;
  assign n7399 = ( n7394 & n7397 ) | ( n7394 & ~n7398 ) | ( n7397 & ~n7398 ) ;
  assign n7400 = x40 & x59 ;
  assign n7401 = x44 & x55 ;
  assign n7402 = x41 & x58 ;
  assign n7403 = ( ~n7400 & n7401 ) | ( ~n7400 & n7402 ) | ( n7401 & n7402 ) ;
  assign n7404 = ( n7400 & n7401 ) | ( n7400 & n7402 ) | ( n7401 & n7402 ) ;
  assign n7405 = ( n7400 & n7403 ) | ( n7400 & ~n7404 ) | ( n7403 & ~n7404 ) ;
  assign n7406 = x45 & x54 ;
  assign n7407 = x47 & x52 ;
  assign n7408 = x46 & x53 ;
  assign n7409 = ( ~n7406 & n7407 ) | ( ~n7406 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7410 = ( n7406 & n7407 ) | ( n7406 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7411 = ( n7406 & n7409 ) | ( n7406 & ~n7410 ) | ( n7409 & ~n7410 ) ;
  assign n7412 = ( ~n7399 & n7405 ) | ( ~n7399 & n7411 ) | ( n7405 & n7411 ) ;
  assign n7413 = ( n7399 & n7405 ) | ( n7399 & n7411 ) | ( n7405 & n7411 ) ;
  assign n7414 = ( n7399 & n7412 ) | ( n7399 & ~n7413 ) | ( n7412 & ~n7413 ) ;
  assign n7415 = ( n7336 & n7339 ) | ( n7336 & n7414 ) | ( n7339 & n7414 ) ;
  assign n7416 = ( ~n7336 & n7339 ) | ( ~n7336 & n7414 ) | ( n7339 & n7414 ) ;
  assign n7417 = ( n7336 & ~n7415 ) | ( n7336 & n7416 ) | ( ~n7415 & n7416 ) ;
  assign n7418 = ( n7342 & n7393 ) | ( n7342 & n7417 ) | ( n7393 & n7417 ) ;
  assign n7419 = ( ~n7342 & n7393 ) | ( ~n7342 & n7417 ) | ( n7393 & n7417 ) ;
  assign n7420 = ( n7342 & ~n7418 ) | ( n7342 & n7419 ) | ( ~n7418 & n7419 ) ;
  assign n7421 = ( ~n7363 & n7366 ) | ( ~n7363 & n7420 ) | ( n7366 & n7420 ) ;
  assign n7422 = ( n7363 & n7366 ) | ( n7363 & n7420 ) | ( n7366 & n7420 ) ;
  assign n7423 = ( n7363 & n7421 ) | ( n7363 & ~n7422 ) | ( n7421 & ~n7422 ) ;
  assign n7424 = ( ~n7383 & n7404 ) | ( ~n7383 & n7410 ) | ( n7404 & n7410 ) ;
  assign n7425 = ( n7383 & n7404 ) | ( n7383 & n7410 ) | ( n7404 & n7410 ) ;
  assign n7426 = ( n7383 & n7424 ) | ( n7383 & ~n7425 ) | ( n7424 & ~n7425 ) ;
  assign n7427 = x37 & x63 ;
  assign n7428 = ( n7370 & n7398 ) | ( n7370 & n7427 ) | ( n7398 & n7427 ) ;
  assign n7429 = ( n7370 & ~n7398 ) | ( n7370 & n7427 ) | ( ~n7398 & n7427 ) ;
  assign n7430 = ( n7398 & ~n7428 ) | ( n7398 & n7429 ) | ( ~n7428 & n7429 ) ;
  assign n7431 = ( ~n7413 & n7426 ) | ( ~n7413 & n7430 ) | ( n7426 & n7430 ) ;
  assign n7432 = ( n7413 & n7426 ) | ( n7413 & n7430 ) | ( n7426 & n7430 ) ;
  assign n7433 = ( n7413 & n7431 ) | ( n7413 & ~n7432 ) | ( n7431 & ~n7432 ) ;
  assign n7434 = x47 & x53 ;
  assign n7435 = x49 & x51 ;
  assign n7436 = x48 & x52 ;
  assign n7437 = ( ~n7434 & n7435 ) | ( ~n7434 & n7436 ) | ( n7435 & n7436 ) ;
  assign n7438 = ( n7434 & n7435 ) | ( n7434 & n7436 ) | ( n7435 & n7436 ) ;
  assign n7439 = ( n7434 & n7437 ) | ( n7434 & ~n7438 ) | ( n7437 & ~n7438 ) ;
  assign n7440 = ( ~n7377 & n7386 ) | ( ~n7377 & n7439 ) | ( n7386 & n7439 ) ;
  assign n7441 = ( n7377 & n7386 ) | ( n7377 & n7439 ) | ( n7386 & n7439 ) ;
  assign n7442 = ( n7377 & n7440 ) | ( n7377 & ~n7441 ) | ( n7440 & ~n7441 ) ;
  assign n7443 = ( n7415 & n7433 ) | ( n7415 & n7442 ) | ( n7433 & n7442 ) ;
  assign n7444 = ( ~n7415 & n7433 ) | ( ~n7415 & n7442 ) | ( n7433 & n7442 ) ;
  assign n7445 = ( n7415 & ~n7443 ) | ( n7415 & n7444 ) | ( ~n7443 & n7444 ) ;
  assign n7446 = x43 & x57 ;
  assign n7447 = x45 & x55 ;
  assign n7448 = x44 & x56 ;
  assign n7449 = ( ~n7446 & n7447 ) | ( ~n7446 & n7448 ) | ( n7447 & n7448 ) ;
  assign n7450 = ( n7446 & n7447 ) | ( n7446 & n7448 ) | ( n7447 & n7448 ) ;
  assign n7451 = ( n7446 & n7449 ) | ( n7446 & ~n7450 ) | ( n7449 & ~n7450 ) ;
  assign n7452 = x46 & x54 ;
  assign n7453 = x41 & x59 ;
  assign n7454 = x42 & x58 ;
  assign n7455 = ( ~n7452 & n7453 ) | ( ~n7452 & n7454 ) | ( n7453 & n7454 ) ;
  assign n7456 = ( n7452 & n7453 ) | ( n7452 & n7454 ) | ( n7453 & n7454 ) ;
  assign n7457 = ( n7452 & n7455 ) | ( n7452 & ~n7456 ) | ( n7455 & ~n7456 ) ;
  assign n7458 = x38 & x62 ;
  assign n7459 = x39 & x61 ;
  assign n7460 = x40 & x60 ;
  assign n7461 = ( ~n7458 & n7459 ) | ( ~n7458 & n7460 ) | ( n7459 & n7460 ) ;
  assign n7462 = ( n7458 & n7459 ) | ( n7458 & n7460 ) | ( n7459 & n7460 ) ;
  assign n7463 = ( n7458 & n7461 ) | ( n7458 & ~n7462 ) | ( n7461 & ~n7462 ) ;
  assign n7464 = ( ~n7451 & n7457 ) | ( ~n7451 & n7463 ) | ( n7457 & n7463 ) ;
  assign n7465 = ( n7451 & n7457 ) | ( n7451 & n7463 ) | ( n7457 & n7463 ) ;
  assign n7466 = ( n7451 & n7464 ) | ( n7451 & ~n7465 ) | ( n7464 & ~n7465 ) ;
  assign n7467 = ( ~n7374 & n7389 ) | ( ~n7374 & n7466 ) | ( n7389 & n7466 ) ;
  assign n7468 = ( n7374 & n7389 ) | ( n7374 & n7466 ) | ( n7389 & n7466 ) ;
  assign n7469 = ( n7374 & n7467 ) | ( n7374 & ~n7468 ) | ( n7467 & ~n7468 ) ;
  assign n7470 = ( n7392 & n7445 ) | ( n7392 & n7469 ) | ( n7445 & n7469 ) ;
  assign n7471 = ( ~n7392 & n7445 ) | ( ~n7392 & n7469 ) | ( n7445 & n7469 ) ;
  assign n7472 = ( n7392 & ~n7470 ) | ( n7392 & n7471 ) | ( ~n7470 & n7471 ) ;
  assign n7473 = ( ~n7418 & n7422 ) | ( ~n7418 & n7472 ) | ( n7422 & n7472 ) ;
  assign n7474 = ( n7418 & n7422 ) | ( n7418 & n7472 ) | ( n7422 & n7472 ) ;
  assign n7475 = ( n7418 & n7473 ) | ( n7418 & ~n7474 ) | ( n7473 & ~n7474 ) ;
  assign n7476 = x40 & x61 ;
  assign n7477 = x41 & x60 ;
  assign n7478 = ( n7438 & n7476 ) | ( n7438 & n7477 ) | ( n7476 & n7477 ) ;
  assign n7479 = ( ~n7438 & n7476 ) | ( ~n7438 & n7477 ) | ( n7476 & n7477 ) ;
  assign n7480 = ( n7438 & ~n7478 ) | ( n7438 & n7479 ) | ( ~n7478 & n7479 ) ;
  assign n7481 = x50 & x51 ;
  assign n7482 = x39 & x62 ;
  assign n7483 = ( x51 & n7481 ) | ( x51 & n7482 ) | ( n7481 & n7482 ) ;
  assign n7484 = ( x51 & ~n7481 ) | ( x51 & n7482 ) | ( ~n7481 & n7482 ) ;
  assign n7485 = ( n7481 & ~n7483 ) | ( n7481 & n7484 ) | ( ~n7483 & n7484 ) ;
  assign n7486 = ( ~n7428 & n7480 ) | ( ~n7428 & n7485 ) | ( n7480 & n7485 ) ;
  assign n7487 = ( n7428 & n7480 ) | ( n7428 & n7485 ) | ( n7480 & n7485 ) ;
  assign n7488 = ( n7428 & n7486 ) | ( n7428 & ~n7487 ) | ( n7486 & ~n7487 ) ;
  assign n7489 = x48 & x53 ;
  assign n7490 = x49 & x52 ;
  assign n7491 = x44 & x57 ;
  assign n7492 = ( ~n7489 & n7490 ) | ( ~n7489 & n7491 ) | ( n7490 & n7491 ) ;
  assign n7493 = ( n7489 & n7490 ) | ( n7489 & n7491 ) | ( n7490 & n7491 ) ;
  assign n7494 = ( n7489 & n7492 ) | ( n7489 & ~n7493 ) | ( n7492 & ~n7493 ) ;
  assign n7495 = x42 & x59 ;
  assign n7496 = x45 & x56 ;
  assign n7497 = x43 & x58 ;
  assign n7498 = ( ~n7495 & n7496 ) | ( ~n7495 & n7497 ) | ( n7496 & n7497 ) ;
  assign n7499 = ( n7495 & n7496 ) | ( n7495 & n7497 ) | ( n7496 & n7497 ) ;
  assign n7500 = ( n7495 & n7498 ) | ( n7495 & ~n7499 ) | ( n7498 & ~n7499 ) ;
  assign n7501 = x38 & x63 ;
  assign n7502 = x46 & x55 ;
  assign n7503 = x47 & x54 ;
  assign n7504 = ( ~n7501 & n7502 ) | ( ~n7501 & n7503 ) | ( n7502 & n7503 ) ;
  assign n7505 = ( n7501 & n7502 ) | ( n7501 & n7503 ) | ( n7502 & n7503 ) ;
  assign n7506 = ( n7501 & n7504 ) | ( n7501 & ~n7505 ) | ( n7504 & ~n7505 ) ;
  assign n7507 = ( ~n7494 & n7500 ) | ( ~n7494 & n7506 ) | ( n7500 & n7506 ) ;
  assign n7508 = ( n7494 & n7500 ) | ( n7494 & n7506 ) | ( n7500 & n7506 ) ;
  assign n7509 = ( n7494 & n7507 ) | ( n7494 & ~n7508 ) | ( n7507 & ~n7508 ) ;
  assign n7510 = ( n7441 & n7488 ) | ( n7441 & n7509 ) | ( n7488 & n7509 ) ;
  assign n7511 = ( ~n7441 & n7488 ) | ( ~n7441 & n7509 ) | ( n7488 & n7509 ) ;
  assign n7512 = ( n7441 & ~n7510 ) | ( n7441 & n7511 ) | ( ~n7510 & n7511 ) ;
  assign n7513 = ( n7450 & n7456 ) | ( n7450 & n7462 ) | ( n7456 & n7462 ) ;
  assign n7514 = ( ~n7450 & n7456 ) | ( ~n7450 & n7462 ) | ( n7456 & n7462 ) ;
  assign n7515 = ( n7450 & ~n7513 ) | ( n7450 & n7514 ) | ( ~n7513 & n7514 ) ;
  assign n7516 = ( n7425 & n7465 ) | ( n7425 & n7515 ) | ( n7465 & n7515 ) ;
  assign n7517 = ( n7425 & n7465 ) | ( n7425 & ~n7515 ) | ( n7465 & ~n7515 ) ;
  assign n7518 = ( n7515 & ~n7516 ) | ( n7515 & n7517 ) | ( ~n7516 & n7517 ) ;
  assign n7519 = ( ~n7432 & n7468 ) | ( ~n7432 & n7518 ) | ( n7468 & n7518 ) ;
  assign n7520 = ( n7432 & n7468 ) | ( n7432 & n7518 ) | ( n7468 & n7518 ) ;
  assign n7521 = ( n7432 & n7519 ) | ( n7432 & ~n7520 ) | ( n7519 & ~n7520 ) ;
  assign n7522 = ( ~n7443 & n7512 ) | ( ~n7443 & n7521 ) | ( n7512 & n7521 ) ;
  assign n7523 = ( n7443 & n7512 ) | ( n7443 & n7521 ) | ( n7512 & n7521 ) ;
  assign n7524 = ( n7443 & n7522 ) | ( n7443 & ~n7523 ) | ( n7522 & ~n7523 ) ;
  assign n7525 = ( n7470 & n7474 ) | ( n7470 & n7524 ) | ( n7474 & n7524 ) ;
  assign n7526 = ( ~n7470 & n7474 ) | ( ~n7470 & n7524 ) | ( n7474 & n7524 ) ;
  assign n7527 = ( n7470 & ~n7525 ) | ( n7470 & n7526 ) | ( ~n7525 & n7526 ) ;
  assign n7528 = ( n7483 & ~n7493 ) | ( n7483 & n7505 ) | ( ~n7493 & n7505 ) ;
  assign n7529 = ( n7483 & n7493 ) | ( n7483 & n7505 ) | ( n7493 & n7505 ) ;
  assign n7530 = ( n7493 & n7528 ) | ( n7493 & ~n7529 ) | ( n7528 & ~n7529 ) ;
  assign n7531 = ( ~n7508 & n7513 ) | ( ~n7508 & n7530 ) | ( n7513 & n7530 ) ;
  assign n7532 = ( n7508 & n7513 ) | ( n7508 & n7530 ) | ( n7513 & n7530 ) ;
  assign n7533 = ( n7508 & n7531 ) | ( n7508 & ~n7532 ) | ( n7531 & ~n7532 ) ;
  assign n7534 = ( ~n7510 & n7516 ) | ( ~n7510 & n7533 ) | ( n7516 & n7533 ) ;
  assign n7535 = ( n7510 & n7516 ) | ( n7510 & n7533 ) | ( n7516 & n7533 ) ;
  assign n7536 = ( n7510 & n7534 ) | ( n7510 & ~n7535 ) | ( n7534 & ~n7535 ) ;
  assign n7537 = x39 & x63 ;
  assign n7538 = x41 & x61 ;
  assign n7539 = x42 & x60 ;
  assign n7540 = ( ~n7537 & n7538 ) | ( ~n7537 & n7539 ) | ( n7538 & n7539 ) ;
  assign n7541 = ( n7537 & n7538 ) | ( n7537 & n7539 ) | ( n7538 & n7539 ) ;
  assign n7542 = ( n7537 & n7540 ) | ( n7537 & ~n7541 ) | ( n7540 & ~n7541 ) ;
  assign n7543 = ( n7478 & n7499 ) | ( n7478 & n7542 ) | ( n7499 & n7542 ) ;
  assign n7544 = ( n7478 & n7499 ) | ( n7478 & ~n7542 ) | ( n7499 & ~n7542 ) ;
  assign n7545 = ( n7542 & ~n7543 ) | ( n7542 & n7544 ) | ( ~n7543 & n7544 ) ;
  assign n7546 = x45 & x57 ;
  assign n7547 = x47 & x55 ;
  assign n7548 = x46 & x56 ;
  assign n7549 = ( ~n7546 & n7547 ) | ( ~n7546 & n7548 ) | ( n7547 & n7548 ) ;
  assign n7550 = ( n7546 & n7547 ) | ( n7546 & n7548 ) | ( n7547 & n7548 ) ;
  assign n7551 = ( n7546 & n7549 ) | ( n7546 & ~n7550 ) | ( n7549 & ~n7550 ) ;
  assign n7552 = x48 & x54 ;
  assign n7553 = x50 & x52 ;
  assign n7554 = x49 & x53 ;
  assign n7555 = ( ~n7552 & n7553 ) | ( ~n7552 & n7554 ) | ( n7553 & n7554 ) ;
  assign n7556 = ( n7552 & n7553 ) | ( n7552 & n7554 ) | ( n7553 & n7554 ) ;
  assign n7557 = ( n7552 & n7555 ) | ( n7552 & ~n7556 ) | ( n7555 & ~n7556 ) ;
  assign n7558 = x40 & x62 ;
  assign n7559 = x44 & x58 ;
  assign n7560 = x43 & x59 ;
  assign n7561 = ( ~n7558 & n7559 ) | ( ~n7558 & n7560 ) | ( n7559 & n7560 ) ;
  assign n7562 = ( n7558 & n7559 ) | ( n7558 & n7560 ) | ( n7559 & n7560 ) ;
  assign n7563 = ( n7558 & n7561 ) | ( n7558 & ~n7562 ) | ( n7561 & ~n7562 ) ;
  assign n7564 = ( ~n7551 & n7557 ) | ( ~n7551 & n7563 ) | ( n7557 & n7563 ) ;
  assign n7565 = ( n7551 & n7557 ) | ( n7551 & n7563 ) | ( n7557 & n7563 ) ;
  assign n7566 = ( n7551 & n7564 ) | ( n7551 & ~n7565 ) | ( n7564 & ~n7565 ) ;
  assign n7567 = ( ~n7487 & n7545 ) | ( ~n7487 & n7566 ) | ( n7545 & n7566 ) ;
  assign n7568 = ( n7487 & n7545 ) | ( n7487 & n7566 ) | ( n7545 & n7566 ) ;
  assign n7569 = ( n7487 & n7567 ) | ( n7487 & ~n7568 ) | ( n7567 & ~n7568 ) ;
  assign n7570 = ( n7520 & n7536 ) | ( n7520 & n7569 ) | ( n7536 & n7569 ) ;
  assign n7571 = ( ~n7520 & n7536 ) | ( ~n7520 & n7569 ) | ( n7536 & n7569 ) ;
  assign n7572 = ( n7520 & ~n7570 ) | ( n7520 & n7571 ) | ( ~n7570 & n7571 ) ;
  assign n7573 = ( n7523 & n7525 ) | ( n7523 & n7572 ) | ( n7525 & n7572 ) ;
  assign n7574 = ( ~n7523 & n7525 ) | ( ~n7523 & n7572 ) | ( n7525 & n7572 ) ;
  assign n7575 = ( n7523 & ~n7573 ) | ( n7523 & n7574 ) | ( ~n7573 & n7574 ) ;
  assign n7576 = x40 & x63 ;
  assign n7577 = ( n7550 & n7556 ) | ( n7550 & n7576 ) | ( n7556 & n7576 ) ;
  assign n7578 = ( ~n7550 & n7556 ) | ( ~n7550 & n7576 ) | ( n7556 & n7576 ) ;
  assign n7579 = ( n7550 & ~n7577 ) | ( n7550 & n7578 ) | ( ~n7577 & n7578 ) ;
  assign n7580 = x51 & x52 ;
  assign n7581 = x41 & x62 ;
  assign n7582 = ( x52 & n7580 ) | ( x52 & n7581 ) | ( n7580 & n7581 ) ;
  assign n7583 = ( x52 & ~n7580 ) | ( x52 & n7581 ) | ( ~n7580 & n7581 ) ;
  assign n7584 = ( n7580 & ~n7582 ) | ( n7580 & n7583 ) | ( ~n7582 & n7583 ) ;
  assign n7585 = x48 & x55 ;
  assign n7586 = x50 & x53 ;
  assign n7587 = x49 & x54 ;
  assign n7588 = ( ~n7585 & n7586 ) | ( ~n7585 & n7587 ) | ( n7586 & n7587 ) ;
  assign n7589 = ( n7585 & n7586 ) | ( n7585 & n7587 ) | ( n7586 & n7587 ) ;
  assign n7590 = ( n7585 & n7588 ) | ( n7585 & ~n7589 ) | ( n7588 & ~n7589 ) ;
  assign n7591 = x43 & x60 ;
  assign n7592 = x47 & x56 ;
  assign n7593 = x46 & x57 ;
  assign n7594 = ( ~n7591 & n7592 ) | ( ~n7591 & n7593 ) | ( n7592 & n7593 ) ;
  assign n7595 = ( n7591 & n7592 ) | ( n7591 & n7593 ) | ( n7592 & n7593 ) ;
  assign n7596 = ( n7591 & n7594 ) | ( n7591 & ~n7595 ) | ( n7594 & ~n7595 ) ;
  assign n7597 = ( n7584 & n7590 ) | ( n7584 & n7596 ) | ( n7590 & n7596 ) ;
  assign n7598 = ( ~n7584 & n7590 ) | ( ~n7584 & n7596 ) | ( n7590 & n7596 ) ;
  assign n7599 = ( n7584 & ~n7597 ) | ( n7584 & n7598 ) | ( ~n7597 & n7598 ) ;
  assign n7600 = x42 & x61 ;
  assign n7601 = x45 & x58 ;
  assign n7602 = x44 & x59 ;
  assign n7603 = ( ~n7600 & n7601 ) | ( ~n7600 & n7602 ) | ( n7601 & n7602 ) ;
  assign n7604 = ( n7600 & n7601 ) | ( n7600 & n7602 ) | ( n7601 & n7602 ) ;
  assign n7605 = ( n7600 & n7603 ) | ( n7600 & ~n7604 ) | ( n7603 & ~n7604 ) ;
  assign n7606 = ( ~n7541 & n7562 ) | ( ~n7541 & n7605 ) | ( n7562 & n7605 ) ;
  assign n7607 = ( n7541 & n7562 ) | ( n7541 & n7605 ) | ( n7562 & n7605 ) ;
  assign n7608 = ( n7541 & n7606 ) | ( n7541 & ~n7607 ) | ( n7606 & ~n7607 ) ;
  assign n7609 = ( ~n7579 & n7599 ) | ( ~n7579 & n7608 ) | ( n7599 & n7608 ) ;
  assign n7610 = ( n7579 & n7599 ) | ( n7579 & n7608 ) | ( n7599 & n7608 ) ;
  assign n7611 = ( n7579 & n7609 ) | ( n7579 & ~n7610 ) | ( n7609 & ~n7610 ) ;
  assign n7612 = ( n7529 & ~n7543 ) | ( n7529 & n7565 ) | ( ~n7543 & n7565 ) ;
  assign n7613 = ( n7529 & n7543 ) | ( n7529 & n7565 ) | ( n7543 & n7565 ) ;
  assign n7614 = ( n7543 & n7612 ) | ( n7543 & ~n7613 ) | ( n7612 & ~n7613 ) ;
  assign n7615 = ( n7532 & n7568 ) | ( n7532 & n7614 ) | ( n7568 & n7614 ) ;
  assign n7616 = ( ~n7532 & n7568 ) | ( ~n7532 & n7614 ) | ( n7568 & n7614 ) ;
  assign n7617 = ( n7532 & ~n7615 ) | ( n7532 & n7616 ) | ( ~n7615 & n7616 ) ;
  assign n7618 = ( n7535 & n7611 ) | ( n7535 & n7617 ) | ( n7611 & n7617 ) ;
  assign n7619 = ( ~n7535 & n7611 ) | ( ~n7535 & n7617 ) | ( n7611 & n7617 ) ;
  assign n7620 = ( n7535 & ~n7618 ) | ( n7535 & n7619 ) | ( ~n7618 & n7619 ) ;
  assign n7621 = ( n7570 & n7573 ) | ( n7570 & n7620 ) | ( n7573 & n7620 ) ;
  assign n7622 = ( ~n7570 & n7573 ) | ( ~n7570 & n7620 ) | ( n7573 & n7620 ) ;
  assign n7623 = ( n7570 & ~n7621 ) | ( n7570 & n7622 ) | ( ~n7621 & n7622 ) ;
  assign n7624 = x42 & x62 ;
  assign n7625 = x41 & x63 ;
  assign n7626 = ( ~n7582 & n7624 ) | ( ~n7582 & n7625 ) | ( n7624 & n7625 ) ;
  assign n7627 = ( n7582 & n7624 ) | ( n7582 & n7625 ) | ( n7624 & n7625 ) ;
  assign n7628 = ( n7582 & n7626 ) | ( n7582 & ~n7627 ) | ( n7626 & ~n7627 ) ;
  assign n7629 = ( n7577 & n7607 ) | ( n7577 & n7628 ) | ( n7607 & n7628 ) ;
  assign n7630 = ( ~n7577 & n7607 ) | ( ~n7577 & n7628 ) | ( n7607 & n7628 ) ;
  assign n7631 = ( n7577 & ~n7629 ) | ( n7577 & n7630 ) | ( ~n7629 & n7630 ) ;
  assign n7632 = ( n7610 & n7613 ) | ( n7610 & n7631 ) | ( n7613 & n7631 ) ;
  assign n7633 = ( ~n7610 & n7613 ) | ( ~n7610 & n7631 ) | ( n7613 & n7631 ) ;
  assign n7634 = ( n7610 & ~n7632 ) | ( n7610 & n7633 ) | ( ~n7632 & n7633 ) ;
  assign n7635 = ( ~n7589 & n7595 ) | ( ~n7589 & n7604 ) | ( n7595 & n7604 ) ;
  assign n7636 = ( n7589 & n7595 ) | ( n7589 & n7604 ) | ( n7595 & n7604 ) ;
  assign n7637 = ( n7589 & n7635 ) | ( n7589 & ~n7636 ) | ( n7635 & ~n7636 ) ;
  assign n7638 = x49 & x55 ;
  assign n7639 = x50 & x54 ;
  assign n7640 = x51 & x53 ;
  assign n7641 = ( ~n7638 & n7639 ) | ( ~n7638 & n7640 ) | ( n7639 & n7640 ) ;
  assign n7642 = ( n7638 & n7639 ) | ( n7638 & n7640 ) | ( n7639 & n7640 ) ;
  assign n7643 = ( n7638 & n7641 ) | ( n7638 & ~n7642 ) | ( n7641 & ~n7642 ) ;
  assign n7644 = x46 & x58 ;
  assign n7645 = x47 & x57 ;
  assign n7646 = x48 & x56 ;
  assign n7647 = ( ~n7644 & n7645 ) | ( ~n7644 & n7646 ) | ( n7645 & n7646 ) ;
  assign n7648 = ( n7644 & n7645 ) | ( n7644 & n7646 ) | ( n7645 & n7646 ) ;
  assign n7649 = ( n7644 & n7647 ) | ( n7644 & ~n7648 ) | ( n7647 & ~n7648 ) ;
  assign n7650 = x44 & x60 ;
  assign n7651 = x45 & x59 ;
  assign n7652 = x43 & x61 ;
  assign n7653 = ( ~n7650 & n7651 ) | ( ~n7650 & n7652 ) | ( n7651 & n7652 ) ;
  assign n7654 = ( n7650 & n7651 ) | ( n7650 & n7652 ) | ( n7651 & n7652 ) ;
  assign n7655 = ( n7650 & n7653 ) | ( n7650 & ~n7654 ) | ( n7653 & ~n7654 ) ;
  assign n7656 = ( ~n7643 & n7649 ) | ( ~n7643 & n7655 ) | ( n7649 & n7655 ) ;
  assign n7657 = ( n7643 & n7649 ) | ( n7643 & n7655 ) | ( n7649 & n7655 ) ;
  assign n7658 = ( n7643 & n7656 ) | ( n7643 & ~n7657 ) | ( n7656 & ~n7657 ) ;
  assign n7659 = ( ~n7597 & n7637 ) | ( ~n7597 & n7658 ) | ( n7637 & n7658 ) ;
  assign n7660 = ( n7597 & n7637 ) | ( n7597 & n7658 ) | ( n7637 & n7658 ) ;
  assign n7661 = ( n7597 & n7659 ) | ( n7597 & ~n7660 ) | ( n7659 & ~n7660 ) ;
  assign n7662 = ( n7615 & n7634 ) | ( n7615 & n7661 ) | ( n7634 & n7661 ) ;
  assign n7663 = ( ~n7615 & n7634 ) | ( ~n7615 & n7661 ) | ( n7634 & n7661 ) ;
  assign n7664 = ( n7615 & ~n7662 ) | ( n7615 & n7663 ) | ( ~n7662 & n7663 ) ;
  assign n7665 = ( ~n7618 & n7621 ) | ( ~n7618 & n7664 ) | ( n7621 & n7664 ) ;
  assign n7666 = ( n7618 & n7621 ) | ( n7618 & n7664 ) | ( n7621 & n7664 ) ;
  assign n7667 = ( n7618 & n7665 ) | ( n7618 & ~n7666 ) | ( n7665 & ~n7666 ) ;
  assign n7668 = x49 & x56 ;
  assign n7669 = x51 & x54 ;
  assign n7670 = x50 & x55 ;
  assign n7671 = ( ~n7668 & n7669 ) | ( ~n7668 & n7670 ) | ( n7669 & n7670 ) ;
  assign n7672 = ( n7668 & n7669 ) | ( n7668 & n7670 ) | ( n7669 & n7670 ) ;
  assign n7673 = ( n7668 & n7671 ) | ( n7668 & ~n7672 ) | ( n7671 & ~n7672 ) ;
  assign n7674 = x52 & x53 ;
  assign n7675 = x43 & x62 ;
  assign n7676 = ( x53 & n7674 ) | ( x53 & n7675 ) | ( n7674 & n7675 ) ;
  assign n7677 = ( x53 & ~n7674 ) | ( x53 & n7675 ) | ( ~n7674 & n7675 ) ;
  assign n7678 = ( n7674 & ~n7676 ) | ( n7674 & n7677 ) | ( ~n7676 & n7677 ) ;
  assign n7679 = ( ~n7636 & n7673 ) | ( ~n7636 & n7678 ) | ( n7673 & n7678 ) ;
  assign n7680 = ( n7636 & n7673 ) | ( n7636 & n7678 ) | ( n7673 & n7678 ) ;
  assign n7681 = ( n7636 & n7679 ) | ( n7636 & ~n7680 ) | ( n7679 & ~n7680 ) ;
  assign n7682 = x46 & x59 ;
  assign n7683 = x48 & x57 ;
  assign n7684 = x47 & x58 ;
  assign n7685 = ( ~n7682 & n7683 ) | ( ~n7682 & n7684 ) | ( n7683 & n7684 ) ;
  assign n7686 = ( n7682 & n7683 ) | ( n7682 & n7684 ) | ( n7683 & n7684 ) ;
  assign n7687 = ( n7682 & n7685 ) | ( n7682 & ~n7686 ) | ( n7685 & ~n7686 ) ;
  assign n7688 = x42 & x63 ;
  assign n7689 = x44 & x61 ;
  assign n7690 = x45 & x60 ;
  assign n7691 = ( ~n7688 & n7689 ) | ( ~n7688 & n7690 ) | ( n7689 & n7690 ) ;
  assign n7692 = ( n7688 & n7689 ) | ( n7688 & n7690 ) | ( n7689 & n7690 ) ;
  assign n7693 = ( n7688 & n7691 ) | ( n7688 & ~n7692 ) | ( n7691 & ~n7692 ) ;
  assign n7694 = ( n7627 & n7687 ) | ( n7627 & n7693 ) | ( n7687 & n7693 ) ;
  assign n7695 = ( ~n7627 & n7687 ) | ( ~n7627 & n7693 ) | ( n7687 & n7693 ) ;
  assign n7696 = ( n7627 & ~n7694 ) | ( n7627 & n7695 ) | ( ~n7694 & n7695 ) ;
  assign n7697 = ( ~n7660 & n7681 ) | ( ~n7660 & n7696 ) | ( n7681 & n7696 ) ;
  assign n7698 = ( n7660 & n7681 ) | ( n7660 & n7696 ) | ( n7681 & n7696 ) ;
  assign n7699 = ( n7660 & n7697 ) | ( n7660 & ~n7698 ) | ( n7697 & ~n7698 ) ;
  assign n7700 = ( ~n7642 & n7648 ) | ( ~n7642 & n7654 ) | ( n7648 & n7654 ) ;
  assign n7701 = ( n7642 & n7648 ) | ( n7642 & n7654 ) | ( n7648 & n7654 ) ;
  assign n7702 = ( n7642 & n7700 ) | ( n7642 & ~n7701 ) | ( n7700 & ~n7701 ) ;
  assign n7703 = ( n7629 & n7657 ) | ( n7629 & n7702 ) | ( n7657 & n7702 ) ;
  assign n7704 = ( n7629 & ~n7657 ) | ( n7629 & n7702 ) | ( ~n7657 & n7702 ) ;
  assign n7705 = ( n7657 & ~n7703 ) | ( n7657 & n7704 ) | ( ~n7703 & n7704 ) ;
  assign n7706 = ( n7632 & n7699 ) | ( n7632 & n7705 ) | ( n7699 & n7705 ) ;
  assign n7707 = ( n7632 & ~n7699 ) | ( n7632 & n7705 ) | ( ~n7699 & n7705 ) ;
  assign n7708 = ( n7699 & ~n7706 ) | ( n7699 & n7707 ) | ( ~n7706 & n7707 ) ;
  assign n7709 = ( ~n7662 & n7666 ) | ( ~n7662 & n7708 ) | ( n7666 & n7708 ) ;
  assign n7710 = ( n7662 & n7666 ) | ( n7662 & n7708 ) | ( n7666 & n7708 ) ;
  assign n7711 = ( n7662 & n7709 ) | ( n7662 & ~n7710 ) | ( n7709 & ~n7710 ) ;
  assign n7712 = x50 & x56 ;
  assign n7713 = x51 & x55 ;
  assign n7714 = x52 & x54 ;
  assign n7715 = ( ~n7712 & n7713 ) | ( ~n7712 & n7714 ) | ( n7713 & n7714 ) ;
  assign n7716 = ( n7712 & n7713 ) | ( n7712 & n7714 ) | ( n7713 & n7714 ) ;
  assign n7717 = ( n7712 & n7715 ) | ( n7712 & ~n7716 ) | ( n7715 & ~n7716 ) ;
  assign n7718 = x47 & x59 ;
  assign n7719 = x49 & x57 ;
  assign n7720 = x48 & x58 ;
  assign n7721 = ( ~n7718 & n7719 ) | ( ~n7718 & n7720 ) | ( n7719 & n7720 ) ;
  assign n7722 = ( n7718 & n7719 ) | ( n7718 & n7720 ) | ( n7719 & n7720 ) ;
  assign n7723 = ( n7718 & n7721 ) | ( n7718 & ~n7722 ) | ( n7721 & ~n7722 ) ;
  assign n7724 = ( ~n7701 & n7717 ) | ( ~n7701 & n7723 ) | ( n7717 & n7723 ) ;
  assign n7725 = ( n7701 & n7717 ) | ( n7701 & n7723 ) | ( n7717 & n7723 ) ;
  assign n7726 = ( n7701 & n7724 ) | ( n7701 & ~n7725 ) | ( n7724 & ~n7725 ) ;
  assign n7727 = x44 & x62 ;
  assign n7728 = x45 & x61 ;
  assign n7729 = x46 & x60 ;
  assign n7730 = ( ~n7727 & n7728 ) | ( ~n7727 & n7729 ) | ( n7728 & n7729 ) ;
  assign n7731 = ( n7727 & n7728 ) | ( n7727 & n7729 ) | ( n7728 & n7729 ) ;
  assign n7732 = ( n7727 & n7730 ) | ( n7727 & ~n7731 ) | ( n7730 & ~n7731 ) ;
  assign n7733 = ( ~n7686 & n7692 ) | ( ~n7686 & n7732 ) | ( n7692 & n7732 ) ;
  assign n7734 = ( n7686 & n7692 ) | ( n7686 & n7732 ) | ( n7692 & n7732 ) ;
  assign n7735 = ( n7686 & n7733 ) | ( n7686 & ~n7734 ) | ( n7733 & ~n7734 ) ;
  assign n7736 = ( n7703 & n7726 ) | ( n7703 & n7735 ) | ( n7726 & n7735 ) ;
  assign n7737 = ( ~n7703 & n7726 ) | ( ~n7703 & n7735 ) | ( n7726 & n7735 ) ;
  assign n7738 = ( n7703 & ~n7736 ) | ( n7703 & n7737 ) | ( ~n7736 & n7737 ) ;
  assign n7739 = x43 & x63 ;
  assign n7740 = ( n7672 & n7676 ) | ( n7672 & n7739 ) | ( n7676 & n7739 ) ;
  assign n7741 = ( ~n7672 & n7676 ) | ( ~n7672 & n7739 ) | ( n7676 & n7739 ) ;
  assign n7742 = ( n7672 & ~n7740 ) | ( n7672 & n7741 ) | ( ~n7740 & n7741 ) ;
  assign n7743 = ( n7680 & n7694 ) | ( n7680 & n7742 ) | ( n7694 & n7742 ) ;
  assign n7744 = ( n7680 & ~n7694 ) | ( n7680 & n7742 ) | ( ~n7694 & n7742 ) ;
  assign n7745 = ( n7694 & ~n7743 ) | ( n7694 & n7744 ) | ( ~n7743 & n7744 ) ;
  assign n7746 = ( n7698 & n7738 ) | ( n7698 & n7745 ) | ( n7738 & n7745 ) ;
  assign n7747 = ( ~n7698 & n7738 ) | ( ~n7698 & n7745 ) | ( n7738 & n7745 ) ;
  assign n7748 = ( n7698 & ~n7746 ) | ( n7698 & n7747 ) | ( ~n7746 & n7747 ) ;
  assign n7749 = ( ~n7706 & n7710 ) | ( ~n7706 & n7748 ) | ( n7710 & n7748 ) ;
  assign n7750 = ( n7706 & n7710 ) | ( n7706 & n7748 ) | ( n7710 & n7748 ) ;
  assign n7751 = ( n7706 & n7749 ) | ( n7706 & ~n7750 ) | ( n7749 & ~n7750 ) ;
  assign n7752 = x46 & x61 ;
  assign n7753 = x47 & x60 ;
  assign n7754 = ( n7716 & n7752 ) | ( n7716 & n7753 ) | ( n7752 & n7753 ) ;
  assign n7755 = ( ~n7716 & n7752 ) | ( ~n7716 & n7753 ) | ( n7752 & n7753 ) ;
  assign n7756 = ( n7716 & ~n7754 ) | ( n7716 & n7755 ) | ( ~n7754 & n7755 ) ;
  assign n7757 = x50 & x57 ;
  assign n7758 = x52 & x55 ;
  assign n7759 = x51 & x56 ;
  assign n7760 = ( ~n7757 & n7758 ) | ( ~n7757 & n7759 ) | ( n7758 & n7759 ) ;
  assign n7761 = ( n7757 & n7758 ) | ( n7757 & n7759 ) | ( n7758 & n7759 ) ;
  assign n7762 = ( n7757 & n7760 ) | ( n7757 & ~n7761 ) | ( n7760 & ~n7761 ) ;
  assign n7763 = x53 & x54 ;
  assign n7764 = x45 & x62 ;
  assign n7765 = ( x54 & n7763 ) | ( x54 & n7764 ) | ( n7763 & n7764 ) ;
  assign n7766 = ( x54 & ~n7763 ) | ( x54 & n7764 ) | ( ~n7763 & n7764 ) ;
  assign n7767 = ( n7763 & ~n7765 ) | ( n7763 & n7766 ) | ( ~n7765 & n7766 ) ;
  assign n7768 = ( ~n7756 & n7762 ) | ( ~n7756 & n7767 ) | ( n7762 & n7767 ) ;
  assign n7769 = ( n7756 & n7762 ) | ( n7756 & n7767 ) | ( n7762 & n7767 ) ;
  assign n7770 = ( n7756 & n7768 ) | ( n7756 & ~n7769 ) | ( n7768 & ~n7769 ) ;
  assign n7771 = x48 & x59 ;
  assign n7772 = x49 & x58 ;
  assign n7773 = x44 & x63 ;
  assign n7774 = ( ~n7771 & n7772 ) | ( ~n7771 & n7773 ) | ( n7772 & n7773 ) ;
  assign n7775 = ( n7771 & n7772 ) | ( n7771 & n7773 ) | ( n7772 & n7773 ) ;
  assign n7776 = ( n7771 & n7774 ) | ( n7771 & ~n7775 ) | ( n7774 & ~n7775 ) ;
  assign n7777 = ( ~n7722 & n7731 ) | ( ~n7722 & n7776 ) | ( n7731 & n7776 ) ;
  assign n7778 = ( n7722 & n7731 ) | ( n7722 & n7776 ) | ( n7731 & n7776 ) ;
  assign n7779 = ( n7722 & n7777 ) | ( n7722 & ~n7778 ) | ( n7777 & ~n7778 ) ;
  assign n7780 = ( n7743 & n7770 ) | ( n7743 & n7779 ) | ( n7770 & n7779 ) ;
  assign n7781 = ( ~n7743 & n7770 ) | ( ~n7743 & n7779 ) | ( n7770 & n7779 ) ;
  assign n7782 = ( n7743 & ~n7780 ) | ( n7743 & n7781 ) | ( ~n7780 & n7781 ) ;
  assign n7783 = ( n7725 & n7734 ) | ( n7725 & n7740 ) | ( n7734 & n7740 ) ;
  assign n7784 = ( ~n7725 & n7734 ) | ( ~n7725 & n7740 ) | ( n7734 & n7740 ) ;
  assign n7785 = ( n7725 & ~n7783 ) | ( n7725 & n7784 ) | ( ~n7783 & n7784 ) ;
  assign n7786 = ( ~n7736 & n7782 ) | ( ~n7736 & n7785 ) | ( n7782 & n7785 ) ;
  assign n7787 = ( n7736 & n7782 ) | ( n7736 & n7785 ) | ( n7782 & n7785 ) ;
  assign n7788 = ( n7736 & n7786 ) | ( n7736 & ~n7787 ) | ( n7786 & ~n7787 ) ;
  assign n7789 = ( ~n7746 & n7750 ) | ( ~n7746 & n7788 ) | ( n7750 & n7788 ) ;
  assign n7790 = ( n7746 & n7750 ) | ( n7746 & n7788 ) | ( n7750 & n7788 ) ;
  assign n7791 = ( n7746 & n7789 ) | ( n7746 & ~n7790 ) | ( n7789 & ~n7790 ) ;
  assign n7792 = x51 & x57 ;
  assign n7793 = x52 & x56 ;
  assign n7794 = x53 & x55 ;
  assign n7795 = ( ~n7792 & n7793 ) | ( ~n7792 & n7794 ) | ( n7793 & n7794 ) ;
  assign n7796 = ( n7792 & n7793 ) | ( n7792 & n7794 ) | ( n7793 & n7794 ) ;
  assign n7797 = ( n7792 & n7795 ) | ( n7792 & ~n7796 ) | ( n7795 & ~n7796 ) ;
  assign n7798 = ( ~n7769 & n7778 ) | ( ~n7769 & n7797 ) | ( n7778 & n7797 ) ;
  assign n7799 = ( n7769 & n7778 ) | ( n7769 & n7797 ) | ( n7778 & n7797 ) ;
  assign n7800 = ( n7769 & n7798 ) | ( n7769 & ~n7799 ) | ( n7798 & ~n7799 ) ;
  assign n7801 = ( ~n7761 & n7765 ) | ( ~n7761 & n7775 ) | ( n7765 & n7775 ) ;
  assign n7802 = ( n7761 & n7765 ) | ( n7761 & n7775 ) | ( n7765 & n7775 ) ;
  assign n7803 = ( n7761 & n7801 ) | ( n7761 & ~n7802 ) | ( n7801 & ~n7802 ) ;
  assign n7804 = x48 & x60 ;
  assign n7805 = x49 & x59 ;
  assign n7806 = x50 & x58 ;
  assign n7807 = ( ~n7804 & n7805 ) | ( ~n7804 & n7806 ) | ( n7805 & n7806 ) ;
  assign n7808 = ( n7804 & n7805 ) | ( n7804 & n7806 ) | ( n7805 & n7806 ) ;
  assign n7809 = ( n7804 & n7807 ) | ( n7804 & ~n7808 ) | ( n7807 & ~n7808 ) ;
  assign n7810 = x45 & x63 ;
  assign n7811 = x47 & x61 ;
  assign n7812 = x46 & x62 ;
  assign n7813 = ( ~n7810 & n7811 ) | ( ~n7810 & n7812 ) | ( n7811 & n7812 ) ;
  assign n7814 = ( n7810 & n7811 ) | ( n7810 & n7812 ) | ( n7811 & n7812 ) ;
  assign n7815 = ( n7810 & n7813 ) | ( n7810 & ~n7814 ) | ( n7813 & ~n7814 ) ;
  assign n7816 = ( n7754 & n7809 ) | ( n7754 & n7815 ) | ( n7809 & n7815 ) ;
  assign n7817 = ( ~n7754 & n7809 ) | ( ~n7754 & n7815 ) | ( n7809 & n7815 ) ;
  assign n7818 = ( n7754 & ~n7816 ) | ( n7754 & n7817 ) | ( ~n7816 & n7817 ) ;
  assign n7819 = ( ~n7783 & n7803 ) | ( ~n7783 & n7818 ) | ( n7803 & n7818 ) ;
  assign n7820 = ( n7783 & n7803 ) | ( n7783 & n7818 ) | ( n7803 & n7818 ) ;
  assign n7821 = ( n7783 & n7819 ) | ( n7783 & ~n7820 ) | ( n7819 & ~n7820 ) ;
  assign n7822 = ( n7780 & n7800 ) | ( n7780 & n7821 ) | ( n7800 & n7821 ) ;
  assign n7823 = ( ~n7780 & n7800 ) | ( ~n7780 & n7821 ) | ( n7800 & n7821 ) ;
  assign n7824 = ( n7780 & ~n7822 ) | ( n7780 & n7823 ) | ( ~n7822 & n7823 ) ;
  assign n7825 = ( n7787 & n7790 ) | ( n7787 & n7824 ) | ( n7790 & n7824 ) ;
  assign n7826 = ( ~n7787 & n7790 ) | ( ~n7787 & n7824 ) | ( n7790 & n7824 ) ;
  assign n7827 = ( n7787 & ~n7825 ) | ( n7787 & n7826 ) | ( ~n7825 & n7826 ) ;
  assign n7828 = x51 & x58 ;
  assign n7829 = x53 & x56 ;
  assign n7830 = x52 & x57 ;
  assign n7831 = ( ~n7828 & n7829 ) | ( ~n7828 & n7830 ) | ( n7829 & n7830 ) ;
  assign n7832 = ( n7828 & n7829 ) | ( n7828 & n7830 ) | ( n7829 & n7830 ) ;
  assign n7833 = ( n7828 & n7831 ) | ( n7828 & ~n7832 ) | ( n7831 & ~n7832 ) ;
  assign n7834 = x48 & x61 ;
  assign n7835 = x50 & x59 ;
  assign n7836 = x49 & x60 ;
  assign n7837 = ( ~n7834 & n7835 ) | ( ~n7834 & n7836 ) | ( n7835 & n7836 ) ;
  assign n7838 = ( n7834 & n7835 ) | ( n7834 & n7836 ) | ( n7835 & n7836 ) ;
  assign n7839 = ( n7834 & n7837 ) | ( n7834 & ~n7838 ) | ( n7837 & ~n7838 ) ;
  assign n7840 = ( n7814 & n7833 ) | ( n7814 & n7839 ) | ( n7833 & n7839 ) ;
  assign n7841 = ( ~n7814 & n7833 ) | ( ~n7814 & n7839 ) | ( n7833 & n7839 ) ;
  assign n7842 = ( n7814 & ~n7840 ) | ( n7814 & n7841 ) | ( ~n7840 & n7841 ) ;
  assign n7843 = x46 & x63 ;
  assign n7844 = ( n7796 & n7808 ) | ( n7796 & n7843 ) | ( n7808 & n7843 ) ;
  assign n7845 = ( ~n7796 & n7808 ) | ( ~n7796 & n7843 ) | ( n7808 & n7843 ) ;
  assign n7846 = ( n7796 & ~n7844 ) | ( n7796 & n7845 ) | ( ~n7844 & n7845 ) ;
  assign n7847 = ( n7799 & n7842 ) | ( n7799 & n7846 ) | ( n7842 & n7846 ) ;
  assign n7848 = ( ~n7799 & n7842 ) | ( ~n7799 & n7846 ) | ( n7842 & n7846 ) ;
  assign n7849 = ( n7799 & ~n7847 ) | ( n7799 & n7848 ) | ( ~n7847 & n7848 ) ;
  assign n7850 = x54 & x55 ;
  assign n7851 = x47 & x62 ;
  assign n7852 = ( x55 & n7850 ) | ( x55 & n7851 ) | ( n7850 & n7851 ) ;
  assign n7853 = ( x55 & ~n7850 ) | ( x55 & n7851 ) | ( ~n7850 & n7851 ) ;
  assign n7854 = ( n7850 & ~n7852 ) | ( n7850 & n7853 ) | ( ~n7852 & n7853 ) ;
  assign n7855 = ( n7802 & n7816 ) | ( n7802 & n7854 ) | ( n7816 & n7854 ) ;
  assign n7856 = ( ~n7802 & n7816 ) | ( ~n7802 & n7854 ) | ( n7816 & n7854 ) ;
  assign n7857 = ( n7802 & ~n7855 ) | ( n7802 & n7856 ) | ( ~n7855 & n7856 ) ;
  assign n7858 = ( n7820 & n7849 ) | ( n7820 & n7857 ) | ( n7849 & n7857 ) ;
  assign n7859 = ( ~n7820 & n7849 ) | ( ~n7820 & n7857 ) | ( n7849 & n7857 ) ;
  assign n7860 = ( n7820 & ~n7858 ) | ( n7820 & n7859 ) | ( ~n7858 & n7859 ) ;
  assign n7861 = ( ~n7822 & n7825 ) | ( ~n7822 & n7860 ) | ( n7825 & n7860 ) ;
  assign n7862 = ( n7822 & n7825 ) | ( n7822 & n7860 ) | ( n7825 & n7860 ) ;
  assign n7863 = ( n7822 & n7861 ) | ( n7822 & ~n7862 ) | ( n7861 & ~n7862 ) ;
  assign n7864 = x49 & x61 ;
  assign n7865 = x50 & x60 ;
  assign n7866 = x51 & x59 ;
  assign n7867 = ( ~n7864 & n7865 ) | ( ~n7864 & n7866 ) | ( n7865 & n7866 ) ;
  assign n7868 = ( n7864 & n7865 ) | ( n7864 & n7866 ) | ( n7865 & n7866 ) ;
  assign n7869 = ( n7864 & n7867 ) | ( n7864 & ~n7868 ) | ( n7867 & ~n7868 ) ;
  assign n7870 = ( ~n7832 & n7838 ) | ( ~n7832 & n7869 ) | ( n7838 & n7869 ) ;
  assign n7871 = ( n7832 & n7838 ) | ( n7832 & n7869 ) | ( n7838 & n7869 ) ;
  assign n7872 = ( n7832 & n7870 ) | ( n7832 & ~n7871 ) | ( n7870 & ~n7871 ) ;
  assign n7873 = ( ~n7840 & n7855 ) | ( ~n7840 & n7872 ) | ( n7855 & n7872 ) ;
  assign n7874 = ( n7840 & n7855 ) | ( n7840 & n7872 ) | ( n7855 & n7872 ) ;
  assign n7875 = ( n7840 & n7873 ) | ( n7840 & ~n7874 ) | ( n7873 & ~n7874 ) ;
  assign n7876 = x48 & x62 ;
  assign n7877 = x47 & x63 ;
  assign n7878 = ( ~n7852 & n7876 ) | ( ~n7852 & n7877 ) | ( n7876 & n7877 ) ;
  assign n7879 = ( n7852 & n7876 ) | ( n7852 & n7877 ) | ( n7876 & n7877 ) ;
  assign n7880 = ( n7852 & n7878 ) | ( n7852 & ~n7879 ) | ( n7878 & ~n7879 ) ;
  assign n7881 = x52 & x58 ;
  assign n7882 = x53 & x57 ;
  assign n7883 = x54 & x56 ;
  assign n7884 = ( ~n7881 & n7882 ) | ( ~n7881 & n7883 ) | ( n7882 & n7883 ) ;
  assign n7885 = ( n7881 & n7882 ) | ( n7881 & n7883 ) | ( n7882 & n7883 ) ;
  assign n7886 = ( n7881 & n7884 ) | ( n7881 & ~n7885 ) | ( n7884 & ~n7885 ) ;
  assign n7887 = ( n7844 & n7880 ) | ( n7844 & n7886 ) | ( n7880 & n7886 ) ;
  assign n7888 = ( ~n7844 & n7880 ) | ( ~n7844 & n7886 ) | ( n7880 & n7886 ) ;
  assign n7889 = ( n7844 & ~n7887 ) | ( n7844 & n7888 ) | ( ~n7887 & n7888 ) ;
  assign n7890 = ( ~n7847 & n7875 ) | ( ~n7847 & n7889 ) | ( n7875 & n7889 ) ;
  assign n7891 = ( n7847 & n7875 ) | ( n7847 & n7889 ) | ( n7875 & n7889 ) ;
  assign n7892 = ( n7847 & n7890 ) | ( n7847 & ~n7891 ) | ( n7890 & ~n7891 ) ;
  assign n7893 = ( ~n7858 & n7862 ) | ( ~n7858 & n7892 ) | ( n7862 & n7892 ) ;
  assign n7894 = ( n7858 & n7862 ) | ( n7858 & n7892 ) | ( n7862 & n7892 ) ;
  assign n7895 = ( n7858 & n7893 ) | ( n7858 & ~n7894 ) | ( n7893 & ~n7894 ) ;
  assign n7896 = x55 & x56 ;
  assign n7897 = x49 & x62 ;
  assign n7898 = ( x56 & n7896 ) | ( x56 & n7897 ) | ( n7896 & n7897 ) ;
  assign n7899 = ( x56 & ~n7896 ) | ( x56 & n7897 ) | ( ~n7896 & n7897 ) ;
  assign n7900 = ( n7896 & ~n7898 ) | ( n7896 & n7899 ) | ( ~n7898 & n7899 ) ;
  assign n7901 = x52 & x59 ;
  assign n7902 = x54 & x57 ;
  assign n7903 = x53 & x58 ;
  assign n7904 = ( ~n7901 & n7902 ) | ( ~n7901 & n7903 ) | ( n7902 & n7903 ) ;
  assign n7905 = ( n7901 & n7902 ) | ( n7901 & n7903 ) | ( n7902 & n7903 ) ;
  assign n7906 = ( n7901 & n7904 ) | ( n7901 & ~n7905 ) | ( n7904 & ~n7905 ) ;
  assign n7907 = x48 & x63 ;
  assign n7908 = x51 & x60 ;
  assign n7909 = x50 & x61 ;
  assign n7910 = ( ~n7907 & n7908 ) | ( ~n7907 & n7909 ) | ( n7908 & n7909 ) ;
  assign n7911 = ( n7907 & n7908 ) | ( n7907 & n7909 ) | ( n7908 & n7909 ) ;
  assign n7912 = ( n7907 & n7910 ) | ( n7907 & ~n7911 ) | ( n7910 & ~n7911 ) ;
  assign n7913 = ( n7900 & n7906 ) | ( n7900 & n7912 ) | ( n7906 & n7912 ) ;
  assign n7914 = ( ~n7900 & n7906 ) | ( ~n7900 & n7912 ) | ( n7906 & n7912 ) ;
  assign n7915 = ( n7900 & ~n7913 ) | ( n7900 & n7914 ) | ( ~n7913 & n7914 ) ;
  assign n7916 = ( n7868 & ~n7879 ) | ( n7868 & n7885 ) | ( ~n7879 & n7885 ) ;
  assign n7917 = ( n7868 & n7879 ) | ( n7868 & n7885 ) | ( n7879 & n7885 ) ;
  assign n7918 = ( n7879 & n7916 ) | ( n7879 & ~n7917 ) | ( n7916 & ~n7917 ) ;
  assign n7919 = ( n7871 & n7887 ) | ( n7871 & n7918 ) | ( n7887 & n7918 ) ;
  assign n7920 = ( ~n7871 & n7887 ) | ( ~n7871 & n7918 ) | ( n7887 & n7918 ) ;
  assign n7921 = ( n7871 & ~n7919 ) | ( n7871 & n7920 ) | ( ~n7919 & n7920 ) ;
  assign n7922 = ( n7874 & n7915 ) | ( n7874 & n7921 ) | ( n7915 & n7921 ) ;
  assign n7923 = ( n7874 & ~n7915 ) | ( n7874 & n7921 ) | ( ~n7915 & n7921 ) ;
  assign n7924 = ( n7915 & ~n7922 ) | ( n7915 & n7923 ) | ( ~n7922 & n7923 ) ;
  assign n7925 = ( n7891 & n7894 ) | ( n7891 & n7924 ) | ( n7894 & n7924 ) ;
  assign n7926 = ( ~n7891 & n7894 ) | ( ~n7891 & n7924 ) | ( n7894 & n7924 ) ;
  assign n7927 = ( n7891 & ~n7925 ) | ( n7891 & n7926 ) | ( ~n7925 & n7926 ) ;
  assign n7928 = x53 & x59 ;
  assign n7929 = x54 & x58 ;
  assign n7930 = x55 & x57 ;
  assign n7931 = ( ~n7928 & n7929 ) | ( ~n7928 & n7930 ) | ( n7929 & n7930 ) ;
  assign n7932 = ( n7928 & n7929 ) | ( n7928 & n7930 ) | ( n7929 & n7930 ) ;
  assign n7933 = ( n7928 & n7931 ) | ( n7928 & ~n7932 ) | ( n7931 & ~n7932 ) ;
  assign n7934 = x49 & x63 ;
  assign n7935 = x51 & x61 ;
  assign n7936 = x52 & x60 ;
  assign n7937 = ( ~n7934 & n7935 ) | ( ~n7934 & n7936 ) | ( n7935 & n7936 ) ;
  assign n7938 = ( n7934 & n7935 ) | ( n7934 & n7936 ) | ( n7935 & n7936 ) ;
  assign n7939 = ( n7934 & n7937 ) | ( n7934 & ~n7938 ) | ( n7937 & ~n7938 ) ;
  assign n7940 = ( n7911 & n7933 ) | ( n7911 & n7939 ) | ( n7933 & n7939 ) ;
  assign n7941 = ( ~n7911 & n7933 ) | ( ~n7911 & n7939 ) | ( n7933 & n7939 ) ;
  assign n7942 = ( n7911 & ~n7940 ) | ( n7911 & n7941 ) | ( ~n7940 & n7941 ) ;
  assign n7943 = x50 & x62 ;
  assign n7944 = ( n7898 & n7905 ) | ( n7898 & n7943 ) | ( n7905 & n7943 ) ;
  assign n7945 = ( n7898 & ~n7905 ) | ( n7898 & n7943 ) | ( ~n7905 & n7943 ) ;
  assign n7946 = ( n7905 & ~n7944 ) | ( n7905 & n7945 ) | ( ~n7944 & n7945 ) ;
  assign n7947 = ( n7913 & n7917 ) | ( n7913 & n7946 ) | ( n7917 & n7946 ) ;
  assign n7948 = ( ~n7913 & n7917 ) | ( ~n7913 & n7946 ) | ( n7917 & n7946 ) ;
  assign n7949 = ( n7913 & ~n7947 ) | ( n7913 & n7948 ) | ( ~n7947 & n7948 ) ;
  assign n7950 = ( n7919 & n7942 ) | ( n7919 & n7949 ) | ( n7942 & n7949 ) ;
  assign n7951 = ( ~n7919 & n7942 ) | ( ~n7919 & n7949 ) | ( n7942 & n7949 ) ;
  assign n7952 = ( n7919 & ~n7950 ) | ( n7919 & n7951 ) | ( ~n7950 & n7951 ) ;
  assign n7953 = ( ~n7922 & n7925 ) | ( ~n7922 & n7952 ) | ( n7925 & n7952 ) ;
  assign n7954 = ( n7922 & n7925 ) | ( n7922 & n7952 ) | ( n7925 & n7952 ) ;
  assign n7955 = ( n7922 & n7953 ) | ( n7922 & ~n7954 ) | ( n7953 & ~n7954 ) ;
  assign n7956 = x52 & x61 ;
  assign n7957 = x53 & x60 ;
  assign n7958 = ( n7932 & n7956 ) | ( n7932 & n7957 ) | ( n7956 & n7957 ) ;
  assign n7959 = ( ~n7932 & n7956 ) | ( ~n7932 & n7957 ) | ( n7956 & n7957 ) ;
  assign n7960 = ( n7932 & ~n7958 ) | ( n7932 & n7959 ) | ( ~n7958 & n7959 ) ;
  assign n7961 = ( ~n7940 & n7944 ) | ( ~n7940 & n7960 ) | ( n7944 & n7960 ) ;
  assign n7962 = ( n7940 & n7944 ) | ( n7940 & n7960 ) | ( n7944 & n7960 ) ;
  assign n7963 = ( n7940 & n7961 ) | ( n7940 & ~n7962 ) | ( n7961 & ~n7962 ) ;
  assign n7964 = x50 & x63 ;
  assign n7965 = x55 & x58 ;
  assign n7966 = x54 & x59 ;
  assign n7967 = ( ~n7964 & n7965 ) | ( ~n7964 & n7966 ) | ( n7965 & n7966 ) ;
  assign n7968 = ( n7964 & n7965 ) | ( n7964 & n7966 ) | ( n7965 & n7966 ) ;
  assign n7969 = ( n7964 & n7967 ) | ( n7964 & ~n7968 ) | ( n7967 & ~n7968 ) ;
  assign n7970 = x56 & x57 ;
  assign n7971 = x51 & x62 ;
  assign n7972 = ( x57 & n7970 ) | ( x57 & n7971 ) | ( n7970 & n7971 ) ;
  assign n7973 = ( x57 & ~n7970 ) | ( x57 & n7971 ) | ( ~n7970 & n7971 ) ;
  assign n7974 = ( n7970 & ~n7972 ) | ( n7970 & n7973 ) | ( ~n7972 & n7973 ) ;
  assign n7975 = ( ~n7938 & n7969 ) | ( ~n7938 & n7974 ) | ( n7969 & n7974 ) ;
  assign n7976 = ( n7938 & n7969 ) | ( n7938 & n7974 ) | ( n7969 & n7974 ) ;
  assign n7977 = ( n7938 & n7975 ) | ( n7938 & ~n7976 ) | ( n7975 & ~n7976 ) ;
  assign n7978 = ( ~n7947 & n7963 ) | ( ~n7947 & n7977 ) | ( n7963 & n7977 ) ;
  assign n7979 = ( n7947 & n7963 ) | ( n7947 & n7977 ) | ( n7963 & n7977 ) ;
  assign n7980 = ( n7947 & n7978 ) | ( n7947 & ~n7979 ) | ( n7978 & ~n7979 ) ;
  assign n7981 = ( ~n7950 & n7954 ) | ( ~n7950 & n7980 ) | ( n7954 & n7980 ) ;
  assign n7982 = ( n7950 & n7954 ) | ( n7950 & n7980 ) | ( n7954 & n7980 ) ;
  assign n7983 = ( n7950 & n7981 ) | ( n7950 & ~n7982 ) | ( n7981 & ~n7982 ) ;
  assign n7984 = ( ~n7958 & n7968 ) | ( ~n7958 & n7972 ) | ( n7968 & n7972 ) ;
  assign n7985 = ( n7958 & n7968 ) | ( n7958 & n7972 ) | ( n7968 & n7972 ) ;
  assign n7986 = ( n7958 & n7984 ) | ( n7958 & ~n7985 ) | ( n7984 & ~n7985 ) ;
  assign n7987 = x54 & x60 ;
  assign n7988 = x55 & x59 ;
  assign n7989 = x56 & x58 ;
  assign n7990 = ( ~n7987 & n7988 ) | ( ~n7987 & n7989 ) | ( n7988 & n7989 ) ;
  assign n7991 = ( n7987 & n7988 ) | ( n7987 & n7989 ) | ( n7988 & n7989 ) ;
  assign n7992 = ( n7987 & n7990 ) | ( n7987 & ~n7991 ) | ( n7990 & ~n7991 ) ;
  assign n7993 = x51 & x63 ;
  assign n7994 = x53 & x61 ;
  assign n7995 = x52 & x62 ;
  assign n7996 = ( ~n7993 & n7994 ) | ( ~n7993 & n7995 ) | ( n7994 & n7995 ) ;
  assign n7997 = ( n7993 & n7994 ) | ( n7993 & n7995 ) | ( n7994 & n7995 ) ;
  assign n7998 = ( n7993 & n7996 ) | ( n7993 & ~n7997 ) | ( n7996 & ~n7997 ) ;
  assign n7999 = ( n7976 & n7992 ) | ( n7976 & n7998 ) | ( n7992 & n7998 ) ;
  assign n8000 = ( ~n7976 & n7992 ) | ( ~n7976 & n7998 ) | ( n7992 & n7998 ) ;
  assign n8001 = ( n7976 & ~n7999 ) | ( n7976 & n8000 ) | ( ~n7999 & n8000 ) ;
  assign n8002 = ( ~n7962 & n7986 ) | ( ~n7962 & n8001 ) | ( n7986 & n8001 ) ;
  assign n8003 = ( n7962 & n7986 ) | ( n7962 & n8001 ) | ( n7986 & n8001 ) ;
  assign n8004 = ( n7962 & n8002 ) | ( n7962 & ~n8003 ) | ( n8002 & ~n8003 ) ;
  assign n8005 = ( n7979 & n7982 ) | ( n7979 & n8004 ) | ( n7982 & n8004 ) ;
  assign n8006 = ( ~n7979 & n7982 ) | ( ~n7979 & n8004 ) | ( n7982 & n8004 ) ;
  assign n8007 = ( n7979 & ~n8005 ) | ( n7979 & n8006 ) | ( ~n8005 & n8006 ) ;
  assign n8008 = x54 & x61 ;
  assign n8009 = x56 & x59 ;
  assign n8010 = x55 & x60 ;
  assign n8011 = ( ~n8008 & n8009 ) | ( ~n8008 & n8010 ) | ( n8009 & n8010 ) ;
  assign n8012 = ( n8008 & n8009 ) | ( n8008 & n8010 ) | ( n8009 & n8010 ) ;
  assign n8013 = ( n8008 & n8011 ) | ( n8008 & ~n8012 ) | ( n8011 & ~n8012 ) ;
  assign n8014 = x57 & x58 ;
  assign n8015 = x53 & x62 ;
  assign n8016 = ( x58 & n8014 ) | ( x58 & n8015 ) | ( n8014 & n8015 ) ;
  assign n8017 = ( x58 & ~n8014 ) | ( x58 & n8015 ) | ( ~n8014 & n8015 ) ;
  assign n8018 = ( n8014 & ~n8016 ) | ( n8014 & n8017 ) | ( ~n8016 & n8017 ) ;
  assign n8019 = ( ~n7985 & n8013 ) | ( ~n7985 & n8018 ) | ( n8013 & n8018 ) ;
  assign n8020 = ( n7985 & n8013 ) | ( n7985 & n8018 ) | ( n8013 & n8018 ) ;
  assign n8021 = ( n7985 & n8019 ) | ( n7985 & ~n8020 ) | ( n8019 & ~n8020 ) ;
  assign n8022 = x52 & x63 ;
  assign n8023 = ( ~n7991 & n7997 ) | ( ~n7991 & n8022 ) | ( n7997 & n8022 ) ;
  assign n8024 = ( n7991 & n7997 ) | ( n7991 & n8022 ) | ( n7997 & n8022 ) ;
  assign n8025 = ( n7991 & n8023 ) | ( n7991 & ~n8024 ) | ( n8023 & ~n8024 ) ;
  assign n8026 = ( ~n7999 & n8021 ) | ( ~n7999 & n8025 ) | ( n8021 & n8025 ) ;
  assign n8027 = ( n7999 & n8021 ) | ( n7999 & n8025 ) | ( n8021 & n8025 ) ;
  assign n8028 = ( n7999 & n8026 ) | ( n7999 & ~n8027 ) | ( n8026 & ~n8027 ) ;
  assign n8029 = ( n8003 & n8005 ) | ( n8003 & n8028 ) | ( n8005 & n8028 ) ;
  assign n8030 = ( ~n8003 & n8005 ) | ( ~n8003 & n8028 ) | ( n8005 & n8028 ) ;
  assign n8031 = ( n8003 & ~n8029 ) | ( n8003 & n8030 ) | ( ~n8029 & n8030 ) ;
  assign n8032 = x54 & x62 ;
  assign n8033 = x53 & x63 ;
  assign n8034 = ( ~n8016 & n8032 ) | ( ~n8016 & n8033 ) | ( n8032 & n8033 ) ;
  assign n8035 = ( n8016 & n8032 ) | ( n8016 & n8033 ) | ( n8032 & n8033 ) ;
  assign n8036 = ( n8016 & n8034 ) | ( n8016 & ~n8035 ) | ( n8034 & ~n8035 ) ;
  assign n8037 = x55 & x61 ;
  assign n8038 = x56 & x60 ;
  assign n8039 = x57 & x59 ;
  assign n8040 = ( ~n8037 & n8038 ) | ( ~n8037 & n8039 ) | ( n8038 & n8039 ) ;
  assign n8041 = ( n8037 & n8038 ) | ( n8037 & n8039 ) | ( n8038 & n8039 ) ;
  assign n8042 = ( n8037 & n8040 ) | ( n8037 & ~n8041 ) | ( n8040 & ~n8041 ) ;
  assign n8043 = ( ~n8012 & n8036 ) | ( ~n8012 & n8042 ) | ( n8036 & n8042 ) ;
  assign n8044 = ( n8012 & n8036 ) | ( n8012 & n8042 ) | ( n8036 & n8042 ) ;
  assign n8045 = ( n8012 & n8043 ) | ( n8012 & ~n8044 ) | ( n8043 & ~n8044 ) ;
  assign n8046 = ( ~n8020 & n8024 ) | ( ~n8020 & n8045 ) | ( n8024 & n8045 ) ;
  assign n8047 = ( n8020 & n8024 ) | ( n8020 & n8045 ) | ( n8024 & n8045 ) ;
  assign n8048 = ( n8020 & n8046 ) | ( n8020 & ~n8047 ) | ( n8046 & ~n8047 ) ;
  assign n8049 = ( n8027 & n8029 ) | ( n8027 & n8048 ) | ( n8029 & n8048 ) ;
  assign n8050 = ( ~n8027 & n8029 ) | ( ~n8027 & n8048 ) | ( n8029 & n8048 ) ;
  assign n8051 = ( n8027 & ~n8049 ) | ( n8027 & n8050 ) | ( ~n8049 & n8050 ) ;
  assign n8052 = x54 & x63 ;
  assign n8053 = x57 & x60 ;
  assign n8054 = x56 & x61 ;
  assign n8055 = ( ~n8052 & n8053 ) | ( ~n8052 & n8054 ) | ( n8053 & n8054 ) ;
  assign n8056 = ( n8052 & n8053 ) | ( n8052 & n8054 ) | ( n8053 & n8054 ) ;
  assign n8057 = ( n8052 & n8055 ) | ( n8052 & ~n8056 ) | ( n8055 & ~n8056 ) ;
  assign n8058 = ( ~n8035 & n8041 ) | ( ~n8035 & n8057 ) | ( n8041 & n8057 ) ;
  assign n8059 = ( n8035 & n8041 ) | ( n8035 & n8057 ) | ( n8041 & n8057 ) ;
  assign n8060 = ( n8035 & n8058 ) | ( n8035 & ~n8059 ) | ( n8058 & ~n8059 ) ;
  assign n8061 = x58 & x59 ;
  assign n8062 = x55 & x62 ;
  assign n8063 = ( x59 & n8061 ) | ( x59 & n8062 ) | ( n8061 & n8062 ) ;
  assign n8064 = ( x59 & ~n8061 ) | ( x59 & n8062 ) | ( ~n8061 & n8062 ) ;
  assign n8065 = ( n8061 & ~n8063 ) | ( n8061 & n8064 ) | ( ~n8063 & n8064 ) ;
  assign n8066 = ( ~n8044 & n8060 ) | ( ~n8044 & n8065 ) | ( n8060 & n8065 ) ;
  assign n8067 = ( n8044 & n8060 ) | ( n8044 & n8065 ) | ( n8060 & n8065 ) ;
  assign n8068 = ( n8044 & n8066 ) | ( n8044 & ~n8067 ) | ( n8066 & ~n8067 ) ;
  assign n8069 = ( ~n8047 & n8049 ) | ( ~n8047 & n8068 ) | ( n8049 & n8068 ) ;
  assign n8070 = ( n8047 & n8049 ) | ( n8047 & n8068 ) | ( n8049 & n8068 ) ;
  assign n8071 = ( n8047 & n8069 ) | ( n8047 & ~n8070 ) | ( n8069 & ~n8070 ) ;
  assign n8072 = x55 & x63 ;
  assign n8073 = ( n8056 & n8063 ) | ( n8056 & n8072 ) | ( n8063 & n8072 ) ;
  assign n8074 = ( ~n8056 & n8063 ) | ( ~n8056 & n8072 ) | ( n8063 & n8072 ) ;
  assign n8075 = ( n8056 & ~n8073 ) | ( n8056 & n8074 ) | ( ~n8073 & n8074 ) ;
  assign n8076 = x56 & x62 ;
  assign n8077 = x57 & x61 ;
  assign n8078 = x58 & x60 ;
  assign n8079 = ( ~n8076 & n8077 ) | ( ~n8076 & n8078 ) | ( n8077 & n8078 ) ;
  assign n8080 = ( n8076 & n8077 ) | ( n8076 & n8078 ) | ( n8077 & n8078 ) ;
  assign n8081 = ( n8076 & n8079 ) | ( n8076 & ~n8080 ) | ( n8079 & ~n8080 ) ;
  assign n8082 = ( ~n8059 & n8075 ) | ( ~n8059 & n8081 ) | ( n8075 & n8081 ) ;
  assign n8083 = ( n8059 & n8075 ) | ( n8059 & n8081 ) | ( n8075 & n8081 ) ;
  assign n8084 = ( n8059 & n8082 ) | ( n8059 & ~n8083 ) | ( n8082 & ~n8083 ) ;
  assign n8085 = ( n8067 & n8070 ) | ( n8067 & n8084 ) | ( n8070 & n8084 ) ;
  assign n8086 = ( ~n8067 & n8070 ) | ( ~n8067 & n8084 ) | ( n8070 & n8084 ) ;
  assign n8087 = ( n8067 & ~n8085 ) | ( n8067 & n8086 ) | ( ~n8085 & n8086 ) ;
  assign n8088 = x58 & x61 ;
  assign n8089 = x56 & x63 ;
  assign n8090 = ( n8080 & n8088 ) | ( n8080 & n8089 ) | ( n8088 & n8089 ) ;
  assign n8091 = ( ~n8080 & n8088 ) | ( ~n8080 & n8089 ) | ( n8088 & n8089 ) ;
  assign n8092 = ( n8080 & ~n8090 ) | ( n8080 & n8091 ) | ( ~n8090 & n8091 ) ;
  assign n8093 = x59 & x60 ;
  assign n8094 = x57 & x62 ;
  assign n8095 = ( x60 & n8093 ) | ( x60 & n8094 ) | ( n8093 & n8094 ) ;
  assign n8096 = ( x60 & ~n8093 ) | ( x60 & n8094 ) | ( ~n8093 & n8094 ) ;
  assign n8097 = ( n8093 & ~n8095 ) | ( n8093 & n8096 ) | ( ~n8095 & n8096 ) ;
  assign n8098 = ( ~n8073 & n8092 ) | ( ~n8073 & n8097 ) | ( n8092 & n8097 ) ;
  assign n8099 = ( n8073 & n8092 ) | ( n8073 & n8097 ) | ( n8092 & n8097 ) ;
  assign n8100 = ( n8073 & n8098 ) | ( n8073 & ~n8099 ) | ( n8098 & ~n8099 ) ;
  assign n8101 = ( n8083 & n8085 ) | ( n8083 & n8100 ) | ( n8085 & n8100 ) ;
  assign n8102 = ( ~n8083 & n8085 ) | ( ~n8083 & n8100 ) | ( n8085 & n8100 ) ;
  assign n8103 = ( n8083 & ~n8101 ) | ( n8083 & n8102 ) | ( ~n8101 & n8102 ) ;
  assign n8104 = x57 & x63 ;
  assign n8105 = x59 & x61 ;
  assign n8106 = x58 & x62 ;
  assign n8107 = ( ~n8104 & n8105 ) | ( ~n8104 & n8106 ) | ( n8105 & n8106 ) ;
  assign n8108 = ( n8104 & n8105 ) | ( n8104 & n8106 ) | ( n8105 & n8106 ) ;
  assign n8109 = ( n8104 & n8107 ) | ( n8104 & ~n8108 ) | ( n8107 & ~n8108 ) ;
  assign n8110 = ( n8090 & n8095 ) | ( n8090 & n8109 ) | ( n8095 & n8109 ) ;
  assign n8111 = ( ~n8090 & n8095 ) | ( ~n8090 & n8109 ) | ( n8095 & n8109 ) ;
  assign n8112 = ( n8090 & ~n8110 ) | ( n8090 & n8111 ) | ( ~n8110 & n8111 ) ;
  assign n8113 = ( n8099 & n8101 ) | ( n8099 & n8112 ) | ( n8101 & n8112 ) ;
  assign n8114 = ( ~n8099 & n8101 ) | ( ~n8099 & n8112 ) | ( n8101 & n8112 ) ;
  assign n8115 = ( n8099 & ~n8113 ) | ( n8099 & n8114 ) | ( ~n8113 & n8114 ) ;
  assign n8116 = x58 & x63 ;
  assign n8117 = x60 & x61 ;
  assign n8118 = x59 & x62 ;
  assign n8119 = ( x61 & n8117 ) | ( x61 & n8118 ) | ( n8117 & n8118 ) ;
  assign n8120 = ( x61 & ~n8117 ) | ( x61 & n8118 ) | ( ~n8117 & n8118 ) ;
  assign n8121 = ( n8117 & ~n8119 ) | ( n8117 & n8120 ) | ( ~n8119 & n8120 ) ;
  assign n8122 = ( n8108 & n8116 ) | ( n8108 & n8121 ) | ( n8116 & n8121 ) ;
  assign n8123 = ( ~n8108 & n8116 ) | ( ~n8108 & n8121 ) | ( n8116 & n8121 ) ;
  assign n8124 = ( n8108 & ~n8122 ) | ( n8108 & n8123 ) | ( ~n8122 & n8123 ) ;
  assign n8125 = ( ~n8110 & n8113 ) | ( ~n8110 & n8124 ) | ( n8113 & n8124 ) ;
  assign n8126 = ( n8110 & n8113 ) | ( n8110 & n8124 ) | ( n8113 & n8124 ) ;
  assign n8127 = ( n8110 & n8125 ) | ( n8110 & ~n8126 ) | ( n8125 & ~n8126 ) ;
  assign n8128 = x60 & x62 ;
  assign n8129 = x59 & x63 ;
  assign n8130 = ( ~n8119 & n8128 ) | ( ~n8119 & n8129 ) | ( n8128 & n8129 ) ;
  assign n8131 = ( n8119 & n8128 ) | ( n8119 & n8129 ) | ( n8128 & n8129 ) ;
  assign n8132 = ( n8119 & n8130 ) | ( n8119 & ~n8131 ) | ( n8130 & ~n8131 ) ;
  assign n8133 = ( n8122 & n8126 ) | ( n8122 & n8132 ) | ( n8126 & n8132 ) ;
  assign n8134 = ( ~n8122 & n8126 ) | ( ~n8122 & n8132 ) | ( n8126 & n8132 ) ;
  assign n8135 = ( n8122 & ~n8133 ) | ( n8122 & n8134 ) | ( ~n8133 & n8134 ) ;
  assign n8136 = ~x61 & x62 ;
  assign n8137 = x60 & x63 ;
  assign n8138 = n8136 & n8137 ;
  assign n8139 = n8136 | n8137 ;
  assign n8140 = ~n8138 & n8139 ;
  assign n8141 = ( n8131 & n8133 ) | ( n8131 & n8140 ) | ( n8133 & n8140 ) ;
  assign n8142 = ( ~n8131 & n8133 ) | ( ~n8131 & n8140 ) | ( n8133 & n8140 ) ;
  assign n8143 = ( n8131 & ~n8141 ) | ( n8131 & n8142 ) | ( ~n8141 & n8142 ) ;
  assign n8144 = x62 | x63 ;
  assign n8145 = ( ~x61 & x62 ) | ( ~x61 & x63 ) | ( x62 & x63 ) ;
  assign n8146 = ( n8138 & n8144 ) | ( n8138 & ~n8145 ) | ( n8144 & ~n8145 ) ;
  assign n8147 = n8141 | n8146 ;
  assign n8148 = n8141 & n8146 ;
  assign n8149 = n8147 & ~n8148 ;
  assign n8150 = ( x63 & ~n8136 ) | ( x63 & n8148 ) | ( ~n8136 & n8148 ) ;
  assign n8151 = ~x62 & n8148 ;
  assign n8152 = n8150 & ~n8151 ;
  assign n8153 = ( x62 & x63 ) | ( x62 & n8151 ) | ( x63 & n8151 ) ;
  assign y0 = x0 ;
  assign y1 = 1'b0 ;
  assign y2 = n65 ;
  assign y3 = n68 ;
  assign y4 = n72 ;
  assign y5 = n84 ;
  assign y6 = n95 ;
  assign y7 = n107 ;
  assign y8 = n123 ;
  assign y9 = n142 ;
  assign y10 = n162 ;
  assign y11 = n182 ;
  assign y12 = n211 ;
  assign y13 = n236 ;
  assign y14 = n263 ;
  assign y15 = n294 ;
  assign y16 = n325 ;
  assign y17 = n355 ;
  assign y18 = n390 ;
  assign y19 = n427 ;
  assign y20 = n469 ;
  assign y21 = n509 ;
  assign y22 = n553 ;
  assign y23 = n597 ;
  assign y24 = n648 ;
  assign y25 = n696 ;
  assign y26 = n744 ;
  assign y27 = n798 ;
  assign y28 = n854 ;
  assign y29 = n911 ;
  assign y30 = n974 ;
  assign y31 = n1035 ;
  assign y32 = n1096 ;
  assign y33 = n1162 ;
  assign y34 = n1230 ;
  assign y35 = n1298 ;
  assign y36 = n1370 ;
  assign y37 = n1443 ;
  assign y38 = n1520 ;
  assign y39 = n1599 ;
  assign y40 = n1679 ;
  assign y41 = n1758 ;
  assign y42 = n1845 ;
  assign y43 = n1930 ;
  assign y44 = n2017 ;
  assign y45 = n2108 ;
  assign y46 = n2200 ;
  assign y47 = n2292 ;
  assign y48 = n2388 ;
  assign y49 = n2485 ;
  assign y50 = n2586 ;
  assign y51 = n2686 ;
  assign y52 = n2790 ;
  assign y53 = n2893 ;
  assign y54 = n3001 ;
  assign y55 = n3110 ;
  assign y56 = n3225 ;
  assign y57 = n3340 ;
  assign y58 = n3456 ;
  assign y59 = n3570 ;
  assign y60 = n3693 ;
  assign y61 = n3813 ;
  assign y62 = n3934 ;
  assign y63 = n4060 ;
  assign y64 = n4188 ;
  assign y65 = n4313 ;
  assign y66 = n4437 ;
  assign y67 = n4557 ;
  assign y68 = n4676 ;
  assign y69 = n4792 ;
  assign y70 = n4908 ;
  assign y71 = n5019 ;
  assign y72 = n5131 ;
  assign y73 = n5239 ;
  assign y74 = n5347 ;
  assign y75 = n5451 ;
  assign y76 = n5555 ;
  assign y77 = n5655 ;
  assign y78 = n5755 ;
  assign y79 = n5851 ;
  assign y80 = n5946 ;
  assign y81 = n6038 ;
  assign y82 = n6130 ;
  assign y83 = n6217 ;
  assign y84 = n6305 ;
  assign y85 = n6389 ;
  assign y86 = n6473 ;
  assign y87 = n6553 ;
  assign y88 = n6633 ;
  assign y89 = n6708 ;
  assign y90 = n6784 ;
  assign y91 = n6856 ;
  assign y92 = n6928 ;
  assign y93 = n6996 ;
  assign y94 = n7064 ;
  assign y95 = n7127 ;
  assign y96 = n7191 ;
  assign y97 = n7251 ;
  assign y98 = n7311 ;
  assign y99 = n7367 ;
  assign y100 = n7423 ;
  assign y101 = n7475 ;
  assign y102 = n7527 ;
  assign y103 = n7575 ;
  assign y104 = n7623 ;
  assign y105 = n7667 ;
  assign y106 = n7711 ;
  assign y107 = n7751 ;
  assign y108 = n7791 ;
  assign y109 = n7827 ;
  assign y110 = n7863 ;
  assign y111 = n7895 ;
  assign y112 = n7927 ;
  assign y113 = n7955 ;
  assign y114 = n7983 ;
  assign y115 = n8007 ;
  assign y116 = n8031 ;
  assign y117 = n8051 ;
  assign y118 = n8071 ;
  assign y119 = n8087 ;
  assign y120 = n8103 ;
  assign y121 = n8115 ;
  assign y122 = n8127 ;
  assign y123 = n8135 ;
  assign y124 = n8143 ;
  assign y125 = n8149 ;
  assign y126 = n8152 ;
  assign y127 = n8153 ;
endmodule
