module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 ;
  assign n11 = x4 | x7 ;
  assign n12 = x5 | x9 ;
  assign n13 = x8 | n12 ;
  assign n14 = x8 & x9 ;
  assign n15 = x5 | x6 ;
  assign n16 = n14 & n15 ;
  assign n17 = n13 & ~n16 ;
  assign n18 = ~x6 & x9 ;
  assign n19 = x1 & ~x3 ;
  assign n20 = ~n18 & n19 ;
  assign n21 = n17 & n20 ;
  assign n22 = ~x6 & x8 ;
  assign n23 = x5 & ~n22 ;
  assign n24 = ~x1 & x5 ;
  assign n25 = ~x9 & n22 ;
  assign n26 = x8 & ~x9 ;
  assign n27 = x1 & n26 ;
  assign n28 = n25 | n27 ;
  assign n29 = x2 & n28 ;
  assign n30 = ~x5 & n29 ;
  assign n31 = ( x1 & x2 ) | ( x1 & n24 ) | ( x2 & n24 ) ;
  assign n32 = ( n24 & n30 ) | ( n24 & n31 ) | ( n30 & n31 ) ;
  assign n33 = ( x2 & n23 ) | ( x2 & n32 ) | ( n23 & n32 ) ;
  assign n34 = n21 | n33 ;
  assign n35 = ~x2 & x3 ;
  assign n36 = ( x5 & x8 ) | ( x5 & x9 ) | ( x8 & x9 ) ;
  assign n37 = x6 | n36 ;
  assign n38 = ( ~n27 & n36 ) | ( ~n27 & n37 ) | ( n36 & n37 ) ;
  assign n39 = n35 & n38 ;
  assign n40 = ( ~x0 & n34 ) | ( ~x0 & n39 ) | ( n34 & n39 ) ;
  assign n41 = x2 | x3 ;
  assign n42 = ~x1 & x9 ;
  assign n43 = x0 & ~x5 ;
  assign n44 = ( n41 & ~n42 ) | ( n41 & n43 ) | ( ~n42 & n43 ) ;
  assign n45 = ~n41 & n44 ;
  assign n46 = x1 & ~x9 ;
  assign n47 = x6 & ~x8 ;
  assign n48 = n46 & ~n47 ;
  assign n49 = n22 | n46 ;
  assign n50 = ( n45 & n48 ) | ( n45 & ~n49 ) | ( n48 & ~n49 ) ;
  assign n51 = x3 & ~x5 ;
  assign n52 = x0 & n51 ;
  assign n53 = x1 & x6 ;
  assign n54 = x3 & ~x9 ;
  assign n55 = ( ~x8 & n53 ) | ( ~x8 & n54 ) | ( n53 & n54 ) ;
  assign n56 = x8 | n55 ;
  assign n57 = ~x2 & x6 ;
  assign n58 = ~x8 & n57 ;
  assign n59 = ( n52 & ~n56 ) | ( n52 & n58 ) | ( ~n56 & n58 ) ;
  assign n60 = n52 & ~n59 ;
  assign n61 = x6 & ~n12 ;
  assign n62 = ( ~x0 & x3 ) | ( ~x0 & n61 ) | ( x3 & n61 ) ;
  assign n63 = ~n56 & n62 ;
  assign n64 = ( ~n29 & n60 ) | ( ~n29 & n63 ) | ( n60 & n63 ) ;
  assign n65 = n50 | n64 ;
  assign n66 = n40 | n65 ;
  assign n67 = x0 | x3 ;
  assign n68 = x1 & x5 ;
  assign n69 = ( ~x1 & x8 ) | ( ~x1 & n68 ) | ( x8 & n68 ) ;
  assign n70 = ( x9 & n24 ) | ( x9 & n69 ) | ( n24 & n69 ) ;
  assign n71 = n67 | n70 ;
  assign n72 = x2 & x3 ;
  assign n73 = ( x3 & n12 ) | ( x3 & n72 ) | ( n12 & n72 ) ;
  assign n74 = x1 | n73 ;
  assign n75 = ( x5 & x8 ) | ( x5 & ~x9 ) | ( x8 & ~x9 ) ;
  assign n76 = ( x2 & ~n26 ) | ( x2 & n75 ) | ( ~n26 & n75 ) ;
  assign n77 = ( x2 & n74 ) | ( x2 & n76 ) | ( n74 & n76 ) ;
  assign n78 = x6 | n11 ;
  assign n79 = n77 & ~n78 ;
  assign n80 = x1 & ~n13 ;
  assign n81 = ( ~n14 & n72 ) | ( ~n14 & n80 ) | ( n72 & n80 ) ;
  assign n82 = x0 & ~x3 ;
  assign n83 = x0 & ~x1 ;
  assign n84 = ( ~n81 & n82 ) | ( ~n81 & n83 ) | ( n82 & n83 ) ;
  assign n85 = ( ~n71 & n79 ) | ( ~n71 & n84 ) | ( n79 & n84 ) ;
  assign n86 = ( ~n11 & n66 ) | ( ~n11 & n85 ) | ( n66 & n85 ) ;
  assign n87 = x2 | n14 ;
  assign n88 = x1 & ~n43 ;
  assign n89 = ( x1 & n87 ) | ( x1 & n88 ) | ( n87 & n88 ) ;
  assign n90 = x9 & ~n89 ;
  assign n91 = ~x0 & x8 ;
  assign n92 = x3 | x4 ;
  assign n93 = n15 | n92 ;
  assign n94 = x2 | n93 ;
  assign n95 = n91 | n94 ;
  assign n96 = ( ~x9 & n89 ) | ( ~x9 & n95 ) | ( n89 & n95 ) ;
  assign n97 = x0 | x1 ;
  assign n98 = n41 | n97 ;
  assign n99 = ( ~x6 & x9 ) | ( ~x6 & n98 ) | ( x9 & n98 ) ;
  assign n100 = x4 & ~x7 ;
  assign n101 = ~n98 & n100 ;
  assign n102 = ~x5 & x6 ;
  assign n103 = x5 & ~x6 ;
  assign n104 = ( n101 & n102 ) | ( n101 & n103 ) | ( n102 & n103 ) ;
  assign n105 = ( n99 & n101 ) | ( n99 & n104 ) | ( n101 & n104 ) ;
  assign n106 = ~x8 & n105 ;
  assign n107 = ( n90 & n96 ) | ( n90 & ~n106 ) | ( n96 & ~n106 ) ;
  assign n108 = n86 | n107 ;
  assign n109 = ~x0 & x3 ;
  assign n110 = x2 & ~x5 ;
  assign n111 = x8 | x9 ;
  assign n112 = x2 | n111 ;
  assign n113 = ( x1 & ~n110 ) | ( x1 & n112 ) | ( ~n110 & n112 ) ;
  assign n114 = n109 | n113 ;
  assign n115 = n58 & n109 ;
  assign n116 = x2 & x9 ;
  assign n117 = ( ~x5 & x8 ) | ( ~x5 & n116 ) | ( x8 & n116 ) ;
  assign n118 = ( ~x8 & n115 ) | ( ~x8 & n117 ) | ( n115 & n117 ) ;
  assign n119 = ~x0 & x9 ;
  assign n120 = ( x8 & ~n54 ) | ( x8 & n119 ) | ( ~n54 & n119 ) ;
  assign n121 = x5 & x6 ;
  assign n122 = n67 & n121 ;
  assign n123 = ( ~n119 & n120 ) | ( ~n119 & n122 ) | ( n120 & n122 ) ;
  assign n124 = ( n114 & ~n118 ) | ( n114 & n123 ) | ( ~n118 & n123 ) ;
  assign n125 = x2 & ~x3 ;
  assign n126 = x0 & ~x9 ;
  assign n127 = n125 | n126 ;
  assign n128 = x1 & ~n51 ;
  assign n129 = ~n127 & n128 ;
  assign n130 = x1 | x2 ;
  assign n131 = x3 & ~n130 ;
  assign n132 = ( n119 & n125 ) | ( n119 & n131 ) | ( n125 & n131 ) ;
  assign n133 = x5 | n132 ;
  assign n134 = x0 | x2 ;
  assign n135 = ~x0 & x5 ;
  assign n136 = x3 | n134 ;
  assign n137 = ( n41 & ~n42 ) | ( n41 & n136 ) | ( ~n42 & n136 ) ;
  assign n138 = ( n134 & n135 ) | ( n134 & n137 ) | ( n135 & n137 ) ;
  assign n139 = ( n132 & n133 ) | ( n132 & n138 ) | ( n133 & n138 ) ;
  assign n140 = ( x8 & n22 ) | ( x8 & ~n139 ) | ( n22 & ~n139 ) ;
  assign n141 = x5 & ~n35 ;
  assign n142 = x6 & ~x9 ;
  assign n143 = ( ~n119 & n141 ) | ( ~n119 & n142 ) | ( n141 & n142 ) ;
  assign n144 = n129 & ~n143 ;
  assign n145 = ( ~n129 & n140 ) | ( ~n129 & n144 ) | ( n140 & n144 ) ;
  assign n146 = x1 & ~x5 ;
  assign n147 = ~n82 & n146 ;
  assign n148 = x2 | x9 ;
  assign n149 = x0 & ~n148 ;
  assign n150 = x3 & ~n24 ;
  assign n151 = ( n116 & n149 ) | ( n116 & n150 ) | ( n149 & n150 ) ;
  assign n152 = x6 | n151 ;
  assign n153 = ( x2 & ~n97 ) | ( x2 & n116 ) | ( ~n97 & n116 ) ;
  assign n154 = n74 | n153 ;
  assign n155 = ( n147 & ~n152 ) | ( n147 & n154 ) | ( ~n152 & n154 ) ;
  assign n156 = x8 | n155 ;
  assign n157 = ( n124 & n145 ) | ( n124 & ~n156 ) | ( n145 & ~n156 ) ;
  assign n158 = ~n11 & n157 ;
  assign n159 = ( x7 & n11 ) | ( x7 & n98 ) | ( n11 & n98 ) ;
  assign n160 = n121 & ~n159 ;
  assign n161 = x2 & ~n97 ;
  assign n162 = n14 | n93 ;
  assign n163 = n161 & ~n162 ;
  assign n164 = ( x8 & n160 ) | ( x8 & n163 ) | ( n160 & n163 ) ;
  assign n165 = n11 & ~n164 ;
  assign n166 = ( n108 & n158 ) | ( n108 & n165 ) | ( n158 & n165 ) ;
  assign n167 = ~x8 & x9 ;
  assign n168 = x3 | x5 ;
  assign n169 = ( x9 & n167 ) | ( x9 & n168 ) | ( n167 & n168 ) ;
  assign n170 = x1 & x3 ;
  assign n171 = x2 | n170 ;
  assign n172 = ( ~x5 & n14 ) | ( ~x5 & n47 ) | ( n14 & n47 ) ;
  assign n173 = ( x2 & n170 ) | ( x2 & ~n172 ) | ( n170 & ~n172 ) ;
  assign n174 = ( n138 & ~n171 ) | ( n138 & n173 ) | ( ~n171 & n173 ) ;
  assign n175 = ( x6 & ~n169 ) | ( x6 & n174 ) | ( ~n169 & n174 ) ;
  assign n176 = ( x2 & ~n111 ) | ( x2 & n130 ) | ( ~n111 & n130 ) ;
  assign n177 = x5 & ~n176 ;
  assign n178 = x5 & ~x9 ;
  assign n179 = x0 & x1 ;
  assign n180 = n178 & n179 ;
  assign n181 = ~x5 & x8 ;
  assign n182 = ~x3 & n70 ;
  assign n183 = ( x3 & ~n181 ) | ( x3 & n182 ) | ( ~n181 & n182 ) ;
  assign n184 = n83 & ~n183 ;
  assign n185 = ( ~n177 & n180 ) | ( ~n177 & n184 ) | ( n180 & n184 ) ;
  assign n186 = ( x6 & ~n169 ) | ( x6 & n185 ) | ( ~n169 & n185 ) ;
  assign n187 = n175 & ~n186 ;
  assign n188 = ( x3 & n89 ) | ( x3 & ~n102 ) | ( n89 & ~n102 ) ;
  assign n189 = ( x3 & n26 ) | ( x3 & n89 ) | ( n26 & n89 ) ;
  assign n190 = ~n188 & n189 ;
  assign n191 = n11 | n103 ;
  assign n192 = ( n11 & n20 ) | ( n11 & n191 ) | ( n20 & n191 ) ;
  assign n193 = x2 | n12 ;
  assign n194 = x6 | x8 ;
  assign n195 = ~x1 & n194 ;
  assign n196 = ( n147 & ~n193 ) | ( n147 & n195 ) | ( ~n193 & n195 ) ;
  assign n197 = x9 & n68 ;
  assign n198 = ( n72 & ~n136 ) | ( n72 & n197 ) | ( ~n136 & n197 ) ;
  assign n199 = n196 | n198 ;
  assign n200 = ( x8 & n22 ) | ( x8 & ~n134 ) | ( n22 & ~n134 ) ;
  assign n201 = ~n54 & n200 ;
  assign n202 = n199 & ~n201 ;
  assign n203 = ( ~n190 & n192 ) | ( ~n190 & n202 ) | ( n192 & n202 ) ;
  assign n204 = n190 | n203 ;
  assign n205 = x5 | n194 ;
  assign n206 = ( ~x0 & n114 ) | ( ~x0 & n205 ) | ( n114 & n205 ) ;
  assign n207 = ~n17 & n83 ;
  assign n208 = ( n25 & n125 ) | ( n25 & n207 ) | ( n125 & n207 ) ;
  assign n209 = ( ~n114 & n206 ) | ( ~n114 & n208 ) | ( n206 & n208 ) ;
  assign n210 = n204 | n209 ;
  assign n211 = n187 | n210 ;
  assign n212 = n66 & ~n94 ;
  assign n213 = ( n13 & n99 ) | ( n13 & n142 ) | ( n99 & n142 ) ;
  assign n214 = ( x4 & ~n13 ) | ( x4 & n213 ) | ( ~n13 & n213 ) ;
  assign n215 = x7 & ~n163 ;
  assign n216 = n214 | n215 ;
  assign n217 = n211 & ~n216 ;
  assign n218 = ( n211 & n212 ) | ( n211 & n217 ) | ( n212 & n217 ) ;
  assign n219 = x0 & x7 ;
  assign n220 = n89 & n219 ;
  assign n221 = ( x0 & x8 ) | ( x0 & x9 ) | ( x8 & x9 ) ;
  assign n222 = ( x0 & n46 ) | ( x0 & ~n221 ) | ( n46 & ~n221 ) ;
  assign n223 = ~n179 & n222 ;
  assign n224 = ( ~n94 & n220 ) | ( ~n94 & n223 ) | ( n220 & n223 ) ;
  assign n225 = n101 & ~n172 ;
  assign n226 = ( n86 & ~n224 ) | ( n86 & n225 ) | ( ~n224 & n225 ) ;
  assign n227 = n224 | n226 ;
  assign n228 = ( x8 & n57 ) | ( x8 & n91 ) | ( n57 & n91 ) ;
  assign n229 = ( x1 & n111 ) | ( x1 & n228 ) | ( n111 & n228 ) ;
  assign n230 = ( x0 & x2 ) | ( x0 & x9 ) | ( x2 & x9 ) ;
  assign n231 = ( x9 & ~n15 ) | ( x9 & n230 ) | ( ~n15 & n230 ) ;
  assign n232 = ( ~x2 & n43 ) | ( ~x2 & n126 ) | ( n43 & n126 ) ;
  assign n233 = ( ~n88 & n231 ) | ( ~n88 & n232 ) | ( n231 & n232 ) ;
  assign n234 = ( ~n111 & n229 ) | ( ~n111 & n233 ) | ( n229 & n233 ) ;
  assign n235 = ( n11 & ~n121 ) | ( n11 & n159 ) | ( ~n121 & n159 ) ;
  assign n236 = ( n159 & ~n234 ) | ( n159 & n235 ) | ( ~n234 & n235 ) ;
  assign n237 = x0 & ~x6 ;
  assign n238 = n148 | n194 ;
  assign n239 = ~n128 & n238 ;
  assign n240 = ( x2 & ~x8 ) | ( x2 & n181 ) | ( ~x8 & n181 ) ;
  assign n241 = ( ~x3 & n14 ) | ( ~x3 & n116 ) | ( n14 & n116 ) ;
  assign n242 = ( n177 & n240 ) | ( n177 & ~n241 ) | ( n240 & ~n241 ) ;
  assign n243 = n237 & n242 ;
  assign n244 = ( n237 & n239 ) | ( n237 & ~n243 ) | ( n239 & ~n243 ) ;
  assign n245 = x6 & n17 ;
  assign n246 = ( x2 & ~n13 ) | ( x2 & n16 ) | ( ~n13 & n16 ) ;
  assign n247 = ( ~n23 & n245 ) | ( ~n23 & n246 ) | ( n245 & n246 ) ;
  assign n248 = x0 | n247 ;
  assign n249 = ~n244 & n248 ;
  assign n250 = n26 & n72 ;
  assign n251 = ( ~x1 & n201 ) | ( ~x1 & n250 ) | ( n201 & n250 ) ;
  assign n252 = ( x6 & ~x9 ) | ( x6 & n116 ) | ( ~x9 & n116 ) ;
  assign n253 = x3 | n252 ;
  assign n254 = ( n121 & ~n251 ) | ( n121 & n253 ) | ( ~n251 & n253 ) ;
  assign n255 = ( x2 & x3 ) | ( x2 & x6 ) | ( x3 & x6 ) ;
  assign n256 = ( n18 & n24 ) | ( n18 & n237 ) | ( n24 & n237 ) ;
  assign n257 = ( x0 & n68 ) | ( x0 & ~n256 ) | ( n68 & ~n256 ) ;
  assign n258 = ( x4 & n255 ) | ( x4 & ~n257 ) | ( n255 & ~n257 ) ;
  assign n259 = x1 & x2 ;
  assign n260 = ~n26 & n259 ;
  assign n261 = ( n121 & n254 ) | ( n121 & n260 ) | ( n254 & n260 ) ;
  assign n262 = ( n254 & n258 ) | ( n254 & ~n261 ) | ( n258 & ~n261 ) ;
  assign n263 = ~n236 & n262 ;
  assign n264 = ( ~n236 & n249 ) | ( ~n236 & n263 ) | ( n249 & n263 ) ;
  assign n265 = n35 & ~n97 ;
  assign n266 = ( x2 & n101 ) | ( x2 & ~n161 ) | ( n101 & ~n161 ) ;
  assign n267 = ( n160 & n265 ) | ( n160 & n266 ) | ( n265 & n266 ) ;
  assign n268 = n92 & ~n265 ;
  assign n269 = n160 & n268 ;
  assign n286 = x2 & n36 ;
  assign n287 = ~n237 & n286 ;
  assign n288 = n57 | n111 ;
  assign n289 = n24 | n288 ;
  assign n290 = ( ~n111 & n287 ) | ( ~n111 & n289 ) | ( n287 & n289 ) ;
  assign n291 = n179 & n182 ;
  assign n292 = ( ~x3 & n290 ) | ( ~x3 & n291 ) | ( n290 & n291 ) ;
  assign n270 = n25 & n82 ;
  assign n271 = n43 | n47 ;
  assign n272 = x9 | n130 ;
  assign n273 = n271 & ~n272 ;
  assign n274 = ( ~n31 & n270 ) | ( ~n31 & n273 ) | ( n270 & n273 ) ;
  assign n275 = n111 & n194 ;
  assign n276 = x2 & n135 ;
  assign n277 = ( n57 & ~n275 ) | ( n57 & n276 ) | ( ~n275 & n276 ) ;
  assign n278 = n18 & ~n41 ;
  assign n279 = n277 | n278 ;
  assign n280 = ~x3 & n237 ;
  assign n281 = ( x3 & n13 ) | ( x3 & ~n280 ) | ( n13 & ~n280 ) ;
  assign n282 = ( n89 & n279 ) | ( n89 & n281 ) | ( n279 & n281 ) ;
  assign n283 = ( n201 & n279 ) | ( n201 & n281 ) | ( n279 & n281 ) ;
  assign n284 = n282 & ~n283 ;
  assign n285 = n73 & n234 ;
  assign n293 = ( n284 & n285 ) | ( n284 & ~n292 ) | ( n285 & ~n292 ) ;
  assign n294 = ( n274 & ~n292 ) | ( n274 & n293 ) | ( ~n292 & n293 ) ;
  assign n295 = n292 | n294 ;
  assign n296 = x8 | n93 ;
  assign n297 = x7 & ~n148 ;
  assign n298 = ( n161 & ~n296 ) | ( n161 & n297 ) | ( ~n296 & n297 ) ;
  assign n299 = n101 | n298 ;
  assign n300 = x7 | n121 ;
  assign n301 = ( ~n215 & n299 ) | ( ~n215 & n300 ) | ( n299 & n300 ) ;
  assign n302 = n224 | n301 ;
  assign n303 = n11 & ~n302 ;
  assign n304 = ( n295 & n302 ) | ( n295 & ~n303 ) | ( n302 & ~n303 ) ;
  assign n305 = ( n26 & ~n97 ) | ( n26 & n167 ) | ( ~n97 & n167 ) ;
  assign n306 = n134 & n272 ;
  assign n307 = ( n223 & ~n305 ) | ( n223 & n306 ) | ( ~n305 & n306 ) ;
  assign n308 = n93 | n307 ;
  assign n309 = x2 | n219 ;
  assign n310 = ~n308 & n309 ;
  assign n311 = ( ~n15 & n101 ) | ( ~n15 & n310 ) | ( n101 & n310 ) ;
  assign n312 = ( x6 & n75 ) | ( x6 & n167 ) | ( n75 & n167 ) ;
  assign n313 = n19 & n69 ;
  assign n314 = ( n51 & ~n312 ) | ( n51 & n313 ) | ( ~n312 & n313 ) ;
  assign n315 = ( ~x6 & n87 ) | ( ~x6 & n97 ) | ( n87 & n97 ) ;
  assign n316 = ~x6 & n97 ;
  assign n317 = n40 & ~n316 ;
  assign n318 = ( ~n40 & n315 ) | ( ~n40 & n317 ) | ( n315 & n317 ) ;
  assign n319 = n147 | n195 ;
  assign n320 = ( x2 & x9 ) | ( x2 & n319 ) | ( x9 & n319 ) ;
  assign n321 = ( n230 & ~n314 ) | ( n230 & n320 ) | ( ~n314 & n320 ) ;
  assign n322 = n230 & ~n321 ;
  assign n323 = ( n314 & ~n318 ) | ( n314 & n322 ) | ( ~n318 & n322 ) ;
  assign n324 = ( x0 & x1 ) | ( x0 & ~n221 ) | ( x1 & ~n221 ) ;
  assign n325 = ( x9 & ~n97 ) | ( x9 & n111 ) | ( ~n97 & n111 ) ;
  assign n326 = ~x2 & n325 ;
  assign n327 = ~n324 & n326 ;
  assign n328 = ~n15 & n72 ;
  assign n329 = n324 & n328 ;
  assign n330 = ( ~x6 & n111 ) | ( ~x6 & n259 ) | ( n111 & n259 ) ;
  assign n331 = ~x1 & x8 ;
  assign n332 = x2 | n97 ;
  assign n333 = ~x3 & x9 ;
  assign n334 = ( ~x1 & x8 ) | ( ~x1 & n333 ) | ( x8 & n333 ) ;
  assign n335 = ( n331 & n332 ) | ( n331 & ~n334 ) | ( n332 & ~n334 ) ;
  assign n336 = ( ~n111 & n330 ) | ( ~n111 & n335 ) | ( n330 & n335 ) ;
  assign n337 = ( x5 & ~n329 ) | ( x5 & n336 ) | ( ~n329 & n336 ) ;
  assign n338 = n327 | n337 ;
  assign n339 = ~x6 & n68 ;
  assign n340 = ~n14 & n35 ;
  assign n341 = ( ~x0 & n241 ) | ( ~x0 & n260 ) | ( n241 & n260 ) ;
  assign n342 = ~n334 & n341 ;
  assign n343 = ( n339 & n340 ) | ( n339 & n342 ) | ( n340 & n342 ) ;
  assign n344 = ( n14 & ~n111 ) | ( n14 & n134 ) | ( ~n111 & n134 ) ;
  assign n345 = ( x2 & x3 ) | ( x2 & n344 ) | ( x3 & n344 ) ;
  assign n346 = ( x6 & n24 ) | ( x6 & ~n345 ) | ( n24 & ~n345 ) ;
  assign n347 = x1 & ~n12 ;
  assign n348 = ( n91 & n253 ) | ( n91 & n347 ) | ( n253 & n347 ) ;
  assign n349 = n347 & ~n348 ;
  assign n350 = ( n24 & ~n346 ) | ( n24 & n349 ) | ( ~n346 & n349 ) ;
  assign n351 = ( ~n323 & n343 ) | ( ~n323 & n350 ) | ( n343 & n350 ) ;
  assign n352 = ( n323 & n338 ) | ( n323 & ~n351 ) | ( n338 & ~n351 ) ;
  assign n353 = ~n323 & n352 ;
  assign n354 = n11 & ~n311 ;
  assign n355 = ( ~n311 & n353 ) | ( ~n311 & n354 ) | ( n353 & n354 ) ;
  assign n356 = ~x5 & n101 ;
  assign n357 = x6 & ~n51 ;
  assign n358 = ( x6 & n327 ) | ( x6 & n357 ) | ( n327 & n357 ) ;
  assign n359 = n11 & n308 ;
  assign n360 = n358 | n359 ;
  assign n361 = x6 | n329 ;
  assign n362 = ( x3 & ~n24 ) | ( x3 & n54 ) | ( ~n24 & n54 ) ;
  assign n363 = n91 & ~n362 ;
  assign n364 = x1 & ~x8 ;
  assign n365 = ( x5 & n70 ) | ( x5 & ~n364 ) | ( n70 & ~n364 ) ;
  assign n366 = x3 & ~n365 ;
  assign n367 = n363 | n366 ;
  assign n368 = x2 | n333 ;
  assign n369 = n222 | n368 ;
  assign n370 = x1 & ~n193 ;
  assign n371 = ( n367 & n369 ) | ( n367 & ~n370 ) | ( n369 & ~n370 ) ;
  assign n372 = ( x3 & n347 ) | ( x3 & ~n363 ) | ( n347 & ~n363 ) ;
  assign n373 = n119 & n364 ;
  assign n374 = ( x2 & ~n70 ) | ( x2 & n373 ) | ( ~n70 & n373 ) ;
  assign n375 = ~n372 & n374 ;
  assign n376 = ( n361 & n371 ) | ( n361 & ~n375 ) | ( n371 & ~n375 ) ;
  assign n377 = ~n361 & n376 ;
  assign n378 = ~n360 & n377 ;
  assign n379 = ( ~n356 & n360 ) | ( ~n356 & n378 ) | ( n360 & n378 ) ;
  assign n380 = ( x2 & ~n182 ) | ( x2 & n372 ) | ( ~n182 & n372 ) ;
  assign n381 = ~n360 & n380 ;
  assign n382 = ( n104 & ~n329 ) | ( n104 & n381 ) | ( ~n329 & n381 ) ;
  assign n383 = ~n11 & n329 ;
  assign n384 = ( ~n15 & n101 ) | ( ~n15 & n383 ) | ( n101 & n383 ) ;
  assign y0 = ~n166 ;
  assign y1 = n218 ;
  assign y2 = n227 ;
  assign y3 = n264 ;
  assign y4 = n267 ;
  assign y5 = n269 ;
  assign y6 = ~n304 ;
  assign y7 = n355 ;
  assign y8 = n379 ;
  assign y9 = n382 ;
  assign y10 = n384 ;
endmodule
