module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , x1001 , x1002 , x1003 , x1004 , x1005 , x1006 , x1007 , x1008 , x1009 , x1010 , x1011 , x1012 , x1013 , x1014 , x1015 , x1016 , x1017 , x1018 , x1019 , x1020 , x1021 , x1022 , x1023 , x1024 , x1025 , x1026 , x1027 , x1028 , x1029 , x1030 , x1031 , x1032 , x1033 , x1034 , x1035 , x1036 , x1037 , x1038 , x1039 , x1040 , x1041 , x1042 , x1043 , x1044 , x1045 , x1046 , x1047 , x1048 , x1049 , x1050 , x1051 , x1052 , x1053 , x1054 , x1055 , x1056 , x1057 , x1058 , x1059 , x1060 , x1061 , x1062 , x1063 , x1064 , x1065 , x1066 , x1067 , x1068 , x1069 , x1070 , x1071 , x1072 , x1073 , x1074 , x1075 , x1076 , x1077 , x1078 , x1079 , x1080 , x1081 , x1082 , x1083 , x1084 , x1085 , x1086 , x1087 , x1088 , x1089 , x1090 , x1091 , x1092 , x1093 , x1094 , x1095 , x1096 , x1097 , x1098 , x1099 , x1100 , x1101 , x1102 , x1103 , x1104 , x1105 , x1106 , x1107 , x1108 , x1109 , x1110 , x1111 , x1112 , x1113 , x1114 , x1115 , x1116 , x1117 , x1118 , x1119 , x1120 , x1121 , x1122 , x1123 , x1124 , x1125 , x1126 , x1127 , x1128 , x1129 , x1130 , x1131 , x1132 , x1133 , x1134 , x1135 , x1136 , x1137 , x1138 , x1139 , x1140 , x1141 , x1142 , x1143 , x1144 , x1145 , x1146 , x1147 , x1148 , x1149 , x1150 , x1151 , x1152 , x1153 , x1154 , x1155 , x1156 , x1157 , x1158 , x1159 , x1160 , x1161 , x1162 , x1163 , x1164 , x1165 , x1166 , x1167 , x1168 , x1169 , x1170 , x1171 , x1172 , x1173 , x1174 , x1175 , x1176 , x1177 , x1178 , x1179 , x1180 , x1181 , x1182 , x1183 , x1184 , x1185 , x1186 , x1187 , x1188 , x1189 , x1190 , x1191 , x1192 , x1193 , x1194 , x1195 , x1196 , x1197 , x1198 , x1199 , x1200 , x1201 , x1202 , x1203 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 ;
  wire n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 ;
  assign n1205 = x57 | x59 ;
  assign n1206 = x56 | x62 ;
  assign n1207 = n1205 | n1206 ;
  assign n1208 = x55 | n1207 ;
  assign n1209 = x38 | x39 ;
  assign n1210 = x75 | x87 ;
  assign n1211 = n1209 | n1210 ;
  assign n1212 = x54 | x74 ;
  assign n1213 = x92 | n1212 ;
  assign n1214 = n1211 | n1213 ;
  assign n1215 = x100 | n1214 ;
  assign n1216 = ( x55 & x56 ) | ( x55 & x62 ) | ( x56 & x62 ) ;
  assign n1217 = n1205 | n1216 ;
  assign n1218 = ( n1208 & n1215 ) | ( n1208 & n1217 ) | ( n1215 & n1217 ) ;
  assign n1219 = x73 | x82 ;
  assign n1220 = x85 | n1219 ;
  assign n1221 = x66 | n1220 ;
  assign n1222 = x68 | x84 ;
  assign n1223 = x61 & x76 ;
  assign n1224 = x49 & x89 ;
  assign n1225 = ( ~n1222 & n1223 ) | ( ~n1222 & n1224 ) | ( n1223 & n1224 ) ;
  assign n1226 = x45 & x48 ;
  assign n1227 = ( ~n1222 & n1225 ) | ( ~n1222 & n1226 ) | ( n1225 & n1226 ) ;
  assign n1228 = n1222 | n1227 ;
  assign n1229 = x45 | x48 ;
  assign n1230 = x111 & n1229 ;
  assign n1231 = ( ~n1221 & n1228 ) | ( ~n1221 & n1230 ) | ( n1228 & n1230 ) ;
  assign n1232 = n1221 | n1231 ;
  assign n1233 = x111 | n1229 ;
  assign n1234 = x49 | x89 ;
  assign n1235 = x106 | n1234 ;
  assign n1236 = n1233 | n1235 ;
  assign n1237 = x61 | x76 ;
  assign n1238 = x104 | n1237 ;
  assign n1239 = n1236 | n1238 ;
  assign n1240 = n1232 | n1239 ;
  assign n1241 = x36 | x67 ;
  assign n1242 = x63 | x64 ;
  assign n1243 = x65 | n1242 ;
  assign n1244 = ( x103 & x107 ) | ( x103 & n1243 ) | ( x107 & n1243 ) ;
  assign n1245 = ( x63 & x64 ) | ( x63 & x65 ) | ( x64 & x65 ) ;
  assign n1246 = ( ~n1241 & n1244 ) | ( ~n1241 & n1245 ) | ( n1244 & n1245 ) ;
  assign n1247 = n1241 | n1246 ;
  assign n1248 = n1240 | n1247 ;
  assign n1249 = x103 | x107 ;
  assign n1250 = n1243 | n1249 ;
  assign n1251 = x69 | x71 ;
  assign n1252 = x83 | n1251 ;
  assign n1253 = n1250 | n1252 ;
  assign n1254 = n1248 | n1253 ;
  assign n1255 = x50 | x53 ;
  assign n1256 = x60 | n1255 ;
  assign n1257 = x77 | x86 ;
  assign n1258 = x94 | n1257 ;
  assign n1259 = n1256 | n1258 ;
  assign n1260 = x88 | x98 ;
  assign n1261 = n1259 | n1260 ;
  assign n1262 = x97 | x108 ;
  assign n1263 = ( x81 & ~x97 ) | ( x81 & x102 ) | ( ~x97 & x102 ) ;
  assign n1264 = n1262 | n1263 ;
  assign n1265 = x46 | n1264 ;
  assign n1266 = n1261 | n1265 ;
  assign n1267 = n1254 | n1266 ;
  assign n1268 = x47 | x109 ;
  assign n1269 = x110 | n1268 ;
  assign n1270 = x91 | n1269 ;
  assign n1271 = n1267 | n1270 ;
  assign n1272 = x70 | x93 ;
  assign n1273 = x58 | x90 ;
  assign n1274 = n1272 | n1273 ;
  assign n1275 = x35 | x51 ;
  assign n1276 = n1274 | n1275 ;
  assign n1277 = n1271 | n1276 ;
  assign n1278 = x40 | x72 ;
  assign n1279 = x96 | n1278 ;
  assign n1280 = x95 | n1279 ;
  assign n1281 = x32 | n1280 ;
  assign n1282 = n1277 | n1281 ;
  assign n1283 = x215 | x221 ;
  assign n1284 = x216 | n1283 ;
  assign n1285 = x228 | n1284 ;
  assign n1286 = n1282 | n1285 ;
  assign n1287 = n1218 | n1286 ;
  assign n1288 = ~x216 & x833 ;
  assign n1289 = ~x215 & x221 ;
  assign n1290 = n1288 & n1289 ;
  assign n1291 = ~x929 & n1290 ;
  assign n1292 = x153 & ~x216 ;
  assign n1293 = x216 & x265 ;
  assign n1294 = ( ~n1283 & n1292 ) | ( ~n1283 & n1293 ) | ( n1292 & n1293 ) ;
  assign n1295 = ( x215 & n1283 ) | ( x215 & ~n1288 ) | ( n1283 & ~n1288 ) ;
  assign n1296 = ~x1144 & n1295 ;
  assign n1297 = ( ~n1291 & n1294 ) | ( ~n1291 & n1296 ) | ( n1294 & n1296 ) ;
  assign n1298 = n1291 | n1297 ;
  assign n1299 = x105 & x228 ;
  assign n1300 = ~n1284 & n1299 ;
  assign n1301 = x95 & ~x479 ;
  assign n1302 = x234 & n1301 ;
  assign n1303 = n1300 & ~n1302 ;
  assign n1304 = n1300 & n1302 ;
  assign n1305 = ( n1298 & n1303 ) | ( n1298 & ~n1304 ) | ( n1303 & ~n1304 ) ;
  assign n1306 = n1287 & ~n1305 ;
  assign n1307 = ~x332 & n1208 ;
  assign n1308 = ~n1306 & n1307 ;
  assign n1309 = n1208 | n1215 ;
  assign n1310 = x74 | x75 ;
  assign n1311 = x100 | n1211 ;
  assign n1312 = x87 | x100 ;
  assign n1313 = n1209 | n1312 ;
  assign n1314 = ( x74 & n1311 ) | ( x74 & n1313 ) | ( n1311 & n1313 ) ;
  assign n1315 = ( x92 & n1310 ) | ( x92 & n1314 ) | ( n1310 & n1314 ) ;
  assign n1316 = x54 | n1315 ;
  assign n1317 = x92 | n1313 ;
  assign n1318 = ( n1310 & n1316 ) | ( n1310 & n1317 ) | ( n1316 & n1317 ) ;
  assign n1319 = x75 | x100 ;
  assign n1320 = x74 | n1319 ;
  assign n1321 = x39 | x87 ;
  assign n1322 = x92 | n1321 ;
  assign n1323 = n1206 | n1322 ;
  assign n1324 = n1320 | n1323 ;
  assign n1325 = x57 & x59 ;
  assign n1326 = x38 | x54 ;
  assign n1327 = x55 | n1326 ;
  assign n1328 = ( ~n1324 & n1325 ) | ( ~n1324 & n1327 ) | ( n1325 & n1327 ) ;
  assign n1329 = n1324 | n1328 ;
  assign n1330 = n1218 & n1329 ;
  assign n1331 = ( n1318 & n1329 ) | ( n1318 & n1330 ) | ( n1329 & n1330 ) ;
  assign n1332 = n1282 | n1331 ;
  assign n1333 = n1309 & n1332 ;
  assign n1334 = x38 | x87 ;
  assign n1335 = ( x38 & x100 ) | ( x38 & n1334 ) | ( x100 & n1334 ) ;
  assign n1336 = ( x39 & n1312 ) | ( x39 & n1335 ) | ( n1312 & n1335 ) ;
  assign n1337 = n1333 | n1336 ;
  assign n1338 = ~x105 & x228 ;
  assign n1339 = n1284 | n1338 ;
  assign n1340 = x55 | n1206 ;
  assign n1341 = x228 | n1340 ;
  assign n1342 = ( x55 & x137 ) | ( x55 & n1341 ) | ( x137 & n1341 ) ;
  assign n1343 = ( n1337 & n1339 ) | ( n1337 & n1342 ) | ( n1339 & n1342 ) ;
  assign n1344 = n1308 & ~n1342 ;
  assign n1345 = ( n1308 & n1343 ) | ( n1308 & n1344 ) | ( n1343 & n1344 ) ;
  assign n1346 = x32 | x40 ;
  assign n1347 = x32 | x96 ;
  assign n1348 = ( x72 & n1346 ) | ( x72 & n1347 ) | ( n1346 & n1347 ) ;
  assign n1349 = ( x95 & n1279 ) | ( x95 & n1348 ) | ( n1279 & n1348 ) ;
  assign n1350 = n1277 | n1349 ;
  assign n1351 = x35 | x58 ;
  assign n1352 = x90 | n1351 ;
  assign n1353 = x35 | x70 ;
  assign n1354 = x90 | n1272 ;
  assign n1355 = ( x58 & x93 ) | ( x58 & n1354 ) | ( x93 & n1354 ) ;
  assign n1356 = ( n1352 & n1353 ) | ( n1352 & n1355 ) | ( n1353 & n1355 ) ;
  assign n1357 = ( x51 & n1274 ) | ( x51 & n1356 ) | ( n1274 & n1356 ) ;
  assign n1358 = ( n1271 & n1276 ) | ( n1271 & n1357 ) | ( n1276 & n1357 ) ;
  assign n1359 = n1281 | n1358 ;
  assign n1360 = n1350 & n1359 ;
  assign n1361 = x91 & ~n1269 ;
  assign n1362 = ~n1267 & n1361 ;
  assign n1363 = n1276 | n1281 ;
  assign n1364 = n1362 | n1363 ;
  assign n1365 = x94 | n1260 ;
  assign n1366 = x50 & x53 ;
  assign n1367 = x77 & x86 ;
  assign n1368 = ( ~n1365 & n1366 ) | ( ~n1365 & n1367 ) | ( n1366 & n1367 ) ;
  assign n1369 = n1365 | n1368 ;
  assign n1370 = ( x60 & n1255 ) | ( x60 & n1257 ) | ( n1255 & n1257 ) ;
  assign n1371 = n1265 | n1370 ;
  assign n1372 = n1369 | n1371 ;
  assign n1373 = x46 | n1257 ;
  assign n1374 = n1256 | n1373 ;
  assign n1375 = ( x81 & x97 ) | ( x81 & x102 ) | ( x97 & x102 ) ;
  assign n1376 = ( x97 & x108 ) | ( x97 & n1263 ) | ( x108 & n1263 ) ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = ( x88 & x94 ) | ( x88 & x98 ) | ( x94 & x98 ) ;
  assign n1379 = ( n1264 & n1365 ) | ( n1264 & n1378 ) | ( n1365 & n1378 ) ;
  assign n1380 = ( ~n1374 & n1377 ) | ( ~n1374 & n1379 ) | ( n1377 & n1379 ) ;
  assign n1381 = n1374 | n1380 ;
  assign n1382 = n1372 & ~n1381 ;
  assign n1383 = ( n1269 & ~n1372 ) | ( n1269 & n1381 ) | ( ~n1372 & n1381 ) ;
  assign n1384 = ( ~n1254 & n1382 ) | ( ~n1254 & n1383 ) | ( n1382 & n1383 ) ;
  assign n1385 = ( x47 & x109 ) | ( x47 & x110 ) | ( x109 & x110 ) ;
  assign n1386 = ( n1267 & n1269 ) | ( n1267 & n1385 ) | ( n1269 & n1385 ) ;
  assign n1387 = x91 | n1386 ;
  assign n1388 = ( x106 & n1233 ) | ( x106 & n1234 ) | ( n1233 & n1234 ) ;
  assign n1389 = n1239 & ~n1388 ;
  assign n1390 = x67 | x84 ;
  assign n1391 = ( x73 & x82 ) | ( x73 & x85 ) | ( x82 & x85 ) ;
  assign n1392 = ( x66 & n1390 ) | ( x66 & ~n1391 ) | ( n1390 & ~n1391 ) ;
  assign n1393 = ~n1220 & n1392 ;
  assign n1394 = ( n1220 & ~n1391 ) | ( n1220 & n1392 ) | ( ~n1391 & n1392 ) ;
  assign n1395 = ( ~x66 & n1393 ) | ( ~x66 & n1394 ) | ( n1393 & n1394 ) ;
  assign n1396 = x68 | n1395 ;
  assign n1397 = ( x68 & x84 ) | ( x68 & n1221 ) | ( x84 & n1221 ) ;
  assign n1398 = n1239 | n1397 ;
  assign n1399 = n1396 & ~n1398 ;
  assign n1400 = ( x104 & n1236 ) | ( x104 & n1237 ) | ( n1236 & n1237 ) ;
  assign n1401 = ( n1232 & n1239 ) | ( n1232 & n1400 ) | ( n1239 & n1400 ) ;
  assign n1402 = ( n1389 & n1399 ) | ( n1389 & ~n1401 ) | ( n1399 & ~n1401 ) ;
  assign n1403 = ~x36 & n1402 ;
  assign n1404 = n1240 & n1247 ;
  assign n1405 = n1266 | n1404 ;
  assign n1406 = ( x69 & x71 ) | ( x69 & x83 ) | ( x71 & x83 ) ;
  assign n1407 = n1248 | n1406 ;
  assign n1408 = ( n1250 & n1252 ) | ( n1250 & n1407 ) | ( n1252 & n1407 ) ;
  assign n1409 = n1405 | n1408 ;
  assign n1410 = ( x36 & n1253 ) | ( x36 & ~n1402 ) | ( n1253 & ~n1402 ) ;
  assign n1411 = ( n1403 & ~n1409 ) | ( n1403 & n1410 ) | ( ~n1409 & n1410 ) ;
  assign n1412 = ~n1387 & n1411 ;
  assign n1413 = ( n1384 & ~n1387 ) | ( n1384 & n1412 ) | ( ~n1387 & n1412 ) ;
  assign n1414 = n1364 | n1413 ;
  assign n1415 = ~n1360 & n1414 ;
  assign n1416 = x228 | n1415 ;
  assign n1417 = x153 & ~n1416 ;
  assign n1418 = x299 & ~x332 ;
  assign n1419 = ~n1339 & n1418 ;
  assign n1420 = x53 | x60 ;
  assign n1421 = ~x32 & x137 ;
  assign n1422 = x35 | n1421 ;
  assign n1423 = n1420 | n1422 ;
  assign n1424 = n1301 | n1347 ;
  assign n1425 = n1423 | n1424 ;
  assign n1426 = ~x1091 & x1093 ;
  assign n1427 = x829 & x1092 ;
  assign n1428 = ~n1426 & n1427 ;
  assign n1429 = x950 & n1428 ;
  assign n1430 = x1092 & x1093 ;
  assign n1431 = x1091 & n1430 ;
  assign n1432 = ~x833 & x957 ;
  assign n1433 = n1431 & n1432 ;
  assign n1434 = n1429 & ~n1433 ;
  assign n1435 = x1093 & n1434 ;
  assign n1436 = x152 | x161 ;
  assign n1437 = x166 | n1436 ;
  assign n1438 = ~x146 & n1437 ;
  assign n1439 = x210 | n1438 ;
  assign n1440 = x97 & ~n1439 ;
  assign n1441 = n1435 & n1440 ;
  assign n1442 = n1425 | n1441 ;
  assign n1443 = x32 & ~x841 ;
  assign n1444 = ( x210 & n1280 ) | ( x210 & n1443 ) | ( n1280 & n1443 ) ;
  assign n1445 = n1443 & ~n1444 ;
  assign n1446 = x96 | n1301 ;
  assign n1447 = ~x234 & n1446 ;
  assign n1448 = ( n1442 & n1445 ) | ( n1442 & n1447 ) | ( n1445 & n1447 ) ;
  assign n1449 = ( n1416 & ~n1442 ) | ( n1416 & n1448 ) | ( ~n1442 & n1448 ) ;
  assign n1450 = ( n1417 & n1419 ) | ( n1417 & n1449 ) | ( n1419 & n1449 ) ;
  assign n1451 = n1339 & n1418 ;
  assign n1452 = n1298 & n1451 ;
  assign n1453 = n1309 | n1452 ;
  assign n1454 = ~x224 & x833 ;
  assign n1455 = x222 | x223 ;
  assign n1456 = ( x223 & ~n1454 ) | ( x223 & n1455 ) | ( ~n1454 & n1455 ) ;
  assign n1457 = x1144 & n1456 ;
  assign n1458 = x299 | x332 ;
  assign n1459 = x222 & ~x223 ;
  assign n1460 = n1454 & n1459 ;
  assign n1461 = x929 | n1458 ;
  assign n1462 = ( n1458 & n1460 ) | ( n1458 & n1461 ) | ( n1460 & n1461 ) ;
  assign n1463 = x224 & ~n1455 ;
  assign n1464 = ~x265 & n1463 ;
  assign n1465 = ( ~n1457 & n1462 ) | ( ~n1457 & n1464 ) | ( n1462 & n1464 ) ;
  assign n1466 = n1457 | n1465 ;
  assign n1467 = x224 | n1455 ;
  assign n1468 = ~x198 & n1443 ;
  assign n1469 = n1467 | n1468 ;
  assign n1470 = n1447 | n1469 ;
  assign n1471 = ~x142 & x189 ;
  assign n1472 = x144 | x174 ;
  assign n1473 = ( ~x142 & n1471 ) | ( ~x142 & n1472 ) | ( n1471 & n1472 ) ;
  assign n1474 = x198 | n1473 ;
  assign n1475 = x97 | n1474 ;
  assign n1476 = ( ~n1435 & n1474 ) | ( ~n1435 & n1475 ) | ( n1474 & n1475 ) ;
  assign n1477 = ( n1425 & n1475 ) | ( n1425 & ~n1476 ) | ( n1475 & ~n1476 ) ;
  assign n1478 = ~n1470 & n1477 ;
  assign n1479 = n1466 | n1478 ;
  assign n1480 = ~n1360 & n1479 ;
  assign n1481 = n1266 & ~n1381 ;
  assign n1482 = x46 & ~n1264 ;
  assign n1483 = ~n1261 & n1482 ;
  assign n1484 = ( ~n1254 & n1481 ) | ( ~n1254 & n1483 ) | ( n1481 & n1483 ) ;
  assign n1485 = n1411 | n1484 ;
  assign n1486 = n1269 & ~n1387 ;
  assign n1487 = ( ~n1387 & n1485 ) | ( ~n1387 & n1486 ) | ( n1485 & n1486 ) ;
  assign n1488 = n1413 | n1487 ;
  assign n1489 = x51 | x93 ;
  assign n1490 = ( n1273 & n1279 ) | ( n1273 & ~n1489 ) | ( n1279 & ~n1489 ) ;
  assign n1491 = n1489 | n1490 ;
  assign n1492 = x32 | x35 ;
  assign n1493 = x225 & n1492 ;
  assign n1494 = ( ~n1362 & n1491 ) | ( ~n1362 & n1493 ) | ( n1491 & n1493 ) ;
  assign n1495 = n1362 | n1494 ;
  assign n1496 = n1488 | n1495 ;
  assign n1497 = x95 & ~n1453 ;
  assign n1498 = ( ~n1453 & n1496 ) | ( ~n1453 & n1497 ) | ( n1496 & n1497 ) ;
  assign n1499 = n1480 & n1498 ;
  assign n1500 = ~n1301 & n1419 ;
  assign n1501 = n1466 & ~n1500 ;
  assign n1502 = ( ~n1416 & n1466 ) | ( ~n1416 & n1501 ) | ( n1466 & n1501 ) ;
  assign n1503 = ( ~n1453 & n1499 ) | ( ~n1453 & n1502 ) | ( n1499 & n1502 ) ;
  assign n1504 = ~n1450 & n1503 ;
  assign n1505 = ( x39 & n1312 ) | ( x39 & ~n1335 ) | ( n1312 & ~n1335 ) ;
  assign n1506 = ~n1336 & n1505 ;
  assign n1507 = ( x75 & n1211 ) | ( x75 & ~n1506 ) | ( n1211 & ~n1506 ) ;
  assign n1508 = n1212 | n1507 ;
  assign n1509 = x100 & x252 ;
  assign n1510 = n1438 | n1509 ;
  assign n1511 = ( ~n1438 & n1508 ) | ( ~n1438 & n1510 ) | ( n1508 & n1510 ) ;
  assign n1512 = n1318 | n1511 ;
  assign n1513 = n1286 | n1512 ;
  assign n1514 = ~n1305 & n1513 ;
  assign n1515 = x100 & ~n1214 ;
  assign n1516 = ~x228 & x299 ;
  assign n1517 = x75 & ~n1516 ;
  assign n1518 = n1515 | n1517 ;
  assign n1519 = ( n1282 & n1318 ) | ( n1282 & n1518 ) | ( n1318 & n1518 ) ;
  assign n1520 = n1518 & ~n1519 ;
  assign n1521 = ( x137 & n1418 ) | ( x137 & ~n1439 ) | ( n1418 & ~n1439 ) ;
  assign n1522 = ( n1418 & n1451 ) | ( n1418 & ~n1521 ) | ( n1451 & ~n1521 ) ;
  assign n1523 = ~x228 & x252 ;
  assign n1524 = ( n1418 & n1438 ) | ( n1418 & n1523 ) | ( n1438 & n1523 ) ;
  assign n1525 = ( ~n1438 & n1522 ) | ( ~n1438 & n1524 ) | ( n1522 & n1524 ) ;
  assign n1526 = ( n1418 & ~n1520 ) | ( n1418 & n1525 ) | ( ~n1520 & n1525 ) ;
  assign n1527 = ~n1514 & n1526 ;
  assign n1528 = x137 | n1302 ;
  assign n1529 = n1474 & ~n1528 ;
  assign n1530 = ( n1302 & n1520 ) | ( n1302 & ~n1529 ) | ( n1520 & ~n1529 ) ;
  assign n1531 = n1215 & n1466 ;
  assign n1532 = n1467 & ~n1531 ;
  assign n1533 = ( n1530 & n1531 ) | ( n1530 & ~n1532 ) | ( n1531 & ~n1532 ) ;
  assign n1534 = ~n1527 & n1533 ;
  assign n1535 = n1208 | n1534 ;
  assign n1536 = ( n1211 & n1213 ) | ( n1211 & ~n1336 ) | ( n1213 & ~n1336 ) ;
  assign n1537 = ~n1318 & n1536 ;
  assign n1538 = n1277 | n1280 ;
  assign n1539 = n1421 & ~n1538 ;
  assign n1540 = ~n1467 & n1539 ;
  assign n1541 = n1466 & n1537 ;
  assign n1542 = ( n1537 & n1540 ) | ( n1537 & n1541 ) | ( n1540 & n1541 ) ;
  assign n1543 = ( n1300 & n1302 ) | ( n1300 & n1539 ) | ( n1302 & n1539 ) ;
  assign n1544 = x299 | n1543 ;
  assign n1545 = x137 | n1286 ;
  assign n1546 = ( n1286 & n1298 ) | ( n1286 & n1300 ) | ( n1298 & n1300 ) ;
  assign n1547 = ( x332 & n1545 ) | ( x332 & ~n1546 ) | ( n1545 & ~n1546 ) ;
  assign n1548 = ~n1508 & n1547 ;
  assign n1549 = ( n1543 & n1544 ) | ( n1543 & n1548 ) | ( n1544 & n1548 ) ;
  assign n1550 = ( n1542 & ~n1544 ) | ( n1542 & n1549 ) | ( ~n1544 & n1549 ) ;
  assign n1551 = n1535 | n1550 ;
  assign n1552 = ( ~n1345 & n1504 ) | ( ~n1345 & n1551 ) | ( n1504 & n1551 ) ;
  assign n1553 = x299 | n1208 ;
  assign n1554 = ( n1218 & n1309 ) | ( n1218 & n1513 ) | ( n1309 & n1513 ) ;
  assign n1555 = n1553 & n1554 ;
  assign n1556 = n1339 | n1555 ;
  assign n1557 = n1317 | n1340 ;
  assign n1558 = ~x228 & n1415 ;
  assign n1559 = ( n1301 & ~n1350 ) | ( n1301 & n1446 ) | ( ~n1350 & n1446 ) ;
  assign n1560 = ( n1299 & n1558 ) | ( n1299 & ~n1559 ) | ( n1558 & ~n1559 ) ;
  assign n1561 = n1557 | n1560 ;
  assign n1562 = x216 | x221 ;
  assign n1563 = x299 & ~n1562 ;
  assign n1564 = ( n1340 & n1561 ) | ( n1340 & n1563 ) | ( n1561 & n1563 ) ;
  assign n1565 = ~n1556 & n1564 ;
  assign n1566 = x939 & n1460 ;
  assign n1567 = x276 & n1463 ;
  assign n1568 = n1566 | n1567 ;
  assign n1569 = x1146 & n1456 ;
  assign n1570 = ( ~n1553 & n1568 ) | ( ~n1553 & n1569 ) | ( n1568 & n1569 ) ;
  assign n1571 = x299 & n1215 ;
  assign n1572 = x299 & ~n1446 ;
  assign n1573 = n1339 | n1350 ;
  assign n1574 = ( x299 & n1572 ) | ( x299 & n1573 ) | ( n1572 & n1573 ) ;
  assign n1575 = n1571 | n1574 ;
  assign n1576 = n1208 | n1575 ;
  assign n1577 = x939 & n1290 ;
  assign n1578 = x216 & ~n1283 ;
  assign n1579 = x216 & ~x276 ;
  assign n1580 = ( n1577 & n1578 ) | ( n1577 & ~n1579 ) | ( n1578 & ~n1579 ) ;
  assign n1581 = n1284 | n1299 ;
  assign n1582 = x1146 & n1295 ;
  assign n1583 = x154 & ~n1581 ;
  assign n1584 = ( n1581 & ~n1582 ) | ( n1581 & n1583 ) | ( ~n1582 & n1583 ) ;
  assign n1585 = ( ~n1570 & n1580 ) | ( ~n1570 & n1584 ) | ( n1580 & n1584 ) ;
  assign n1586 = ~n1580 & n1585 ;
  assign n1587 = ( n1570 & n1576 ) | ( n1570 & ~n1586 ) | ( n1576 & ~n1586 ) ;
  assign n1588 = n1300 & n1301 ;
  assign n1589 = n1576 & ~n1588 ;
  assign n1590 = ( ~n1215 & n1301 ) | ( ~n1215 & n1559 ) | ( n1301 & n1559 ) ;
  assign n1591 = ~n1467 & n1590 ;
  assign n1592 = n1553 | n1591 ;
  assign n1593 = ~n1589 & n1592 ;
  assign n1594 = ~x239 & n1593 ;
  assign n1595 = ( n1587 & n1593 ) | ( n1587 & ~n1594 ) | ( n1593 & ~n1594 ) ;
  assign n1596 = ~n1565 & n1595 ;
  assign n1597 = x235 & n1593 ;
  assign n1598 = ~x235 & n1593 ;
  assign n1599 = n1460 & ~n1553 ;
  assign n1600 = n1290 & n1553 ;
  assign n1601 = ( x927 & n1599 ) | ( x927 & n1600 ) | ( n1599 & n1600 ) ;
  assign n1602 = n1599 | n1600 ;
  assign n1603 = n1455 | n1553 ;
  assign n1604 = ~n1283 & n1553 ;
  assign n1605 = n1603 & ~n1604 ;
  assign n1606 = ~n1602 & n1605 ;
  assign n1607 = n1463 & ~n1553 ;
  assign n1608 = n1553 & n1578 ;
  assign n1609 = ( ~x274 & n1607 ) | ( ~x274 & n1608 ) | ( n1607 & n1608 ) ;
  assign n1610 = x1145 | n1609 ;
  assign n1611 = ( n1606 & n1609 ) | ( n1606 & n1610 ) | ( n1609 & n1610 ) ;
  assign n1612 = n1601 | n1611 ;
  assign n1613 = x151 | n1309 ;
  assign n1614 = ~x215 & n1563 ;
  assign n1615 = ( ~n1560 & n1613 ) | ( ~n1560 & n1614 ) | ( n1613 & n1614 ) ;
  assign n1616 = ~n1613 & n1615 ;
  assign n1617 = n1555 & ~n1581 ;
  assign n1618 = ( ~x151 & n1616 ) | ( ~x151 & n1617 ) | ( n1616 & n1617 ) ;
  assign n1619 = n1612 | n1618 ;
  assign n1620 = ( n1597 & ~n1598 ) | ( n1597 & n1619 ) | ( ~n1598 & n1619 ) ;
  assign n1621 = n1575 & ~n1588 ;
  assign n1622 = x299 | n1591 ;
  assign n1623 = ~n1621 & n1622 ;
  assign n1624 = ~x238 & n1623 ;
  assign n1625 = ~x1143 & n1295 ;
  assign n1626 = ~x944 & n1290 ;
  assign n1627 = x216 & ~x264 ;
  assign n1628 = ( n1578 & n1626 ) | ( n1578 & ~n1627 ) | ( n1626 & ~n1627 ) ;
  assign n1629 = n1625 | n1628 ;
  assign n1630 = n1300 & ~n1301 ;
  assign n1631 = x284 & n1630 ;
  assign n1632 = x146 & ~n1581 ;
  assign n1633 = ( n1581 & ~n1631 ) | ( n1581 & n1632 ) | ( ~n1631 & n1632 ) ;
  assign n1634 = ~n1629 & n1633 ;
  assign n1635 = n1513 & ~n1634 ;
  assign n1636 = x284 & ~n1513 ;
  assign n1637 = ( n1571 & n1635 ) | ( n1571 & n1636 ) | ( n1635 & n1636 ) ;
  assign n1638 = x944 & ~n1208 ;
  assign n1639 = ( n1208 & n1599 ) | ( n1208 & ~n1638 ) | ( n1599 & ~n1638 ) ;
  assign n1640 = n1637 | n1639 ;
  assign n1641 = ~x1143 & n1456 ;
  assign n1642 = x224 & x264 ;
  assign n1643 = ~x224 & x284 ;
  assign n1644 = ( ~n1455 & n1642 ) | ( ~n1455 & n1643 ) | ( n1642 & n1643 ) ;
  assign n1645 = ( ~n1622 & n1641 ) | ( ~n1622 & n1644 ) | ( n1641 & n1644 ) ;
  assign n1646 = n1640 | n1645 ;
  assign n1647 = n1624 | n1646 ;
  assign n1648 = x238 & n1208 ;
  assign n1649 = ( n1208 & ~n1588 ) | ( n1208 & n1648 ) | ( ~n1588 & n1648 ) ;
  assign n1650 = x284 | n1287 ;
  assign n1651 = n1287 & n1634 ;
  assign n1652 = ( n1649 & ~n1650 ) | ( n1649 & n1651 ) | ( ~n1650 & n1651 ) ;
  assign n1653 = ~n1285 & n1415 ;
  assign n1654 = x284 & n1653 ;
  assign n1655 = ~n1215 & n1574 ;
  assign n1656 = n1634 | n1653 ;
  assign n1657 = ( n1654 & n1655 ) | ( n1654 & ~n1656 ) | ( n1655 & ~n1656 ) ;
  assign n1658 = ~n1652 & n1657 ;
  assign n1659 = ( n1647 & ~n1652 ) | ( n1647 & n1658 ) | ( ~n1652 & n1658 ) ;
  assign n1660 = ( x249 & n1589 ) | ( x249 & n1592 ) | ( n1589 & n1592 ) ;
  assign n1661 = x932 & n1460 ;
  assign n1662 = x277 & n1463 ;
  assign n1663 = ( ~x1142 & n1455 ) | ( ~x1142 & n1460 ) | ( n1455 & n1460 ) ;
  assign n1664 = ( ~n1661 & n1662 ) | ( ~n1661 & n1663 ) | ( n1662 & n1663 ) ;
  assign n1665 = n1592 | n1664 ;
  assign n1666 = n1467 | n1553 ;
  assign n1667 = n1590 & ~n1666 ;
  assign n1668 = ( ~n1565 & n1666 ) | ( ~n1565 & n1667 ) | ( n1666 & n1667 ) ;
  assign n1669 = x262 & ~n1668 ;
  assign n1670 = ( ~n1660 & n1665 ) | ( ~n1660 & n1669 ) | ( n1665 & n1669 ) ;
  assign n1671 = ~x1142 & n1295 ;
  assign n1672 = ~x932 & n1290 ;
  assign n1673 = x262 | n1672 ;
  assign n1674 = ( n1630 & n1672 ) | ( n1630 & n1673 ) | ( n1672 & n1673 ) ;
  assign n1675 = n1671 | n1674 ;
  assign n1676 = n1576 & n1675 ;
  assign n1677 = x172 & ~n1581 ;
  assign n1678 = x216 & x277 ;
  assign n1679 = ( ~n1565 & n1677 ) | ( ~n1565 & n1678 ) | ( n1677 & n1678 ) ;
  assign n1680 = ~n1283 & n1679 ;
  assign n1681 = ( n1576 & n1676 ) | ( n1576 & n1680 ) | ( n1676 & n1680 ) ;
  assign n1682 = n1670 | n1681 ;
  assign n1683 = x861 & n1565 ;
  assign n1684 = x216 & ~x270 ;
  assign n1685 = ~x935 & n1290 ;
  assign n1686 = ( n1578 & ~n1684 ) | ( n1578 & n1685 ) | ( ~n1684 & n1685 ) ;
  assign n1687 = x171 & ~n1581 ;
  assign n1688 = ~x1141 & n1295 ;
  assign n1689 = ( ~n1686 & n1687 ) | ( ~n1686 & n1688 ) | ( n1687 & n1688 ) ;
  assign n1690 = n1686 | n1689 ;
  assign n1691 = x861 | n1301 ;
  assign n1692 = n1300 & ~n1691 ;
  assign n1693 = n1690 | n1692 ;
  assign n1694 = n1207 & n1693 ;
  assign n1695 = ( n1207 & ~n1287 ) | ( n1207 & n1694 ) | ( ~n1287 & n1694 ) ;
  assign n1696 = x241 & ~n1695 ;
  assign n1697 = ( n1593 & n1695 ) | ( n1593 & ~n1696 ) | ( n1695 & ~n1696 ) ;
  assign n1698 = x55 | x299 ;
  assign n1699 = ~n1467 & n1691 ;
  assign n1700 = ~x270 & n1463 ;
  assign n1701 = n1699 | n1700 ;
  assign n1702 = ~x935 & n1460 ;
  assign n1703 = ( x1141 & n1455 ) | ( x1141 & n1460 ) | ( n1455 & n1460 ) ;
  assign n1704 = ~n1702 & n1703 ;
  assign n1705 = ( ~n1698 & n1701 ) | ( ~n1698 & n1704 ) | ( n1701 & n1704 ) ;
  assign n1706 = ~n1697 & n1705 ;
  assign n1707 = x55 | n1215 ;
  assign n1708 = n1622 & ~n1707 ;
  assign n1709 = ~n1284 & n1560 ;
  assign n1710 = n1708 & ~n1709 ;
  assign n1711 = n1555 & ~n1693 ;
  assign n1712 = n1574 & n1690 ;
  assign n1713 = ( n1710 & n1711 ) | ( n1710 & ~n1712 ) | ( n1711 & ~n1712 ) ;
  assign n1714 = ( ~n1697 & n1706 ) | ( ~n1697 & n1713 ) | ( n1706 & n1713 ) ;
  assign n1715 = n1683 | n1714 ;
  assign n1716 = x170 | n1299 ;
  assign n1717 = x869 & n1299 ;
  assign n1718 = ( n1284 & n1716 ) | ( n1284 & ~n1717 ) | ( n1716 & ~n1717 ) ;
  assign n1719 = n1589 & ~n1718 ;
  assign n1720 = ~n1565 & n1719 ;
  assign n1721 = ( ~x282 & n1607 ) | ( ~x282 & n1608 ) | ( n1607 & n1608 ) ;
  assign n1722 = x1140 | n1721 ;
  assign n1723 = ( n1606 & n1721 ) | ( n1606 & n1722 ) | ( n1721 & n1722 ) ;
  assign n1724 = ( x921 & n1599 ) | ( x921 & n1600 ) | ( n1599 & n1600 ) ;
  assign n1725 = x248 | n1724 ;
  assign n1726 = ( n1593 & n1724 ) | ( n1593 & n1725 ) | ( n1724 & n1725 ) ;
  assign n1727 = n1723 | n1726 ;
  assign n1728 = x869 | n1727 ;
  assign n1729 = ( ~n1668 & n1727 ) | ( ~n1668 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1730 = n1720 | n1729 ;
  assign n1731 = ~x920 & n1290 ;
  assign n1732 = x216 & ~x281 ;
  assign n1733 = ( n1578 & n1731 ) | ( n1578 & ~n1732 ) | ( n1731 & ~n1732 ) ;
  assign n1734 = ~x1139 & n1295 ;
  assign n1735 = x148 & ~n1581 ;
  assign n1736 = ( ~n1733 & n1734 ) | ( ~n1733 & n1735 ) | ( n1734 & n1735 ) ;
  assign n1737 = ( n1589 & n1733 ) | ( n1589 & n1736 ) | ( n1733 & n1736 ) ;
  assign n1738 = ~n1565 & n1737 ;
  assign n1739 = ( ~x1139 & n1455 ) | ( ~x1139 & n1460 ) | ( n1455 & n1460 ) ;
  assign n1740 = x281 & n1463 ;
  assign n1741 = x920 & n1460 ;
  assign n1742 = ( n1739 & n1740 ) | ( n1739 & ~n1741 ) | ( n1740 & ~n1741 ) ;
  assign n1743 = ~n1592 & n1742 ;
  assign n1744 = ~x247 & n1593 ;
  assign n1745 = n1743 | n1744 ;
  assign n1746 = n1738 | n1745 ;
  assign n1747 = ~x862 & n1630 ;
  assign n1748 = n1576 & n1747 ;
  assign n1749 = ( x862 & n1668 ) | ( x862 & ~n1748 ) | ( n1668 & ~n1748 ) ;
  assign n1750 = ~n1746 & n1749 ;
  assign n1751 = ~x55 & n1571 ;
  assign n1752 = x55 | x62 ;
  assign n1753 = ~n1215 & n1752 ;
  assign n1754 = ( ~n1512 & n1751 ) | ( ~n1512 & n1753 ) | ( n1751 & n1753 ) ;
  assign n1755 = x877 & n1754 ;
  assign n1756 = x56 | n1755 ;
  assign n1757 = ~n1286 & n1756 ;
  assign n1758 = ~x877 & n1630 ;
  assign n1759 = x169 | n1299 ;
  assign n1760 = ( ~n1581 & n1758 ) | ( ~n1581 & n1759 ) | ( n1758 & n1759 ) ;
  assign n1761 = x216 & ~x269 ;
  assign n1762 = ~x940 & n1290 ;
  assign n1763 = ( n1578 & ~n1761 ) | ( n1578 & n1762 ) | ( ~n1761 & n1762 ) ;
  assign n1764 = ~x1138 & n1295 ;
  assign n1765 = ( ~n1760 & n1763 ) | ( ~n1760 & n1764 ) | ( n1763 & n1764 ) ;
  assign n1766 = n1760 | n1765 ;
  assign n1767 = n1574 & n1766 ;
  assign n1768 = ( n1653 & ~n1757 ) | ( n1653 & n1767 ) | ( ~n1757 & n1767 ) ;
  assign n1769 = ~n1653 & n1768 ;
  assign n1770 = n1555 & n1766 ;
  assign n1771 = n1301 & ~n1467 ;
  assign n1772 = x224 | x299 ;
  assign n1773 = ~x223 & x877 ;
  assign n1774 = n1772 | n1773 ;
  assign n1775 = x222 | x224 ;
  assign n1776 = ( x269 & n1455 ) | ( x269 & n1775 ) | ( n1455 & n1775 ) ;
  assign n1777 = n1774 & ~n1776 ;
  assign n1778 = x1138 & n1456 ;
  assign n1779 = x299 | x940 ;
  assign n1780 = ( x299 & n1460 ) | ( x299 & n1779 ) | ( n1460 & n1779 ) ;
  assign n1781 = ( ~n1777 & n1778 ) | ( ~n1777 & n1780 ) | ( n1778 & n1780 ) ;
  assign n1782 = n1777 | n1781 ;
  assign n1783 = ( ~x299 & n1215 ) | ( ~x299 & n1771 ) | ( n1215 & n1771 ) ;
  assign n1784 = ( n1771 & n1782 ) | ( n1771 & n1783 ) | ( n1782 & n1783 ) ;
  assign n1785 = n1555 | n1784 ;
  assign n1786 = x299 & ~x877 ;
  assign n1787 = n1653 & n1786 ;
  assign n1788 = n1559 & n1782 ;
  assign n1789 = ( n1782 & ~n1787 ) | ( n1782 & n1788 ) | ( ~n1787 & n1788 ) ;
  assign n1790 = x96 & ~n1350 ;
  assign n1791 = ~n1467 & n1790 ;
  assign n1792 = ~n1707 & n1791 ;
  assign n1793 = ( ~n1707 & n1789 ) | ( ~n1707 & n1792 ) | ( n1789 & n1792 ) ;
  assign n1794 = ( ~n1770 & n1785 ) | ( ~n1770 & n1793 ) | ( n1785 & n1793 ) ;
  assign n1795 = ( n1757 & ~n1769 ) | ( n1757 & n1794 ) | ( ~n1769 & n1794 ) ;
  assign n1796 = ( ~x246 & n1589 ) | ( ~x246 & n1592 ) | ( n1589 & n1592 ) ;
  assign n1797 = n1287 & n1766 ;
  assign n1798 = x877 | n1287 ;
  assign n1799 = ( n1207 & n1797 ) | ( n1207 & ~n1798 ) | ( n1797 & ~n1798 ) ;
  assign n1800 = ( ~n1589 & n1796 ) | ( ~n1589 & n1799 ) | ( n1796 & n1799 ) ;
  assign n1801 = n1795 & ~n1800 ;
  assign n1802 = x280 & n1578 ;
  assign n1803 = x168 & ~n1299 ;
  assign n1804 = ~x878 & n1299 ;
  assign n1805 = ( ~n1284 & n1803 ) | ( ~n1284 & n1804 ) | ( n1803 & n1804 ) ;
  assign n1806 = ~x1137 & n1295 ;
  assign n1807 = ~x933 & n1290 ;
  assign n1808 = ( ~n1802 & n1806 ) | ( ~n1802 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1809 = ( ~n1802 & n1805 ) | ( ~n1802 & n1808 ) | ( n1805 & n1808 ) ;
  assign n1810 = n1802 | n1809 ;
  assign n1811 = x55 & ~n1810 ;
  assign n1812 = ( n1512 & ~n1810 ) | ( n1512 & n1811 ) | ( ~n1810 & n1811 ) ;
  assign n1813 = n1215 & n1812 ;
  assign n1814 = ~x280 & n1463 ;
  assign n1815 = ( x878 & ~n1467 ) | ( x878 & n1771 ) | ( ~n1467 & n1771 ) ;
  assign n1816 = n1814 | n1815 ;
  assign n1817 = x933 & n1460 ;
  assign n1818 = ( ~n1553 & n1816 ) | ( ~n1553 & n1817 ) | ( n1816 & n1817 ) ;
  assign n1819 = x1137 & n1456 ;
  assign n1820 = ( ~n1553 & n1818 ) | ( ~n1553 & n1819 ) | ( n1818 & n1819 ) ;
  assign n1821 = n1553 | n1820 ;
  assign n1822 = ( ~n1207 & n1588 ) | ( ~n1207 & n1698 ) | ( n1588 & n1698 ) ;
  assign n1823 = ( ~n1588 & n1813 ) | ( ~n1588 & n1822 ) | ( n1813 & n1822 ) ;
  assign n1824 = ( n1813 & n1821 ) | ( n1813 & ~n1823 ) | ( n1821 & ~n1823 ) ;
  assign n1825 = n1754 | n1824 ;
  assign n1826 = n1287 & n1810 ;
  assign n1827 = x878 | n1287 ;
  assign n1828 = ( n1588 & ~n1826 ) | ( n1588 & n1827 ) | ( ~n1826 & n1827 ) ;
  assign n1829 = ( n1824 & n1825 ) | ( n1824 & n1828 ) | ( n1825 & n1828 ) ;
  assign n1830 = n1708 | n1829 ;
  assign n1831 = ~n1653 & n1810 ;
  assign n1832 = ~x878 & n1653 ;
  assign n1833 = ( n1574 & n1831 ) | ( n1574 & n1832 ) | ( n1831 & n1832 ) ;
  assign n1834 = ( n1829 & n1830 ) | ( n1829 & ~n1833 ) | ( n1830 & ~n1833 ) ;
  assign n1835 = ( ~x240 & n1589 ) | ( ~x240 & n1592 ) | ( n1589 & n1592 ) ;
  assign n1836 = n1207 & ~n1828 ;
  assign n1837 = ( ~n1589 & n1835 ) | ( ~n1589 & n1836 ) | ( n1835 & n1836 ) ;
  assign n1838 = n1834 & ~n1837 ;
  assign n1839 = ~x928 & n1460 ;
  assign n1840 = x266 & n1463 ;
  assign n1841 = ( x1136 & n1455 ) | ( x1136 & n1460 ) | ( n1455 & n1460 ) ;
  assign n1842 = ( ~n1839 & n1840 ) | ( ~n1839 & n1841 ) | ( n1840 & n1841 ) ;
  assign n1843 = ~n1592 & n1842 ;
  assign n1844 = x245 | n1843 ;
  assign n1845 = ( n1593 & n1843 ) | ( n1593 & n1844 ) | ( n1843 & n1844 ) ;
  assign n1846 = x266 & n1578 ;
  assign n1847 = x928 & n1290 ;
  assign n1848 = x1136 & n1295 ;
  assign n1849 = ( ~n1846 & n1847 ) | ( ~n1846 & n1848 ) | ( n1847 & n1848 ) ;
  assign n1850 = n1846 | n1849 ;
  assign n1851 = x875 & n1630 ;
  assign n1852 = x166 & ~n1581 ;
  assign n1853 = ( ~n1850 & n1851 ) | ( ~n1850 & n1852 ) | ( n1851 & n1852 ) ;
  assign n1854 = n1850 | n1853 ;
  assign n1855 = n1576 & n1854 ;
  assign n1856 = n1668 & ~n1855 ;
  assign n1857 = x875 | n1668 ;
  assign n1858 = ( n1845 & ~n1856 ) | ( n1845 & n1857 ) | ( ~n1856 & n1857 ) ;
  assign n1859 = x879 | n1301 ;
  assign n1860 = n1300 & ~n1859 ;
  assign n1861 = n1208 & ~n1860 ;
  assign n1862 = ~x244 & n1588 ;
  assign n1863 = n1861 & ~n1862 ;
  assign n1864 = x161 | n1581 ;
  assign n1865 = ~x279 & n1578 ;
  assign n1866 = ~x938 & n1290 ;
  assign n1867 = n1865 | n1866 ;
  assign n1868 = n1864 & ~n1867 ;
  assign n1869 = ~x1135 & n1295 ;
  assign n1870 = n1868 & ~n1869 ;
  assign n1871 = n1287 & n1870 ;
  assign n1872 = x879 & ~n1287 ;
  assign n1873 = ( n1863 & n1871 ) | ( n1863 & n1872 ) | ( n1871 & n1872 ) ;
  assign n1874 = x299 & ~x879 ;
  assign n1875 = n1320 | n1326 ;
  assign n1876 = x92 & ~n1321 ;
  assign n1877 = ~n1875 & n1876 ;
  assign n1878 = ~n1874 & n1877 ;
  assign n1879 = ( ~n1286 & n1877 ) | ( ~n1286 & n1878 ) | ( n1877 & n1878 ) ;
  assign n1880 = ( n1208 & ~n1878 ) | ( n1208 & n1879 ) | ( ~n1878 & n1879 ) ;
  assign n1881 = x244 & ~n1880 ;
  assign n1882 = ( n1623 & n1880 ) | ( n1623 & ~n1881 ) | ( n1880 & ~n1881 ) ;
  assign n1883 = ~n1873 & n1882 ;
  assign n1884 = x299 | x938 ;
  assign n1885 = ( x299 & n1460 ) | ( x299 & n1884 ) | ( n1460 & n1884 ) ;
  assign n1886 = x1135 & n1456 ;
  assign n1887 = ~n1467 & n1859 ;
  assign n1888 = ( ~n1885 & n1886 ) | ( ~n1885 & n1887 ) | ( n1886 & n1887 ) ;
  assign n1889 = x279 & n1463 ;
  assign n1890 = ( ~n1885 & n1888 ) | ( ~n1885 & n1889 ) | ( n1888 & n1889 ) ;
  assign n1891 = n1885 | n1890 ;
  assign n1892 = n1215 & ~n1891 ;
  assign n1893 = ( x299 & n1860 ) | ( x299 & ~n1870 ) | ( n1860 & ~n1870 ) ;
  assign n1894 = n1282 & n1893 ;
  assign n1895 = ( n1215 & n1892 ) | ( n1215 & n1894 ) | ( n1892 & n1894 ) ;
  assign n1896 = n1513 | n1874 ;
  assign n1897 = n1513 & ~n1893 ;
  assign n1898 = ( n1215 & ~n1896 ) | ( n1215 & n1897 ) | ( ~n1896 & n1897 ) ;
  assign n1899 = ~n1895 & n1898 ;
  assign n1900 = ~n1339 & n1415 ;
  assign n1901 = n1893 | n1900 ;
  assign n1902 = ~n1559 & n1874 ;
  assign n1903 = n1900 & ~n1902 ;
  assign n1904 = ~n1313 & n1891 ;
  assign n1905 = ( ~n1313 & n1791 ) | ( ~n1313 & n1904 ) | ( n1791 & n1904 ) ;
  assign n1906 = ( ~n1901 & n1903 ) | ( ~n1901 & n1905 ) | ( n1903 & n1905 ) ;
  assign n1907 = ( ~n1895 & n1899 ) | ( ~n1895 & n1906 ) | ( n1899 & n1906 ) ;
  assign n1908 = ( n1873 & ~n1883 ) | ( n1873 & n1907 ) | ( ~n1883 & n1907 ) ;
  assign n1909 = ~x846 & n1564 ;
  assign n1910 = x152 & x299 ;
  assign n1911 = ( n1285 & n1415 ) | ( n1285 & n1910 ) | ( n1415 & n1910 ) ;
  assign n1912 = n1910 & ~n1911 ;
  assign n1913 = ~x930 & n1460 ;
  assign n1914 = x224 | x846 ;
  assign n1915 = x224 & ~x278 ;
  assign n1916 = ( n1455 & n1914 ) | ( n1455 & ~n1915 ) | ( n1914 & ~n1915 ) ;
  assign n1917 = ~n1913 & n1916 ;
  assign n1918 = ~n1622 & n1917 ;
  assign n1919 = ( n1564 & ~n1912 ) | ( n1564 & n1918 ) | ( ~n1912 & n1918 ) ;
  assign n1920 = n1912 | n1919 ;
  assign n1921 = x299 & n1285 ;
  assign n1922 = x152 | n1283 ;
  assign n1923 = ( n1283 & ~n1581 ) | ( n1283 & n1922 ) | ( ~n1581 & n1922 ) ;
  assign n1924 = x216 & x278 ;
  assign n1925 = ~x930 & n1290 ;
  assign n1926 = ( n1923 & n1924 ) | ( n1923 & ~n1925 ) | ( n1924 & ~n1925 ) ;
  assign n1927 = n1921 & n1926 ;
  assign n1928 = x242 | n1927 ;
  assign n1929 = ( n1623 & n1927 ) | ( n1623 & n1928 ) | ( n1927 & n1928 ) ;
  assign n1930 = n1555 | n1929 ;
  assign n1931 = ( ~n1909 & n1920 ) | ( ~n1909 & n1930 ) | ( n1920 & n1930 ) ;
  assign n1932 = x242 & n1301 ;
  assign n1933 = x846 & ~n1301 ;
  assign n1934 = ( n1300 & n1932 ) | ( n1300 & n1933 ) | ( n1932 & n1933 ) ;
  assign n1935 = n1926 | n1934 ;
  assign n1936 = n1555 & ~n1935 ;
  assign n1937 = x1134 & n1606 ;
  assign n1938 = ( n1606 & n1936 ) | ( n1606 & ~n1937 ) | ( n1936 & ~n1937 ) ;
  assign n1939 = n1931 & ~n1938 ;
  assign n1940 = n1337 | n1360 ;
  assign n1941 = x42 | x44 ;
  assign n1942 = x41 | x101 ;
  assign n1943 = x99 | n1942 ;
  assign n1944 = x113 | n1943 ;
  assign n1945 = x116 | n1944 ;
  assign n1946 = x115 | n1945 ;
  assign n1947 = ( x114 & ~n1941 ) | ( x114 & n1946 ) | ( ~n1941 & n1946 ) ;
  assign n1948 = n1941 | n1947 ;
  assign n1949 = x43 | x52 ;
  assign n1950 = n1948 | n1949 ;
  assign n1951 = x299 & n1438 ;
  assign n1952 = ~x299 & n1473 ;
  assign n1953 = n1951 | n1952 ;
  assign n1954 = n1950 & n1953 ;
  assign n1955 = x129 & x250 ;
  assign n1956 = ~x129 & x250 ;
  assign n1957 = x950 & x1092 ;
  assign n1958 = x824 & n1957 ;
  assign n1959 = ( x950 & n1428 ) | ( x950 & n1958 ) | ( n1428 & n1958 ) ;
  assign n1960 = ~x1093 & n1959 ;
  assign n1961 = ( ~n1955 & n1956 ) | ( ~n1955 & n1960 ) | ( n1956 & n1960 ) ;
  assign n1962 = x683 & ~n1961 ;
  assign n1963 = n1954 & n1962 ;
  assign n1964 = x57 | x74 ;
  assign n1965 = n1206 | n1964 ;
  assign n1966 = n1334 | n1965 ;
  assign n1967 = x252 & ~n1953 ;
  assign n1968 = ( x100 & n1963 ) | ( x100 & ~n1967 ) | ( n1963 & ~n1967 ) ;
  assign n1969 = ( ~n1963 & n1966 ) | ( ~n1963 & n1968 ) | ( n1966 & n1968 ) ;
  assign n1970 = x39 | x51 ;
  assign n1971 = x93 & ~x841 ;
  assign n1972 = n1281 | n1352 ;
  assign n1973 = ( ~n1487 & n1971 ) | ( ~n1487 & n1972 ) | ( n1971 & n1972 ) ;
  assign n1974 = ( ~n1487 & n1970 ) | ( ~n1487 & n1973 ) | ( n1970 & n1973 ) ;
  assign n1975 = n1487 | n1974 ;
  assign n1976 = x215 & x299 ;
  assign n1977 = x223 & ~x299 ;
  assign n1978 = n1976 | n1977 ;
  assign n1979 = x614 | x616 ;
  assign n1980 = x603 & ~x642 ;
  assign n1981 = ~n1979 & n1980 ;
  assign n1982 = x332 | x468 ;
  assign n1983 = x661 | x662 ;
  assign n1984 = x680 & ~x681 ;
  assign n1985 = ~n1983 & n1984 ;
  assign n1986 = n1982 & ~n1985 ;
  assign n1987 = ~n1981 & n1986 ;
  assign n1988 = ~x287 & x835 ;
  assign n1989 = x252 | x1001 ;
  assign n1990 = x979 | x984 ;
  assign n1991 = ( n1988 & ~n1989 ) | ( n1988 & n1990 ) | ( ~n1989 & n1990 ) ;
  assign n1992 = n1988 & ~n1991 ;
  assign n1993 = ~n1987 & n1992 ;
  assign n1994 = x39 & n1993 ;
  assign n1995 = ~n1433 & n1959 ;
  assign n1996 = x971 | x974 ;
  assign n1997 = x602 | x961 ;
  assign n1998 = x967 | x969 ;
  assign n1999 = x299 | x587 ;
  assign n2000 = ( ~n1997 & n1998 ) | ( ~n1997 & n1999 ) | ( n1998 & n1999 ) ;
  assign n2001 = n1997 | n2000 ;
  assign n2002 = ( x977 & ~n1996 ) | ( x977 & n2001 ) | ( ~n1996 & n2001 ) ;
  assign n2003 = n1996 | n2002 ;
  assign n2004 = x975 | x978 ;
  assign n2005 = x970 | x972 ;
  assign n2006 = x960 | x963 ;
  assign n2007 = x907 | x947 ;
  assign n2008 = ( ~n2004 & n2006 ) | ( ~n2004 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2009 = ( ~n2004 & n2005 ) | ( ~n2004 & n2008 ) | ( n2005 & n2008 ) ;
  assign n2010 = n2004 | n2009 ;
  assign n2011 = x299 & ~n2010 ;
  assign n2012 = ( n1982 & n2003 ) | ( n1982 & ~n2011 ) | ( n2003 & ~n2011 ) ;
  assign n2013 = ( n1987 & n1995 ) | ( n1987 & ~n2012 ) | ( n1995 & ~n2012 ) ;
  assign n2014 = n1995 & ~n2013 ;
  assign n2015 = n1994 & n2014 ;
  assign n2016 = n1978 & n2015 ;
  assign n2017 = n1435 & n2012 ;
  assign n2018 = n1994 & n2017 ;
  assign n2019 = ~x299 & n1459 ;
  assign n2020 = x224 & n2019 ;
  assign n2021 = x299 & n1289 ;
  assign n2022 = x216 & n2021 ;
  assign n2023 = n2020 | n2022 ;
  assign n2024 = n2018 & n2023 ;
  assign n2025 = x210 & x299 ;
  assign n2026 = x198 & ~x299 ;
  assign n2027 = n2025 | n2026 ;
  assign n2028 = n1443 & ~n2027 ;
  assign n2029 = ( ~n2016 & n2024 ) | ( ~n2016 & n2028 ) | ( n2024 & n2028 ) ;
  assign n2030 = n2016 | n2029 ;
  assign n2031 = ~n1969 & n2030 ;
  assign n2032 = ( n1969 & n1975 ) | ( n1969 & ~n2031 ) | ( n1975 & ~n2031 ) ;
  assign n2033 = ~n1940 & n2032 ;
  assign n2034 = ~x907 & n1553 ;
  assign n2035 = x602 | n1553 ;
  assign n2036 = ( n1982 & ~n2034 ) | ( n1982 & n2035 ) | ( ~n2034 & n2035 ) ;
  assign n2037 = ~n1986 & n2036 ;
  assign n2038 = n1301 | n2028 ;
  assign n2039 = ~n1350 & n2038 ;
  assign n2040 = x39 & x1093 ;
  assign n2041 = ( n1992 & n1995 ) | ( n1992 & ~n2040 ) | ( n1995 & ~n2040 ) ;
  assign n2042 = n2040 & n2041 ;
  assign n2043 = ~x216 & n2021 ;
  assign n2044 = n1459 & ~n1772 ;
  assign n2045 = x829 & x1091 ;
  assign n2046 = ( n2043 & n2044 ) | ( n2043 & ~n2045 ) | ( n2044 & ~n2045 ) ;
  assign n2047 = ( n2023 & n2042 ) | ( n2023 & n2046 ) | ( n2042 & n2046 ) ;
  assign n2048 = x40 | n1347 ;
  assign n2049 = x95 | n1276 ;
  assign n2050 = ( n1271 & ~n2048 ) | ( n1271 & n2049 ) | ( ~n2048 & n2049 ) ;
  assign n2051 = n2048 | n2050 ;
  assign n2052 = x72 & ~n2051 ;
  assign n2053 = ( ~n2039 & n2047 ) | ( ~n2039 & n2052 ) | ( n2047 & n2052 ) ;
  assign n2054 = n2039 | n2053 ;
  assign n2055 = x90 | n1362 ;
  assign n2056 = n1266 & ~n1372 ;
  assign n2057 = ( ~n1254 & n1483 ) | ( ~n1254 & n2056 ) | ( n1483 & n2056 ) ;
  assign n2058 = ~n1387 & n2057 ;
  assign n2059 = x103 & ~x314 ;
  assign n2060 = x109 | n1272 ;
  assign n2061 = x81 | x83 ;
  assign n2062 = ( n1251 & n1399 ) | ( n1251 & ~n2061 ) | ( n1399 & ~n2061 ) ;
  assign n2063 = n2061 | n2062 ;
  assign n2064 = ( ~n2059 & n2060 ) | ( ~n2059 & n2063 ) | ( n2060 & n2063 ) ;
  assign n2065 = n1485 | n2060 ;
  assign n2066 = ( n2059 & n2064 ) | ( n2059 & n2065 ) | ( n2064 & n2065 ) ;
  assign n2067 = ( ~n1387 & n2058 ) | ( ~n1387 & n2066 ) | ( n2058 & n2066 ) ;
  assign n2068 = n2055 | n2067 ;
  assign n2069 = x109 | n1971 ;
  assign n2070 = x109 & ~x197 ;
  assign n2071 = x158 & x159 ;
  assign n2072 = x232 & ~n1982 ;
  assign n2073 = x299 & n2072 ;
  assign n2074 = x160 & n2073 ;
  assign n2075 = n2071 & n2074 ;
  assign n2076 = ( x109 & n2070 ) | ( x109 & ~n2075 ) | ( n2070 & ~n2075 ) ;
  assign n2077 = x145 & x180 ;
  assign n2078 = x181 & n2077 ;
  assign n2079 = ~x299 & n2072 ;
  assign n2080 = x182 & n2079 ;
  assign n2081 = n2078 & n2080 ;
  assign n2082 = n2076 & ~n2081 ;
  assign n2083 = ( n1359 & n2069 ) | ( n1359 & ~n2082 ) | ( n2069 & ~n2082 ) ;
  assign n2084 = n2068 & ~n2083 ;
  assign n2085 = n2054 | n2084 ;
  assign n2086 = ( x55 & n1215 ) | ( x55 & ~n1312 ) | ( n1215 & ~n1312 ) ;
  assign n2087 = n1205 | n2086 ;
  assign n2088 = ~x39 & n2087 ;
  assign n2089 = ( n1515 & n1963 ) | ( n1515 & n1967 ) | ( n1963 & n1967 ) ;
  assign n2090 = n2088 | n2089 ;
  assign n2091 = ~n1333 & n2090 ;
  assign n2092 = n1213 | n1319 ;
  assign n2093 = n1334 | n2092 ;
  assign n2094 = ( n1333 & n2085 ) | ( n1333 & n2093 ) | ( n2085 & n2093 ) ;
  assign n2095 = ( n2085 & n2091 ) | ( n2085 & ~n2094 ) | ( n2091 & ~n2094 ) ;
  assign n2096 = ~x30 & x228 ;
  assign n2097 = x30 & x228 ;
  assign n2098 = ( n2095 & ~n2096 ) | ( n2095 & n2097 ) | ( ~n2096 & n2097 ) ;
  assign n2099 = n2037 & n2098 ;
  assign n2100 = ~n1982 & n1999 ;
  assign n2101 = ( n1208 & ~n1982 ) | ( n1208 & n2100 ) | ( ~n1982 & n2100 ) ;
  assign n2102 = n1981 & n1982 ;
  assign n2103 = x947 | n1982 ;
  assign n2104 = n1553 & ~n2103 ;
  assign n2105 = ( n2101 & n2102 ) | ( n2101 & ~n2104 ) | ( n2102 & ~n2104 ) ;
  assign n2106 = n2098 & n2105 ;
  assign n2107 = x970 & n1553 ;
  assign n2108 = ~n1982 & n2098 ;
  assign n2109 = x967 & ~n1553 ;
  assign n2110 = ( n2107 & n2108 ) | ( n2107 & n2109 ) | ( n2108 & n2109 ) ;
  assign n2111 = x972 & n1553 ;
  assign n2112 = x961 & ~n1553 ;
  assign n2113 = ( n2108 & n2111 ) | ( n2108 & n2112 ) | ( n2111 & n2112 ) ;
  assign n2114 = x977 & ~n1553 ;
  assign n2115 = x960 & n1553 ;
  assign n2116 = ( n2108 & n2114 ) | ( n2108 & n2115 ) | ( n2114 & n2115 ) ;
  assign n2117 = x969 & ~n1553 ;
  assign n2118 = x963 & n1553 ;
  assign n2119 = ( n2108 & n2117 ) | ( n2108 & n2118 ) | ( n2117 & n2118 ) ;
  assign n2120 = x971 & ~n1553 ;
  assign n2121 = x975 & n1553 ;
  assign n2122 = ( n2108 & n2120 ) | ( n2108 & n2121 ) | ( n2120 & n2121 ) ;
  assign n2123 = x974 & ~n1553 ;
  assign n2124 = x978 & n1553 ;
  assign n2125 = ( n2108 & n2123 ) | ( n2108 & n2124 ) | ( n2123 & n2124 ) ;
  assign n2126 = x24 & x954 ;
  assign n2127 = ~x24 & x954 ;
  assign n2128 = x39 & ~x287 ;
  assign n2129 = ~x979 & n2128 ;
  assign n2130 = x835 & x984 ;
  assign n2131 = n2129 & ~n2130 ;
  assign n2132 = n1989 & n2131 ;
  assign n2133 = ( x1093 & ~n1976 ) | ( x1093 & n1977 ) | ( ~n1976 & n1977 ) ;
  assign n2134 = ( x835 & n1976 ) | ( x835 & n2133 ) | ( n1976 & n2133 ) ;
  assign n2135 = n2014 & n2134 ;
  assign n2136 = n2132 & ~n2135 ;
  assign n2137 = n1336 | n2136 ;
  assign n2138 = ( n1333 & n2085 ) | ( n1333 & n2137 ) | ( n2085 & n2137 ) ;
  assign n2139 = ( n2085 & n2091 ) | ( n2085 & ~n2138 ) | ( n2091 & ~n2138 ) ;
  assign n2140 = ( ~n2126 & n2127 ) | ( ~n2126 & n2139 ) | ( n2127 & n2139 ) ;
  assign n2141 = ~n1309 & n1415 ;
  assign n2142 = ( x55 & x92 ) | ( x55 & n1321 ) | ( x92 & n1321 ) ;
  assign n2143 = ( x55 & x92 ) | ( x55 & ~n1206 ) | ( x92 & ~n1206 ) ;
  assign n2144 = x91 | x110 ;
  assign n2145 = x65 | x71 ;
  assign n2146 = x47 | x64 ;
  assign n2147 = ( ~n2144 & n2145 ) | ( ~n2144 & n2146 ) | ( n2145 & n2146 ) ;
  assign n2148 = n2144 | n2147 ;
  assign n2149 = n1266 | n2148 ;
  assign n2150 = x72 | n1347 ;
  assign n2151 = x67 | x103 ;
  assign n2152 = x109 | n2151 ;
  assign n2153 = x36 | x69 ;
  assign n2154 = x83 | n2153 ;
  assign n2155 = ( ~n2150 & n2152 ) | ( ~n2150 & n2154 ) | ( n2152 & n2154 ) ;
  assign n2156 = n2150 | n2155 ;
  assign n2157 = n1240 | n2156 ;
  assign n2158 = n2149 | n2157 ;
  assign n2159 = n2049 | n2158 ;
  assign n2160 = ( n2142 & n2143 ) | ( n2142 & ~n2159 ) | ( n2143 & ~n2159 ) ;
  assign n2161 = ~n2142 & n2160 ;
  assign n2162 = n1206 | n1506 ;
  assign n2163 = ~x100 & n2162 ;
  assign n2164 = ( ~n1967 & n2162 ) | ( ~n1967 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2165 = n2161 | n2164 ;
  assign n2166 = ~n1332 & n2165 ;
  assign n2167 = n2141 | n2166 ;
  assign n2168 = ( n1299 & ~n1338 ) | ( n1299 & n2167 ) | ( ~n1338 & n2167 ) ;
  assign n2169 = x119 & ~x1056 ;
  assign n2170 = ~x119 & n1523 ;
  assign n2171 = ( ~x468 & n2169 ) | ( ~x468 & n2170 ) | ( n2169 & n2170 ) ;
  assign n2172 = x119 & ~x1077 ;
  assign n2173 = ( ~x468 & n2170 ) | ( ~x468 & n2172 ) | ( n2170 & n2172 ) ;
  assign n2174 = x119 & ~x1073 ;
  assign n2175 = ( ~x468 & n2170 ) | ( ~x468 & n2174 ) | ( n2170 & n2174 ) ;
  assign n2176 = x119 & ~x1041 ;
  assign n2177 = ( ~x468 & n2170 ) | ( ~x468 & n2176 ) | ( n2170 & n2176 ) ;
  assign n2178 = ~x31 & n1430 ;
  assign n2179 = x1161 | x1162 ;
  assign n2180 = x1163 | n2179 ;
  assign n2181 = ~x98 & x567 ;
  assign n2182 = n1430 & ~n2181 ;
  assign n2183 = x591 | x592 ;
  assign n2184 = x588 & ~x590 ;
  assign n2185 = ~n2183 & n2184 ;
  assign n2186 = ( x418 & x431 ) | ( x418 & x437 ) | ( x431 & x437 ) ;
  assign n2187 = ( ~x418 & x431 ) | ( ~x418 & x437 ) | ( x431 & x437 ) ;
  assign n2188 = ( x418 & ~n2186 ) | ( x418 & n2187 ) | ( ~n2186 & n2187 ) ;
  assign n2189 = ( ~x417 & x438 ) | ( ~x417 & n2188 ) | ( x438 & n2188 ) ;
  assign n2190 = ( x417 & x438 ) | ( x417 & n2188 ) | ( x438 & n2188 ) ;
  assign n2191 = ( x417 & n2189 ) | ( x417 & ~n2190 ) | ( n2189 & ~n2190 ) ;
  assign n2192 = x415 | x416 ;
  assign n2193 = ~x415 & x416 ;
  assign n2194 = ( ~x416 & n2192 ) | ( ~x416 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2195 = ( x453 & x464 ) | ( x453 & n2194 ) | ( x464 & n2194 ) ;
  assign n2196 = ( x453 & x464 ) | ( x453 & ~n2194 ) | ( x464 & ~n2194 ) ;
  assign n2197 = ( n2194 & ~n2195 ) | ( n2194 & n2196 ) | ( ~n2195 & n2196 ) ;
  assign n2198 = ( x1197 & n2191 ) | ( x1197 & n2197 ) | ( n2191 & n2197 ) ;
  assign n2199 = ( ~x1197 & n2191 ) | ( ~x1197 & n2197 ) | ( n2191 & n2197 ) ;
  assign n2200 = n2198 & ~n2199 ;
  assign n2201 = x419 | x421 ;
  assign n2202 = ~x419 & x421 ;
  assign n2203 = ( ~x421 & n2201 ) | ( ~x421 & n2202 ) | ( n2201 & n2202 ) ;
  assign n2204 = ( x423 & x425 ) | ( x423 & ~n2203 ) | ( x425 & ~n2203 ) ;
  assign n2205 = ( x423 & x425 ) | ( x423 & n2203 ) | ( x425 & n2203 ) ;
  assign n2206 = ( n2203 & n2204 ) | ( n2203 & ~n2205 ) | ( n2204 & ~n2205 ) ;
  assign n2207 = ( x432 & x454 ) | ( x432 & x459 ) | ( x454 & x459 ) ;
  assign n2208 = ( ~x432 & x454 ) | ( ~x432 & x459 ) | ( x454 & x459 ) ;
  assign n2209 = ( x432 & ~n2207 ) | ( x432 & n2208 ) | ( ~n2207 & n2208 ) ;
  assign n2210 = ( ~x420 & x424 ) | ( ~x420 & n2209 ) | ( x424 & n2209 ) ;
  assign n2211 = ( x420 & x424 ) | ( x420 & n2209 ) | ( x424 & n2209 ) ;
  assign n2212 = ( x420 & n2210 ) | ( x420 & ~n2211 ) | ( n2210 & ~n2211 ) ;
  assign n2213 = n2206 & n2212 ;
  assign n2214 = ( x1198 & n2206 ) | ( x1198 & n2212 ) | ( n2206 & n2212 ) ;
  assign n2215 = ( n2200 & ~n2213 ) | ( n2200 & n2214 ) | ( ~n2213 & n2214 ) ;
  assign n2216 = x427 | x428 ;
  assign n2217 = ~x427 & x428 ;
  assign n2218 = ( ~x428 & n2216 ) | ( ~x428 & n2217 ) | ( n2216 & n2217 ) ;
  assign n2219 = ( x430 & x451 ) | ( x430 & n2218 ) | ( x451 & n2218 ) ;
  assign n2220 = ( x430 & x451 ) | ( x430 & ~n2218 ) | ( x451 & ~n2218 ) ;
  assign n2221 = ( n2218 & ~n2219 ) | ( n2218 & n2220 ) | ( ~n2219 & n2220 ) ;
  assign n2222 = x433 | x445 ;
  assign n2223 = ~x433 & x445 ;
  assign n2224 = ( ~x445 & n2222 ) | ( ~x445 & n2223 ) | ( n2222 & n2223 ) ;
  assign n2225 = ( x448 & x449 ) | ( x448 & n2224 ) | ( x449 & n2224 ) ;
  assign n2226 = ( x448 & x449 ) | ( x448 & ~n2224 ) | ( x449 & ~n2224 ) ;
  assign n2227 = ( n2224 & ~n2225 ) | ( n2224 & n2226 ) | ( ~n2225 & n2226 ) ;
  assign n2228 = ( x426 & n2221 ) | ( x426 & n2227 ) | ( n2221 & n2227 ) ;
  assign n2229 = ( ~x426 & n2221 ) | ( ~x426 & n2227 ) | ( n2221 & n2227 ) ;
  assign n2230 = ( x426 & ~n2228 ) | ( x426 & n2229 ) | ( ~n2228 & n2229 ) ;
  assign n2231 = x1199 & n2230 ;
  assign n2232 = ( x435 & x436 ) | ( x435 & x443 ) | ( x436 & x443 ) ;
  assign n2233 = ( ~x435 & x436 ) | ( ~x435 & x443 ) | ( x436 & x443 ) ;
  assign n2234 = ( x435 & ~n2232 ) | ( x435 & n2233 ) | ( ~n2232 & n2233 ) ;
  assign n2235 = ( ~x414 & x429 ) | ( ~x414 & n2234 ) | ( x429 & n2234 ) ;
  assign n2236 = ( x414 & x429 ) | ( x414 & n2234 ) | ( x429 & n2234 ) ;
  assign n2237 = ( x414 & n2235 ) | ( x414 & ~n2236 ) | ( n2235 & ~n2236 ) ;
  assign n2238 = x422 | x434 ;
  assign n2239 = ~x422 & x434 ;
  assign n2240 = ( ~x434 & n2238 ) | ( ~x434 & n2239 ) | ( n2238 & n2239 ) ;
  assign n2241 = ( x444 & x446 ) | ( x444 & n2240 ) | ( x446 & n2240 ) ;
  assign n2242 = ( x444 & x446 ) | ( x444 & ~n2240 ) | ( x446 & ~n2240 ) ;
  assign n2243 = ( n2240 & ~n2241 ) | ( n2240 & n2242 ) | ( ~n2241 & n2242 ) ;
  assign n2244 = n2237 & n2243 ;
  assign n2245 = ( x1196 & n2237 ) | ( x1196 & n2243 ) | ( n2237 & n2243 ) ;
  assign n2246 = ( n2231 & ~n2244 ) | ( n2231 & n2245 ) | ( ~n2244 & n2245 ) ;
  assign n2247 = n2215 | n2246 ;
  assign n2248 = n2185 & n2247 ;
  assign n2249 = x318 | x325 ;
  assign n2250 = ~x318 & x325 ;
  assign n2251 = ( ~x325 & n2249 ) | ( ~x325 & n2250 ) | ( n2249 & n2250 ) ;
  assign n2252 = ( x405 & x409 ) | ( x405 & n2251 ) | ( x409 & n2251 ) ;
  assign n2253 = ( x405 & x409 ) | ( x405 & ~n2251 ) | ( x409 & ~n2251 ) ;
  assign n2254 = ( n2251 & ~n2252 ) | ( n2251 & n2253 ) | ( ~n2252 & n2253 ) ;
  assign n2255 = ~x401 & x402 ;
  assign n2256 = x401 | x402 ;
  assign n2257 = ( ~x402 & n2255 ) | ( ~x402 & n2256 ) | ( n2255 & n2256 ) ;
  assign n2258 = ( x403 & x406 ) | ( x403 & ~n2257 ) | ( x406 & ~n2257 ) ;
  assign n2259 = ( x403 & x406 ) | ( x403 & n2257 ) | ( x406 & n2257 ) ;
  assign n2260 = ( n2257 & n2258 ) | ( n2257 & ~n2259 ) | ( n2258 & ~n2259 ) ;
  assign n2261 = ( x326 & n2254 ) | ( x326 & n2260 ) | ( n2254 & n2260 ) ;
  assign n2262 = ( ~x326 & n2254 ) | ( ~x326 & n2260 ) | ( n2254 & n2260 ) ;
  assign n2263 = ( x326 & ~n2261 ) | ( x326 & n2262 ) | ( ~n2261 & n2262 ) ;
  assign n2264 = x1199 & n2263 ;
  assign n2265 = ( x324 & x390 ) | ( x324 & x410 ) | ( x390 & x410 ) ;
  assign n2266 = ( ~x324 & x390 ) | ( ~x324 & x410 ) | ( x390 & x410 ) ;
  assign n2267 = ( x324 & ~n2265 ) | ( x324 & n2266 ) | ( ~n2265 & n2266 ) ;
  assign n2268 = ( x319 & x456 ) | ( x319 & n2267 ) | ( x456 & n2267 ) ;
  assign n2269 = ( ~x319 & x456 ) | ( ~x319 & n2267 ) | ( x456 & n2267 ) ;
  assign n2270 = ( x319 & ~n2268 ) | ( x319 & n2269 ) | ( ~n2268 & n2269 ) ;
  assign n2271 = x397 | x404 ;
  assign n2272 = ~x397 & x404 ;
  assign n2273 = ( ~x404 & n2271 ) | ( ~x404 & n2272 ) | ( n2271 & n2272 ) ;
  assign n2274 = ( x411 & x412 ) | ( x411 & ~n2273 ) | ( x412 & ~n2273 ) ;
  assign n2275 = ( x411 & x412 ) | ( x411 & n2273 ) | ( x412 & n2273 ) ;
  assign n2276 = ( n2273 & n2274 ) | ( n2273 & ~n2275 ) | ( n2274 & ~n2275 ) ;
  assign n2277 = n2270 & n2276 ;
  assign n2278 = ( x1196 & n2270 ) | ( x1196 & n2276 ) | ( n2270 & n2276 ) ;
  assign n2279 = ( n2264 & ~n2277 ) | ( n2264 & n2278 ) | ( ~n2277 & n2278 ) ;
  assign n2280 = x394 | x395 ;
  assign n2281 = ~x394 & x395 ;
  assign n2282 = ( ~x395 & n2280 ) | ( ~x395 & n2281 ) | ( n2280 & n2281 ) ;
  assign n2283 = ( x399 & x400 ) | ( x399 & n2282 ) | ( x400 & n2282 ) ;
  assign n2284 = ( x399 & x400 ) | ( x399 & ~n2282 ) | ( x400 & ~n2282 ) ;
  assign n2285 = ( n2282 & ~n2283 ) | ( n2282 & n2284 ) | ( ~n2283 & n2284 ) ;
  assign n2286 = x328 | x396 ;
  assign n2287 = ~x328 & x396 ;
  assign n2288 = ( ~x396 & n2286 ) | ( ~x396 & n2287 ) | ( n2286 & n2287 ) ;
  assign n2289 = ( x398 & x408 ) | ( x398 & n2288 ) | ( x408 & n2288 ) ;
  assign n2290 = ( x398 & x408 ) | ( x398 & ~n2288 ) | ( x408 & ~n2288 ) ;
  assign n2291 = ( n2288 & ~n2289 ) | ( n2288 & n2290 ) | ( ~n2289 & n2290 ) ;
  assign n2292 = ( x329 & n2285 ) | ( x329 & n2291 ) | ( n2285 & n2291 ) ;
  assign n2293 = ( ~x329 & n2285 ) | ( ~x329 & n2291 ) | ( n2285 & n2291 ) ;
  assign n2294 = ( x329 & ~n2292 ) | ( x329 & n2293 ) | ( ~n2292 & n2293 ) ;
  assign n2295 = x1198 & n2294 ;
  assign n2296 = ~x391 & x393 ;
  assign n2297 = x391 | x393 ;
  assign n2298 = ( ~x393 & n2296 ) | ( ~x393 & n2297 ) | ( n2296 & n2297 ) ;
  assign n2299 = ( x407 & x413 ) | ( x407 & ~n2298 ) | ( x413 & ~n2298 ) ;
  assign n2300 = ( x407 & x413 ) | ( x407 & n2298 ) | ( x413 & n2298 ) ;
  assign n2301 = ( n2298 & n2299 ) | ( n2298 & ~n2300 ) | ( n2299 & ~n2300 ) ;
  assign n2302 = ( ~x335 & x392 ) | ( ~x335 & x463 ) | ( x392 & x463 ) ;
  assign n2303 = ( x335 & x392 ) | ( x335 & x463 ) | ( x392 & x463 ) ;
  assign n2304 = ( x335 & n2302 ) | ( x335 & ~n2303 ) | ( n2302 & ~n2303 ) ;
  assign n2305 = ( ~x333 & x334 ) | ( ~x333 & n2304 ) | ( x334 & n2304 ) ;
  assign n2306 = ( x333 & x334 ) | ( x333 & n2304 ) | ( x334 & n2304 ) ;
  assign n2307 = ( x333 & n2305 ) | ( x333 & ~n2306 ) | ( n2305 & ~n2306 ) ;
  assign n2308 = n2301 & n2307 ;
  assign n2309 = ( x1197 & n2301 ) | ( x1197 & n2307 ) | ( n2301 & n2307 ) ;
  assign n2310 = ( n2295 & ~n2308 ) | ( n2295 & n2309 ) | ( ~n2308 & n2309 ) ;
  assign n2311 = n2279 | n2310 ;
  assign n2312 = x588 | x590 ;
  assign n2313 = x591 & ~x592 ;
  assign n2314 = ~n2312 & n2313 ;
  assign n2315 = n2311 & n2314 ;
  assign n2316 = n2248 | n2315 ;
  assign n2317 = ( ~x317 & x378 ) | ( ~x317 & x381 ) | ( x378 & x381 ) ;
  assign n2318 = ( x317 & x378 ) | ( x317 & x381 ) | ( x378 & x381 ) ;
  assign n2319 = ( x317 & n2317 ) | ( x317 & ~n2318 ) | ( n2317 & ~n2318 ) ;
  assign n2320 = ( x377 & x385 ) | ( x377 & n2319 ) | ( x385 & n2319 ) ;
  assign n2321 = ( ~x377 & x385 ) | ( ~x377 & n2319 ) | ( x385 & n2319 ) ;
  assign n2322 = ( x377 & ~n2320 ) | ( x377 & n2321 ) | ( ~n2320 & n2321 ) ;
  assign n2323 = ~x376 & x379 ;
  assign n2324 = x376 | x379 ;
  assign n2325 = ( ~x379 & n2323 ) | ( ~x379 & n2324 ) | ( n2323 & n2324 ) ;
  assign n2326 = ( x382 & x439 ) | ( x382 & ~n2325 ) | ( x439 & ~n2325 ) ;
  assign n2327 = ( x382 & x439 ) | ( x382 & n2325 ) | ( x439 & n2325 ) ;
  assign n2328 = ( n2325 & n2326 ) | ( n2325 & ~n2327 ) | ( n2326 & ~n2327 ) ;
  assign n2329 = ( ~x1199 & n2322 ) | ( ~x1199 & n2328 ) | ( n2322 & n2328 ) ;
  assign n2330 = ( x1199 & n2322 ) | ( x1199 & n2328 ) | ( n2322 & n2328 ) ;
  assign n2331 = ~n2329 & n2330 ;
  assign n2332 = ~x369 & x371 ;
  assign n2333 = x369 | x371 ;
  assign n2334 = ( ~x371 & n2332 ) | ( ~x371 & n2333 ) | ( n2332 & n2333 ) ;
  assign n2335 = ( x373 & x442 ) | ( x373 & n2334 ) | ( x442 & n2334 ) ;
  assign n2336 = ( x373 & x442 ) | ( x373 & ~n2334 ) | ( x442 & ~n2334 ) ;
  assign n2337 = ( n2334 & ~n2335 ) | ( n2334 & n2336 ) | ( ~n2335 & n2336 ) ;
  assign n2338 = ( ~x374 & x384 ) | ( ~x374 & n2337 ) | ( x384 & n2337 ) ;
  assign n2339 = ( x374 & x384 ) | ( x374 & n2337 ) | ( x384 & n2337 ) ;
  assign n2340 = ( x374 & n2338 ) | ( x374 & ~n2339 ) | ( n2338 & ~n2339 ) ;
  assign n2341 = ( ~x370 & x375 ) | ( ~x370 & x440 ) | ( x375 & x440 ) ;
  assign n2342 = ( x370 & x375 ) | ( x370 & x440 ) | ( x375 & x440 ) ;
  assign n2343 = ( x370 & n2341 ) | ( x370 & ~n2342 ) | ( n2341 & ~n2342 ) ;
  assign n2344 = n2340 & n2343 ;
  assign n2345 = ( x1198 & n2340 ) | ( x1198 & n2343 ) | ( n2340 & n2343 ) ;
  assign n2346 = ( n2331 & ~n2344 ) | ( n2331 & n2345 ) | ( ~n2344 & n2345 ) ;
  assign n2347 = ( ~x363 & x372 ) | ( ~x363 & x380 ) | ( x372 & x380 ) ;
  assign n2348 = ( x363 & x372 ) | ( x363 & x380 ) | ( x372 & x380 ) ;
  assign n2349 = ( x363 & n2347 ) | ( x363 & ~n2348 ) | ( n2347 & ~n2348 ) ;
  assign n2350 = ( x337 & x386 ) | ( x337 & n2349 ) | ( x386 & n2349 ) ;
  assign n2351 = ( ~x337 & x386 ) | ( ~x337 & n2349 ) | ( x386 & n2349 ) ;
  assign n2352 = ( x337 & ~n2350 ) | ( x337 & n2351 ) | ( ~n2350 & n2351 ) ;
  assign n2353 = ~x338 & x339 ;
  assign n2354 = x338 | x339 ;
  assign n2355 = ( ~x339 & n2353 ) | ( ~x339 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2356 = ( x387 & x388 ) | ( x387 & ~n2355 ) | ( x388 & ~n2355 ) ;
  assign n2357 = ( x387 & x388 ) | ( x387 & n2355 ) | ( x388 & n2355 ) ;
  assign n2358 = ( n2355 & n2356 ) | ( n2355 & ~n2357 ) | ( n2356 & ~n2357 ) ;
  assign n2359 = ( x1196 & n2352 ) | ( x1196 & n2358 ) | ( n2352 & n2358 ) ;
  assign n2360 = ( ~x1196 & n2352 ) | ( ~x1196 & n2358 ) | ( n2352 & n2358 ) ;
  assign n2361 = n2359 & ~n2360 ;
  assign n2362 = ( x367 & x383 ) | ( x367 & x389 ) | ( x383 & x389 ) ;
  assign n2363 = ( ~x367 & x383 ) | ( ~x367 & x389 ) | ( x383 & x389 ) ;
  assign n2364 = ( x367 & ~n2362 ) | ( x367 & n2363 ) | ( ~n2362 & n2363 ) ;
  assign n2365 = x364 | x365 ;
  assign n2366 = ~x364 & x365 ;
  assign n2367 = ( ~x365 & n2365 ) | ( ~x365 & n2366 ) | ( n2365 & n2366 ) ;
  assign n2368 = ( x368 & x447 ) | ( x368 & n2367 ) | ( x447 & n2367 ) ;
  assign n2369 = ( x368 & x447 ) | ( x368 & ~n2367 ) | ( x447 & ~n2367 ) ;
  assign n2370 = ( n2367 & ~n2368 ) | ( n2367 & n2369 ) | ( ~n2368 & n2369 ) ;
  assign n2371 = ( ~x336 & x366 ) | ( ~x336 & n2370 ) | ( x366 & n2370 ) ;
  assign n2372 = ( x336 & x366 ) | ( x336 & n2370 ) | ( x366 & n2370 ) ;
  assign n2373 = ( x336 & n2371 ) | ( x336 & ~n2372 ) | ( n2371 & ~n2372 ) ;
  assign n2374 = n2364 & n2373 ;
  assign n2375 = ( x1197 & n2364 ) | ( x1197 & n2373 ) | ( n2364 & n2373 ) ;
  assign n2376 = ( n2361 & ~n2374 ) | ( n2361 & n2375 ) | ( ~n2374 & n2375 ) ;
  assign n2377 = n2346 | n2376 ;
  assign n2378 = ~x591 & x592 ;
  assign n2379 = ~x590 & n2378 ;
  assign n2380 = n2377 & n2379 ;
  assign n2381 = x590 & ~n2183 ;
  assign n2382 = ( ~x353 & x357 ) | ( ~x353 & x462 ) | ( x357 & x462 ) ;
  assign n2383 = ( x353 & x357 ) | ( x353 & x462 ) | ( x357 & x462 ) ;
  assign n2384 = ( x353 & n2382 ) | ( x353 & ~n2383 ) | ( n2382 & ~n2383 ) ;
  assign n2385 = ( ~x351 & x352 ) | ( ~x351 & n2384 ) | ( x352 & n2384 ) ;
  assign n2386 = ( x351 & x352 ) | ( x351 & n2384 ) | ( x352 & n2384 ) ;
  assign n2387 = ( x351 & n2385 ) | ( x351 & ~n2386 ) | ( n2385 & ~n2386 ) ;
  assign n2388 = ~x354 & x356 ;
  assign n2389 = x354 | x356 ;
  assign n2390 = ( ~x356 & n2388 ) | ( ~x356 & n2389 ) | ( n2388 & n2389 ) ;
  assign n2391 = ( x360 & x461 ) | ( x360 & n2390 ) | ( x461 & n2390 ) ;
  assign n2392 = ( x360 & x461 ) | ( x360 & ~n2390 ) | ( x461 & ~n2390 ) ;
  assign n2393 = ( n2390 & ~n2391 ) | ( n2390 & n2392 ) | ( ~n2391 & n2392 ) ;
  assign n2394 = ( ~x1199 & n2387 ) | ( ~x1199 & n2393 ) | ( n2387 & n2393 ) ;
  assign n2395 = ( x1199 & n2387 ) | ( x1199 & n2393 ) | ( n2387 & n2393 ) ;
  assign n2396 = ~n2394 & n2395 ;
  assign n2397 = ( x321 & x347 ) | ( x321 & x359 ) | ( x347 & x359 ) ;
  assign n2398 = ( ~x321 & x347 ) | ( ~x321 & x359 ) | ( x347 & x359 ) ;
  assign n2399 = ( x321 & ~n2397 ) | ( x321 & n2398 ) | ( ~n2397 & n2398 ) ;
  assign n2400 = ( ~x315 & x316 ) | ( ~x315 & n2399 ) | ( x316 & n2399 ) ;
  assign n2401 = ( x315 & x316 ) | ( x315 & n2399 ) | ( x316 & n2399 ) ;
  assign n2402 = ( x315 & n2400 ) | ( x315 & ~n2401 ) | ( n2400 & ~n2401 ) ;
  assign n2403 = x322 | x348 ;
  assign n2404 = ~x322 & x348 ;
  assign n2405 = ( ~x348 & n2403 ) | ( ~x348 & n2404 ) | ( n2403 & n2404 ) ;
  assign n2406 = ( x349 & x350 ) | ( x349 & n2405 ) | ( x350 & n2405 ) ;
  assign n2407 = ( x349 & x350 ) | ( x349 & ~n2405 ) | ( x350 & ~n2405 ) ;
  assign n2408 = ( n2405 & ~n2406 ) | ( n2405 & n2407 ) | ( ~n2406 & n2407 ) ;
  assign n2409 = n2402 & n2408 ;
  assign n2410 = ( x1198 & n2402 ) | ( x1198 & n2408 ) | ( n2402 & n2408 ) ;
  assign n2411 = ( n2396 & ~n2409 ) | ( n2396 & n2410 ) | ( ~n2409 & n2410 ) ;
  assign n2412 = ( ~x320 & x452 ) | ( ~x320 & x458 ) | ( x452 & x458 ) ;
  assign n2413 = ( x320 & x452 ) | ( x320 & x458 ) | ( x452 & x458 ) ;
  assign n2414 = ( x320 & n2412 ) | ( x320 & ~n2413 ) | ( n2412 & ~n2413 ) ;
  assign n2415 = ( ~x342 & x361 ) | ( ~x342 & x460 ) | ( x361 & x460 ) ;
  assign n2416 = ( x342 & x361 ) | ( x342 & x460 ) | ( x361 & x460 ) ;
  assign n2417 = ( x342 & n2415 ) | ( x342 & ~n2416 ) | ( n2415 & ~n2416 ) ;
  assign n2418 = ( ~x355 & x441 ) | ( ~x355 & x455 ) | ( x441 & x455 ) ;
  assign n2419 = ( x355 & x441 ) | ( x355 & x455 ) | ( x441 & x455 ) ;
  assign n2420 = ( x355 & n2418 ) | ( x355 & ~n2419 ) | ( n2418 & ~n2419 ) ;
  assign n2421 = ( ~n2414 & n2417 ) | ( ~n2414 & n2420 ) | ( n2417 & n2420 ) ;
  assign n2422 = ( n2414 & n2417 ) | ( n2414 & n2420 ) | ( n2417 & n2420 ) ;
  assign n2423 = ( n2414 & n2421 ) | ( n2414 & ~n2422 ) | ( n2421 & ~n2422 ) ;
  assign n2424 = x1196 & n2423 ;
  assign n2425 = x323 | x346 ;
  assign n2426 = ~x323 & x346 ;
  assign n2427 = ( ~x346 & n2425 ) | ( ~x346 & n2426 ) | ( n2425 & n2426 ) ;
  assign n2428 = ( x358 & x362 ) | ( x358 & n2427 ) | ( x362 & n2427 ) ;
  assign n2429 = ( x358 & x362 ) | ( x358 & ~n2427 ) | ( x362 & ~n2427 ) ;
  assign n2430 = ( n2427 & ~n2428 ) | ( n2427 & n2429 ) | ( ~n2428 & n2429 ) ;
  assign n2431 = ( x344 & x345 ) | ( x344 & x450 ) | ( x345 & x450 ) ;
  assign n2432 = ( ~x344 & x345 ) | ( ~x344 & x450 ) | ( x345 & x450 ) ;
  assign n2433 = ( x344 & ~n2431 ) | ( x344 & n2432 ) | ( ~n2431 & n2432 ) ;
  assign n2434 = ( ~x327 & x343 ) | ( ~x327 & n2433 ) | ( x343 & n2433 ) ;
  assign n2435 = ( x327 & x343 ) | ( x327 & n2433 ) | ( x343 & n2433 ) ;
  assign n2436 = ( x327 & n2434 ) | ( x327 & ~n2435 ) | ( n2434 & ~n2435 ) ;
  assign n2437 = n2430 & n2436 ;
  assign n2438 = ( x1197 & n2430 ) | ( x1197 & n2436 ) | ( n2430 & n2436 ) ;
  assign n2439 = ( n2424 & ~n2437 ) | ( n2424 & n2438 ) | ( ~n2437 & n2438 ) ;
  assign n2440 = n2381 & n2439 ;
  assign n2441 = ( n2381 & n2411 ) | ( n2381 & n2440 ) | ( n2411 & n2440 ) ;
  assign n2442 = ( ~x588 & n2380 ) | ( ~x588 & n2441 ) | ( n2380 & n2441 ) ;
  assign n2443 = n2316 | n2442 ;
  assign n2444 = x88 | n1259 ;
  assign n2445 = n1426 & n1958 ;
  assign n2446 = ~n1265 & n2445 ;
  assign n2447 = ~n2444 & n2446 ;
  assign n2448 = ( x51 & ~n1353 ) | ( x51 & n1354 ) | ( ~n1353 & n1354 ) ;
  assign n2449 = x51 | x841 ;
  assign n2450 = ( x90 & n1272 ) | ( x90 & n2449 ) | ( n1272 & n2449 ) ;
  assign n2451 = n2448 & ~n2450 ;
  assign n2452 = x87 | n2451 ;
  assign n2453 = n2447 & n2452 ;
  assign n2454 = x58 | n1270 ;
  assign n2455 = n1205 | n1326 ;
  assign n2456 = n1319 | n2455 ;
  assign n2457 = n1213 | n1340 ;
  assign n2458 = n2456 | n2457 ;
  assign n2459 = x39 | n2458 ;
  assign n2460 = n2454 | n2459 ;
  assign n2461 = n1275 | n1354 ;
  assign n2462 = n1281 | n2461 ;
  assign n2463 = ( x87 & n1281 ) | ( x87 & n2462 ) | ( n1281 & n2462 ) ;
  assign n2464 = n2460 | n2463 ;
  assign n2465 = n1254 | n2464 ;
  assign n2466 = n2453 & ~n2465 ;
  assign n2467 = ~x122 & n2445 ;
  assign n2468 = x286 | x288 ;
  assign n2469 = x285 | x289 ;
  assign n2470 = n2468 | n2469 ;
  assign n2471 = n2467 & n2470 ;
  assign n2472 = ~x217 & n2471 ;
  assign n2473 = ( ~x217 & n2466 ) | ( ~x217 & n2472 ) | ( n2466 & n2472 ) ;
  assign n2474 = n2182 | n2473 ;
  assign n2475 = ( n2182 & n2443 ) | ( n2182 & n2474 ) | ( n2443 & n2474 ) ;
  assign n2476 = n2180 | n2475 ;
  assign n2477 = x166 & x299 ;
  assign n2478 = x189 & ~x299 ;
  assign n2479 = n2477 | n2478 ;
  assign n2480 = ~x161 & x299 ;
  assign n2481 = x144 | x299 ;
  assign n2482 = ( n2072 & n2480 ) | ( n2072 & ~n2481 ) | ( n2480 & ~n2481 ) ;
  assign n2483 = ~n2479 & n2482 ;
  assign n2484 = x174 & ~x299 ;
  assign n2485 = n1910 | n2484 ;
  assign n2486 = n2483 & ~n2485 ;
  assign n2487 = n1950 & ~n2486 ;
  assign n2488 = x252 & n2487 ;
  assign n2489 = x24 | x122 ;
  assign n2490 = n1313 & ~n2489 ;
  assign n2491 = ( n1507 & n2489 ) | ( n1507 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2492 = ( ~n1435 & n1507 ) | ( ~n1435 & n2491 ) | ( n1507 & n2491 ) ;
  assign n2493 = ( n1507 & ~n2488 ) | ( n1507 & n2492 ) | ( ~n2488 & n2492 ) ;
  assign n2494 = n1213 | n2493 ;
  assign n2495 = ~x39 & n1995 ;
  assign n2496 = ( n1993 & n2043 ) | ( n1993 & n2044 ) | ( n2043 & n2044 ) ;
  assign n2497 = n2017 & n2496 ;
  assign n2498 = ( n1995 & n2495 ) | ( n1995 & n2497 ) | ( n2495 & n2497 ) ;
  assign n2499 = ~n2494 & n2498 ;
  assign n2500 = ~n1337 & n2499 ;
  assign n2501 = x72 | x122 ;
  assign n2502 = ( n1346 & n2049 ) | ( n1346 & ~n2501 ) | ( n2049 & ~n2501 ) ;
  assign n2503 = n2501 | n2502 ;
  assign n2504 = ~x96 & x1093 ;
  assign n2505 = x841 & ~n2504 ;
  assign n2506 = ( n1271 & ~n2504 ) | ( n1271 & n2505 ) | ( ~n2504 & n2505 ) ;
  assign n2507 = n1434 & ~n2506 ;
  assign n2508 = ( n1254 & n1381 ) | ( n1254 & ~n2454 ) | ( n1381 & ~n2454 ) ;
  assign n2509 = n2454 | n2508 ;
  assign n2510 = x97 & ~n2509 ;
  assign n2511 = x96 | n2510 ;
  assign n2512 = n2507 & n2511 ;
  assign n2513 = ~x24 & n1362 ;
  assign n2514 = ( n2507 & n2512 ) | ( n2507 & n2513 ) | ( n2512 & n2513 ) ;
  assign n2515 = ~n2503 & n2514 ;
  assign n2516 = ~n1254 & n1481 ;
  assign n2517 = ( ~x98 & n1387 ) | ( ~x98 & n2516 ) | ( n1387 & n2516 ) ;
  assign n2518 = n2516 & ~n2517 ;
  assign n2519 = ~n1359 & n2451 ;
  assign n2520 = ( ~n1359 & n2518 ) | ( ~n1359 & n2519 ) | ( n2518 & n2519 ) ;
  assign n2521 = n2515 | n2520 ;
  assign n2522 = x100 & n2501 ;
  assign n2523 = ( x100 & ~n1435 ) | ( x100 & n2522 ) | ( ~n1435 & n2522 ) ;
  assign n2524 = x228 & ~n2051 ;
  assign n2525 = n2487 & n2524 ;
  assign n2526 = ( x100 & n2523 ) | ( x100 & ~n2525 ) | ( n2523 & ~n2525 ) ;
  assign n2527 = ( n1311 & n2521 ) | ( n1311 & ~n2526 ) | ( n2521 & ~n2526 ) ;
  assign n2528 = n2471 | n2527 ;
  assign n2529 = ( n2471 & n2500 ) | ( n2471 & n2528 ) | ( n2500 & n2528 ) ;
  assign n2530 = ~n2476 & n2529 ;
  assign n2531 = x1161 & x1162 ;
  assign n2532 = ~x1163 & n2531 ;
  assign n2533 = n2178 & ~n2532 ;
  assign n2534 = ( n2178 & n2530 ) | ( n2178 & ~n2533 ) | ( n2530 & ~n2533 ) ;
  assign n2535 = ~n1434 & n2470 ;
  assign n2536 = x137 | n2027 ;
  assign n2537 = n2535 | n2536 ;
  assign n2538 = x252 & ~n2487 ;
  assign n2539 = ~x24 & x75 ;
  assign n2540 = ~n1313 & n2539 ;
  assign n2541 = n1434 & n2540 ;
  assign n2542 = n2538 & n2541 ;
  assign n2543 = ~n1434 & n2540 ;
  assign n2544 = ( ~n1954 & n2542 ) | ( ~n1954 & n2543 ) | ( n2542 & n2543 ) ;
  assign n2545 = ~n2538 & n2544 ;
  assign n2546 = x100 & ~n1211 ;
  assign n2547 = ~n1954 & n2546 ;
  assign n2548 = ( ~x250 & n1951 ) | ( ~x250 & n1952 ) | ( n1951 & n1952 ) ;
  assign n2549 = ~n1960 & n2548 ;
  assign n2550 = x129 & ~n2548 ;
  assign n2551 = ( n2547 & n2549 ) | ( n2547 & n2550 ) | ( n2549 & n2550 ) ;
  assign n2552 = n1953 | n2538 ;
  assign n2553 = ( x137 & n2551 ) | ( x137 & ~n2552 ) | ( n2551 & ~n2552 ) ;
  assign n2554 = n2551 & ~n2553 ;
  assign n2555 = ( ~x137 & n2545 ) | ( ~x137 & n2554 ) | ( n2545 & n2554 ) ;
  assign n2556 = n1208 | n1282 ;
  assign n2557 = n1213 | n2556 ;
  assign n2558 = n2555 & ~n2557 ;
  assign n2559 = n1309 | n2462 ;
  assign n2560 = n2454 | n2559 ;
  assign n2561 = n1409 | n2560 ;
  assign n2562 = x76 & ~n1401 ;
  assign n2563 = ~n2561 & n2562 ;
  assign n2564 = n2537 | n2563 ;
  assign n2565 = ( ~n2537 & n2558 ) | ( ~n2537 & n2564 ) | ( n2558 & n2564 ) ;
  assign n2566 = ~x24 & x50 ;
  assign n2567 = ( ~x841 & n2025 ) | ( ~x841 & n2026 ) | ( n2025 & n2026 ) ;
  assign n2568 = ( x24 & x841 ) | ( x24 & ~n2567 ) | ( x841 & ~n2567 ) ;
  assign n2569 = x32 & n2568 ;
  assign n2570 = ( ~n2565 & n2566 ) | ( ~n2565 & n2569 ) | ( n2566 & n2569 ) ;
  assign n2571 = n2565 | n2570 ;
  assign n2572 = n1313 | n1415 ;
  assign n2573 = ~n1337 & n2572 ;
  assign n2574 = ( n2565 & n2571 ) | ( n2565 & n2573 ) | ( n2571 & n2573 ) ;
  assign n2575 = ~x33 & x954 ;
  assign n2576 = n1205 | n1875 ;
  assign n2577 = x40 | x63 ;
  assign n2578 = x107 | n2577 ;
  assign n2579 = n2576 | n2578 ;
  assign n2580 = n2161 | n2579 ;
  assign n2581 = n1254 | n1372 ;
  assign n2582 = n2454 | n2581 ;
  assign n2583 = x70 | n1420 ;
  assign n2584 = x50 | n2583 ;
  assign n2585 = ~n1359 & n2584 ;
  assign n2586 = ~n2582 & n2585 ;
  assign n2587 = n2039 | n2586 ;
  assign n2588 = x73 & ~n1359 ;
  assign n2589 = n1487 & n2588 ;
  assign n2590 = n1278 | n1347 ;
  assign n2591 = x90 & ~x841 ;
  assign n2592 = ( x58 & ~x95 ) | ( x58 & n2591 ) | ( ~x95 & n2591 ) ;
  assign n2593 = ~x51 & n2592 ;
  assign n2594 = ~n1356 & n2593 ;
  assign n2595 = ( ~n1271 & n2590 ) | ( ~n1271 & n2594 ) | ( n2590 & n2594 ) ;
  assign n2596 = ~n2590 & n2595 ;
  assign n2597 = n2589 | n2596 ;
  assign n2598 = n2587 | n2597 ;
  assign n2599 = n2024 | n2598 ;
  assign n2600 = n2043 | n2044 ;
  assign n2601 = ( x39 & n2019 ) | ( x39 & n2021 ) | ( n2019 & n2021 ) ;
  assign n2602 = ~n1266 & n2601 ;
  assign n2603 = n1272 | n2454 ;
  assign n2604 = n1972 | n2603 ;
  assign n2605 = n1221 | n1239 ;
  assign n2606 = n1250 | n2154 ;
  assign n2607 = n2605 | n2606 ;
  assign n2608 = ( n2602 & n2604 ) | ( n2602 & n2607 ) | ( n2604 & n2607 ) ;
  assign n2609 = n2602 & ~n2608 ;
  assign n2610 = ~n2600 & n2609 ;
  assign n2611 = x1093 & n1992 ;
  assign n2612 = n2014 & n2611 ;
  assign n2613 = x110 | n2045 ;
  assign n2614 = n2601 & ~n2613 ;
  assign n2615 = n2612 & n2614 ;
  assign n2616 = n2610 & n2615 ;
  assign n2617 = x73 & ~n2610 ;
  assign n2618 = ~n1312 & n2573 ;
  assign n2619 = ( n2616 & n2617 ) | ( n2616 & n2618 ) | ( n2617 & n2618 ) ;
  assign n2620 = ( ~n1337 & n2599 ) | ( ~n1337 & n2619 ) | ( n2599 & n2619 ) ;
  assign n2621 = n2580 | n2620 ;
  assign n2622 = x139 | x195 ;
  assign n2623 = ( ~x118 & x138 ) | ( ~x118 & x196 ) | ( x138 & x196 ) ;
  assign n2624 = ( ~x118 & n2622 ) | ( ~x118 & n2623 ) | ( n2622 & n2623 ) ;
  assign n2625 = x118 | n2624 ;
  assign n2626 = x33 | x34 ;
  assign n2627 = x79 | n2626 ;
  assign n2628 = n2625 | n2627 ;
  assign n2629 = ( ~x33 & x954 ) | ( ~x33 & n2628 ) | ( x954 & n2628 ) ;
  assign n2630 = ( ~n2575 & n2621 ) | ( ~n2575 & n2629 ) | ( n2621 & n2629 ) ;
  assign n2631 = n1319 & n2072 ;
  assign n2632 = ( x149 & x157 ) | ( x149 & ~n2631 ) | ( x157 & ~n2631 ) ;
  assign n2633 = x149 | x157 ;
  assign n2634 = ~n2079 & n2633 ;
  assign n2635 = ~n2632 & n2634 ;
  assign n2636 = x178 | x183 ;
  assign n2637 = n1319 & n2079 ;
  assign n2638 = ( x178 & x183 ) | ( x178 & ~n2637 ) | ( x183 & ~n2637 ) ;
  assign n2639 = ( n2635 & n2636 ) | ( n2635 & ~n2638 ) | ( n2636 & ~n2638 ) ;
  assign n2640 = ~n1208 & n2639 ;
  assign n2641 = x38 & n1322 ;
  assign n2642 = ( x38 & n1282 ) | ( x38 & n2641 ) | ( n1282 & n2641 ) ;
  assign n2643 = x54 | n2642 ;
  assign n2644 = x191 & ~x299 ;
  assign n2645 = x169 & x299 ;
  assign n2646 = ( n2072 & n2644 ) | ( n2072 & n2645 ) | ( n2644 & n2645 ) ;
  assign n2647 = ( n1319 & n1320 ) | ( n1319 & n2646 ) | ( n1320 & n2646 ) ;
  assign n2648 = x154 & x299 ;
  assign n2649 = x176 & ~x299 ;
  assign n2650 = n2648 | n2649 ;
  assign n2651 = n1435 & n2650 ;
  assign n2652 = ( x39 & n2020 ) | ( x39 & n2022 ) | ( n2020 & n2022 ) ;
  assign n2653 = ~n2093 & n2652 ;
  assign n2654 = n1992 & n2072 ;
  assign n2655 = ( ~n2003 & n2011 ) | ( ~n2003 & n2654 ) | ( n2011 & n2654 ) ;
  assign n2656 = n2654 & ~n2655 ;
  assign n2657 = n2653 & n2656 ;
  assign n2658 = ~n1433 & n1958 ;
  assign n2659 = ~x1093 & n1958 ;
  assign n2660 = ( n1429 & ~n1433 ) | ( n1429 & n2659 ) | ( ~n1433 & n2659 ) ;
  assign n2661 = n2658 & ~n2660 ;
  assign n2662 = ~n2485 & n2661 ;
  assign n2663 = ( n2651 & n2657 ) | ( n2651 & n2662 ) | ( n2657 & n2662 ) ;
  assign n2664 = n2072 & n2650 ;
  assign n2665 = n1877 & n2664 ;
  assign n2666 = ( ~n2647 & n2663 ) | ( ~n2647 & n2665 ) | ( n2663 & n2665 ) ;
  assign n2667 = n2647 | n2666 ;
  assign n2668 = ( ~n1282 & n2647 ) | ( ~n1282 & n2667 ) | ( n2647 & n2667 ) ;
  assign n2669 = x164 & x299 ;
  assign n2670 = x186 & ~x299 ;
  assign n2671 = ( ~x74 & n2669 ) | ( ~x74 & n2670 ) | ( n2669 & n2670 ) ;
  assign n2672 = n2072 & n2671 ;
  assign n2673 = n2668 | n2672 ;
  assign n2674 = ( n2643 & n2668 ) | ( n2643 & n2673 ) | ( n2668 & n2673 ) ;
  assign n2675 = ( n1208 & ~n2640 ) | ( n1208 & n2674 ) | ( ~n2640 & n2674 ) ;
  assign n2676 = ~n1215 & n2072 ;
  assign n2677 = ( n2485 & ~n2589 ) | ( n2485 & n2676 ) | ( ~n2589 & n2676 ) ;
  assign n2678 = n2676 & ~n2677 ;
  assign n2679 = ~n1277 & n1445 ;
  assign n2680 = n2586 | n2679 ;
  assign n2681 = x149 & x299 ;
  assign n2682 = n2680 & n2681 ;
  assign n2683 = ~n1276 & n1301 ;
  assign n2684 = x158 & x299 ;
  assign n2685 = x180 & ~x299 ;
  assign n2686 = ( ~n2590 & n2684 ) | ( ~n2590 & n2685 ) | ( n2684 & n2685 ) ;
  assign n2687 = n2683 & n2686 ;
  assign n2688 = x193 & ~x299 ;
  assign n2689 = x172 & x299 ;
  assign n2690 = ( n2594 & n2688 ) | ( n2594 & n2689 ) | ( n2688 & n2689 ) ;
  assign n2691 = ( ~n2590 & n2687 ) | ( ~n2590 & n2690 ) | ( n2687 & n2690 ) ;
  assign n2692 = ~n1271 & n2691 ;
  assign n2693 = n1468 & ~n1538 ;
  assign n2694 = x183 & ~x299 ;
  assign n2695 = ( n2586 & n2693 ) | ( n2586 & n2694 ) | ( n2693 & n2694 ) ;
  assign n2696 = n2692 | n2695 ;
  assign n2697 = n2682 | n2696 ;
  assign n2698 = ( n2676 & n2678 ) | ( n2676 & n2697 ) | ( n2678 & n2697 ) ;
  assign n2699 = n2675 | n2698 ;
  assign n2700 = x169 & n1320 ;
  assign n2701 = ~x74 & n2455 ;
  assign n2702 = x164 & n2701 ;
  assign n2703 = ( n2072 & n2700 ) | ( n2072 & n2702 ) | ( n2700 & n2702 ) ;
  assign n2704 = n1319 | n2703 ;
  assign n2705 = ( n2632 & ~n2633 ) | ( n2632 & n2704 ) | ( ~n2633 & n2704 ) ;
  assign n2706 = n1207 & ~n2705 ;
  assign n2707 = x149 & ~n1282 ;
  assign n2708 = x55 & ~n2676 ;
  assign n2709 = ( x55 & ~n2707 ) | ( x55 & n2708 ) | ( ~n2707 & n2708 ) ;
  assign n2710 = ( ~n2705 & n2706 ) | ( ~n2705 & n2709 ) | ( n2706 & n2709 ) ;
  assign n2711 = ( n2630 & ~n2699 ) | ( n2630 & n2710 ) | ( ~n2699 & n2710 ) ;
  assign n2712 = ~n2158 & n2683 ;
  assign n2713 = x73 & x161 ;
  assign n2714 = x146 | n2713 ;
  assign n2715 = ( n2594 & n2713 ) | ( n2594 & n2714 ) | ( n2713 & n2714 ) ;
  assign n2716 = n2073 & ~n2715 ;
  assign n2717 = x159 & n2716 ;
  assign n2718 = ( ~n2712 & n2716 ) | ( ~n2712 & n2717 ) | ( n2716 & n2717 ) ;
  assign n2719 = x162 & n2718 ;
  assign n2720 = ( ~n2680 & n2718 ) | ( ~n2680 & n2719 ) | ( n2718 & n2719 ) ;
  assign n2721 = ( n1317 & n2598 ) | ( n1317 & ~n2720 ) | ( n2598 & ~n2720 ) ;
  assign n2722 = ~x142 & n1273 ;
  assign n2723 = x140 & ~n1273 ;
  assign n2724 = ( ~x73 & n2722 ) | ( ~x73 & n2723 ) | ( n2722 & n2723 ) ;
  assign n2725 = n2712 | n2724 ;
  assign n2726 = x73 & ~x144 ;
  assign n2727 = ~x181 & n2712 ;
  assign n2728 = ( n2725 & n2726 ) | ( n2725 & ~n2727 ) | ( n2726 & ~n2727 ) ;
  assign n2729 = n2079 & n2728 ;
  assign n2730 = ( n1317 & n2721 ) | ( n1317 & ~n2729 ) | ( n2721 & ~n2729 ) ;
  assign n2731 = ~n1317 & n2730 ;
  assign n2732 = n1207 | n1212 ;
  assign n2733 = x162 & n2072 ;
  assign n2734 = ( n1317 & ~n2732 ) | ( n1317 & n2733 ) | ( ~n2732 & n2733 ) ;
  assign n2735 = n2732 | n2734 ;
  assign n2736 = n2159 | n2735 ;
  assign n2737 = ( x140 & x145 ) | ( x140 & n2636 ) | ( x145 & n2636 ) ;
  assign n2738 = ( ~x140 & x145 ) | ( ~x140 & n2636 ) | ( x145 & n2636 ) ;
  assign n2739 = ( x140 & ~n2737 ) | ( x140 & n2738 ) | ( ~n2737 & n2738 ) ;
  assign n2740 = ~n1553 & n2739 ;
  assign n2741 = ( ~x162 & x197 ) | ( ~x162 & n2633 ) | ( x197 & n2633 ) ;
  assign n2742 = ( x162 & x197 ) | ( x162 & n2633 ) | ( x197 & n2633 ) ;
  assign n2743 = ( x162 & n2741 ) | ( x162 & ~n2742 ) | ( n2741 & ~n2742 ) ;
  assign n2744 = n1553 & n2743 ;
  assign n2745 = ( n1319 & n2740 ) | ( n1319 & n2744 ) | ( n2740 & n2744 ) ;
  assign n2746 = x188 & ~x299 ;
  assign n2747 = x54 & ~x74 ;
  assign n2748 = x167 & x299 ;
  assign n2749 = ( n2746 & n2747 ) | ( n2746 & n2748 ) | ( n2747 & n2748 ) ;
  assign n2750 = x148 & x299 ;
  assign n2751 = x141 & ~x299 ;
  assign n2752 = ( x74 & n2750 ) | ( x74 & n2751 ) | ( n2750 & n2751 ) ;
  assign n2753 = ( ~n1208 & n2749 ) | ( ~n1208 & n2752 ) | ( n2749 & n2752 ) ;
  assign n2754 = ( n1208 & ~n1319 ) | ( n1208 & n2753 ) | ( ~n1319 & n2753 ) ;
  assign n2755 = n2745 | n2754 ;
  assign n2756 = ( n2736 & n2745 ) | ( n2736 & n2755 ) | ( n2745 & n2755 ) ;
  assign n2757 = x68 | x71 ;
  assign n2758 = n1390 | n2757 ;
  assign n2759 = x51 | x87 ;
  assign n2760 = n2758 | n2759 ;
  assign n2761 = n2610 & ~n2760 ;
  assign n2762 = n2612 & n2761 ;
  assign n2763 = x155 & x299 ;
  assign n2764 = x177 & ~x299 ;
  assign n2765 = ( n2072 & n2763 ) | ( n2072 & n2764 ) | ( n2763 & n2764 ) ;
  assign n2766 = n1435 & ~n2765 ;
  assign n2767 = n1435 | n2482 ;
  assign n2768 = ( x92 & ~n2766 ) | ( x92 & n2767 ) | ( ~n2766 & n2767 ) ;
  assign n2769 = n2762 & ~n2768 ;
  assign n2770 = ~n1327 & n2765 ;
  assign n2771 = n1876 & ~n2159 ;
  assign n2772 = ( n1327 & ~n2770 ) | ( n1327 & n2771 ) | ( ~n2770 & n2771 ) ;
  assign n2773 = n2769 | n2772 ;
  assign n2774 = ( n2642 & n2746 ) | ( n2642 & n2748 ) | ( n2746 & n2748 ) ;
  assign n2775 = ( n1320 & n2773 ) | ( n1320 & ~n2774 ) | ( n2773 & ~n2774 ) ;
  assign n2776 = ~n2756 & n2775 ;
  assign n2777 = ( n2731 & ~n2756 ) | ( n2731 & n2776 ) | ( ~n2756 & n2776 ) ;
  assign n2778 = x167 & n1208 ;
  assign n2779 = ( ~n1208 & n2701 ) | ( ~n1208 & n2778 ) | ( n2701 & n2778 ) ;
  assign n2780 = ~x148 & n1208 ;
  assign n2781 = ( n1319 & n1320 ) | ( n1319 & ~n2780 ) | ( n1320 & ~n2780 ) ;
  assign n2782 = n2779 | n2781 ;
  assign n2783 = ~n2072 & n2579 ;
  assign n2784 = ( n2579 & ~n2782 ) | ( n2579 & n2783 ) | ( ~n2782 & n2783 ) ;
  assign n2785 = n2777 | n2784 ;
  assign n2786 = x33 | x954 ;
  assign n2787 = ( x34 & n2628 ) | ( x34 & ~n2786 ) | ( n2628 & ~n2786 ) ;
  assign n2788 = n2628 & ~n2786 ;
  assign n2789 = ( x34 & n2621 ) | ( x34 & n2788 ) | ( n2621 & n2788 ) ;
  assign n2790 = ( n2785 & n2787 ) | ( n2785 & ~n2789 ) | ( n2787 & ~n2789 ) ;
  assign n2791 = x683 & n2658 ;
  assign n2792 = n2488 & ~n2791 ;
  assign n2793 = n2551 & ~n2792 ;
  assign n2794 = ~n1965 & n2793 ;
  assign n2795 = x38 & ~n1336 ;
  assign n2796 = ~x24 & n2732 ;
  assign n2797 = ( ~x24 & n2795 ) | ( ~x24 & n2796 ) | ( n2795 & n2796 ) ;
  assign n2798 = n2544 | n2797 ;
  assign n2799 = ( ~n1965 & n2794 ) | ( ~n1965 & n2798 ) | ( n2794 & n2798 ) ;
  assign n2800 = ( n1332 & n2555 ) | ( n1332 & n2799 ) | ( n2555 & n2799 ) ;
  assign n2801 = n2799 & ~n2800 ;
  assign n2802 = x35 & ~x841 ;
  assign n2803 = ~n1538 & n2028 ;
  assign n2804 = ~x24 & n2803 ;
  assign n2805 = ~x93 & x841 ;
  assign n2806 = x93 | n1351 ;
  assign n2807 = x40 & x1082 ;
  assign n2808 = x76 & ~x122 ;
  assign n2809 = ( n1960 & ~n2536 ) | ( n1960 & n2808 ) | ( ~n2536 & n2808 ) ;
  assign n2810 = n2808 & ~n2809 ;
  assign n2811 = n2535 & ~n2807 ;
  assign n2812 = ( n2807 & n2810 ) | ( n2807 & ~n2811 ) | ( n2810 & ~n2811 ) ;
  assign n2813 = n2806 | n2812 ;
  assign n2814 = x35 | x841 ;
  assign n2815 = ( n2805 & n2813 ) | ( n2805 & ~n2814 ) | ( n2813 & ~n2814 ) ;
  assign n2816 = ( ~n2802 & n2804 ) | ( ~n2802 & n2815 ) | ( n2804 & n2815 ) ;
  assign n2817 = n2801 | n2816 ;
  assign n2818 = ( n2141 & n2801 ) | ( n2141 & n2817 ) | ( n2801 & n2817 ) ;
  assign n2819 = x58 | n2559 ;
  assign n2820 = x36 & n1412 ;
  assign n2821 = ( n2513 & ~n2819 ) | ( n2513 & n2820 ) | ( ~n2819 & n2820 ) ;
  assign n2822 = n1960 & n2821 ;
  assign n2823 = n1487 & ~n2819 ;
  assign n2824 = x89 & x332 ;
  assign n2825 = x64 & ~x841 ;
  assign n2826 = ( ~x841 & n2824 ) | ( ~x841 & n2825 ) | ( n2824 & n2825 ) ;
  assign n2827 = n2823 & n2826 ;
  assign n2828 = x24 & ~n1324 ;
  assign n2829 = x46 | x97 ;
  assign n2830 = ( x108 & n2560 ) | ( x108 & ~n2829 ) | ( n2560 & ~n2829 ) ;
  assign n2831 = n2829 | n2830 ;
  assign n2832 = ( n2557 & n2828 ) | ( n2557 & ~n2831 ) | ( n2828 & ~n2831 ) ;
  assign n2833 = n2828 & ~n2832 ;
  assign n2834 = n2827 | n2833 ;
  assign n2835 = x786 & ~x1082 ;
  assign n2836 = ( n2015 & ~n2132 ) | ( n2015 & n2835 ) | ( ~n2132 & n2835 ) ;
  assign n2837 = n2835 & ~n2836 ;
  assign n2838 = ( x48 & ~x841 ) | ( x48 & n2802 ) | ( ~x841 & n2802 ) ;
  assign n2839 = x47 | n2838 ;
  assign n2840 = x108 & x314 ;
  assign n2841 = x986 | n1960 ;
  assign n2842 = ~x252 & n2840 ;
  assign n2843 = ( n2840 & ~n2841 ) | ( n2840 & n2842 ) | ( ~n2841 & n2842 ) ;
  assign n2844 = ( ~x47 & n2136 ) | ( ~x47 & n2843 ) | ( n2136 & n2843 ) ;
  assign n2845 = ~n2837 & n2844 ;
  assign n2846 = ( ~n2837 & n2839 ) | ( ~n2837 & n2845 ) | ( n2839 & n2845 ) ;
  assign n2847 = ( n1280 & n1359 ) | ( n1280 & ~n2567 ) | ( n1359 & ~n2567 ) ;
  assign n2848 = ( n1359 & n2846 ) | ( n1359 & ~n2847 ) | ( n2846 & ~n2847 ) ;
  assign n2849 = n2618 & n2848 ;
  assign n2850 = x40 | x102 ;
  assign n2851 = ( ~n2573 & n2807 ) | ( ~n2573 & n2850 ) | ( n2807 & n2850 ) ;
  assign n2852 = n2850 & ~n2851 ;
  assign n2853 = x39 & ~x72 ;
  assign n2854 = ( x41 & x72 ) | ( x41 & ~n2853 ) | ( x72 & ~n2853 ) ;
  assign n2855 = x39 & ~x152 ;
  assign n2856 = ~x161 & n2855 ;
  assign n2857 = ~x166 & n2072 ;
  assign n2858 = x287 & ~n2093 ;
  assign n2859 = ~n2051 & n2858 ;
  assign n2860 = ( n1208 & n1553 ) | ( n1208 & ~n2859 ) | ( n1553 & ~n2859 ) ;
  assign n2861 = n2857 & n2860 ;
  assign n2862 = ( n2855 & n2856 ) | ( n2855 & n2861 ) | ( n2856 & n2861 ) ;
  assign n2863 = ( n2854 & ~n2856 ) | ( n2854 & n2862 ) | ( ~n2856 & n2862 ) ;
  assign n2864 = ~x189 & n2079 ;
  assign n2865 = ~n1208 & n2864 ;
  assign n2866 = ~n2859 & n2865 ;
  assign n2867 = ~x144 & n2866 ;
  assign n2868 = x144 & x174 ;
  assign n2869 = x39 & ~n2868 ;
  assign n2870 = ( n2866 & n2867 ) | ( n2866 & n2869 ) | ( n2867 & n2869 ) ;
  assign n2871 = ( n2863 & ~n2867 ) | ( n2863 & n2870 ) | ( ~n2867 & n2870 ) ;
  assign n2872 = x101 & n2871 ;
  assign n2873 = x44 | n1208 ;
  assign n2874 = ~x72 & n1210 ;
  assign n2875 = ( n2494 & ~n2524 ) | ( n2494 & n2874 ) | ( ~n2524 & n2874 ) ;
  assign n2876 = n2874 & ~n2875 ;
  assign n2877 = ~n2526 & n2876 ;
  assign n2878 = x228 & n2521 ;
  assign n2879 = ( ~n1214 & n1515 ) | ( ~n1214 & n2878 ) | ( n1515 & n2878 ) ;
  assign n2880 = x901 & ~x959 ;
  assign n2881 = x94 & ~n2509 ;
  assign n2882 = ~x250 & x252 ;
  assign n2883 = ( ~n2880 & n2881 ) | ( ~n2880 & n2882 ) | ( n2881 & n2882 ) ;
  assign n2884 = n2880 & n2883 ;
  assign n2885 = x110 & ~x480 ;
  assign n2886 = ~x949 & n2885 ;
  assign n2887 = ( n2884 & n2885 ) | ( n2884 & ~n2886 ) | ( n2885 & ~n2886 ) ;
  assign n2888 = ( n1214 & n1558 ) | ( n1214 & ~n2887 ) | ( n1558 & ~n2887 ) ;
  assign n2889 = ( n1558 & n2879 ) | ( n1558 & ~n2888 ) | ( n2879 & ~n2888 ) ;
  assign n2890 = ( ~n2526 & n2877 ) | ( ~n2526 & n2889 ) | ( n2877 & n2889 ) ;
  assign n2891 = ~n2873 & n2890 ;
  assign n2892 = ( ~x101 & n2871 ) | ( ~x101 & n2891 ) | ( n2871 & n2891 ) ;
  assign n2893 = n2871 & n2891 ;
  assign n2894 = ( n2872 & n2892 ) | ( n2872 & ~n2893 ) | ( n2892 & ~n2893 ) ;
  assign n2895 = x39 | x72 ;
  assign n2896 = x42 & ~n2895 ;
  assign n2897 = ~n1946 & n2891 ;
  assign n2898 = ~x114 & n2897 ;
  assign n2899 = n2896 & ~n2898 ;
  assign n2900 = ~n1948 & n2890 ;
  assign n2901 = ~n1208 & n2900 ;
  assign n2902 = n2853 & ~n2861 ;
  assign n2903 = x207 & x208 ;
  assign n2904 = x199 | x200 ;
  assign n2905 = ( x199 & n2903 ) | ( x199 & n2904 ) | ( n2903 & n2904 ) ;
  assign n2906 = n1553 | n2905 ;
  assign n2907 = x211 | x219 ;
  assign n2908 = x212 & x214 ;
  assign n2909 = ( x219 & n2907 ) | ( x219 & n2908 ) | ( n2907 & n2908 ) ;
  assign n2910 = n1553 & ~n2909 ;
  assign n2911 = n2906 & ~n2910 ;
  assign n2912 = ~n2866 & n2911 ;
  assign n2913 = n2902 & ~n2912 ;
  assign n2914 = ( n2901 & n2902 ) | ( n2901 & ~n2913 ) | ( n2902 & ~n2913 ) ;
  assign n2915 = n2899 | n2914 ;
  assign n2916 = ~x39 & x43 ;
  assign n2917 = x211 & ~n2908 ;
  assign n2918 = ~n2907 & n2908 ;
  assign n2919 = ( x39 & n2917 ) | ( x39 & n2918 ) | ( n2917 & n2918 ) ;
  assign n2920 = ~n2857 & n2919 ;
  assign n2921 = ( n1208 & n2916 ) | ( n1208 & ~n2920 ) | ( n2916 & ~n2920 ) ;
  assign n2922 = ( x72 & ~n2916 ) | ( x72 & n2921 ) | ( ~n2916 & n2921 ) ;
  assign n2923 = x43 & n2900 ;
  assign n2924 = n2900 | n2916 ;
  assign n2925 = x200 & ~n2903 ;
  assign n2926 = n2903 & ~n2904 ;
  assign n2927 = ( ~x299 & n2925 ) | ( ~x299 & n2926 ) | ( n2925 & n2926 ) ;
  assign n2928 = ( x299 & n2917 ) | ( x299 & n2918 ) | ( n2917 & n2918 ) ;
  assign n2929 = ( x39 & n2927 ) | ( x39 & n2928 ) | ( n2927 & n2928 ) ;
  assign n2930 = n1208 | n2929 ;
  assign n2931 = n2072 & ~n2479 ;
  assign n2932 = ~n2859 & n2931 ;
  assign n2933 = ( n1208 & n2930 ) | ( n1208 & ~n2932 ) | ( n2930 & ~n2932 ) ;
  assign n2934 = ( ~n2923 & n2924 ) | ( ~n2923 & n2933 ) | ( n2924 & n2933 ) ;
  assign n2935 = ~n2922 & n2934 ;
  assign n2936 = x39 | x44 ;
  assign n2937 = x39 & ~n2486 ;
  assign n2938 = ( x39 & n2859 ) | ( x39 & n2937 ) | ( n2859 & n2937 ) ;
  assign n2939 = ( n1208 & n2936 ) | ( n1208 & ~n2938 ) | ( n2936 & ~n2938 ) ;
  assign n2940 = ~n2890 & n2939 ;
  assign n2941 = ~x72 & n2940 ;
  assign n2942 = ~n1437 & n2072 ;
  assign n2943 = x39 & ~n2942 ;
  assign n2944 = ( n1208 & ~n2936 ) | ( n1208 & n2943 ) | ( ~n2936 & n2943 ) ;
  assign n2945 = ( n1208 & ~n2873 ) | ( n1208 & n2890 ) | ( ~n2873 & n2890 ) ;
  assign n2946 = ( n2941 & ~n2944 ) | ( n2941 & n2945 ) | ( ~n2944 & n2945 ) ;
  assign n2947 = ~n1337 & n2128 ;
  assign n2948 = x979 & n2947 ;
  assign n2949 = x61 & x841 ;
  assign n2950 = x24 & n1483 ;
  assign n2951 = ( x61 & ~n2949 ) | ( x61 & n2950 ) | ( ~n2949 & n2950 ) ;
  assign n2952 = n2823 & n2951 ;
  assign n2953 = ~n2660 & n2821 ;
  assign n2954 = x88 | x104 ;
  assign n2955 = ~n2658 & n2954 ;
  assign n2956 = n2823 & ~n2955 ;
  assign n2957 = ( n2823 & n2953 ) | ( n2823 & ~n2956 ) | ( n2953 & ~n2956 ) ;
  assign n2958 = x48 & x841 ;
  assign n2959 = n2823 & n2958 ;
  assign n2960 = x49 & x841 ;
  assign n2961 = n2823 & n2960 ;
  assign n2962 = n1557 | n2456 ;
  assign n2963 = n1282 | n2962 ;
  assign n2964 = n2797 & ~n2963 ;
  assign n2965 = n2961 | n2964 ;
  assign n2966 = n1257 | n1260 ;
  assign n2967 = ( n1265 & n1420 ) | ( n1265 & ~n2966 ) | ( n1420 & ~n2966 ) ;
  assign n2968 = n2966 | n2967 ;
  assign n2969 = ( n1254 & n2560 ) | ( n1254 & ~n2968 ) | ( n2560 & ~n2968 ) ;
  assign n2970 = n2968 | n2969 ;
  assign n2971 = x24 & ~x94 ;
  assign n2972 = x252 & n1434 ;
  assign n2973 = ~x252 & n2487 ;
  assign n2974 = ( ~x50 & n2972 ) | ( ~x50 & n2973 ) | ( n2972 & n2973 ) ;
  assign n2975 = n2971 | n2974 ;
  assign n2976 = ~n2970 & n2975 ;
  assign n2977 = n2557 & ~n2976 ;
  assign n2978 = n1515 & n1963 ;
  assign n2979 = ( n1954 & n2543 ) | ( n1954 & n2978 ) | ( n2543 & n2978 ) ;
  assign n2980 = n2557 | n2979 ;
  assign n2981 = ~n2977 & n2980 ;
  assign n2982 = n1411 & ~n2560 ;
  assign n2983 = x82 & n2982 ;
  assign n2984 = ~x43 & n2901 ;
  assign n2985 = x52 & ~n2895 ;
  assign n2986 = ( n1553 & n2907 ) | ( n1553 & n2918 ) | ( n2907 & n2918 ) ;
  assign n2987 = ( ~n1553 & n2904 ) | ( ~n1553 & n2926 ) | ( n2904 & n2926 ) ;
  assign n2988 = n2986 | n2987 ;
  assign n2989 = ( ~n2866 & n2902 ) | ( ~n2866 & n2988 ) | ( n2902 & n2988 ) ;
  assign n2990 = ~n2988 & n2989 ;
  assign n2991 = ( ~n2984 & n2985 ) | ( ~n2984 & n2990 ) | ( n2985 & n2990 ) ;
  assign n2992 = n2984 & n2985 ;
  assign n2993 = ( n2984 & n2991 ) | ( n2984 & ~n2992 ) | ( n2991 & ~n2992 ) ;
  assign n2994 = x24 & x53 ;
  assign n2995 = n2560 | n2581 ;
  assign n2996 = n2994 & ~n2995 ;
  assign n2997 = n2129 & n2130 ;
  assign n2998 = n2093 & n2997 ;
  assign n2999 = ( n2556 & n2997 ) | ( n2556 & n2998 ) | ( n2997 & n2998 ) ;
  assign n3000 = ( n2996 & n2997 ) | ( n2996 & ~n2999 ) | ( n2997 & ~n2999 ) ;
  assign n3001 = x106 & n2982 ;
  assign n3002 = ~x841 & n3001 ;
  assign n3003 = x54 & ~n1332 ;
  assign n3004 = x24 & n3003 ;
  assign n3005 = n3002 | n3004 ;
  assign n3006 = x45 & ~n2819 ;
  assign n3007 = n1412 & n3006 ;
  assign n3008 = x24 & ~x92 ;
  assign n3009 = ~n2576 & n3008 ;
  assign n3010 = x55 | x59 ;
  assign n3011 = ~n1332 & n3010 ;
  assign n3012 = n3009 & n3011 ;
  assign n3013 = n3007 | n3012 ;
  assign n3014 = x56 & x841 ;
  assign n3015 = ~x24 & x55 ;
  assign n3016 = n3014 | n3015 ;
  assign n3017 = ~n1337 & n3016 ;
  assign n3018 = x62 & ~x924 ;
  assign n3019 = ( x56 & ~x841 ) | ( x56 & n3018 ) | ( ~x841 & n3018 ) ;
  assign n3020 = ~n1217 & n3019 ;
  assign n3021 = x24 & x57 ;
  assign n3022 = ( x59 & n1340 ) | ( x59 & n3021 ) | ( n1340 & n3021 ) ;
  assign n3023 = n3021 & ~n3022 ;
  assign n3024 = ( ~n1215 & n3020 ) | ( ~n1215 & n3023 ) | ( n3020 & n3023 ) ;
  assign n3025 = ~n1282 & n3024 ;
  assign n3026 = ~n2464 & n2594 ;
  assign n3027 = ~n1267 & n3026 ;
  assign n3028 = x62 & ~x841 ;
  assign n3029 = ~x59 & x924 ;
  assign n3030 = n3028 & n3029 ;
  assign n3031 = x24 & ~x62 ;
  assign n3032 = x59 & n3031 ;
  assign n3033 = x55 | x56 ;
  assign n3034 = x57 | n3033 ;
  assign n3035 = ( n3030 & n3032 ) | ( n3030 & ~n3034 ) | ( n3032 & ~n3034 ) ;
  assign n3036 = ~n1215 & n3035 ;
  assign n3037 = ~n1282 & n3036 ;
  assign n3038 = ~n1989 & n2131 ;
  assign n3039 = ~n1337 & n3038 ;
  assign n3040 = x60 & ~n2995 ;
  assign n3041 = ~x24 & n3040 ;
  assign n3042 = ( n3039 & n3040 ) | ( n3039 & ~n3041 ) | ( n3040 & ~n3041 ) ;
  assign n3043 = ( n1487 & n2819 ) | ( n1487 & n2949 ) | ( n2819 & n2949 ) ;
  assign n3044 = ( ~n2819 & n3041 ) | ( ~n2819 & n3043 ) | ( n3041 & n3043 ) ;
  assign n3045 = ~x24 & x57 ;
  assign n3046 = ( x62 & ~n3028 ) | ( x62 & n3045 ) | ( ~n3028 & n3045 ) ;
  assign n3047 = ~n1333 & n3046 ;
  assign n3048 = ~n1254 & n1483 ;
  assign n3049 = ( x24 & n2560 ) | ( x24 & n3048 ) | ( n2560 & n3048 ) ;
  assign n3050 = x63 & x999 ;
  assign n3051 = ~n2561 & n3050 ;
  assign n3052 = ( n3048 & ~n3049 ) | ( n3048 & n3051 ) | ( ~n3049 & n3051 ) ;
  assign n3053 = x64 & x841 ;
  assign n3054 = ~x64 & x107 ;
  assign n3055 = ( ~n2561 & n3053 ) | ( ~n2561 & n3054 ) | ( n3053 & n3054 ) ;
  assign n3056 = ~n1337 & n2837 ;
  assign n3057 = ~x102 & x314 ;
  assign n3058 = ( n1261 & n2831 ) | ( n1261 & n3057 ) | ( n2831 & n3057 ) ;
  assign n3059 = n3057 & ~n3058 ;
  assign n3060 = x199 & ~n1553 ;
  assign n3061 = x219 & n1553 ;
  assign n3062 = n3060 | n3061 ;
  assign n3063 = n2516 & n3062 ;
  assign n3064 = n3059 & n3063 ;
  assign n3065 = x81 | n1404 ;
  assign n3066 = ( ~n1408 & n3059 ) | ( ~n1408 & n3065 ) | ( n3059 & n3065 ) ;
  assign n3067 = ~n3065 & n3066 ;
  assign n3068 = x83 & n3067 ;
  assign n3069 = ( n1607 & n1608 ) | ( n1607 & ~n2660 ) | ( n1608 & ~n2660 ) ;
  assign n3070 = ( n2015 & n2618 ) | ( n2015 & ~n3069 ) | ( n2618 & ~n3069 ) ;
  assign n3071 = n3069 & n3070 ;
  assign n3072 = x69 & ~x314 ;
  assign n3073 = ( x71 & ~n2560 ) | ( x71 & n3072 ) | ( ~n2560 & n3072 ) ;
  assign n3074 = ~n1409 & n3073 ;
  assign n3075 = x39 & x287 ;
  assign n3076 = x299 | n1775 ;
  assign n3077 = x1093 & ~n1978 ;
  assign n3078 = ( n1563 & ~n3076 ) | ( n1563 & n3077 ) | ( ~n3076 & n3077 ) ;
  assign n3079 = n2015 & n3078 ;
  assign n3080 = ( x589 & n2025 ) | ( x589 & n2026 ) | ( n2025 & n2026 ) ;
  assign n3081 = n3079 & n3080 ;
  assign n3082 = x593 & ~n3075 ;
  assign n3083 = ( n3075 & n3081 ) | ( n3075 & ~n3082 ) | ( n3081 & ~n3082 ) ;
  assign n3084 = ~n1266 & n2586 ;
  assign n3085 = ~x24 & n3084 ;
  assign n3086 = ( n3083 & n3084 ) | ( n3083 & ~n3085 ) | ( n3084 & ~n3085 ) ;
  assign n3087 = n2618 & n3086 ;
  assign n3088 = x85 & n3067 ;
  assign n3089 = x211 & n1553 ;
  assign n3090 = x200 & ~n1553 ;
  assign n3091 = n3089 | n3090 ;
  assign n3092 = ~n3062 & n3091 ;
  assign n3093 = ~n1254 & n3092 ;
  assign n3094 = ( n3059 & n3088 ) | ( n3059 & n3093 ) | ( n3088 & n3093 ) ;
  assign n3095 = n2063 & n3094 ;
  assign n3096 = x88 & x1093 ;
  assign n3097 = n2658 & n3096 ;
  assign n3098 = x1093 & n2046 ;
  assign n3099 = n2015 & n3098 ;
  assign n3100 = x24 | n3099 ;
  assign n3101 = ( n2052 & n3099 ) | ( n2052 & n3100 ) | ( n3099 & n3100 ) ;
  assign n3102 = n3097 | n3101 ;
  assign n3103 = n2573 & n3102 ;
  assign n3104 = ~x314 & x1050 ;
  assign n3105 = x39 | n3104 ;
  assign n3106 = n2619 & n3105 ;
  assign n3107 = x479 | x841 ;
  assign n3108 = n1790 & ~n3107 ;
  assign n3109 = x74 | n1434 ;
  assign n3110 = ( n2962 & n2963 ) | ( n2962 & n3109 ) | ( n2963 & n3109 ) ;
  assign n3111 = ( x479 & n2025 ) | ( x479 & n2026 ) | ( n2025 & n2026 ) ;
  assign n3112 = n1960 | n3111 ;
  assign n3113 = ( ~n2462 & n2510 ) | ( ~n2462 & n3112 ) | ( n2510 & n3112 ) ;
  assign n3114 = n3112 & n3113 ;
  assign n3115 = x24 & n1310 ;
  assign n3116 = ~n1316 & n3115 ;
  assign n3117 = ( n3113 & ~n3114 ) | ( n3113 & n3116 ) | ( ~n3114 & n3116 ) ;
  assign n3118 = ~n3110 & n3117 ;
  assign n3119 = ( n3108 & ~n3110 ) | ( n3108 & n3118 ) | ( ~n3110 & n3118 ) ;
  assign n3120 = ~x74 & n3116 ;
  assign n3121 = n2512 | n3120 ;
  assign n3122 = ~n1940 & n3121 ;
  assign n3123 = ~n2487 & n2881 ;
  assign n3124 = ( ~n2559 & n2972 ) | ( ~n2559 & n3123 ) | ( n2972 & n3123 ) ;
  assign n3125 = ( n2535 & n2536 ) | ( n2535 & ~n2810 ) | ( n2536 & ~n2810 ) ;
  assign n3126 = n2563 & n3125 ;
  assign n3127 = ( ~n2972 & n3124 ) | ( ~n2972 & n3126 ) | ( n3124 & n3126 ) ;
  assign n3128 = ( x86 & ~x314 ) | ( x86 & n1257 ) | ( ~x314 & n1257 ) ;
  assign n3129 = ~n2995 & n3128 ;
  assign n3130 = x119 & x232 ;
  assign n3131 = ~x468 & n3130 ;
  assign n3132 = x163 & n2742 ;
  assign n3133 = x163 | n2742 ;
  assign n3134 = ~n3132 & n3133 ;
  assign n3135 = n2631 & n3134 ;
  assign n3136 = x40 | n2455 ;
  assign n3137 = x147 & n2072 ;
  assign n3138 = n2455 & ~n3137 ;
  assign n3139 = ( n1320 & n3136 ) | ( n1320 & ~n3138 ) | ( n3136 & ~n3138 ) ;
  assign n3140 = ~n3135 & n3139 ;
  assign n3141 = n1207 & ~n3140 ;
  assign n3142 = ( n1282 & ~n1323 ) | ( n1282 & n1875 ) | ( ~n1323 & n1875 ) ;
  assign n3143 = n1323 | n3142 ;
  assign n3144 = x55 & n3143 ;
  assign n3145 = x163 & n2072 ;
  assign n3146 = ( x55 & n3144 ) | ( x55 & ~n3145 ) | ( n3144 & ~n3145 ) ;
  assign n3147 = ( ~n3140 & n3141 ) | ( ~n3140 & n3146 ) | ( n3141 & n3146 ) ;
  assign n3148 = x156 & x299 ;
  assign n3149 = x179 & ~x299 ;
  assign n3150 = n3148 | n3149 ;
  assign n3151 = n1876 & n2072 ;
  assign n3152 = ~n3150 & n3151 ;
  assign n3153 = ( ~n1282 & n3151 ) | ( ~n1282 & n3152 ) | ( n3151 & n3152 ) ;
  assign n3154 = ( x40 & ~n3152 ) | ( x40 & n3153 ) | ( ~n3152 & n3153 ) ;
  assign n3155 = ~n1326 & n3154 ;
  assign n3156 = n1320 | n3155 ;
  assign n3157 = x187 & n2079 ;
  assign n3158 = ~n2079 & n3137 ;
  assign n3159 = ( n2643 & n3157 ) | ( n2643 & n3158 ) | ( n3157 & n3158 ) ;
  assign n3160 = n3156 | n3159 ;
  assign n3161 = ~n2479 & n2661 ;
  assign n3162 = n1435 & n3150 ;
  assign n3163 = ( ~n2049 & n3161 ) | ( ~n2049 & n3162 ) | ( n3161 & n3162 ) ;
  assign n3164 = n2657 & n3163 ;
  assign n3165 = x175 & n2594 ;
  assign n3166 = ~n1215 & n2079 ;
  assign n3167 = x182 & n2683 ;
  assign n3168 = n3166 & n3167 ;
  assign n3169 = ( n3165 & n3166 ) | ( n3165 & n3168 ) | ( n3166 & n3168 ) ;
  assign n3170 = n3164 | n3169 ;
  assign n3171 = ~n1208 & n2156 ;
  assign n3172 = ( n1208 & n3170 ) | ( n1208 & ~n3171 ) | ( n3170 & ~n3171 ) ;
  assign n3173 = ( n1208 & ~n1271 ) | ( n1208 & n3172 ) | ( ~n1271 & n3172 ) ;
  assign n3174 = x184 | n2737 ;
  assign n3175 = x299 & n2631 ;
  assign n3176 = n3134 & n3175 ;
  assign n3177 = ( x184 & ~n2637 ) | ( x184 & n2737 ) | ( ~n2637 & n2737 ) ;
  assign n3178 = ( n3174 & n3176 ) | ( n3174 & ~n3177 ) | ( n3176 & ~n3177 ) ;
  assign n3179 = ~n3173 & n3178 ;
  assign n3180 = ( n3160 & n3173 ) | ( n3160 & ~n3179 ) | ( n3173 & ~n3179 ) ;
  assign n3181 = ~n3147 & n3180 ;
  assign n3182 = x184 & ~x299 ;
  assign n3183 = ( n2586 & n2693 ) | ( n2586 & n3182 ) | ( n2693 & n3182 ) ;
  assign n3184 = ~n2479 & n2589 ;
  assign n3185 = n1271 | n1279 ;
  assign n3186 = ~x32 & x153 ;
  assign n3187 = n2594 & n3186 ;
  assign n3188 = x160 | n3187 ;
  assign n3189 = ( n2712 & n3187 ) | ( n2712 & n3188 ) | ( n3187 & n3188 ) ;
  assign n3190 = ~n3185 & n3189 ;
  assign n3191 = x163 & x299 ;
  assign n3192 = ( n2586 & n2679 ) | ( n2586 & n3191 ) | ( n2679 & n3191 ) ;
  assign n3193 = ( x299 & n3190 ) | ( x299 & n3192 ) | ( n3190 & n3192 ) ;
  assign n3194 = ( ~n3183 & n3184 ) | ( ~n3183 & n3193 ) | ( n3184 & n3193 ) ;
  assign n3195 = ( n2676 & n3183 ) | ( n2676 & n3194 ) | ( n3183 & n3194 ) ;
  assign n3196 = ( ~n3147 & n3181 ) | ( ~n3147 & n3195 ) | ( n3181 & n3195 ) ;
  assign n3197 = x954 | n2626 ;
  assign n3198 = x79 & ~n3197 ;
  assign n3199 = ( n2625 & n3197 ) | ( n2625 & ~n3198 ) | ( n3197 & ~n3198 ) ;
  assign n3200 = ( ~x79 & n3197 ) | ( ~x79 & n3198 ) | ( n3197 & n3198 ) ;
  assign n3201 = ( n2621 & n3199 ) | ( n2621 & ~n3200 ) | ( n3199 & ~n3200 ) ;
  assign n3202 = ~n3196 & n3201 ;
  assign n3203 = x80 | n2180 ;
  assign n3204 = n2475 & ~n3203 ;
  assign n3205 = n1485 & ~n2831 ;
  assign n3206 = x81 & ~x314 ;
  assign n3207 = x68 | n3206 ;
  assign n3208 = n3205 & n3207 ;
  assign n3209 = ( x66 & x69 ) | ( x66 & ~n3072 ) | ( x69 & ~n3072 ) ;
  assign n3210 = n2982 & n3209 ;
  assign n3211 = x83 & ~x314 ;
  assign n3212 = x84 | n3211 ;
  assign n3213 = n2982 & n3212 ;
  assign n3214 = n3062 | n3091 ;
  assign n3215 = ( n2516 & n3059 ) | ( n2516 & n3214 ) | ( n3059 & n3214 ) ;
  assign n3216 = ~n3214 & n3215 ;
  assign n3217 = x85 & x314 ;
  assign n3218 = ( x67 & x85 ) | ( x67 & ~n3217 ) | ( x85 & ~n3217 ) ;
  assign n3219 = n2982 & n3218 ;
  assign n3220 = ( n1607 & n1608 ) | ( n1607 & n2018 ) | ( n1608 & n2018 ) ;
  assign n3221 = ~n1337 & n3220 ;
  assign n3222 = x103 & n3067 ;
  assign n3223 = x104 & ~n2470 ;
  assign n3224 = ( x88 & ~n3096 ) | ( x88 & n3223 ) | ( ~n3096 & n3223 ) ;
  assign n3225 = ( n2658 & n2823 ) | ( n2658 & ~n3224 ) | ( n2823 & ~n3224 ) ;
  assign n3226 = n3224 & n3225 ;
  assign n3227 = x24 | n1309 ;
  assign n3228 = n3084 & ~n3227 ;
  assign n3229 = x89 & x841 ;
  assign n3230 = ~n2823 & n3229 ;
  assign n3231 = ( n3228 & n3229 ) | ( n3228 & ~n3230 ) | ( n3229 & ~n3230 ) ;
  assign n3232 = x73 & ~x1050 ;
  assign n3233 = ( x90 & ~n2591 ) | ( x90 & n3232 ) | ( ~n2591 & n3232 ) ;
  assign n3234 = n2573 & n3233 ;
  assign n3235 = ~n1282 & n2497 ;
  assign n3236 = x24 & ~x36 ;
  assign n3237 = n1435 | n3236 ;
  assign n3238 = ( ~n2559 & n3235 ) | ( ~n2559 & n3237 ) | ( n3235 & n3237 ) ;
  assign n3239 = ~x58 & n3238 ;
  assign n3240 = ~n1337 & n3239 ;
  assign n3241 = x39 | n2820 ;
  assign n3242 = x58 & n2820 ;
  assign n3243 = ( n1362 & n3241 ) | ( n1362 & ~n3242 ) | ( n3241 & ~n3242 ) ;
  assign n3244 = n3240 & n3243 ;
  assign n3245 = n2024 & ~n2093 ;
  assign n3246 = n1877 & n3104 ;
  assign n3247 = n3245 | n3246 ;
  assign n3248 = ~n2556 & n3247 ;
  assign n3249 = ~x1050 & n1877 ;
  assign n3250 = ( x93 & ~n1971 ) | ( x93 & n3249 ) | ( ~n1971 & n3249 ) ;
  assign n3251 = ~n1940 & n3250 ;
  assign n3252 = ~n1434 & n2488 ;
  assign n3253 = n2881 & n3252 ;
  assign n3254 = ( x49 & ~n2960 ) | ( x49 & n3253 ) | ( ~n2960 & n3253 ) ;
  assign n3255 = n2823 & n3254 ;
  assign n3256 = x24 & x95 ;
  assign n3257 = ( n1309 & n1350 ) | ( n1309 & n3256 ) | ( n1350 & n3256 ) ;
  assign n3258 = n3256 & ~n3257 ;
  assign n3259 = x841 & ~n3258 ;
  assign n3260 = x89 & ~x332 ;
  assign n3261 = n2823 & n3260 ;
  assign n3262 = ( n3258 & ~n3259 ) | ( n3258 & n3261 ) | ( ~n3259 & n3261 ) ;
  assign n3263 = n3079 & ~n3080 ;
  assign n3264 = n2618 & n3263 ;
  assign n3265 = n3262 | n3264 ;
  assign n3266 = ~x24 & x95 ;
  assign n3267 = ( x841 & ~n1434 ) | ( x841 & n3107 ) | ( ~n1434 & n3107 ) ;
  assign n3268 = x96 & n3267 ;
  assign n3269 = ( ~n1309 & n3266 ) | ( ~n1309 & n3268 ) | ( n3266 & n3268 ) ;
  assign n3270 = ~n1350 & n3269 ;
  assign n3271 = x97 & ~n1435 ;
  assign n3272 = n3112 & n3271 ;
  assign n3273 = x593 | n3272 ;
  assign n3274 = ( n3081 & n3272 ) | ( n3081 & n3273 ) | ( n3272 & n3273 ) ;
  assign n3275 = n2618 & n3274 ;
  assign n3276 = x92 | n2589 ;
  assign n3277 = x314 & x1050 ;
  assign n3278 = ~n1333 & n3277 ;
  assign n3279 = n3276 & n3278 ;
  assign n3280 = ( ~x72 & x99 ) | ( ~x72 & n2853 ) | ( x99 & n2853 ) ;
  assign n3281 = x152 & x161 ;
  assign n3282 = n2861 & n3281 ;
  assign n3283 = ( x39 & ~n2866 ) | ( x39 & n2869 ) | ( ~n2866 & n2869 ) ;
  assign n3284 = n3280 & ~n3283 ;
  assign n3285 = ( n3280 & n3282 ) | ( n3280 & n3284 ) | ( n3282 & n3284 ) ;
  assign n3286 = n1942 & ~n3285 ;
  assign n3287 = n2891 & ~n3285 ;
  assign n3288 = ( n1942 & ~n2891 ) | ( n1942 & n3285 ) | ( ~n2891 & n3285 ) ;
  assign n3289 = ( ~n3286 & n3287 ) | ( ~n3286 & n3288 ) | ( n3287 & n3288 ) ;
  assign n3290 = ~n1963 & n2546 ;
  assign n3291 = ~n2793 & n3290 ;
  assign n3292 = ( n2541 & ~n2542 ) | ( n2541 & n3291 ) | ( ~n2542 & n3291 ) ;
  assign n3293 = ~n2557 & n3292 ;
  assign n3294 = x287 & n2618 ;
  assign n3295 = x101 & ~n2895 ;
  assign n3296 = n2891 & n3295 ;
  assign n3297 = ~x161 & n2853 ;
  assign n3298 = x152 & n1208 ;
  assign n3299 = ( n2857 & ~n3297 ) | ( n2857 & n3298 ) | ( ~n3297 & n3298 ) ;
  assign n3300 = n3297 & n3299 ;
  assign n3301 = ~n1208 & n2485 ;
  assign n3302 = ( n2483 & ~n2853 ) | ( n2483 & n3301 ) | ( ~n2853 & n3301 ) ;
  assign n3303 = ( n2853 & n3300 ) | ( n2853 & n3302 ) | ( n3300 & n3302 ) ;
  assign n3304 = ( n3294 & ~n3296 ) | ( n3294 & n3303 ) | ( ~n3296 & n3303 ) ;
  assign n3305 = n2891 | n3295 ;
  assign n3306 = ~n3296 & n3305 ;
  assign n3307 = ( ~n3294 & n3304 ) | ( ~n3294 & n3306 ) | ( n3304 & n3306 ) ;
  assign n3308 = x65 & ~n2561 ;
  assign n3309 = n2561 & n2823 ;
  assign n3310 = n2059 & ~n2561 ;
  assign n3311 = ( ~n2149 & n3309 ) | ( ~n2149 & n3310 ) | ( n3309 & n3310 ) ;
  assign n3312 = x104 & n2470 ;
  assign n3313 = n2658 & n3312 ;
  assign n3314 = n2487 & n2658 ;
  assign n3315 = x110 & n3314 ;
  assign n3316 = ( x110 & n3313 ) | ( x110 & ~n3315 ) | ( n3313 & ~n3315 ) ;
  assign n3317 = n2823 & n3316 ;
  assign n3318 = ~x24 & x53 ;
  assign n3319 = ~n2995 & n3318 ;
  assign n3320 = ( n3001 & ~n3002 ) | ( n3001 & n3319 ) | ( ~n3002 & n3319 ) ;
  assign n3321 = x63 & ~x999 ;
  assign n3322 = ~n2561 & n3321 ;
  assign n3323 = x51 | x98 ;
  assign n3324 = x100 & ~x108 ;
  assign n3325 = ( ~x108 & n1282 ) | ( ~x108 & n3324 ) | ( n1282 & n3324 ) ;
  assign n3326 = n1209 & ~n3323 ;
  assign n3327 = ( ~n3323 & n3325 ) | ( ~n3323 & n3326 ) | ( n3325 & n3326 ) ;
  assign n3328 = n2573 & ~n2843 ;
  assign n3329 = ~n3327 & n3328 ;
  assign n3330 = x77 & x314 ;
  assign n3331 = ~n2995 & n3330 ;
  assign n3332 = x111 & ~x314 ;
  assign n3333 = ( x111 & n3315 ) | ( x111 & ~n3332 ) | ( n3315 & ~n3332 ) ;
  assign n3334 = n2823 & n3333 ;
  assign n3335 = n2823 & n3332 ;
  assign n3336 = n2052 | n3227 ;
  assign n3337 = ( ~n3227 & n3335 ) | ( ~n3227 & n3336 ) | ( n3335 & n3336 ) ;
  assign n3338 = x124 & ~x468 ;
  assign n3339 = x113 & ~n2895 ;
  assign n3340 = n2891 & ~n3339 ;
  assign n3341 = n1943 & ~n3339 ;
  assign n3342 = ( n1943 & ~n2891 ) | ( n1943 & n3339 ) | ( ~n2891 & n3339 ) ;
  assign n3343 = ( n3340 & ~n3341 ) | ( n3340 & n3342 ) | ( ~n3341 & n3342 ) ;
  assign n3344 = x114 & n2897 ;
  assign n3345 = x114 & ~n2895 ;
  assign n3346 = ( n2898 & ~n3344 ) | ( n2898 & n3345 ) | ( ~n3344 & n3345 ) ;
  assign n3347 = ~n1945 & n2891 ;
  assign n3348 = ( x115 & n2895 ) | ( x115 & n3347 ) | ( n2895 & n3347 ) ;
  assign n3349 = ( x115 & n2897 ) | ( x115 & ~n3348 ) | ( n2897 & ~n3348 ) ;
  assign n3350 = x116 & ~n2895 ;
  assign n3351 = n1944 & ~n3350 ;
  assign n3352 = n2891 & ~n3350 ;
  assign n3353 = ( n1944 & ~n2891 ) | ( n1944 & n3350 ) | ( ~n2891 & n3350 ) ;
  assign n3354 = ( ~n3351 & n3352 ) | ( ~n3351 & n3353 ) | ( n3352 & n3353 ) ;
  assign n3355 = x79 | n3197 ;
  assign n3356 = x118 & ~n3355 ;
  assign n3357 = ( x118 & n2625 ) | ( x118 & ~n3355 ) | ( n2625 & ~n3355 ) ;
  assign n3358 = ( n2161 & ~n3356 ) | ( n2161 & n3357 ) | ( ~n3356 & n3357 ) ;
  assign n3359 = ~n2456 & n2578 ;
  assign n3360 = ( n2456 & n3358 ) | ( n2456 & ~n3359 ) | ( n3358 & ~n3359 ) ;
  assign n3361 = n1333 & ~n3360 ;
  assign n3362 = n2762 | n2803 ;
  assign n3363 = ( n2586 & n2597 ) | ( n2586 & ~n3362 ) | ( n2597 & ~n3362 ) ;
  assign n3364 = n3362 | n3363 ;
  assign n3365 = ( n3360 & ~n3361 ) | ( n3360 & n3364 ) | ( ~n3361 & n3364 ) ;
  assign n3366 = x150 & n3133 ;
  assign n3367 = ( x150 & n2631 ) | ( x150 & n3133 ) | ( n2631 & n3133 ) ;
  assign n3368 = x165 & n2072 ;
  assign n3369 = n2455 & n3368 ;
  assign n3370 = n1208 & n1320 ;
  assign n3371 = ( n1208 & n3369 ) | ( n1208 & n3370 ) | ( n3369 & n3370 ) ;
  assign n3372 = ( n3366 & ~n3367 ) | ( n3366 & n3371 ) | ( ~n3367 & n3371 ) ;
  assign n3373 = ~n1320 & n1326 ;
  assign n3374 = x165 & n2073 ;
  assign n3375 = x143 & n2079 ;
  assign n3376 = ( n3373 & n3374 ) | ( n3373 & n3375 ) | ( n3374 & n3375 ) ;
  assign n3377 = ( x55 & n3373 ) | ( x55 & ~n3376 ) | ( n3373 & ~n3376 ) ;
  assign n3378 = ( x150 & n3133 ) | ( x150 & n3175 ) | ( n3133 & n3175 ) ;
  assign n3379 = ( ~n3366 & n3377 ) | ( ~n3366 & n3378 ) | ( n3377 & n3378 ) ;
  assign n3380 = n1215 & n3379 ;
  assign n3381 = ( n1282 & n3379 ) | ( n1282 & n3380 ) | ( n3379 & n3380 ) ;
  assign n3382 = x185 & n3174 ;
  assign n3383 = ( x185 & n2637 ) | ( x185 & n3174 ) | ( n2637 & n3174 ) ;
  assign n3384 = ( n1207 & ~n3382 ) | ( n1207 & n3383 ) | ( ~n3382 & n3383 ) ;
  assign n3385 = x92 & ~n1875 ;
  assign n3386 = x178 & ~x299 ;
  assign n3387 = x157 & x299 ;
  assign n3388 = ( ~n1321 & n3386 ) | ( ~n1321 & n3387 ) | ( n3386 & n3387 ) ;
  assign n3389 = ( ~n2072 & n2159 ) | ( ~n2072 & n3388 ) | ( n2159 & n3388 ) ;
  assign n3390 = n3388 & ~n3389 ;
  assign n3391 = n3385 & ~n3390 ;
  assign n3392 = ( ~n3381 & n3384 ) | ( ~n3381 & n3391 ) | ( n3384 & n3391 ) ;
  assign n3393 = n3381 | n3392 ;
  assign n3394 = ( n1435 & n3386 ) | ( n1435 & n3387 ) | ( n3386 & n3387 ) ;
  assign n3395 = x168 & x299 ;
  assign n3396 = x190 & ~x299 ;
  assign n3397 = ( n2661 & n3395 ) | ( n2661 & n3396 ) | ( n3395 & n3396 ) ;
  assign n3398 = n3394 | n3397 ;
  assign n3399 = ( n2656 & n2761 ) | ( n2656 & ~n3398 ) | ( n2761 & ~n3398 ) ;
  assign n3400 = x55 & x150 ;
  assign n3401 = ~n2072 & n3400 ;
  assign n3402 = ( n2092 & n3400 ) | ( n2092 & ~n3401 ) | ( n3400 & ~n3401 ) ;
  assign n3403 = ~n3398 & n3399 ;
  assign n3404 = ( n3399 & n3402 ) | ( n3399 & ~n3403 ) | ( n3402 & ~n3403 ) ;
  assign n3405 = n2642 | n3404 ;
  assign n3406 = ~n3393 & n3405 ;
  assign n3407 = ( n3365 & n3372 ) | ( n3365 & n3406 ) | ( n3372 & n3406 ) ;
  assign n3408 = n3365 & ~n3407 ;
  assign n3409 = ( x150 & n2586 ) | ( x150 & n2679 ) | ( n2586 & n2679 ) ;
  assign n3410 = n2597 | n3409 ;
  assign n3411 = x73 & ~x168 ;
  assign n3412 = ~x151 & n1273 ;
  assign n3413 = ( n2073 & n3411 ) | ( n2073 & n3412 ) | ( n3411 & n3412 ) ;
  assign n3414 = n2073 & ~n3413 ;
  assign n3415 = n2712 | n3414 ;
  assign n3416 = ( n2712 & n3410 ) | ( n2712 & n3415 ) | ( n3410 & n3415 ) ;
  assign n3417 = x173 & n1273 ;
  assign n3418 = x73 & x190 ;
  assign n3419 = ~x73 & x185 ;
  assign n3420 = ( ~n1273 & n3418 ) | ( ~n1273 & n3419 ) | ( n3418 & n3419 ) ;
  assign n3421 = ( n2079 & n3417 ) | ( n2079 & n3420 ) | ( n3417 & n3420 ) ;
  assign n3422 = ( n2586 & ~n2597 ) | ( n2586 & n2693 ) | ( ~n2597 & n2693 ) ;
  assign n3423 = ( n2597 & n3421 ) | ( n2597 & n3422 ) | ( n3421 & n3422 ) ;
  assign n3424 = ~n3416 & n3423 ;
  assign n3425 = ( ~n1309 & n3416 ) | ( ~n1309 & n3424 ) | ( n3416 & n3424 ) ;
  assign n3426 = n3408 & ~n3425 ;
  assign n3427 = ~x128 & x228 ;
  assign n3428 = x128 & x228 ;
  assign n3429 = x92 | n1319 ;
  assign n3430 = n1978 & ~n3429 ;
  assign n3431 = ~n1563 & n3076 ;
  assign n3432 = n2018 & n3431 ;
  assign n3433 = ( n3429 & ~n3430 ) | ( n3429 & n3432 ) | ( ~n3430 & n3432 ) ;
  assign n3434 = x91 | x93 ;
  assign n3435 = ( n1257 & n2082 ) | ( n1257 & ~n3434 ) | ( n2082 & ~n3434 ) ;
  assign n3436 = n3434 | n3435 ;
  assign n3437 = x36 | x97 ;
  assign n3438 = n1435 & n3437 ;
  assign n3439 = ( ~n3433 & n3436 ) | ( ~n3433 & n3438 ) | ( n3436 & n3438 ) ;
  assign n3440 = n3433 | n3439 ;
  assign n3441 = ( n1415 & n3433 ) | ( n1415 & n3440 ) | ( n3433 & n3440 ) ;
  assign n3442 = ~n1337 & n3441 ;
  assign n3443 = ( ~n3427 & n3428 ) | ( ~n3427 & n3442 ) | ( n3428 & n3442 ) ;
  assign n3444 = x951 & x982 ;
  assign n3445 = ( ~n1430 & n2180 ) | ( ~n1430 & n3444 ) | ( n2180 & n3444 ) ;
  assign n3446 = n3444 & ~n3445 ;
  assign n3447 = x31 | x80 ;
  assign n3448 = x818 & ~n3447 ;
  assign n3449 = ( x1093 & n3446 ) | ( x1093 & n3448 ) | ( n3446 & n3448 ) ;
  assign n3450 = x120 | n3449 ;
  assign n3451 = ~n2529 & n3450 ;
  assign n3452 = ( ~x161 & n1208 ) | ( ~x161 & n2480 ) | ( n1208 & n2480 ) ;
  assign n3453 = ~x51 & n2758 ;
  assign n3454 = n1208 | n2481 ;
  assign n3455 = ( n3452 & n3453 ) | ( n3452 & ~n3454 ) | ( n3453 & ~n3454 ) ;
  assign n3456 = ~x146 & n1553 ;
  assign n3457 = x142 | n1553 ;
  assign n3458 = ( x51 & n3456 ) | ( x51 & ~n3457 ) | ( n3456 & ~n3457 ) ;
  assign n3459 = ( ~x87 & n3455 ) | ( ~x87 & n3458 ) | ( n3455 & n3458 ) ;
  assign n3460 = ~n1208 & n3182 ;
  assign n3461 = ( x163 & n1208 ) | ( x163 & n3191 ) | ( n1208 & n3191 ) ;
  assign n3462 = ( x87 & n3460 ) | ( x87 & n3461 ) | ( n3460 & n3461 ) ;
  assign n3463 = n3459 | n3462 ;
  assign n3464 = ~x24 & x77 ;
  assign n3465 = x314 & n3464 ;
  assign n3466 = ( n2684 & n2685 ) | ( n2684 & n3465 ) | ( n2685 & n3465 ) ;
  assign n3467 = ( x77 & x86 ) | ( x77 & ~n3464 ) | ( x86 & ~n3464 ) ;
  assign n3468 = n3150 & n3467 ;
  assign n3469 = ( n3463 & ~n3466 ) | ( n3463 & n3468 ) | ( ~n3466 & n3468 ) ;
  assign n3470 = n3466 | n3469 ;
  assign n3471 = ( ~n2995 & n3463 ) | ( ~n2995 & n3470 ) | ( n3463 & n3470 ) ;
  assign n3472 = x159 & x299 ;
  assign n3473 = x181 & ~x299 ;
  assign n3474 = n3472 | n3473 ;
  assign n3475 = ( n2020 & n2022 ) | ( n2020 & n3474 ) | ( n2022 & n3474 ) ;
  assign n3476 = n3471 | n3475 ;
  assign n3477 = ( n2947 & n3471 ) | ( n2947 & n3476 ) | ( n3471 & n3476 ) ;
  assign n3478 = n2072 & n3477 ;
  assign n3479 = n1209 | n2092 ;
  assign n3480 = n3330 | n3467 ;
  assign n3481 = ~n2604 & n3480 ;
  assign n3482 = ( n2582 & n3479 ) | ( n2582 & n3481 ) | ( n3479 & n3481 ) ;
  assign n3483 = n3481 & ~n3482 ;
  assign n3484 = ( n2052 & ~n3479 ) | ( n2052 & n3483 ) | ( ~n3479 & n3483 ) ;
  assign n3485 = ~n1208 & n3484 ;
  assign n3486 = ~n2458 & n2609 ;
  assign n3487 = n3485 | n3486 ;
  assign n3488 = x125 | x133 ;
  assign n3489 = ~x121 & n3488 ;
  assign n3490 = x121 | n3488 ;
  assign n3491 = x126 | n3490 ;
  assign n3492 = x132 | n3491 ;
  assign n3493 = x130 | n3492 ;
  assign n3494 = x136 | n3493 ;
  assign n3495 = x135 | n3494 ;
  assign n3496 = x134 | n3495 ;
  assign n3497 = ( ~x121 & n3488 ) | ( ~x121 & n3496 ) | ( n3488 & n3496 ) ;
  assign n3498 = ( n2760 & ~n3489 ) | ( n2760 & n3497 ) | ( ~n3489 & n3497 ) ;
  assign n3499 = ~n3487 & n3498 ;
  assign n3500 = ( ~n3478 & n3487 ) | ( ~n3478 & n3499 ) | ( n3487 & n3499 ) ;
  assign n3501 = x82 & ~x111 ;
  assign n3502 = x90 | n2063 ;
  assign n3503 = ( x111 & ~n3501 ) | ( x111 & n3502 ) | ( ~n3501 & n3502 ) ;
  assign n3504 = ~n1215 & n3503 ;
  assign n3505 = ( ~n1215 & n2052 ) | ( ~n1215 & n3504 ) | ( n2052 & n3504 ) ;
  assign n3506 = n1415 & n3505 ;
  assign n3507 = ~x39 & x110 ;
  assign n3508 = ~n2942 & n3507 ;
  assign n3509 = n1950 & n3508 ;
  assign n3510 = n1982 | n2010 ;
  assign n3511 = ( n1993 & n2613 ) | ( n1993 & ~n3510 ) | ( n2613 & ~n3510 ) ;
  assign n3512 = n1289 & n2040 ;
  assign n3513 = ( n1993 & n3511 ) | ( n1993 & ~n3512 ) | ( n3511 & ~n3512 ) ;
  assign n3514 = n1993 & ~n3513 ;
  assign n3515 = ( n2658 & n3509 ) | ( n2658 & n3514 ) | ( n3509 & n3514 ) ;
  assign n3516 = n1208 & ~n3515 ;
  assign n3517 = n1208 | n3507 ;
  assign n3518 = ( n1208 & n3314 ) | ( n1208 & n3517 ) | ( n3314 & n3517 ) ;
  assign n3519 = ~n1208 & n2615 ;
  assign n3520 = ( ~n3506 & n3518 ) | ( ~n3506 & n3519 ) | ( n3518 & n3519 ) ;
  assign n3521 = ( n3506 & ~n3516 ) | ( n3506 & n3520 ) | ( ~n3516 & n3520 ) ;
  assign n3522 = ~x162 & n1553 ;
  assign n3523 = x140 | n1553 ;
  assign n3524 = ( x87 & n3522 ) | ( x87 & ~n3523 ) | ( n3522 & ~n3523 ) ;
  assign n3525 = x87 & n2072 ;
  assign n3526 = ( n3298 & ~n3301 ) | ( n3298 & n3453 ) | ( ~n3301 & n3453 ) ;
  assign n3527 = ~n1208 & n2688 ;
  assign n3528 = ( x172 & n1208 ) | ( x172 & n2689 ) | ( n1208 & n2689 ) ;
  assign n3529 = ( x51 & n3527 ) | ( x51 & n3528 ) | ( n3527 & n3528 ) ;
  assign n3530 = ( ~n3298 & n3526 ) | ( ~n3298 & n3529 ) | ( n3526 & n3529 ) ;
  assign n3531 = ( n2072 & n3525 ) | ( n2072 & n3530 ) | ( n3525 & n3530 ) ;
  assign n3532 = ~n3524 & n3531 ;
  assign n3533 = n2760 & ~n3532 ;
  assign n3534 = ~x287 & n2072 ;
  assign n3535 = ( n2684 & n2685 ) | ( n2684 & n3534 ) | ( n2685 & n3534 ) ;
  assign n3536 = n2600 | n3535 ;
  assign n3537 = n3486 & n3536 ;
  assign n3538 = ~x125 & x133 ;
  assign n3539 = ~n2600 & n3486 ;
  assign n3540 = n1372 | n2607 ;
  assign n3541 = n3481 & ~n3540 ;
  assign n3542 = ~n1309 & n3541 ;
  assign n3543 = n3539 | n3542 ;
  assign n3544 = ( ~x125 & x133 ) | ( ~x125 & n3496 ) | ( x133 & n3496 ) ;
  assign n3545 = ( ~n3538 & n3543 ) | ( ~n3538 & n3544 ) | ( n3543 & n3544 ) ;
  assign n3546 = ~n3537 & n3545 ;
  assign n3547 = x197 & x299 ;
  assign n3548 = x145 & ~x299 ;
  assign n3549 = ( n2072 & n3547 ) | ( n2072 & n3548 ) | ( n3547 & n3548 ) ;
  assign n3550 = n3464 & ~n3549 ;
  assign n3551 = n2765 | n3464 ;
  assign n3552 = ( n2052 & ~n3550 ) | ( n2052 & n3551 ) | ( ~n3550 & n3551 ) ;
  assign n3553 = n3546 & ~n3552 ;
  assign n3554 = ( ~n3485 & n3546 ) | ( ~n3485 & n3553 ) | ( n3546 & n3553 ) ;
  assign n3555 = ( ~n3532 & n3533 ) | ( ~n3532 & n3554 ) | ( n3533 & n3554 ) ;
  assign n3556 = ~n2072 & n2760 ;
  assign n3557 = ( x39 & n1282 ) | ( x39 & ~n2023 ) | ( n1282 & ~n2023 ) ;
  assign n3558 = ( ~x287 & n2074 ) | ( ~x287 & n2080 ) | ( n2074 & n2080 ) ;
  assign n3559 = ( x39 & n3557 ) | ( x39 & n3558 ) | ( n3557 & n3558 ) ;
  assign n3560 = x39 & ~n3559 ;
  assign n3561 = ( x126 & ~n3490 ) | ( x126 & n3496 ) | ( ~n3490 & n3496 ) ;
  assign n3562 = x51 | n2758 ;
  assign n3563 = ( x126 & ~n3490 ) | ( x126 & n3562 ) | ( ~n3490 & n3562 ) ;
  assign n3564 = n3561 & ~n3563 ;
  assign n3565 = ~n3541 & n3564 ;
  assign n3566 = ~n2072 & n3541 ;
  assign n3567 = ( ~n2052 & n3565 ) | ( ~n2052 & n3566 ) | ( n3565 & n3566 ) ;
  assign n3568 = n3386 | n3387 ;
  assign n3569 = n3467 & ~n3568 ;
  assign n3570 = n3465 & ~n3474 ;
  assign n3571 = ( ~n2462 & n3569 ) | ( ~n2462 & n3570 ) | ( n3569 & n3570 ) ;
  assign n3572 = ( x39 & n2582 ) | ( x39 & n3571 ) | ( n2582 & n3571 ) ;
  assign n3573 = n3571 & ~n3572 ;
  assign n3574 = ( ~x39 & n3567 ) | ( ~x39 & n3573 ) | ( n3567 & n3573 ) ;
  assign n3575 = ( ~n2458 & n3560 ) | ( ~n2458 & n3574 ) | ( n3560 & n3574 ) ;
  assign n3576 = n2459 & n3564 ;
  assign n3577 = ~n1208 & n2478 ;
  assign n3578 = ( x166 & n1208 ) | ( x166 & n2477 ) | ( n1208 & n2477 ) ;
  assign n3579 = ( n3453 & n3577 ) | ( n3453 & n3578 ) | ( n3577 & n3578 ) ;
  assign n3580 = x87 | n3579 ;
  assign n3581 = ~x153 & n1553 ;
  assign n3582 = x175 | n1553 ;
  assign n3583 = ( x51 & n3581 ) | ( x51 & ~n3582 ) | ( n3581 & ~n3582 ) ;
  assign n3584 = n3580 | n3583 ;
  assign n3585 = n3486 & ~n3584 ;
  assign n3586 = ( n3576 & n3584 ) | ( n3576 & ~n3585 ) | ( n3584 & ~n3585 ) ;
  assign n3587 = n3575 | n3586 ;
  assign n3588 = x185 & ~n1553 ;
  assign n3589 = x150 & n1553 ;
  assign n3590 = ( x87 & n3588 ) | ( x87 & n3589 ) | ( n3588 & n3589 ) ;
  assign n3591 = ~n3556 & n3590 ;
  assign n3592 = ( n3556 & n3587 ) | ( n3556 & ~n3591 ) | ( n3587 & ~n3591 ) ;
  assign n3593 = ~x63 & x129 ;
  assign n3594 = x250 & n2488 ;
  assign n3595 = n1960 & n3594 ;
  assign n3596 = x127 | n3594 ;
  assign n3597 = ( x94 & n3595 ) | ( x94 & ~n3596 ) | ( n3595 & ~n3596 ) ;
  assign n3598 = n3593 & ~n3597 ;
  assign n3599 = n1309 | n1364 ;
  assign n3600 = ~n1940 & n3599 ;
  assign n3601 = n1488 & ~n1940 ;
  assign n3602 = n3600 | n3601 ;
  assign n3603 = n3598 & n3602 ;
  assign n3604 = n2487 & n2882 ;
  assign n3605 = n1960 & n3604 ;
  assign n3606 = x129 | n3604 ;
  assign n3607 = ( x75 & n3605 ) | ( x75 & ~n3606 ) | ( n3605 & ~n3606 ) ;
  assign n3608 = x100 & n1961 ;
  assign n3609 = ( n2141 & n3600 ) | ( n2141 & ~n3608 ) | ( n3600 & ~n3608 ) ;
  assign n3610 = ~n3607 & n3609 ;
  assign n3611 = ( ~n1208 & n2746 ) | ( ~n1208 & n2748 ) | ( n2746 & n2748 ) ;
  assign n3612 = ( n2072 & n2778 ) | ( n2072 & n3611 ) | ( n2778 & n3611 ) ;
  assign n3613 = x87 & ~n3612 ;
  assign n3614 = ( x169 & n1208 ) | ( x169 & n2645 ) | ( n1208 & n2645 ) ;
  assign n3615 = ~n1208 & n2644 ;
  assign n3616 = n2072 & n2758 ;
  assign n3617 = ( n3614 & n3615 ) | ( n3614 & n3616 ) | ( n3615 & n3616 ) ;
  assign n3618 = n2759 | n3617 ;
  assign n3619 = ~x130 & n3492 ;
  assign n3620 = ~n3487 & n3496 ;
  assign n3621 = ( ~x130 & n3492 ) | ( ~x130 & n3620 ) | ( n3492 & n3620 ) ;
  assign n3622 = x162 & x299 ;
  assign n3623 = x140 & ~x299 ;
  assign n3624 = ( ~n2758 & n3622 ) | ( ~n2758 & n3623 ) | ( n3622 & n3623 ) ;
  assign n3625 = n3534 & n3624 ;
  assign n3626 = ( n2758 & n3539 ) | ( n2758 & ~n3625 ) | ( n3539 & ~n3625 ) ;
  assign n3627 = ( ~n3619 & n3621 ) | ( ~n3619 & n3626 ) | ( n3621 & n3626 ) ;
  assign n3628 = ~n3618 & n3627 ;
  assign n3629 = n3613 | n3628 ;
  assign n3630 = ( x164 & n1208 ) | ( x164 & n2669 ) | ( n1208 & n2669 ) ;
  assign n3631 = ~n1208 & n2670 ;
  assign n3632 = ( n3525 & n3630 ) | ( n3525 & n3631 ) | ( n3630 & n3631 ) ;
  assign n3633 = x51 & x151 ;
  assign n3634 = x168 | n3633 ;
  assign n3635 = ( n3453 & n3633 ) | ( n3453 & n3634 ) | ( n3633 & n3634 ) ;
  assign n3636 = ~x132 & n3491 ;
  assign n3637 = ( ~x132 & n3491 ) | ( ~x132 & n3496 ) | ( n3491 & n3496 ) ;
  assign n3638 = ( n3562 & ~n3636 ) | ( n3562 & n3637 ) | ( ~n3636 & n3637 ) ;
  assign n3639 = ( n1208 & n3635 ) | ( n1208 & n3638 ) | ( n3635 & n3638 ) ;
  assign n3640 = ( x87 & ~n3635 ) | ( x87 & n3639 ) | ( ~n3635 & n3639 ) ;
  assign n3641 = ( n2074 & n2080 ) | ( n2074 & n3464 ) | ( n2080 & n3464 ) ;
  assign n3642 = ( x51 & n3464 ) | ( x51 & ~n3641 ) | ( n3464 & ~n3641 ) ;
  assign n3643 = n3484 & ~n3642 ;
  assign n3644 = ( n2681 & n2694 ) | ( n2681 & n3534 ) | ( n2694 & n3534 ) ;
  assign n3645 = n2600 | n3644 ;
  assign n3646 = n3486 & n3645 ;
  assign n3647 = n1282 | n3646 ;
  assign n3648 = n3543 | n3638 ;
  assign n3649 = x190 & n3453 ;
  assign n3650 = x51 & x173 ;
  assign n3651 = ( ~x299 & n3649 ) | ( ~x299 & n3650 ) | ( n3649 & n3650 ) ;
  assign n3652 = n2072 & n3651 ;
  assign n3653 = n1553 & n3635 ;
  assign n3654 = ( n2072 & n3652 ) | ( n2072 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3655 = n1282 & ~n3654 ;
  assign n3656 = ( ~n3647 & n3648 ) | ( ~n3647 & n3655 ) | ( n3648 & n3655 ) ;
  assign n3657 = n3640 | n3656 ;
  assign n3658 = ( n3640 & ~n3643 ) | ( n3640 & n3657 ) | ( ~n3643 & n3657 ) ;
  assign n3659 = ~n3632 & n3658 ;
  assign n3660 = n2560 | n3540 ;
  assign n3661 = ~n2664 & n3467 ;
  assign n3662 = n2760 | n3661 ;
  assign n3663 = ( n2760 & ~n3660 ) | ( n2760 & n3662 ) | ( ~n3660 & n3662 ) ;
  assign n3664 = ~x287 & n3549 ;
  assign n3665 = n3539 | n3663 ;
  assign n3666 = ( n3663 & ~n3664 ) | ( n3663 & n3665 ) | ( ~n3664 & n3665 ) ;
  assign n3667 = x133 & ~n3666 ;
  assign n3668 = ( n3620 & n3666 ) | ( n3620 & ~n3667 ) | ( n3666 & ~n3667 ) ;
  assign n3669 = ~n1208 & n2694 ;
  assign n3670 = ( x149 & n1208 ) | ( x149 & n2681 ) | ( n1208 & n2681 ) ;
  assign n3671 = ( n3525 & n3669 ) | ( n3525 & n3670 ) | ( n3669 & n3670 ) ;
  assign n3672 = n3668 & ~n3671 ;
  assign n3673 = ( x39 & n2043 ) | ( x39 & n2044 ) | ( n2043 & n2044 ) ;
  assign n3674 = ( n1282 & n2458 ) | ( n1282 & n3673 ) | ( n2458 & n3673 ) ;
  assign n3675 = n3673 & ~n3674 ;
  assign n3676 = n3485 | n3675 ;
  assign n3677 = ( n2669 & n2670 ) | ( n2669 & ~n2758 ) | ( n2670 & ~n2758 ) ;
  assign n3678 = n3534 & n3677 ;
  assign n3679 = ( n2758 & n3486 ) | ( n2758 & ~n3678 ) | ( n3486 & ~n3678 ) ;
  assign n3680 = x134 & ~n2760 ;
  assign n3681 = ( ~n3495 & n3539 ) | ( ~n3495 & n3680 ) | ( n3539 & n3680 ) ;
  assign n3682 = n3680 & ~n3681 ;
  assign n3683 = x192 & ~x299 ;
  assign n3684 = x171 & x299 ;
  assign n3685 = ( n2072 & n3683 ) | ( n2072 & n3684 ) | ( n3683 & n3684 ) ;
  assign n3686 = ( n1208 & n2072 ) | ( n1208 & n3685 ) | ( n2072 & n3685 ) ;
  assign n3687 = x171 & n2758 ;
  assign n3688 = ( ~n1208 & n2758 ) | ( ~n1208 & n3687 ) | ( n2758 & n3687 ) ;
  assign n3689 = n3686 & n3688 ;
  assign n3690 = ( n2759 & n3679 ) | ( n2759 & n3689 ) | ( n3679 & n3689 ) ;
  assign n3691 = ( n3679 & n3682 ) | ( n3679 & ~n3690 ) | ( n3682 & ~n3690 ) ;
  assign n3692 = ~n3676 & n3691 ;
  assign n3693 = n3484 | n3675 ;
  assign n3694 = x170 & x299 ;
  assign n3695 = x194 & ~x299 ;
  assign n3696 = ( n2072 & n3694 ) | ( n2072 & n3695 ) | ( n3694 & n3695 ) ;
  assign n3697 = n2758 & ~n3696 ;
  assign n3698 = x134 & ~x135 ;
  assign n3699 = ~n3494 & n3698 ;
  assign n3700 = x135 & n3494 ;
  assign n3701 = ( ~n3539 & n3699 ) | ( ~n3539 & n3700 ) | ( n3699 & n3700 ) ;
  assign n3702 = x185 & n2079 ;
  assign n3703 = x150 & n2073 ;
  assign n3704 = ( ~x287 & n3702 ) | ( ~x287 & n3703 ) | ( n3702 & n3703 ) ;
  assign n3705 = n3539 & ~n3704 ;
  assign n3706 = ( ~n2758 & n3701 ) | ( ~n2758 & n3705 ) | ( n3701 & n3705 ) ;
  assign n3707 = ( ~n1208 & n3697 ) | ( ~n1208 & n3706 ) | ( n3697 & n3706 ) ;
  assign n3708 = ~n3693 & n3707 ;
  assign n3709 = x170 & n2072 ;
  assign n3710 = n2758 & ~n3709 ;
  assign n3711 = ( ~n2758 & n3699 ) | ( ~n2758 & n3700 ) | ( n3699 & n3700 ) ;
  assign n3712 = ( n1208 & n3710 ) | ( n1208 & n3711 ) | ( n3710 & n3711 ) ;
  assign n3713 = ( ~n2759 & n3708 ) | ( ~n2759 & n3712 ) | ( n3708 & n3712 ) ;
  assign n3714 = ( n2072 & n2750 ) | ( n2072 & n2751 ) | ( n2750 & n2751 ) ;
  assign n3715 = ( n1208 & n2072 ) | ( n1208 & n3714 ) | ( n2072 & n3714 ) ;
  assign n3716 = n2759 | n3715 ;
  assign n3717 = n2758 & ~n2780 ;
  assign n3718 = ( n2759 & n3716 ) | ( n2759 & n3717 ) | ( n3716 & n3717 ) ;
  assign n3719 = ( n3182 & n3191 ) | ( n3182 & n3534 ) | ( n3191 & n3534 ) ;
  assign n3720 = n3486 & n3719 ;
  assign n3721 = ~x136 & n3493 ;
  assign n3722 = ( ~x136 & n3493 ) | ( ~x136 & n3496 ) | ( n3493 & n3496 ) ;
  assign n3723 = ( n3486 & ~n3721 ) | ( n3486 & n3722 ) | ( ~n3721 & n3722 ) ;
  assign n3724 = ( n2758 & ~n3720 ) | ( n2758 & n3723 ) | ( ~n3720 & n3723 ) ;
  assign n3725 = ~n3718 & n3724 ;
  assign n3726 = ~n3676 & n3725 ;
  assign n3727 = ~x39 & x137 ;
  assign n3728 = n1208 | n2027 ;
  assign n3729 = n2486 & ~n3728 ;
  assign n3730 = ~x210 & n1208 ;
  assign n3731 = n2942 & n3730 ;
  assign n3732 = ( x39 & n3729 ) | ( x39 & n3731 ) | ( n3729 & n3731 ) ;
  assign n3733 = n3727 | n3732 ;
  assign n3734 = ( ~n3294 & n3727 ) | ( ~n3294 & n3733 ) | ( n3727 & n3733 ) ;
  assign n3735 = n2619 & ~n3714 ;
  assign n3736 = x118 | n3355 ;
  assign n3737 = x139 | n3736 ;
  assign n3738 = ( x138 & n2625 ) | ( x138 & ~n3737 ) | ( n2625 & ~n3737 ) ;
  assign n3739 = ( x138 & n2621 ) | ( x138 & ~n3737 ) | ( n2621 & ~n3737 ) ;
  assign n3740 = n3738 & ~n3739 ;
  assign n3741 = n3735 | n3740 ;
  assign n3742 = n2619 & ~n2646 ;
  assign n3743 = ( ~x139 & n2621 ) | ( ~x139 & n3736 ) | ( n2621 & n3736 ) ;
  assign n3744 = ( ~x139 & n2625 ) | ( ~x139 & n3736 ) | ( n2625 & n3736 ) ;
  assign n3745 = n3742 | n3744 ;
  assign n3746 = ( n3742 & ~n3743 ) | ( n3742 & n3745 ) | ( ~n3743 & n3745 ) ;
  assign n3747 = x618 & x1154 ;
  assign n3748 = ( x618 & x781 ) | ( x618 & x1154 ) | ( x781 & x1154 ) ;
  assign n3749 = ( x630 & ~x787 ) | ( x630 & x1157 ) | ( ~x787 & x1157 ) ;
  assign n3750 = ( x630 & x787 ) | ( x630 & x1157 ) | ( x787 & x1157 ) ;
  assign n3751 = ~n3749 & n3750 ;
  assign n3752 = ( ~n3747 & n3748 ) | ( ~n3747 & n3751 ) | ( n3748 & n3751 ) ;
  assign n3753 = ( x608 & ~x778 ) | ( x608 & x1153 ) | ( ~x778 & x1153 ) ;
  assign n3754 = ( x608 & x778 ) | ( x608 & x1153 ) | ( x778 & x1153 ) ;
  assign n3755 = ~n3753 & n3754 ;
  assign n3756 = x609 & x1155 ;
  assign n3757 = ( x609 & x785 ) | ( x609 & x1155 ) | ( x785 & x1155 ) ;
  assign n3758 = ( n3755 & ~n3756 ) | ( n3755 & n3757 ) | ( ~n3756 & n3757 ) ;
  assign n3759 = n3752 | n3758 ;
  assign n3760 = x626 & x1158 ;
  assign n3761 = ( x626 & x788 ) | ( x626 & x1158 ) | ( x788 & x1158 ) ;
  assign n3762 = ( x603 & n3760 ) | ( x603 & ~n3761 ) | ( n3760 & ~n3761 ) ;
  assign n3763 = x619 & x1159 ;
  assign n3764 = ( x644 & ~x790 ) | ( x644 & x1160 ) | ( ~x790 & x1160 ) ;
  assign n3765 = ( x644 & x790 ) | ( x644 & x1160 ) | ( x790 & x1160 ) ;
  assign n3766 = ~n3764 & n3765 ;
  assign n3767 = ( x619 & x789 ) | ( x619 & x1159 ) | ( x789 & x1159 ) ;
  assign n3768 = ( ~n3763 & n3766 ) | ( ~n3763 & n3767 ) | ( n3766 & n3767 ) ;
  assign n3769 = x629 | x1156 ;
  assign n3770 = ( x629 & ~x792 ) | ( x629 & x1156 ) | ( ~x792 & x1156 ) ;
  assign n3771 = ( n3768 & n3769 ) | ( n3768 & ~n3770 ) | ( n3769 & ~n3770 ) ;
  assign n3772 = ( n3759 & n3762 ) | ( n3759 & ~n3771 ) | ( n3762 & ~n3771 ) ;
  assign n3773 = ~n3759 & n3772 ;
  assign n3774 = x621 & x1091 ;
  assign n3775 = n3773 & ~n3774 ;
  assign n3776 = ~x761 & n3775 ;
  assign n3777 = x45 | n1209 ;
  assign n3778 = n2850 | n3777 ;
  assign n3779 = n2802 | n2840 ;
  assign n3780 = ~n1960 & n3779 ;
  assign n3781 = x47 & x252 ;
  assign n3782 = ( x252 & n3780 ) | ( x252 & n3781 ) | ( n3780 & n3781 ) ;
  assign n3783 = x1093 & n1443 ;
  assign n3784 = n2027 & n3783 ;
  assign n3785 = ( n1995 & n3097 ) | ( n1995 & n3784 ) | ( n3097 & n3784 ) ;
  assign n3786 = ( ~n3778 & n3782 ) | ( ~n3778 & n3785 ) | ( n3782 & n3785 ) ;
  assign n3787 = n3778 | n3786 ;
  assign n3788 = ~n2016 & n3787 ;
  assign n3789 = ( ~x120 & n2132 ) | ( ~x120 & n3075 ) | ( n2132 & n3075 ) ;
  assign n3790 = n2612 & n3431 ;
  assign n3791 = n3789 & ~n3790 ;
  assign n3792 = ( n2618 & ~n3788 ) | ( n2618 & n3791 ) | ( ~n3788 & n3791 ) ;
  assign n3793 = n2618 & ~n3792 ;
  assign n3794 = n1430 & n3793 ;
  assign n3795 = ( x832 & n1430 ) | ( x832 & n3794 ) | ( n1430 & n3794 ) ;
  assign n3796 = x140 & ~n3795 ;
  assign n3797 = x648 & x1159 ;
  assign n3798 = ( x628 & ~x792 ) | ( x628 & x1156 ) | ( ~x792 & x1156 ) ;
  assign n3799 = ( x628 & x792 ) | ( x628 & x1156 ) | ( x792 & x1156 ) ;
  assign n3800 = ~n3798 & n3799 ;
  assign n3801 = ( x648 & x789 ) | ( x648 & x1159 ) | ( x789 & x1159 ) ;
  assign n3802 = ( ~n3797 & n3800 ) | ( ~n3797 & n3801 ) | ( n3800 & n3801 ) ;
  assign n3803 = ( x641 & ~x788 ) | ( x641 & x1158 ) | ( ~x788 & x1158 ) ;
  assign n3804 = ( x641 & x788 ) | ( x641 & x1158 ) | ( x788 & x1158 ) ;
  assign n3805 = ~n3803 & n3804 ;
  assign n3806 = x627 & x1154 ;
  assign n3807 = ( x627 & x781 ) | ( x627 & x1154 ) | ( x781 & x1154 ) ;
  assign n3808 = ( n3805 & ~n3806 ) | ( n3805 & n3807 ) | ( ~n3806 & n3807 ) ;
  assign n3809 = n3802 | n3808 ;
  assign n3810 = x660 | x1155 ;
  assign n3811 = ( x660 & ~x785 ) | ( x660 & x1155 ) | ( ~x785 & x1155 ) ;
  assign n3812 = ( x680 & ~n3810 ) | ( x680 & n3811 ) | ( ~n3810 & n3811 ) ;
  assign n3813 = ~n3809 & n3812 ;
  assign n3814 = x647 | x1157 ;
  assign n3815 = x625 & x1153 ;
  assign n3816 = ( x625 & x778 ) | ( x625 & x1153 ) | ( x778 & x1153 ) ;
  assign n3817 = ( x715 & ~x790 ) | ( x715 & x1160 ) | ( ~x790 & x1160 ) ;
  assign n3818 = ( x715 & x790 ) | ( x715 & x1160 ) | ( x790 & x1160 ) ;
  assign n3819 = ~n3817 & n3818 ;
  assign n3820 = ( ~n3815 & n3816 ) | ( ~n3815 & n3819 ) | ( n3816 & n3819 ) ;
  assign n3821 = ( x647 & ~x787 ) | ( x647 & x1157 ) | ( ~x787 & x1157 ) ;
  assign n3822 = ( n3814 & n3820 ) | ( n3814 & ~n3821 ) | ( n3820 & ~n3821 ) ;
  assign n3823 = n3813 & ~n3822 ;
  assign n3824 = x665 & x1091 ;
  assign n3825 = n3823 & ~n3824 ;
  assign n3826 = ~n3775 & n3825 ;
  assign n3827 = ~x738 & n3826 ;
  assign n3828 = ( n3776 & n3795 ) | ( n3776 & ~n3827 ) | ( n3795 & ~n3827 ) ;
  assign n3829 = ( ~n3776 & n3796 ) | ( ~n3776 & n3828 ) | ( n3796 & n3828 ) ;
  assign n3830 = x141 & ~n3795 ;
  assign n3831 = x706 & n3826 ;
  assign n3832 = x749 & n3775 ;
  assign n3833 = ( n3795 & n3831 ) | ( n3795 & ~n3832 ) | ( n3831 & ~n3832 ) ;
  assign n3834 = ( n3830 & ~n3831 ) | ( n3830 & n3833 ) | ( ~n3831 & n3833 ) ;
  assign n3835 = x142 | n3795 ;
  assign n3836 = x735 & n3826 ;
  assign n3837 = x743 & n3775 ;
  assign n3838 = ( n3795 & n3836 ) | ( n3795 & ~n3837 ) | ( n3836 & ~n3837 ) ;
  assign n3839 = ( n3835 & n3836 ) | ( n3835 & ~n3838 ) | ( n3836 & ~n3838 ) ;
  assign n3840 = x143 & ~n3795 ;
  assign n3841 = ~x774 & n3775 ;
  assign n3842 = x687 & n3826 ;
  assign n3843 = ( n3795 & n3841 ) | ( n3795 & ~n3842 ) | ( n3841 & ~n3842 ) ;
  assign n3844 = ( n3840 & ~n3841 ) | ( n3840 & n3843 ) | ( ~n3841 & n3843 ) ;
  assign n3845 = x144 | n3795 ;
  assign n3846 = x758 & n3775 ;
  assign n3847 = x736 & n3826 ;
  assign n3848 = ( n3795 & n3846 ) | ( n3795 & ~n3847 ) | ( n3846 & ~n3847 ) ;
  assign n3849 = ( n3845 & n3846 ) | ( n3845 & ~n3848 ) | ( n3846 & ~n3848 ) ;
  assign n3850 = x145 & ~n3795 ;
  assign n3851 = ~x698 & n3826 ;
  assign n3852 = ~x767 & n3775 ;
  assign n3853 = ( n3795 & n3851 ) | ( n3795 & ~n3852 ) | ( n3851 & ~n3852 ) ;
  assign n3854 = ( n3850 & ~n3851 ) | ( n3850 & n3853 ) | ( ~n3851 & n3853 ) ;
  assign n3855 = x146 & ~n3795 ;
  assign n3856 = ~x743 & x947 ;
  assign n3857 = ( x735 & x947 ) | ( x735 & n2007 ) | ( x947 & n2007 ) ;
  assign n3858 = ( n3795 & n3856 ) | ( n3795 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3859 = ( n3855 & ~n3856 ) | ( n3855 & n3858 ) | ( ~n3856 & n3858 ) ;
  assign n3860 = x147 | n3795 ;
  assign n3861 = ( x726 & x947 ) | ( x726 & n2007 ) | ( x947 & n2007 ) ;
  assign n3862 = x770 & x947 ;
  assign n3863 = ( ~n3795 & n3861 ) | ( ~n3795 & n3862 ) | ( n3861 & n3862 ) ;
  assign n3864 = ( n3860 & ~n3861 ) | ( n3860 & n3863 ) | ( ~n3861 & n3863 ) ;
  assign n3865 = x148 | n3795 ;
  assign n3866 = ( x706 & x947 ) | ( x706 & n2007 ) | ( x947 & n2007 ) ;
  assign n3867 = ~x749 & x947 ;
  assign n3868 = ( ~n3795 & n3866 ) | ( ~n3795 & n3867 ) | ( n3866 & n3867 ) ;
  assign n3869 = ( n3865 & ~n3866 ) | ( n3865 & n3868 ) | ( ~n3866 & n3868 ) ;
  assign n3870 = x149 | n3795 ;
  assign n3871 = ( ~x725 & x947 ) | ( ~x725 & n2007 ) | ( x947 & n2007 ) ;
  assign n3872 = x755 & x947 ;
  assign n3873 = ( ~n3795 & n3871 ) | ( ~n3795 & n3872 ) | ( n3871 & n3872 ) ;
  assign n3874 = ( n3870 & ~n3871 ) | ( n3870 & n3873 ) | ( ~n3871 & n3873 ) ;
  assign n3875 = x150 | n3795 ;
  assign n3876 = x751 & x947 ;
  assign n3877 = ( ~x701 & x947 ) | ( ~x701 & n2007 ) | ( x947 & n2007 ) ;
  assign n3878 = ( n3795 & n3876 ) | ( n3795 & n3877 ) | ( n3876 & n3877 ) ;
  assign n3879 = ( n3875 & n3876 ) | ( n3875 & ~n3878 ) | ( n3876 & ~n3878 ) ;
  assign n3880 = x151 | n3795 ;
  assign n3881 = ( ~x723 & x947 ) | ( ~x723 & n2007 ) | ( x947 & n2007 ) ;
  assign n3882 = x745 & x947 ;
  assign n3883 = ( ~n3795 & n3881 ) | ( ~n3795 & n3882 ) | ( n3881 & n3882 ) ;
  assign n3884 = ( n3880 & ~n3881 ) | ( n3880 & n3883 ) | ( ~n3881 & n3883 ) ;
  assign n3885 = x152 & ~n3795 ;
  assign n3886 = ~x759 & x947 ;
  assign n3887 = ( x696 & x947 ) | ( x696 & n2007 ) | ( x947 & n2007 ) ;
  assign n3888 = ( n3795 & n3886 ) | ( n3795 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3889 = ( n3885 & ~n3886 ) | ( n3885 & n3888 ) | ( ~n3886 & n3888 ) ;
  assign n3890 = x153 | n3795 ;
  assign n3891 = ~x766 & x947 ;
  assign n3892 = ( x700 & x947 ) | ( x700 & n2007 ) | ( x947 & n2007 ) ;
  assign n3893 = ( n3795 & n3891 ) | ( n3795 & n3892 ) | ( n3891 & n3892 ) ;
  assign n3894 = ( n3890 & n3891 ) | ( n3890 & ~n3893 ) | ( n3891 & ~n3893 ) ;
  assign n3895 = x154 | n3795 ;
  assign n3896 = ( ~x704 & x947 ) | ( ~x704 & n2007 ) | ( x947 & n2007 ) ;
  assign n3897 = x742 & x947 ;
  assign n3898 = ( ~n3795 & n3896 ) | ( ~n3795 & n3897 ) | ( n3896 & n3897 ) ;
  assign n3899 = ( n3895 & ~n3896 ) | ( n3895 & n3898 ) | ( ~n3896 & n3898 ) ;
  assign n3900 = x155 | n3795 ;
  assign n3901 = x757 & x947 ;
  assign n3902 = ( ~x686 & x947 ) | ( ~x686 & n2007 ) | ( x947 & n2007 ) ;
  assign n3903 = ( n3795 & n3901 ) | ( n3795 & n3902 ) | ( n3901 & n3902 ) ;
  assign n3904 = ( n3900 & n3901 ) | ( n3900 & ~n3903 ) | ( n3901 & ~n3903 ) ;
  assign n3905 = x156 | n3795 ;
  assign n3906 = ( ~x724 & x947 ) | ( ~x724 & n2007 ) | ( x947 & n2007 ) ;
  assign n3907 = x741 & x947 ;
  assign n3908 = ( ~n3795 & n3906 ) | ( ~n3795 & n3907 ) | ( n3906 & n3907 ) ;
  assign n3909 = ( n3905 & ~n3906 ) | ( n3905 & n3908 ) | ( ~n3906 & n3908 ) ;
  assign n3910 = x157 | n3795 ;
  assign n3911 = ( ~x688 & x947 ) | ( ~x688 & n2007 ) | ( x947 & n2007 ) ;
  assign n3912 = x760 & x947 ;
  assign n3913 = ( ~n3795 & n3911 ) | ( ~n3795 & n3912 ) | ( n3911 & n3912 ) ;
  assign n3914 = ( n3910 & ~n3911 ) | ( n3910 & n3913 ) | ( ~n3911 & n3913 ) ;
  assign n3915 = x158 | n3795 ;
  assign n3916 = ( ~x702 & x947 ) | ( ~x702 & n2007 ) | ( x947 & n2007 ) ;
  assign n3917 = x753 & x947 ;
  assign n3918 = ( ~n3795 & n3916 ) | ( ~n3795 & n3917 ) | ( n3916 & n3917 ) ;
  assign n3919 = ( n3915 & ~n3916 ) | ( n3915 & n3918 ) | ( ~n3916 & n3918 ) ;
  assign n3920 = x159 | n3795 ;
  assign n3921 = ( ~x709 & x947 ) | ( ~x709 & n2007 ) | ( x947 & n2007 ) ;
  assign n3922 = x754 & x947 ;
  assign n3923 = ( ~n3795 & n3921 ) | ( ~n3795 & n3922 ) | ( n3921 & n3922 ) ;
  assign n3924 = ( n3920 & ~n3921 ) | ( n3920 & n3923 ) | ( ~n3921 & n3923 ) ;
  assign n3925 = x160 | n3795 ;
  assign n3926 = ( ~x734 & x947 ) | ( ~x734 & n2007 ) | ( x947 & n2007 ) ;
  assign n3927 = x756 & x947 ;
  assign n3928 = ( ~n3795 & n3926 ) | ( ~n3795 & n3927 ) | ( n3926 & n3927 ) ;
  assign n3929 = ( n3925 & ~n3926 ) | ( n3925 & n3928 ) | ( ~n3926 & n3928 ) ;
  assign n3930 = x161 & ~n3795 ;
  assign n3931 = ( x736 & x947 ) | ( x736 & n2007 ) | ( x947 & n2007 ) ;
  assign n3932 = ~x758 & x947 ;
  assign n3933 = ( ~n3795 & n3931 ) | ( ~n3795 & n3932 ) | ( n3931 & n3932 ) ;
  assign n3934 = ( n3930 & n3931 ) | ( n3930 & ~n3933 ) | ( n3931 & ~n3933 ) ;
  assign n3935 = x162 | n3795 ;
  assign n3936 = x761 & x947 ;
  assign n3937 = ( ~x738 & x947 ) | ( ~x738 & n2007 ) | ( x947 & n2007 ) ;
  assign n3938 = ( n3795 & n3936 ) | ( n3795 & n3937 ) | ( n3936 & n3937 ) ;
  assign n3939 = ( n3935 & n3936 ) | ( n3935 & ~n3938 ) | ( n3936 & ~n3938 ) ;
  assign n3940 = x163 | n3795 ;
  assign n3941 = ( ~x737 & x947 ) | ( ~x737 & n2007 ) | ( x947 & n2007 ) ;
  assign n3942 = x777 & x947 ;
  assign n3943 = ( ~n3795 & n3941 ) | ( ~n3795 & n3942 ) | ( n3941 & n3942 ) ;
  assign n3944 = ( n3940 & ~n3941 ) | ( n3940 & n3943 ) | ( ~n3941 & n3943 ) ;
  assign n3945 = x164 | n3795 ;
  assign n3946 = x752 & x947 ;
  assign n3947 = ( x703 & x947 ) | ( x703 & n2007 ) | ( x947 & n2007 ) ;
  assign n3948 = ( n3795 & n3946 ) | ( n3795 & n3947 ) | ( n3946 & n3947 ) ;
  assign n3949 = ( n3945 & n3946 ) | ( n3945 & ~n3948 ) | ( n3946 & ~n3948 ) ;
  assign n3950 = x165 | n3795 ;
  assign n3951 = ( x687 & x947 ) | ( x687 & n2007 ) | ( x947 & n2007 ) ;
  assign n3952 = x774 & x947 ;
  assign n3953 = ( ~n3795 & n3951 ) | ( ~n3795 & n3952 ) | ( n3951 & n3952 ) ;
  assign n3954 = ( n3950 & ~n3951 ) | ( n3950 & n3953 ) | ( ~n3951 & n3953 ) ;
  assign n3955 = x166 & ~n3795 ;
  assign n3956 = ~x772 & x947 ;
  assign n3957 = ( x727 & x947 ) | ( x727 & n2007 ) | ( x947 & n2007 ) ;
  assign n3958 = ( n3795 & n3956 ) | ( n3795 & n3957 ) | ( n3956 & n3957 ) ;
  assign n3959 = ( n3955 & ~n3956 ) | ( n3955 & n3958 ) | ( ~n3956 & n3958 ) ;
  assign n3960 = x167 | n3795 ;
  assign n3961 = ( x705 & x947 ) | ( x705 & n2007 ) | ( x947 & n2007 ) ;
  assign n3962 = x768 & x947 ;
  assign n3963 = ( ~n3795 & n3961 ) | ( ~n3795 & n3962 ) | ( n3961 & n3962 ) ;
  assign n3964 = ( n3960 & ~n3961 ) | ( n3960 & n3963 ) | ( ~n3961 & n3963 ) ;
  assign n3965 = x168 | n3795 ;
  assign n3966 = ~x763 & x947 ;
  assign n3967 = ( x699 & x947 ) | ( x699 & n2007 ) | ( x947 & n2007 ) ;
  assign n3968 = ( n3795 & n3966 ) | ( n3795 & n3967 ) | ( n3966 & n3967 ) ;
  assign n3969 = ( n3965 & n3966 ) | ( n3965 & ~n3968 ) | ( n3966 & ~n3968 ) ;
  assign n3970 = x169 | n3795 ;
  assign n3971 = ~x746 & x947 ;
  assign n3972 = ( x729 & x947 ) | ( x729 & n2007 ) | ( x947 & n2007 ) ;
  assign n3973 = ( n3795 & n3971 ) | ( n3795 & n3972 ) | ( n3971 & n3972 ) ;
  assign n3974 = ( n3970 & n3971 ) | ( n3970 & ~n3973 ) | ( n3971 & ~n3973 ) ;
  assign n3975 = x170 | n3795 ;
  assign n3976 = ~x748 & x947 ;
  assign n3977 = ( x730 & x947 ) | ( x730 & n2007 ) | ( x947 & n2007 ) ;
  assign n3978 = ( n3795 & n3976 ) | ( n3795 & n3977 ) | ( n3976 & n3977 ) ;
  assign n3979 = ( n3975 & n3976 ) | ( n3975 & ~n3978 ) | ( n3976 & ~n3978 ) ;
  assign n3980 = x171 | n3795 ;
  assign n3981 = ~x764 & x947 ;
  assign n3982 = ( x691 & x947 ) | ( x691 & n2007 ) | ( x947 & n2007 ) ;
  assign n3983 = ( n3795 & n3981 ) | ( n3795 & n3982 ) | ( n3981 & n3982 ) ;
  assign n3984 = ( n3980 & n3981 ) | ( n3980 & ~n3983 ) | ( n3981 & ~n3983 ) ;
  assign n3985 = x172 | n3795 ;
  assign n3986 = ~x739 & x947 ;
  assign n3987 = ( x690 & x947 ) | ( x690 & n2007 ) | ( x947 & n2007 ) ;
  assign n3988 = ( n3795 & n3986 ) | ( n3795 & n3987 ) | ( n3986 & n3987 ) ;
  assign n3989 = ( n3985 & n3986 ) | ( n3985 & ~n3988 ) | ( n3986 & ~n3988 ) ;
  assign n3990 = x173 & ~n3795 ;
  assign n3991 = ~x745 & n3775 ;
  assign n3992 = ~x723 & n3826 ;
  assign n3993 = ( n3795 & n3991 ) | ( n3795 & ~n3992 ) | ( n3991 & ~n3992 ) ;
  assign n3994 = ( n3990 & ~n3991 ) | ( n3990 & n3993 ) | ( ~n3991 & n3993 ) ;
  assign n3995 = x174 | n3795 ;
  assign n3996 = x696 & n3826 ;
  assign n3997 = x759 & n3775 ;
  assign n3998 = ( n3795 & n3996 ) | ( n3795 & ~n3997 ) | ( n3996 & ~n3997 ) ;
  assign n3999 = ( n3995 & n3996 ) | ( n3995 & ~n3998 ) | ( n3996 & ~n3998 ) ;
  assign n4000 = x175 & ~n3795 ;
  assign n4001 = x700 & n3826 ;
  assign n4002 = x766 & n3775 ;
  assign n4003 = ( n3795 & n4001 ) | ( n3795 & ~n4002 ) | ( n4001 & ~n4002 ) ;
  assign n4004 = ( n4000 & ~n4001 ) | ( n4000 & n4003 ) | ( ~n4001 & n4003 ) ;
  assign n4005 = x176 & ~n3795 ;
  assign n4006 = ~x704 & n3826 ;
  assign n4007 = ~x742 & n3775 ;
  assign n4008 = ( n3795 & n4006 ) | ( n3795 & ~n4007 ) | ( n4006 & ~n4007 ) ;
  assign n4009 = ( n4005 & ~n4006 ) | ( n4005 & n4008 ) | ( ~n4006 & n4008 ) ;
  assign n4010 = x177 & ~n3795 ;
  assign n4011 = ~x757 & n3775 ;
  assign n4012 = ~x686 & n3826 ;
  assign n4013 = ( n3795 & n4011 ) | ( n3795 & ~n4012 ) | ( n4011 & ~n4012 ) ;
  assign n4014 = ( n4010 & ~n4011 ) | ( n4010 & n4013 ) | ( ~n4011 & n4013 ) ;
  assign n4015 = x178 & ~n3795 ;
  assign n4016 = ~x760 & n3775 ;
  assign n4017 = ~x688 & n3826 ;
  assign n4018 = ( n3795 & n4016 ) | ( n3795 & ~n4017 ) | ( n4016 & ~n4017 ) ;
  assign n4019 = ( n4015 & ~n4016 ) | ( n4015 & n4018 ) | ( ~n4016 & n4018 ) ;
  assign n4020 = x179 & ~n3795 ;
  assign n4021 = ~x741 & n3775 ;
  assign n4022 = ~x724 & n3826 ;
  assign n4023 = ( n3795 & n4021 ) | ( n3795 & ~n4022 ) | ( n4021 & ~n4022 ) ;
  assign n4024 = ( n4020 & ~n4021 ) | ( n4020 & n4023 ) | ( ~n4021 & n4023 ) ;
  assign n4025 = x180 & ~n3795 ;
  assign n4026 = ~x702 & n3826 ;
  assign n4027 = ~x753 & n3775 ;
  assign n4028 = ( n3795 & n4026 ) | ( n3795 & ~n4027 ) | ( n4026 & ~n4027 ) ;
  assign n4029 = ( n4025 & ~n4026 ) | ( n4025 & n4028 ) | ( ~n4026 & n4028 ) ;
  assign n4030 = x181 & ~n3795 ;
  assign n4031 = ~x709 & n3826 ;
  assign n4032 = ~x754 & n3775 ;
  assign n4033 = ( n3795 & n4031 ) | ( n3795 & ~n4032 ) | ( n4031 & ~n4032 ) ;
  assign n4034 = ( n4030 & ~n4031 ) | ( n4030 & n4033 ) | ( ~n4031 & n4033 ) ;
  assign n4035 = x182 & ~n3795 ;
  assign n4036 = ~x734 & n3826 ;
  assign n4037 = ~x756 & n3775 ;
  assign n4038 = ( n3795 & n4036 ) | ( n3795 & ~n4037 ) | ( n4036 & ~n4037 ) ;
  assign n4039 = ( n4035 & ~n4036 ) | ( n4035 & n4038 ) | ( ~n4036 & n4038 ) ;
  assign n4040 = x183 & ~n3795 ;
  assign n4041 = ~x755 & n3775 ;
  assign n4042 = ~x725 & n3826 ;
  assign n4043 = ( n3795 & n4041 ) | ( n3795 & ~n4042 ) | ( n4041 & ~n4042 ) ;
  assign n4044 = ( n4040 & ~n4041 ) | ( n4040 & n4043 ) | ( ~n4041 & n4043 ) ;
  assign n4045 = x184 & ~n3795 ;
  assign n4046 = ~x777 & n3775 ;
  assign n4047 = ~x737 & n3826 ;
  assign n4048 = ( n3795 & n4046 ) | ( n3795 & ~n4047 ) | ( n4046 & ~n4047 ) ;
  assign n4049 = ( n4045 & ~n4046 ) | ( n4045 & n4048 ) | ( ~n4046 & n4048 ) ;
  assign n4050 = x185 & ~n3795 ;
  assign n4051 = ~x701 & n3826 ;
  assign n4052 = ~x751 & n3775 ;
  assign n4053 = ( n3795 & n4051 ) | ( n3795 & ~n4052 ) | ( n4051 & ~n4052 ) ;
  assign n4054 = ( n4050 & ~n4051 ) | ( n4050 & n4053 ) | ( ~n4051 & n4053 ) ;
  assign n4055 = x186 & ~n3795 ;
  assign n4056 = x703 & n3826 ;
  assign n4057 = ~x752 & n3775 ;
  assign n4058 = ( n3795 & n4056 ) | ( n3795 & ~n4057 ) | ( n4056 & ~n4057 ) ;
  assign n4059 = ( n4055 & ~n4056 ) | ( n4055 & n4058 ) | ( ~n4056 & n4058 ) ;
  assign n4060 = x187 & ~n3795 ;
  assign n4061 = x726 & n3826 ;
  assign n4062 = ~x770 & n3775 ;
  assign n4063 = ( n3795 & n4061 ) | ( n3795 & ~n4062 ) | ( n4061 & ~n4062 ) ;
  assign n4064 = ( n4060 & ~n4061 ) | ( n4060 & n4063 ) | ( ~n4061 & n4063 ) ;
  assign n4065 = x188 & ~n3795 ;
  assign n4066 = ~x768 & n3775 ;
  assign n4067 = x705 & n3826 ;
  assign n4068 = ( n3795 & n4066 ) | ( n3795 & ~n4067 ) | ( n4066 & ~n4067 ) ;
  assign n4069 = ( n4065 & ~n4066 ) | ( n4065 & n4068 ) | ( ~n4066 & n4068 ) ;
  assign n4070 = x189 | n3795 ;
  assign n4071 = x727 & n3826 ;
  assign n4072 = x772 & n3775 ;
  assign n4073 = ( n3795 & n4071 ) | ( n3795 & ~n4072 ) | ( n4071 & ~n4072 ) ;
  assign n4074 = ( n4070 & n4071 ) | ( n4070 & ~n4073 ) | ( n4071 & ~n4073 ) ;
  assign n4075 = x190 & ~n3795 ;
  assign n4076 = x699 & n3826 ;
  assign n4077 = x763 & n3775 ;
  assign n4078 = ( n3795 & n4076 ) | ( n3795 & ~n4077 ) | ( n4076 & ~n4077 ) ;
  assign n4079 = ( n4075 & ~n4076 ) | ( n4075 & n4078 ) | ( ~n4076 & n4078 ) ;
  assign n4080 = x191 & ~n3795 ;
  assign n4081 = x729 & n3826 ;
  assign n4082 = x746 & n3775 ;
  assign n4083 = ( n3795 & n4081 ) | ( n3795 & ~n4082 ) | ( n4081 & ~n4082 ) ;
  assign n4084 = ( n4080 & ~n4081 ) | ( n4080 & n4083 ) | ( ~n4081 & n4083 ) ;
  assign n4085 = x192 & ~n3795 ;
  assign n4086 = x691 & n3826 ;
  assign n4087 = x764 & n3775 ;
  assign n4088 = ( n3795 & n4086 ) | ( n3795 & ~n4087 ) | ( n4086 & ~n4087 ) ;
  assign n4089 = ( n4085 & ~n4086 ) | ( n4085 & n4088 ) | ( ~n4086 & n4088 ) ;
  assign n4090 = x193 & ~n3795 ;
  assign n4091 = x739 & n3775 ;
  assign n4092 = x690 & n3826 ;
  assign n4093 = ( n3795 & n4091 ) | ( n3795 & ~n4092 ) | ( n4091 & ~n4092 ) ;
  assign n4094 = ( n4090 & ~n4091 ) | ( n4090 & n4093 ) | ( ~n4091 & n4093 ) ;
  assign n4095 = x194 & ~n3795 ;
  assign n4096 = x748 & n3775 ;
  assign n4097 = x730 & n3826 ;
  assign n4098 = ( n3795 & n4096 ) | ( n3795 & ~n4097 ) | ( n4096 & ~n4097 ) ;
  assign n4099 = ( n4095 & ~n4096 ) | ( n4095 & n4098 ) | ( ~n4096 & n4098 ) ;
  assign n4100 = x138 | n3737 ;
  assign n4101 = x195 & x196 ;
  assign n4102 = ( x195 & n4100 ) | ( x195 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4103 = ~n2621 & n4102 ;
  assign n4104 = n2619 & ~n3685 ;
  assign n4105 = n4103 | n4104 ;
  assign n4106 = n2619 & ~n3696 ;
  assign n4107 = x195 & ~x196 ;
  assign n4108 = ~n4100 & n4107 ;
  assign n4109 = x196 & n4100 ;
  assign n4110 = ( ~n2621 & n4108 ) | ( ~n2621 & n4109 ) | ( n4108 & n4109 ) ;
  assign n4111 = n4106 | n4110 ;
  assign n4112 = x197 | n3795 ;
  assign n4113 = ( ~x698 & x947 ) | ( ~x698 & n2007 ) | ( x947 & n2007 ) ;
  assign n4114 = x767 & x947 ;
  assign n4115 = ( ~n3795 & n4113 ) | ( ~n3795 & n4114 ) | ( n4113 & n4114 ) ;
  assign n4116 = ( n4112 & ~n4113 ) | ( n4112 & n4115 ) | ( ~n4113 & n4115 ) ;
  assign n4117 = x634 & n3826 ;
  assign n4118 = x633 & n3775 ;
  assign n4119 = ( n3794 & n4117 ) | ( n3794 & ~n4118 ) | ( n4117 & ~n4118 ) ;
  assign n4120 = x198 | n3794 ;
  assign n4121 = ( n4117 & ~n4119 ) | ( n4117 & n4120 ) | ( ~n4119 & n4120 ) ;
  assign n4122 = x199 | n3794 ;
  assign n4123 = x637 & n3826 ;
  assign n4124 = x617 & n3775 ;
  assign n4125 = ( n3794 & n4123 ) | ( n3794 & ~n4124 ) | ( n4123 & ~n4124 ) ;
  assign n4126 = ( n4122 & n4123 ) | ( n4122 & ~n4125 ) | ( n4123 & ~n4125 ) ;
  assign n4127 = x200 | n3794 ;
  assign n4128 = x643 & n3826 ;
  assign n4129 = x606 & n3775 ;
  assign n4130 = ( n3794 & n4128 ) | ( n3794 & ~n4129 ) | ( n4128 & ~n4129 ) ;
  assign n4131 = ( n4127 & n4128 ) | ( n4127 & ~n4130 ) | ( n4128 & ~n4130 ) ;
  assign n4132 = x233 & x237 ;
  assign n4133 = n3728 & ~n3730 ;
  assign n4134 = x96 & n4133 ;
  assign n4135 = n4132 & n4134 ;
  assign n4136 = n2105 & n4135 ;
  assign n4137 = n1420 & ~n2995 ;
  assign n4138 = ( ~n3003 & n3011 ) | ( ~n3003 & n4137 ) | ( n3011 & n4137 ) ;
  assign n4139 = n3003 | n4138 ;
  assign n4140 = ~x32 & x70 ;
  assign n4141 = ~x70 & n1443 ;
  assign n4142 = ( ~n3728 & n3730 ) | ( ~n3728 & n4141 ) | ( n3730 & n4141 ) ;
  assign n4143 = ( n4132 & n4140 ) | ( n4132 & n4142 ) | ( n4140 & n4142 ) ;
  assign n4144 = n4139 | n4143 ;
  assign n4145 = n2105 & n4144 ;
  assign n4146 = x201 | x332 ;
  assign n4147 = ~n4136 & n4146 ;
  assign n4148 = ( ~n4136 & n4145 ) | ( ~n4136 & n4147 ) | ( n4145 & n4147 ) ;
  assign n4149 = ~x233 & x237 ;
  assign n4150 = n4134 & n4149 ;
  assign n4151 = n2105 & n4150 ;
  assign n4152 = ( n4140 & n4142 ) | ( n4140 & n4149 ) | ( n4142 & n4149 ) ;
  assign n4153 = n4139 | n4152 ;
  assign n4154 = n2105 & n4153 ;
  assign n4155 = x202 | x332 ;
  assign n4156 = ~n4151 & n4155 ;
  assign n4157 = ( ~n4151 & n4154 ) | ( ~n4151 & n4156 ) | ( n4154 & n4156 ) ;
  assign n4158 = x233 | x237 ;
  assign n4159 = n4134 & ~n4158 ;
  assign n4160 = n2105 & n4159 ;
  assign n4161 = x203 | x332 ;
  assign n4162 = n2105 | n4161 ;
  assign n4163 = ( n4140 & n4142 ) | ( n4140 & ~n4158 ) | ( n4142 & ~n4158 ) ;
  assign n4164 = n4139 | n4163 ;
  assign n4165 = ( n4161 & n4162 ) | ( n4161 & n4164 ) | ( n4162 & n4164 ) ;
  assign n4166 = ~n4160 & n4165 ;
  assign n4167 = n2037 & n4135 ;
  assign n4168 = x204 | x332 ;
  assign n4169 = n2037 | n4168 ;
  assign n4170 = ( n4144 & n4168 ) | ( n4144 & n4169 ) | ( n4168 & n4169 ) ;
  assign n4171 = ~n4167 & n4170 ;
  assign n4172 = n2037 & n4150 ;
  assign n4173 = x205 | x332 ;
  assign n4174 = n2037 | n4173 ;
  assign n4175 = ( n4153 & n4173 ) | ( n4153 & n4174 ) | ( n4173 & n4174 ) ;
  assign n4176 = ~n4172 & n4175 ;
  assign n4177 = x233 & ~x237 ;
  assign n4178 = n4134 & n4177 ;
  assign n4179 = n2037 & n4178 ;
  assign n4180 = ( n4140 & n4142 ) | ( n4140 & n4177 ) | ( n4142 & n4177 ) ;
  assign n4181 = n4139 | n4180 ;
  assign n4182 = n2037 & n4181 ;
  assign n4183 = x206 | x332 ;
  assign n4184 = ~n4179 & n4183 ;
  assign n4185 = ( ~n4179 & n4182 ) | ( ~n4179 & n4184 ) | ( n4182 & n4184 ) ;
  assign n4186 = x207 & ~n3794 ;
  assign n4187 = x623 & n3775 ;
  assign n4188 = x710 & n3826 ;
  assign n4189 = ( n3794 & n4187 ) | ( n3794 & ~n4188 ) | ( n4187 & ~n4188 ) ;
  assign n4190 = ( n4186 & ~n4187 ) | ( n4186 & n4189 ) | ( ~n4187 & n4189 ) ;
  assign n4191 = x208 & ~n3794 ;
  assign n4192 = x607 & n3775 ;
  assign n4193 = x638 & n3826 ;
  assign n4194 = ( n3794 & n4192 ) | ( n3794 & ~n4193 ) | ( n4192 & ~n4193 ) ;
  assign n4195 = ( n4191 & ~n4192 ) | ( n4191 & n4194 ) | ( ~n4192 & n4194 ) ;
  assign n4196 = x209 & ~n3794 ;
  assign n4197 = x622 & n3775 ;
  assign n4198 = x639 & n3826 ;
  assign n4199 = ( n3794 & n4197 ) | ( n3794 & ~n4198 ) | ( n4197 & ~n4198 ) ;
  assign n4200 = ( n4196 & ~n4197 ) | ( n4196 & n4199 ) | ( ~n4197 & n4199 ) ;
  assign n4201 = x210 & ~n3794 ;
  assign n4202 = ~x633 & x947 ;
  assign n4203 = ( x634 & x947 ) | ( x634 & n2007 ) | ( x947 & n2007 ) ;
  assign n4204 = ( n3794 & n4202 ) | ( n3794 & n4203 ) | ( n4202 & n4203 ) ;
  assign n4205 = ( n4201 & ~n4202 ) | ( n4201 & n4204 ) | ( ~n4202 & n4204 ) ;
  assign n4206 = x211 & ~n3794 ;
  assign n4207 = ~x606 & x947 ;
  assign n4208 = ( x643 & x947 ) | ( x643 & n2007 ) | ( x947 & n2007 ) ;
  assign n4209 = ( n3794 & n4207 ) | ( n3794 & n4208 ) | ( n4207 & n4208 ) ;
  assign n4210 = ( n4206 & ~n4207 ) | ( n4206 & n4209 ) | ( ~n4207 & n4209 ) ;
  assign n4211 = x212 | n3794 ;
  assign n4212 = ~x607 & x947 ;
  assign n4213 = ( x638 & x947 ) | ( x638 & n2007 ) | ( x947 & n2007 ) ;
  assign n4214 = ( n3794 & n4212 ) | ( n3794 & n4213 ) | ( n4212 & n4213 ) ;
  assign n4215 = ( n4211 & n4212 ) | ( n4211 & ~n4214 ) | ( n4212 & ~n4214 ) ;
  assign n4216 = x213 | n3794 ;
  assign n4217 = ( x639 & x947 ) | ( x639 & n2007 ) | ( x947 & n2007 ) ;
  assign n4218 = ~x622 & x947 ;
  assign n4219 = ( ~n3794 & n4217 ) | ( ~n3794 & n4218 ) | ( n4217 & n4218 ) ;
  assign n4220 = ( n4216 & ~n4217 ) | ( n4216 & n4219 ) | ( ~n4217 & n4219 ) ;
  assign n4221 = x214 | n3794 ;
  assign n4222 = ( x710 & x947 ) | ( x710 & n2007 ) | ( x947 & n2007 ) ;
  assign n4223 = ~x623 & x947 ;
  assign n4224 = ( ~n3794 & n4222 ) | ( ~n3794 & n4223 ) | ( n4222 & n4223 ) ;
  assign n4225 = ( n4221 & ~n4222 ) | ( n4221 & n4224 ) | ( ~n4222 & n4224 ) ;
  assign n4226 = x215 & ~n3794 ;
  assign n4227 = ( x681 & x947 ) | ( x681 & n2007 ) | ( x947 & n2007 ) ;
  assign n4228 = ~x642 & x947 ;
  assign n4229 = ( ~n3794 & n4227 ) | ( ~n3794 & n4228 ) | ( n4227 & n4228 ) ;
  assign n4230 = ( n4226 & n4227 ) | ( n4226 & ~n4229 ) | ( n4227 & ~n4229 ) ;
  assign n4231 = x216 & ~n3794 ;
  assign n4232 = ( x662 & x947 ) | ( x662 & n2007 ) | ( x947 & n2007 ) ;
  assign n4233 = ~x614 & x947 ;
  assign n4234 = ( ~n3794 & n4232 ) | ( ~n3794 & n4233 ) | ( n4232 & n4233 ) ;
  assign n4235 = ( n4231 & n4232 ) | ( n4231 & ~n4234 ) | ( n4232 & ~n4234 ) ;
  assign n4236 = x217 & ~n3794 ;
  assign n4237 = ~x695 & n3826 ;
  assign n4238 = x612 & n3775 ;
  assign n4239 = ( n3794 & n4237 ) | ( n3794 & ~n4238 ) | ( n4237 & ~n4238 ) ;
  assign n4240 = ( n4236 & ~n4237 ) | ( n4236 & n4239 ) | ( ~n4237 & n4239 ) ;
  assign n4241 = n2037 & n4159 ;
  assign n4242 = x218 | x332 ;
  assign n4243 = n2037 | n4242 ;
  assign n4244 = ( n4164 & n4242 ) | ( n4164 & n4243 ) | ( n4242 & n4243 ) ;
  assign n4245 = ~n4241 & n4244 ;
  assign n4246 = x219 & ~n3794 ;
  assign n4247 = ~x617 & x947 ;
  assign n4248 = ( x637 & x947 ) | ( x637 & n2007 ) | ( x947 & n2007 ) ;
  assign n4249 = ( n3794 & n4247 ) | ( n3794 & n4248 ) | ( n4247 & n4248 ) ;
  assign n4250 = ( n4246 & ~n4247 ) | ( n4246 & n4249 ) | ( ~n4247 & n4249 ) ;
  assign n4251 = n2105 & n4178 ;
  assign n4252 = x220 | x332 ;
  assign n4253 = n2105 | n4252 ;
  assign n4254 = ( n4181 & n4252 ) | ( n4181 & n4253 ) | ( n4252 & n4253 ) ;
  assign n4255 = ~n4251 & n4254 ;
  assign n4256 = x221 & ~n3794 ;
  assign n4257 = ~x616 & x947 ;
  assign n4258 = ( x661 & x947 ) | ( x661 & n2007 ) | ( x947 & n2007 ) ;
  assign n4259 = ( n3794 & n4257 ) | ( n3794 & n4258 ) | ( n4257 & n4258 ) ;
  assign n4260 = ( n4256 & ~n4257 ) | ( n4256 & n4259 ) | ( ~n4257 & n4259 ) ;
  assign n4261 = x222 | n3794 ;
  assign n4262 = x661 & n3826 ;
  assign n4263 = x616 & n3775 ;
  assign n4264 = ( n3794 & n4262 ) | ( n3794 & ~n4263 ) | ( n4262 & ~n4263 ) ;
  assign n4265 = ( n4261 & n4262 ) | ( n4261 & ~n4264 ) | ( n4262 & ~n4264 ) ;
  assign n4266 = x223 | n3794 ;
  assign n4267 = x642 & n3775 ;
  assign n4268 = x681 & n3826 ;
  assign n4269 = ( n3794 & n4267 ) | ( n3794 & ~n4268 ) | ( n4267 & ~n4268 ) ;
  assign n4270 = ( n4266 & n4267 ) | ( n4266 & ~n4269 ) | ( n4267 & ~n4269 ) ;
  assign n4271 = x224 | n3794 ;
  assign n4272 = x662 & n3826 ;
  assign n4273 = x614 & n3775 ;
  assign n4274 = ( n3794 & n4272 ) | ( n3794 & ~n4273 ) | ( n4272 & ~n4273 ) ;
  assign n4275 = ( n4271 & n4272 ) | ( n4271 & ~n4274 ) | ( n4272 & ~n4274 ) ;
  assign n4276 = ( x841 & ~n1279 ) | ( x841 & n2567 ) | ( ~n1279 & n2567 ) ;
  assign n4277 = n1423 | n4276 ;
  assign n4278 = ( ~n1277 & n1423 ) | ( ~n1277 & n4277 ) | ( n1423 & n4277 ) ;
  assign n4279 = n1953 | n2027 ;
  assign n4280 = ~n4278 & n4279 ;
  assign n4281 = ( n2512 & n4278 ) | ( n2512 & ~n4280 ) | ( n4278 & ~n4280 ) ;
  assign n4282 = n1496 & n4281 ;
  assign n4283 = x95 & x137 ;
  assign n4284 = ( x137 & n1309 ) | ( x137 & n4283 ) | ( n1309 & n4283 ) ;
  assign n4285 = x70 & x332 ;
  assign n4286 = x55 | n4285 ;
  assign n4287 = n1319 & ~n4279 ;
  assign n4288 = n4286 | n4287 ;
  assign n4289 = n4284 | n4288 ;
  assign n4290 = ~n1496 & n4289 ;
  assign n4291 = ( ~n1940 & n4282 ) | ( ~n1940 & n4290 ) | ( n4282 & n4290 ) ;
  assign n4292 = n2038 | n2583 ;
  assign n4293 = n1324 & ~n4292 ;
  assign n4294 = ( n1415 & ~n4292 ) | ( n1415 & n4293 ) | ( ~n4292 & n4293 ) ;
  assign n4295 = ~n1337 & n4294 ;
  assign n4296 = x228 & ~x231 ;
  assign n4297 = x228 & x231 ;
  assign n4298 = ( n4295 & ~n4296 ) | ( n4295 & n4297 ) | ( ~n4296 & n4297 ) ;
  assign n4299 = x47 | x72 ;
  assign n4300 = x36 & ~n2660 ;
  assign n4301 = ( ~n2955 & n4299 ) | ( ~n2955 & n4300 ) | ( n4299 & n4300 ) ;
  assign n4302 = n2955 | n4301 ;
  assign n4303 = n3099 | n4302 ;
  assign n4304 = n1362 | n4303 ;
  assign n4305 = n2573 & n4304 ;
  assign n4306 = ~x39 & x228 ;
  assign n4307 = x96 | x97 ;
  assign n4308 = x1091 & x1093 ;
  assign n4309 = n4307 & n4308 ;
  assign n4310 = ( n1429 & n4307 ) | ( n1429 & n4309 ) | ( n4307 & n4309 ) ;
  assign n4311 = n4306 | n4310 ;
  assign n4312 = ( n2141 & n4306 ) | ( n2141 & n4311 ) | ( n4306 & n4311 ) ;
  assign n4313 = x1091 & n3079 ;
  assign n4314 = n4312 | n4313 ;
  assign n4315 = ( n2618 & n4312 ) | ( n2618 & n4314 ) | ( n4312 & n4314 ) ;
  assign n4316 = x65 | x102 ;
  assign n4317 = n3601 & ~n4316 ;
  assign n4318 = ( ~n2807 & n2837 ) | ( ~n2807 & n3600 ) | ( n2837 & n3600 ) ;
  assign n4319 = ( ~n2837 & n4317 ) | ( ~n2837 & n4318 ) | ( n4317 & n4318 ) ;
  assign n4320 = ~x230 & x233 ;
  assign n4321 = ~x211 & x219 ;
  assign n4322 = x214 & x1153 ;
  assign n4323 = ~x214 & x1154 ;
  assign n4324 = ( n4321 & n4322 ) | ( n4321 & n4323 ) | ( n4322 & n4323 ) ;
  assign n4325 = x212 & ~x213 ;
  assign n4326 = n1553 & n4325 ;
  assign n4327 = x1155 & ~n2908 ;
  assign n4328 = x1154 & n2908 ;
  assign n4329 = ( x211 & n4327 ) | ( x211 & n4328 ) | ( n4327 & n4328 ) ;
  assign n4330 = x1155 & n2908 ;
  assign n4331 = x1156 & ~n2908 ;
  assign n4332 = ( ~x211 & n4330 ) | ( ~x211 & n4331 ) | ( n4330 & n4331 ) ;
  assign n4333 = ( ~x219 & n4329 ) | ( ~x219 & n4332 ) | ( n4329 & n4332 ) ;
  assign n4334 = ( n4324 & n4326 ) | ( n4324 & n4333 ) | ( n4326 & n4333 ) ;
  assign n4335 = x207 | x208 ;
  assign n4336 = x199 & ~x200 ;
  assign n4337 = ( x199 & n1553 ) | ( x199 & ~n4336 ) | ( n1553 & ~n4336 ) ;
  assign n4338 = n4335 & ~n4337 ;
  assign n4339 = ~x199 & x200 ;
  assign n4340 = x1156 & n4339 ;
  assign n4341 = x1157 & ~n2904 ;
  assign n4342 = n4340 | n4341 ;
  assign n4343 = x199 & x1155 ;
  assign n4344 = ( ~n2903 & n4342 ) | ( ~n2903 & n4343 ) | ( n4342 & n4343 ) ;
  assign n4345 = x208 | n4344 ;
  assign n4346 = x1155 & ~n2904 ;
  assign n4347 = x1154 & n4339 ;
  assign n4348 = n4346 | n4347 ;
  assign n4349 = x200 & x1155 ;
  assign n4350 = ~x200 & x1156 ;
  assign n4351 = ( ~x199 & n4349 ) | ( ~x199 & n4350 ) | ( n4349 & n4350 ) ;
  assign n4352 = x1154 & n4336 ;
  assign n4353 = ( ~x209 & n4351 ) | ( ~x209 & n4352 ) | ( n4351 & n4352 ) ;
  assign n4354 = ( x207 & ~x209 ) | ( x207 & n4353 ) | ( ~x209 & n4353 ) ;
  assign n4355 = x199 & x1153 ;
  assign n4356 = ( n2903 & n4348 ) | ( n2903 & ~n4355 ) | ( n4348 & ~n4355 ) ;
  assign n4357 = ( n4348 & n4354 ) | ( n4348 & ~n4356 ) | ( n4354 & ~n4356 ) ;
  assign n4358 = n4345 & n4357 ;
  assign n4359 = ~x1142 & n2905 ;
  assign n4360 = x200 | n2903 ;
  assign n4361 = x1144 | n4360 ;
  assign n4362 = ~x1143 & n4360 ;
  assign n4363 = ( n2905 & n4361 ) | ( n2905 & ~n4362 ) | ( n4361 & ~n4362 ) ;
  assign n4364 = ~n4359 & n4363 ;
  assign n4365 = x209 & n4364 ;
  assign n4366 = ( n4338 & n4358 ) | ( n4338 & n4365 ) | ( n4358 & n4365 ) ;
  assign n4367 = n4334 | n4366 ;
  assign n4368 = x211 & x219 ;
  assign n4369 = x212 | x214 ;
  assign n4370 = ( n1553 & n4368 ) | ( n1553 & ~n4369 ) | ( n4368 & ~n4369 ) ;
  assign n4371 = n1553 & ~n4370 ;
  assign n4372 = ~x1142 & n2909 ;
  assign n4373 = x211 | n2908 ;
  assign n4374 = ~x1143 & n4373 ;
  assign n4375 = x1144 | n4373 ;
  assign n4376 = ( n2909 & ~n4374 ) | ( n2909 & n4375 ) | ( ~n4374 & n4375 ) ;
  assign n4377 = ~n4372 & n4376 ;
  assign n4378 = x213 & n4377 ;
  assign n4379 = x1157 & ~n2908 ;
  assign n4380 = x1156 & n2908 ;
  assign n4381 = ( ~n2907 & n4379 ) | ( ~n2907 & n4380 ) | ( n4379 & n4380 ) ;
  assign n4382 = x212 | x213 ;
  assign n4383 = x219 & x1155 ;
  assign n4384 = ~n2908 & n4383 ;
  assign n4385 = ( x211 & n4330 ) | ( x211 & n4331 ) | ( n4330 & n4331 ) ;
  assign n4386 = n4384 | n4385 ;
  assign n4387 = ( n4381 & ~n4382 ) | ( n4381 & n4386 ) | ( ~n4382 & n4386 ) ;
  assign n4388 = ( n4371 & n4378 ) | ( n4371 & n4387 ) | ( n4378 & n4387 ) ;
  assign n4389 = x230 & ~n4388 ;
  assign n4390 = n4367 | n4389 ;
  assign n4391 = ( n4320 & ~n4367 ) | ( n4320 & n4390 ) | ( ~n4367 & n4390 ) ;
  assign n4392 = x230 | x234 ;
  assign n4393 = x213 & n4371 ;
  assign n4394 = x219 & x1154 ;
  assign n4395 = ( n4333 & n4393 ) | ( n4333 & n4394 ) | ( n4393 & n4394 ) ;
  assign n4396 = ~x209 & x230 ;
  assign n4397 = ( x230 & ~n4335 ) | ( x230 & n4396 ) | ( ~n4335 & n4396 ) ;
  assign n4398 = n2903 & ~n4348 ;
  assign n4399 = n2903 | n4351 ;
  assign n4400 = ( n4352 & ~n4398 ) | ( n4352 & n4399 ) | ( ~n4398 & n4399 ) ;
  assign n4401 = ~n1553 & n4400 ;
  assign n4402 = ( x230 & n4397 ) | ( x230 & ~n4401 ) | ( n4397 & ~n4401 ) ;
  assign n4403 = ~n4395 & n4402 ;
  assign n4404 = x209 & n4338 ;
  assign n4405 = n4393 | n4404 ;
  assign n4406 = ( x230 & n4338 ) | ( x230 & n4371 ) | ( n4338 & n4371 ) ;
  assign n4407 = ~n4405 & n4406 ;
  assign n4408 = x1152 & n2911 ;
  assign n4409 = x1154 | n2988 ;
  assign n4410 = ( ~x1153 & n2986 ) | ( ~x1153 & n2987 ) | ( n2986 & n2987 ) ;
  assign n4411 = ( n2911 & ~n4408 ) | ( n2911 & n4410 ) | ( ~n4408 & n4410 ) ;
  assign n4412 = ( n4408 & n4409 ) | ( n4408 & ~n4411 ) | ( n4409 & ~n4411 ) ;
  assign n4413 = n4407 & n4412 ;
  assign n4414 = ( n4392 & ~n4403 ) | ( n4392 & n4413 ) | ( ~n4403 & n4413 ) ;
  assign n4415 = x230 | x235 ;
  assign n4416 = n2903 & n4351 ;
  assign n4417 = ( x209 & n4344 ) | ( x209 & n4416 ) | ( n4344 & n4416 ) ;
  assign n4418 = n4355 & ~n4360 ;
  assign n4419 = ~x200 & x1154 ;
  assign n4420 = x200 & x1153 ;
  assign n4421 = ( ~x199 & n4419 ) | ( ~x199 & n4420 ) | ( n4419 & n4420 ) ;
  assign n4422 = n2903 & ~n4421 ;
  assign n4423 = ( n4348 & n4398 ) | ( n4348 & ~n4422 ) | ( n4398 & ~n4422 ) ;
  assign n4424 = ( ~x209 & n4418 ) | ( ~x209 & n4423 ) | ( n4418 & n4423 ) ;
  assign n4425 = ( n4338 & n4417 ) | ( n4338 & n4424 ) | ( n4417 & n4424 ) ;
  assign n4426 = ( ~x230 & n4415 ) | ( ~x230 & n4425 ) | ( n4415 & n4425 ) ;
  assign n4427 = ( x213 & n4381 ) | ( x213 & n4386 ) | ( n4381 & n4386 ) ;
  assign n4428 = ( ~n2907 & n4327 ) | ( ~n2907 & n4328 ) | ( n4327 & n4328 ) ;
  assign n4429 = ( x211 & x1153 ) | ( x211 & ~n2908 ) | ( x1153 & ~n2908 ) ;
  assign n4430 = x211 & x1154 ;
  assign n4431 = ~n2908 & n4430 ;
  assign n4432 = ( n2909 & n4429 ) | ( n2909 & n4431 ) | ( n4429 & n4431 ) ;
  assign n4433 = ( ~x213 & n4428 ) | ( ~x213 & n4432 ) | ( n4428 & n4432 ) ;
  assign n4434 = ( n4371 & n4427 ) | ( n4371 & n4433 ) | ( n4427 & n4433 ) ;
  assign n4435 = ( n4415 & n4426 ) | ( n4415 & n4434 ) | ( n4426 & n4434 ) ;
  assign n4436 = ~x1143 & n2911 ;
  assign n4437 = x1145 | n2988 ;
  assign n4438 = ( ~x1144 & n2986 ) | ( ~x1144 & n2987 ) | ( n2986 & n2987 ) ;
  assign n4439 = ( n2911 & n4437 ) | ( n2911 & ~n4438 ) | ( n4437 & ~n4438 ) ;
  assign n4440 = ( n4405 & n4436 ) | ( n4405 & ~n4439 ) | ( n4436 & ~n4439 ) ;
  assign n4441 = x230 | x237 ;
  assign n4442 = n2908 & n4394 ;
  assign n4443 = x213 | n4442 ;
  assign n4444 = x211 & ~x1157 ;
  assign n4445 = x219 | x1158 ;
  assign n4446 = x219 & ~x1156 ;
  assign n4447 = ( x211 & n4445 ) | ( x211 & ~n4446 ) | ( n4445 & ~n4446 ) ;
  assign n4448 = ( x212 & ~n4444 ) | ( x212 & n4447 ) | ( ~n4444 & n4447 ) ;
  assign n4449 = ( ~x212 & n4443 ) | ( ~x212 & n4448 ) | ( n4443 & n4448 ) ;
  assign n4450 = n1553 & ~n4449 ;
  assign n4451 = ( x212 & n4381 ) | ( x212 & n4386 ) | ( n4381 & n4386 ) ;
  assign n4452 = n4450 & ~n4451 ;
  assign n4453 = x1156 & n4336 ;
  assign n4454 = ~x200 & x1158 ;
  assign n4455 = x200 & x1157 ;
  assign n4456 = ( ~x199 & n4454 ) | ( ~x199 & n4455 ) | ( n4454 & n4455 ) ;
  assign n4457 = ( ~x208 & n4453 ) | ( ~x208 & n4456 ) | ( n4453 & n4456 ) ;
  assign n4458 = ( x209 & n1553 ) | ( x209 & ~n4457 ) | ( n1553 & ~n4457 ) ;
  assign n4459 = n4457 | n4458 ;
  assign n4460 = ( n2903 & n4351 ) | ( n2903 & n4352 ) | ( n4351 & n4352 ) ;
  assign n4461 = ( x208 & n4344 ) | ( x208 & n4460 ) | ( n4344 & n4460 ) ;
  assign n4462 = n4459 | n4461 ;
  assign n4463 = ( n4406 & ~n4441 ) | ( n4406 & n4462 ) | ( ~n4441 & n4462 ) ;
  assign n4464 = ( n4441 & n4452 ) | ( n4441 & ~n4463 ) | ( n4452 & ~n4463 ) ;
  assign n4465 = ( n4440 & n4441 ) | ( n4440 & n4464 ) | ( n4441 & n4464 ) ;
  assign n4466 = x230 | x238 ;
  assign n4467 = ~x1152 & n4373 ;
  assign n4468 = x1151 & n2909 ;
  assign n4469 = n2908 | n4429 ;
  assign n4470 = ( ~n2909 & n4468 ) | ( ~n2909 & n4469 ) | ( n4468 & n4469 ) ;
  assign n4471 = ( ~n4467 & n4468 ) | ( ~n4467 & n4470 ) | ( n4468 & n4470 ) ;
  assign n4472 = ~x213 & n4471 ;
  assign n4473 = x1153 & n2909 ;
  assign n4474 = ( n4428 & ~n4431 ) | ( n4428 & n4473 ) | ( ~n4431 & n4473 ) ;
  assign n4475 = ( x213 & n4431 ) | ( x213 & n4474 ) | ( n4431 & n4474 ) ;
  assign n4476 = ( n4371 & n4472 ) | ( n4371 & n4475 ) | ( n4472 & n4475 ) ;
  assign n4477 = x230 & ~n4476 ;
  assign n4478 = ~x1152 & n4360 ;
  assign n4479 = x1151 & n2905 ;
  assign n4480 = x1153 | n4360 ;
  assign n4481 = ( ~n2905 & n4479 ) | ( ~n2905 & n4480 ) | ( n4479 & n4480 ) ;
  assign n4482 = ( ~n4478 & n4479 ) | ( ~n4478 & n4481 ) | ( n4479 & n4481 ) ;
  assign n4483 = ~x209 & n4482 ;
  assign n4484 = x230 & n4338 ;
  assign n4485 = ( x209 & n4355 ) | ( x209 & n4423 ) | ( n4355 & n4423 ) ;
  assign n4486 = ( n4483 & n4484 ) | ( n4483 & n4485 ) | ( n4484 & n4485 ) ;
  assign n4487 = ( n4466 & ~n4477 ) | ( n4466 & n4486 ) | ( ~n4477 & n4486 ) ;
  assign n4488 = x230 | x239 ;
  assign n4489 = x207 & ~x208 ;
  assign n4490 = ~n1553 & n4489 ;
  assign n4491 = ( x209 & n4453 ) | ( x209 & n4456 ) | ( n4453 & n4456 ) ;
  assign n4492 = ( n4353 & n4490 ) | ( n4353 & n4491 ) | ( n4490 & n4491 ) ;
  assign n4493 = ( ~x230 & n4488 ) | ( ~x230 & n4492 ) | ( n4488 & n4492 ) ;
  assign n4494 = ( ~x213 & n4333 ) | ( ~x213 & n4394 ) | ( n4333 & n4394 ) ;
  assign n4495 = ~x212 & n4371 ;
  assign n4496 = x213 & ~n4444 ;
  assign n4497 = n4447 & n4496 ;
  assign n4498 = ( n4494 & n4495 ) | ( n4494 & n4497 ) | ( n4495 & n4497 ) ;
  assign n4499 = ( n4488 & n4493 ) | ( n4488 & n4498 ) | ( n4493 & n4498 ) ;
  assign n4500 = ~n2911 & n2988 ;
  assign n4501 = x1146 & n4500 ;
  assign n4502 = x1145 & n2911 ;
  assign n4503 = x1147 & ~n2988 ;
  assign n4504 = n4502 | n4503 ;
  assign n4505 = ( n4407 & n4501 ) | ( n4407 & n4504 ) | ( n4501 & n4504 ) ;
  assign n4506 = ( x230 & n4393 ) | ( x230 & n4404 ) | ( n4393 & n4404 ) ;
  assign n4507 = x1147 & n2911 ;
  assign n4508 = x1149 & ~n2988 ;
  assign n4509 = n4507 | n4508 ;
  assign n4510 = x1148 & n4500 ;
  assign n4511 = ( n4506 & n4509 ) | ( n4506 & n4510 ) | ( n4509 & n4510 ) ;
  assign n4512 = ~x230 & x240 ;
  assign n4513 = n4511 | n4512 ;
  assign n4514 = n4505 | n4513 ;
  assign n4515 = n4404 & ~n4482 ;
  assign n4516 = ~x1149 & n2911 ;
  assign n4517 = x1151 | n2988 ;
  assign n4518 = ( ~x1150 & n2986 ) | ( ~x1150 & n2987 ) | ( n2986 & n2987 ) ;
  assign n4519 = ( n2911 & n4517 ) | ( n2911 & ~n4518 ) | ( n4517 & ~n4518 ) ;
  assign n4520 = ( n4404 & ~n4516 ) | ( n4404 & n4519 ) | ( ~n4516 & n4519 ) ;
  assign n4521 = ( n4393 & ~n4515 ) | ( n4393 & n4520 ) | ( ~n4515 & n4520 ) ;
  assign n4522 = n4393 & ~n4471 ;
  assign n4523 = ( ~n4406 & n4521 ) | ( ~n4406 & n4522 ) | ( n4521 & n4522 ) ;
  assign n4524 = ~x230 & x241 ;
  assign n4525 = ( n4521 & ~n4523 ) | ( n4521 & n4524 ) | ( ~n4523 & n4524 ) ;
  assign n4526 = ( ~x1145 & n2986 ) | ( ~x1145 & n2987 ) | ( n2986 & n2987 ) ;
  assign n4527 = x1144 & n2911 ;
  assign n4528 = x1146 | n2988 ;
  assign n4529 = ( ~n2911 & n4527 ) | ( ~n2911 & n4528 ) | ( n4527 & n4528 ) ;
  assign n4530 = ( ~n4526 & n4527 ) | ( ~n4526 & n4529 ) | ( n4527 & n4529 ) ;
  assign n4531 = n4405 & n4530 ;
  assign n4532 = ~x209 & n4364 ;
  assign n4533 = n4484 & n4532 ;
  assign n4534 = ( x230 & n4531 ) | ( x230 & n4533 ) | ( n4531 & n4533 ) ;
  assign n4535 = x230 | x242 ;
  assign n4536 = ( ~x230 & n4371 ) | ( ~x230 & n4377 ) | ( n4371 & n4377 ) ;
  assign n4537 = ( x230 & n4393 ) | ( x230 & ~n4536 ) | ( n4393 & ~n4536 ) ;
  assign n4538 = ( n4534 & n4535 ) | ( n4534 & ~n4537 ) | ( n4535 & ~n4537 ) ;
  assign n4539 = ( x83 & n2061 ) | ( x83 & ~n3062 ) | ( n2061 & ~n3062 ) ;
  assign n4540 = ( x314 & n3217 ) | ( x314 & n4539 ) | ( n3217 & n4539 ) ;
  assign n4541 = x802 & n4540 ;
  assign n4542 = x276 & n4541 ;
  assign n4543 = x271 & n4542 ;
  assign n4544 = x273 & n4543 ;
  assign n4545 = x283 & n4544 ;
  assign n4546 = x272 & n4545 ;
  assign n4547 = x275 & n4546 ;
  assign n4548 = x268 & n4547 ;
  assign n4549 = x253 & n4548 ;
  assign n4550 = x254 & n4549 ;
  assign n4551 = x267 & n4550 ;
  assign n4552 = ~x263 & n4551 ;
  assign n4553 = x243 & n4552 ;
  assign n4554 = n3062 & ~n3091 ;
  assign n4555 = ~x211 & x1155 ;
  assign n4556 = x211 & x1156 ;
  assign n4557 = ( ~x219 & n4555 ) | ( ~x219 & n4556 ) | ( n4555 & n4556 ) ;
  assign n4558 = n1553 & ~n4557 ;
  assign n4559 = n4340 | n4346 ;
  assign n4560 = n1553 | n4559 ;
  assign n4561 = x230 | x1091 ;
  assign n4562 = ( n4558 & ~n4560 ) | ( n4558 & n4561 ) | ( ~n4560 & n4561 ) ;
  assign n4563 = ~x1157 & n4562 ;
  assign n4564 = ( ~n4554 & n4562 ) | ( ~n4554 & n4563 ) | ( n4562 & n4563 ) ;
  assign n4565 = ( x243 & n4552 ) | ( x243 & ~n4561 ) | ( n4552 & ~n4561 ) ;
  assign n4566 = ( ~n4553 & n4564 ) | ( ~n4553 & n4565 ) | ( n4564 & n4565 ) ;
  assign n4567 = ~n4436 & n4439 ;
  assign n4568 = n4407 & n4567 ;
  assign n4569 = ~x230 & x244 ;
  assign n4570 = ( n4501 & n4504 ) | ( n4501 & n4506 ) | ( n4504 & n4506 ) ;
  assign n4571 = n4569 | n4570 ;
  assign n4572 = n4568 | n4571 ;
  assign n4573 = n4407 & n4530 ;
  assign n4574 = ~x230 & x245 ;
  assign n4575 = x1146 & n2911 ;
  assign n4576 = ( ~x1147 & n2986 ) | ( ~x1147 & n2987 ) | ( n2986 & n2987 ) ;
  assign n4577 = x1148 | n2988 ;
  assign n4578 = ( ~n2911 & n4575 ) | ( ~n2911 & n4577 ) | ( n4575 & n4577 ) ;
  assign n4579 = ( n4575 & ~n4576 ) | ( n4575 & n4578 ) | ( ~n4576 & n4578 ) ;
  assign n4580 = n4506 & n4579 ;
  assign n4581 = ( ~n4573 & n4574 ) | ( ~n4573 & n4580 ) | ( n4574 & n4580 ) ;
  assign n4582 = n4573 | n4581 ;
  assign n4583 = n4407 & n4579 ;
  assign n4584 = ~x230 & x246 ;
  assign n4585 = x1148 & n2911 ;
  assign n4586 = ( ~x1149 & n2986 ) | ( ~x1149 & n2987 ) | ( n2986 & n2987 ) ;
  assign n4587 = x1150 | n2988 ;
  assign n4588 = ( ~n2911 & n4585 ) | ( ~n2911 & n4587 ) | ( n4585 & n4587 ) ;
  assign n4589 = ( n4585 & ~n4586 ) | ( n4585 & n4588 ) | ( ~n4586 & n4588 ) ;
  assign n4590 = n4506 & n4589 ;
  assign n4591 = ( ~n4583 & n4584 ) | ( ~n4583 & n4590 ) | ( n4584 & n4590 ) ;
  assign n4592 = n4583 | n4591 ;
  assign n4593 = ~x230 & x247 ;
  assign n4594 = ( n4506 & n4516 ) | ( n4506 & n4519 ) | ( n4516 & n4519 ) ;
  assign n4595 = ( ~n4516 & n4593 ) | ( ~n4516 & n4594 ) | ( n4593 & n4594 ) ;
  assign n4596 = ( n4407 & n4509 ) | ( n4407 & n4510 ) | ( n4509 & n4510 ) ;
  assign n4597 = n4595 | n4596 ;
  assign n4598 = n4407 & n4589 ;
  assign n4599 = ~x230 & x248 ;
  assign n4600 = ( ~x1151 & n2986 ) | ( ~x1151 & n2987 ) | ( n2986 & n2987 ) ;
  assign n4601 = x1150 & n2911 ;
  assign n4602 = x1152 | n2988 ;
  assign n4603 = ( ~n2911 & n4601 ) | ( ~n2911 & n4602 ) | ( n4601 & n4602 ) ;
  assign n4604 = ( ~n4600 & n4601 ) | ( ~n4600 & n4603 ) | ( n4601 & n4603 ) ;
  assign n4605 = n4506 & n4604 ;
  assign n4606 = ( ~n4598 & n4599 ) | ( ~n4598 & n4605 ) | ( n4599 & n4605 ) ;
  assign n4607 = n4598 | n4606 ;
  assign n4608 = n4407 & n4604 ;
  assign n4609 = ~x230 & x249 ;
  assign n4610 = n4506 | n4609 ;
  assign n4611 = ( n4412 & n4609 ) | ( n4412 & n4610 ) | ( n4609 & n4610 ) ;
  assign n4612 = n4608 | n4611 ;
  assign n4613 = x250 | n2462 ;
  assign n4614 = n1319 | n2881 ;
  assign n4615 = ~n4613 & n4614 ;
  assign n4616 = ~n1337 & n4615 ;
  assign n4617 = x200 & ~x476 ;
  assign n4618 = ~x200 & x897 ;
  assign n4619 = ( ~x199 & n4617 ) | ( ~x199 & n4618 ) | ( n4617 & n4618 ) ;
  assign n4620 = x251 & ~n4619 ;
  assign n4621 = ~x200 & x1053 ;
  assign n4622 = x200 & x1039 ;
  assign n4623 = ( ~x199 & n4621 ) | ( ~x199 & n4622 ) | ( n4621 & n4622 ) ;
  assign n4624 = n4619 & ~n4623 ;
  assign n4625 = ( n4619 & n4620 ) | ( n4619 & ~n4624 ) | ( n4620 & ~n4624 ) ;
  assign n4626 = ~n1337 & n2015 ;
  assign n4627 = x252 & x1092 ;
  assign n4628 = x1093 & n2180 ;
  assign n4629 = n4627 & ~n4628 ;
  assign n4630 = n4626 | n4629 ;
  assign n4631 = ( x253 & n4548 ) | ( x253 & ~n4561 ) | ( n4548 & ~n4561 ) ;
  assign n4632 = x1153 & n4554 ;
  assign n4633 = ( x1152 & n3089 ) | ( x1152 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4634 = x1151 & ~n3091 ;
  assign n4635 = ( ~n3062 & n4633 ) | ( ~n3062 & n4634 ) | ( n4633 & n4634 ) ;
  assign n4636 = ( n4561 & n4632 ) | ( n4561 & n4635 ) | ( n4632 & n4635 ) ;
  assign n4637 = ( ~n4549 & n4631 ) | ( ~n4549 & n4636 ) | ( n4631 & n4636 ) ;
  assign n4638 = ~x254 & n4549 ;
  assign n4639 = ( x254 & ~n4549 ) | ( x254 & n4561 ) | ( ~n4549 & n4561 ) ;
  assign n4640 = x1153 & n3092 ;
  assign n4641 = x1154 & n4554 ;
  assign n4642 = x1152 & ~n3091 ;
  assign n4643 = ( n3060 & n3061 ) | ( n3060 & n4561 ) | ( n3061 & n4561 ) ;
  assign n4644 = ( n4561 & ~n4642 ) | ( n4561 & n4643 ) | ( ~n4642 & n4643 ) ;
  assign n4645 = ( n4640 & ~n4641 ) | ( n4640 & n4644 ) | ( ~n4641 & n4644 ) ;
  assign n4646 = ~n4640 & n4645 ;
  assign n4647 = ( n4638 & n4639 ) | ( n4638 & ~n4646 ) | ( n4639 & ~n4646 ) ;
  assign n4648 = x255 & ~n4619 ;
  assign n4649 = ~x200 & x1049 ;
  assign n4650 = x200 & x1036 ;
  assign n4651 = ( ~x199 & n4649 ) | ( ~x199 & n4650 ) | ( n4649 & n4650 ) ;
  assign n4652 = n4619 & ~n4651 ;
  assign n4653 = ( n4619 & n4648 ) | ( n4619 & ~n4652 ) | ( n4648 & ~n4652 ) ;
  assign n4654 = ~x200 & x1048 ;
  assign n4655 = x200 & x1070 ;
  assign n4656 = ( ~x199 & n4654 ) | ( ~x199 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4657 = n4619 & ~n4656 ;
  assign n4658 = x256 & ~n4619 ;
  assign n4659 = ( n4619 & ~n4657 ) | ( n4619 & n4658 ) | ( ~n4657 & n4658 ) ;
  assign n4660 = x257 & ~n4619 ;
  assign n4661 = ~x200 & x1084 ;
  assign n4662 = x200 & x1065 ;
  assign n4663 = ( ~x199 & n4661 ) | ( ~x199 & n4662 ) | ( n4661 & n4662 ) ;
  assign n4664 = n4619 & ~n4663 ;
  assign n4665 = ( n4619 & n4660 ) | ( n4619 & ~n4664 ) | ( n4660 & ~n4664 ) ;
  assign n4666 = x258 & ~n4619 ;
  assign n4667 = x200 & x1062 ;
  assign n4668 = ~x200 & x1072 ;
  assign n4669 = ( ~x199 & n4667 ) | ( ~x199 & n4668 ) | ( n4667 & n4668 ) ;
  assign n4670 = n4619 & ~n4669 ;
  assign n4671 = ( n4619 & n4666 ) | ( n4619 & ~n4670 ) | ( n4666 & ~n4670 ) ;
  assign n4672 = x259 & ~n4619 ;
  assign n4673 = x200 & x1069 ;
  assign n4674 = ~x200 & x1059 ;
  assign n4675 = ( ~x199 & n4673 ) | ( ~x199 & n4674 ) | ( n4673 & n4674 ) ;
  assign n4676 = n4619 & ~n4675 ;
  assign n4677 = ( n4619 & n4672 ) | ( n4619 & ~n4676 ) | ( n4672 & ~n4676 ) ;
  assign n4678 = x260 & ~n4619 ;
  assign n4679 = ~x200 & x1044 ;
  assign n4680 = x200 & x1067 ;
  assign n4681 = ( ~x199 & n4679 ) | ( ~x199 & n4680 ) | ( n4679 & n4680 ) ;
  assign n4682 = n4619 & ~n4681 ;
  assign n4683 = ( n4619 & n4678 ) | ( n4619 & ~n4682 ) | ( n4678 & ~n4682 ) ;
  assign n4684 = x261 & ~n4619 ;
  assign n4685 = ~x200 & x1037 ;
  assign n4686 = x200 & x1040 ;
  assign n4687 = ( ~x199 & n4685 ) | ( ~x199 & n4686 ) | ( n4685 & n4686 ) ;
  assign n4688 = n4619 & ~n4687 ;
  assign n4689 = ( n4619 & n4684 ) | ( n4619 & ~n4688 ) | ( n4684 & ~n4688 ) ;
  assign n4690 = ~x123 & x228 ;
  assign n4691 = ~x228 & x1093 ;
  assign n4692 = n4690 | n4691 ;
  assign n4693 = x262 | n4692 ;
  assign n4694 = ( x1142 & ~n2906 ) | ( x1142 & n2910 ) | ( ~n2906 & n2910 ) ;
  assign n4695 = ( n4338 & n4371 ) | ( n4338 & n4692 ) | ( n4371 & n4692 ) ;
  assign n4696 = n4694 & ~n4695 ;
  assign n4697 = ( n4693 & ~n4694 ) | ( n4693 & n4696 ) | ( ~n4694 & n4696 ) ;
  assign n4698 = ( x263 & ~n4551 ) | ( x263 & n4561 ) | ( ~n4551 & n4561 ) ;
  assign n4699 = ( ~x1155 & n3089 ) | ( ~x1155 & n4383 ) | ( n3089 & n4383 ) ;
  assign n4700 = x219 | x1154 ;
  assign n4701 = ( x211 & ~n4446 ) | ( x211 & n4700 ) | ( ~n4446 & n4700 ) ;
  assign n4702 = n1553 & n4701 ;
  assign n4703 = ( ~x199 & n4349 ) | ( ~x199 & n4419 ) | ( n4349 & n4419 ) ;
  assign n4704 = ( ~n1553 & n4453 ) | ( ~n1553 & n4703 ) | ( n4453 & n4703 ) ;
  assign n4705 = ( n4561 & n4702 ) | ( n4561 & n4704 ) | ( n4702 & n4704 ) ;
  assign n4706 = ~n4699 & n4705 ;
  assign n4707 = ( n4552 & n4698 ) | ( n4552 & ~n4706 ) | ( n4698 & ~n4706 ) ;
  assign n4708 = x1142 & n3092 ;
  assign n4709 = ( x1143 & n3060 ) | ( x1143 & n3061 ) | ( n3060 & n3061 ) ;
  assign n4710 = x1141 & ~n3062 ;
  assign n4711 = ( ~n3091 & n4709 ) | ( ~n3091 & n4710 ) | ( n4709 & n4710 ) ;
  assign n4712 = ( n4561 & n4708 ) | ( n4561 & n4711 ) | ( n4708 & n4711 ) ;
  assign n4713 = x796 & n4540 ;
  assign n4714 = x264 | n4540 ;
  assign n4715 = ( n4561 & ~n4713 ) | ( n4561 & n4714 ) | ( ~n4713 & n4714 ) ;
  assign n4716 = ~n4712 & n4715 ;
  assign n4717 = x1144 & ~n3091 ;
  assign n4718 = ( ~x1143 & n3089 ) | ( ~x1143 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4719 = ( n3062 & ~n4717 ) | ( n3062 & n4718 ) | ( ~n4717 & n4718 ) ;
  assign n4720 = x1142 | n3214 ;
  assign n4721 = ( n4561 & n4719 ) | ( n4561 & ~n4720 ) | ( n4719 & ~n4720 ) ;
  assign n4722 = x265 & ~n4540 ;
  assign n4723 = ~x819 & n4540 ;
  assign n4724 = ( ~n4561 & n4722 ) | ( ~n4561 & n4723 ) | ( n4722 & n4723 ) ;
  assign n4725 = n4721 | n4724 ;
  assign n4726 = ( x1136 & n3060 ) | ( x1136 & n3061 ) | ( n3060 & n3061 ) ;
  assign n4727 = x1134 & ~n3062 ;
  assign n4728 = ( ~n3091 & n4726 ) | ( ~n3091 & n4727 ) | ( n4726 & n4727 ) ;
  assign n4729 = x1135 & n3092 ;
  assign n4730 = ( n4561 & n4728 ) | ( n4561 & n4729 ) | ( n4728 & n4729 ) ;
  assign n4731 = x948 & n4540 ;
  assign n4732 = x266 & ~n4540 ;
  assign n4733 = ( ~n4561 & n4731 ) | ( ~n4561 & n4732 ) | ( n4731 & n4732 ) ;
  assign n4734 = n4730 | n4733 ;
  assign n4735 = ~x267 & n4550 ;
  assign n4736 = x1153 & ~n3214 ;
  assign n4737 = ( n1553 & ~n3090 ) | ( n1553 & n4343 ) | ( ~n3090 & n4343 ) ;
  assign n4738 = n4347 | n4737 ;
  assign n4739 = n4383 | n4430 ;
  assign n4740 = ~n4368 & n4739 ;
  assign n4741 = n1553 & ~n4740 ;
  assign n4742 = ( n4561 & ~n4738 ) | ( n4561 & n4741 ) | ( ~n4738 & n4741 ) ;
  assign n4743 = ~n4736 & n4742 ;
  assign n4744 = ( x267 & ~n4550 ) | ( x267 & n4561 ) | ( ~n4550 & n4561 ) ;
  assign n4745 = ( n4735 & ~n4743 ) | ( n4735 & n4744 ) | ( ~n4743 & n4744 ) ;
  assign n4746 = x1150 & n4561 ;
  assign n4747 = ( n3214 & n4561 ) | ( n3214 & n4746 ) | ( n4561 & n4746 ) ;
  assign n4748 = ( ~x1151 & n3089 ) | ( ~x1151 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4749 = ( n3062 & ~n4642 ) | ( n3062 & n4748 ) | ( ~n4642 & n4748 ) ;
  assign n4750 = n4747 & ~n4749 ;
  assign n4751 = ( x268 & n4547 ) | ( x268 & ~n4561 ) | ( n4547 & ~n4561 ) ;
  assign n4752 = ( ~n4548 & n4750 ) | ( ~n4548 & n4751 ) | ( n4750 & n4751 ) ;
  assign n4753 = x1136 & ~n3091 ;
  assign n4754 = ( x1137 & n3089 ) | ( x1137 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4755 = ( ~n3062 & n4753 ) | ( ~n3062 & n4754 ) | ( n4753 & n4754 ) ;
  assign n4756 = x1138 & n4554 ;
  assign n4757 = ( n4561 & n4755 ) | ( n4561 & n4756 ) | ( n4755 & n4756 ) ;
  assign n4758 = x269 | n4540 ;
  assign n4759 = x817 & n4540 ;
  assign n4760 = ( n4561 & n4758 ) | ( n4561 & ~n4759 ) | ( n4758 & ~n4759 ) ;
  assign n4761 = ~n4757 & n4760 ;
  assign n4762 = x1139 & ~n3091 ;
  assign n4763 = ( x1140 & n3089 ) | ( x1140 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4764 = ( ~n3062 & n4762 ) | ( ~n3062 & n4763 ) | ( n4762 & n4763 ) ;
  assign n4765 = x1141 & n4554 ;
  assign n4766 = ( n4561 & n4764 ) | ( n4561 & n4765 ) | ( n4764 & n4765 ) ;
  assign n4767 = x270 | n4540 ;
  assign n4768 = x805 & n4540 ;
  assign n4769 = ( n4561 & n4767 ) | ( n4561 & ~n4768 ) | ( n4767 & ~n4768 ) ;
  assign n4770 = ~n4766 & n4769 ;
  assign n4771 = x1146 & n3092 ;
  assign n4772 = ( x1147 & n3060 ) | ( x1147 & n3061 ) | ( n3060 & n3061 ) ;
  assign n4773 = x1145 & ~n3062 ;
  assign n4774 = ( ~n3091 & n4772 ) | ( ~n3091 & n4773 ) | ( n4772 & n4773 ) ;
  assign n4775 = ( n4561 & n4771 ) | ( n4561 & n4774 ) | ( n4771 & n4774 ) ;
  assign n4776 = ( x271 & n4542 ) | ( x271 & ~n4561 ) | ( n4542 & ~n4561 ) ;
  assign n4777 = ( ~n4543 & n4775 ) | ( ~n4543 & n4776 ) | ( n4775 & n4776 ) ;
  assign n4778 = x1148 & ~n3091 ;
  assign n4779 = ( x1149 & n3089 ) | ( x1149 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4780 = ( ~n3062 & n4778 ) | ( ~n3062 & n4779 ) | ( n4778 & n4779 ) ;
  assign n4781 = x1150 & n4554 ;
  assign n4782 = ( n4561 & n4780 ) | ( n4561 & n4781 ) | ( n4780 & n4781 ) ;
  assign n4783 = ( x272 & n4545 ) | ( x272 & ~n4561 ) | ( n4545 & ~n4561 ) ;
  assign n4784 = ( ~n4546 & n4782 ) | ( ~n4546 & n4783 ) | ( n4782 & n4783 ) ;
  assign n4785 = n3062 & ~n4778 ;
  assign n4786 = x1146 | n3091 ;
  assign n4787 = ( ~x1147 & n3089 ) | ( ~x1147 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4788 = ( n3062 & n4786 ) | ( n3062 & ~n4787 ) | ( n4786 & ~n4787 ) ;
  assign n4789 = ( n4561 & n4785 ) | ( n4561 & ~n4788 ) | ( n4785 & ~n4788 ) ;
  assign n4790 = x273 & ~n4543 ;
  assign n4791 = ( ~x273 & n4543 ) | ( ~x273 & n4561 ) | ( n4543 & n4561 ) ;
  assign n4792 = ( ~n4789 & n4790 ) | ( ~n4789 & n4791 ) | ( n4790 & n4791 ) ;
  assign n4793 = x1145 & n4554 ;
  assign n4794 = x274 & ~n4540 ;
  assign n4795 = ~x659 & n4540 ;
  assign n4796 = ( ~n4561 & n4794 ) | ( ~n4561 & n4795 ) | ( n4794 & n4795 ) ;
  assign n4797 = ~x1143 & n4561 ;
  assign n4798 = ( n3214 & n4561 ) | ( n3214 & n4797 ) | ( n4561 & n4797 ) ;
  assign n4799 = x1144 & n3092 ;
  assign n4800 = ( n4793 & n4798 ) | ( n4793 & ~n4799 ) | ( n4798 & ~n4799 ) ;
  assign n4801 = ( ~n4793 & n4796 ) | ( ~n4793 & n4800 ) | ( n4796 & n4800 ) ;
  assign n4802 = ( x275 & n4546 ) | ( x275 & ~n4561 ) | ( n4546 & ~n4561 ) ;
  assign n4803 = x1149 & ~n3214 ;
  assign n4804 = x1150 & n3092 ;
  assign n4805 = ( n3214 & n4634 ) | ( n3214 & n4804 ) | ( n4634 & n4804 ) ;
  assign n4806 = ( n4561 & n4803 ) | ( n4561 & n4805 ) | ( n4803 & n4805 ) ;
  assign n4807 = ( ~n4547 & n4802 ) | ( ~n4547 & n4806 ) | ( n4802 & n4806 ) ;
  assign n4808 = ( x1145 & n3089 ) | ( x1145 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4809 = ( ~n3062 & n4717 ) | ( ~n3062 & n4808 ) | ( n4717 & n4808 ) ;
  assign n4810 = x1146 & n4554 ;
  assign n4811 = ( n4561 & n4809 ) | ( n4561 & n4810 ) | ( n4809 & n4810 ) ;
  assign n4812 = ( x276 & n4541 ) | ( x276 & ~n4561 ) | ( n4541 & ~n4561 ) ;
  assign n4813 = ( ~n4542 & n4811 ) | ( ~n4542 & n4812 ) | ( n4811 & n4812 ) ;
  assign n4814 = x1141 & n3092 ;
  assign n4815 = ( x1142 & n3060 ) | ( x1142 & n3061 ) | ( n3060 & n3061 ) ;
  assign n4816 = x1140 & ~n3062 ;
  assign n4817 = ( ~n3091 & n4815 ) | ( ~n3091 & n4816 ) | ( n4815 & n4816 ) ;
  assign n4818 = ( n4561 & n4814 ) | ( n4561 & n4817 ) | ( n4814 & n4817 ) ;
  assign n4819 = x277 | n4540 ;
  assign n4820 = x820 & n4540 ;
  assign n4821 = ( n4561 & n4819 ) | ( n4561 & ~n4820 ) | ( n4819 & ~n4820 ) ;
  assign n4822 = ~n4818 & n4821 ;
  assign n4823 = ( x1133 & n3089 ) | ( x1133 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4824 = x1132 & ~n3091 ;
  assign n4825 = ( ~n3062 & n4823 ) | ( ~n3062 & n4824 ) | ( n4823 & n4824 ) ;
  assign n4826 = x1134 & n4554 ;
  assign n4827 = ( n4561 & n4825 ) | ( n4561 & n4826 ) | ( n4825 & n4826 ) ;
  assign n4828 = x278 & ~n4540 ;
  assign n4829 = x976 & n4540 ;
  assign n4830 = ( ~n4561 & n4828 ) | ( ~n4561 & n4829 ) | ( n4828 & n4829 ) ;
  assign n4831 = n4827 | n4830 ;
  assign n4832 = ( x1135 & n3060 ) | ( x1135 & n3061 ) | ( n3060 & n3061 ) ;
  assign n4833 = x1133 & ~n3062 ;
  assign n4834 = ( ~n3091 & n4832 ) | ( ~n3091 & n4833 ) | ( n4832 & n4833 ) ;
  assign n4835 = x1134 & n3092 ;
  assign n4836 = ( n4561 & n4834 ) | ( n4561 & n4835 ) | ( n4834 & n4835 ) ;
  assign n4837 = x279 & ~n4540 ;
  assign n4838 = x958 & n4540 ;
  assign n4839 = ( ~n4561 & n4837 ) | ( ~n4561 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4840 = n4836 | n4839 ;
  assign n4841 = ( x1136 & n3089 ) | ( x1136 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4842 = x1135 & ~n3091 ;
  assign n4843 = ( ~n3062 & n4841 ) | ( ~n3062 & n4842 ) | ( n4841 & n4842 ) ;
  assign n4844 = x1137 & n4554 ;
  assign n4845 = ( n4561 & n4843 ) | ( n4561 & n4844 ) | ( n4843 & n4844 ) ;
  assign n4846 = x914 & n4540 ;
  assign n4847 = x280 | n4540 ;
  assign n4848 = ( n4561 & ~n4846 ) | ( n4561 & n4847 ) | ( ~n4846 & n4847 ) ;
  assign n4849 = ~n4845 & n4848 ;
  assign n4850 = x1137 | n3214 ;
  assign n4851 = ( ~x1138 & n3089 ) | ( ~x1138 & n3090 ) | ( n3089 & n3090 ) ;
  assign n4852 = ( n3062 & ~n4762 ) | ( n3062 & n4851 ) | ( ~n4762 & n4851 ) ;
  assign n4853 = ( n4561 & ~n4850 ) | ( n4561 & n4852 ) | ( ~n4850 & n4852 ) ;
  assign n4854 = x281 & ~n4540 ;
  assign n4855 = ~x830 & n4540 ;
  assign n4856 = ( ~n4561 & n4854 ) | ( ~n4561 & n4855 ) | ( n4854 & n4855 ) ;
  assign n4857 = n4853 | n4856 ;
  assign n4858 = ~x1138 & n4561 ;
  assign n4859 = ( n3214 & n4561 ) | ( n3214 & n4858 ) | ( n4561 & n4858 ) ;
  assign n4860 = x282 & ~n4540 ;
  assign n4861 = ~x836 & n4540 ;
  assign n4862 = ( ~n4561 & n4860 ) | ( ~n4561 & n4861 ) | ( n4860 & n4861 ) ;
  assign n4863 = x1140 & n4554 ;
  assign n4864 = x1139 & n3092 ;
  assign n4865 = ( n4859 & n4863 ) | ( n4859 & n4864 ) | ( n4863 & n4864 ) ;
  assign n4866 = ( n4859 & n4862 ) | ( n4859 & ~n4865 ) | ( n4862 & ~n4865 ) ;
  assign n4867 = ~x283 & n4544 ;
  assign n4868 = ( x283 & ~n4544 ) | ( x283 & n4561 ) | ( ~n4544 & n4561 ) ;
  assign n4869 = x1148 & n3092 ;
  assign n4870 = x1149 & n4554 ;
  assign n4871 = ~x1147 & n4561 ;
  assign n4872 = ( n3214 & n4561 ) | ( n3214 & n4871 ) | ( n4561 & n4871 ) ;
  assign n4873 = ~n4870 & n4872 ;
  assign n4874 = ~n4869 & n4873 ;
  assign n4875 = ( n4867 & n4868 ) | ( n4867 & ~n4874 ) | ( n4868 & ~n4874 ) ;
  assign n4876 = x284 | n4692 ;
  assign n4877 = x1143 & ~n2988 ;
  assign n4878 = n4695 & ~n4877 ;
  assign n4879 = ( ~n4695 & n4876 ) | ( ~n4695 & n4878 ) | ( n4876 & n4878 ) ;
  assign n4880 = n2823 & n2887 ;
  assign n4881 = x286 & x288 ;
  assign n4882 = ~n2467 & n4881 ;
  assign n4883 = n4880 & n4882 ;
  assign n4884 = x289 & n4883 ;
  assign n4885 = ( x285 & ~x793 ) | ( x285 & n4884 ) | ( ~x793 & n4884 ) ;
  assign n4886 = n2467 & ~n2468 ;
  assign n4887 = ~n4880 & n4886 ;
  assign n4888 = ~x289 & n4887 ;
  assign n4889 = x285 | n4887 ;
  assign n4890 = ( n4884 & n4888 ) | ( n4884 & n4889 ) | ( n4888 & n4889 ) ;
  assign n4891 = n4885 & ~n4890 ;
  assign n4892 = ( ~x288 & n2467 ) | ( ~x288 & n4880 ) | ( n2467 & n4880 ) ;
  assign n4893 = ( x286 & n4880 ) | ( x286 & ~n4892 ) | ( n4880 & ~n4892 ) ;
  assign n4894 = ~n4883 & n4893 ;
  assign n4895 = n2469 & n4887 ;
  assign n4896 = ( ~x793 & n4894 ) | ( ~x793 & n4895 ) | ( n4894 & n4895 ) ;
  assign n4897 = ~x287 & x457 ;
  assign n4898 = x332 | n4897 ;
  assign n4899 = ( x288 & n2467 ) | ( x288 & ~n2470 ) | ( n2467 & ~n2470 ) ;
  assign n4900 = ( x288 & n2467 ) | ( x288 & n2470 ) | ( n2467 & n2470 ) ;
  assign n4901 = ~n4899 & n4900 ;
  assign n4902 = ~n4880 & n4901 ;
  assign n4903 = ( x793 & n4880 ) | ( x793 & n4901 ) | ( n4880 & n4901 ) ;
  assign n4904 = ( n4880 & n4902 ) | ( n4880 & ~n4903 ) | ( n4902 & ~n4903 ) ;
  assign n4905 = n4883 | n4887 ;
  assign n4906 = ( x289 & ~n2470 ) | ( x289 & n4905 ) | ( ~n2470 & n4905 ) ;
  assign n4907 = ( x289 & ~x793 ) | ( x289 & n4905 ) | ( ~x793 & n4905 ) ;
  assign n4908 = ~n4906 & n4907 ;
  assign n4909 = x290 & x476 ;
  assign n4910 = ~x476 & x1048 ;
  assign n4911 = n4909 | n4910 ;
  assign n4912 = x291 & x476 ;
  assign n4913 = ~x476 & x1049 ;
  assign n4914 = n4912 | n4913 ;
  assign n4915 = x292 & x476 ;
  assign n4916 = ~x476 & x1084 ;
  assign n4917 = n4915 | n4916 ;
  assign n4918 = x293 & x476 ;
  assign n4919 = ~x476 & x1059 ;
  assign n4920 = n4918 | n4919 ;
  assign n4921 = x294 & x476 ;
  assign n4922 = ~x476 & x1072 ;
  assign n4923 = n4921 | n4922 ;
  assign n4924 = x295 & x476 ;
  assign n4925 = ~x476 & x1053 ;
  assign n4926 = n4924 | n4925 ;
  assign n4927 = x296 & x476 ;
  assign n4928 = ~x476 & x1037 ;
  assign n4929 = n4927 | n4928 ;
  assign n4930 = x297 & x476 ;
  assign n4931 = ~x476 & x1044 ;
  assign n4932 = n4930 | n4931 ;
  assign n4933 = x298 & x478 ;
  assign n4934 = ~x478 & x1044 ;
  assign n4935 = n4933 | n4934 ;
  assign n4936 = x53 | n2997 ;
  assign n4937 = ( ~n2995 & n2997 ) | ( ~n2995 & n4936 ) | ( n2997 & n4936 ) ;
  assign n4938 = n3001 | n4937 ;
  assign n4939 = n3003 | n4938 ;
  assign n4940 = ~x59 & n3045 ;
  assign n4941 = ( x312 & n3143 ) | ( x312 & n4940 ) | ( n3143 & n4940 ) ;
  assign n4942 = n4940 & ~n4941 ;
  assign n4943 = ( x55 & ~x300 ) | ( x55 & n4942 ) | ( ~x300 & n4942 ) ;
  assign n4944 = ( x55 & x300 ) | ( x55 & ~n4942 ) | ( x300 & ~n4942 ) ;
  assign n4945 = n4943 | n4944 ;
  assign n4946 = ( x55 & ~x301 ) | ( x55 & n4943 ) | ( ~x301 & n4943 ) ;
  assign n4947 = ( x55 & x301 ) | ( x55 & ~n4943 ) | ( x301 & ~n4943 ) ;
  assign n4948 = n4946 | n4947 ;
  assign n4949 = ~x1148 & n1606 ;
  assign n4950 = ( ~x937 & n1599 ) | ( ~x937 & n1600 ) | ( n1599 & n1600 ) ;
  assign n4951 = n1607 | n1608 ;
  assign n4952 = ( x237 & ~n1605 ) | ( x237 & n4951 ) | ( ~n1605 & n4951 ) ;
  assign n4953 = n4950 | n4952 ;
  assign n4954 = ( x273 & n1607 ) | ( x273 & n1608 ) | ( n1607 & n1608 ) ;
  assign n4955 = ( n4949 & n4953 ) | ( n4949 & ~n4954 ) | ( n4953 & ~n4954 ) ;
  assign n4956 = x303 & x478 ;
  assign n4957 = ~x478 & x1049 ;
  assign n4958 = n4956 | n4957 ;
  assign n4959 = x304 & x478 ;
  assign n4960 = ~x478 & x1048 ;
  assign n4961 = n4959 | n4960 ;
  assign n4962 = x305 & x478 ;
  assign n4963 = ~x478 & x1084 ;
  assign n4964 = n4962 | n4963 ;
  assign n4965 = x306 & x478 ;
  assign n4966 = ~x478 & x1059 ;
  assign n4967 = n4965 | n4966 ;
  assign n4968 = x307 & x478 ;
  assign n4969 = ~x478 & x1053 ;
  assign n4970 = n4968 | n4969 ;
  assign n4971 = x308 & x478 ;
  assign n4972 = ~x478 & x1037 ;
  assign n4973 = n4971 | n4972 ;
  assign n4974 = x309 & x478 ;
  assign n4975 = ~x478 & x1072 ;
  assign n4976 = n4974 | n4975 ;
  assign n4977 = ( x934 & n1599 ) | ( x934 & n1600 ) | ( n1599 & n1600 ) ;
  assign n4978 = x233 & ~n4951 ;
  assign n4979 = ( ~x271 & n1607 ) | ( ~x271 & n1608 ) | ( n1607 & n1608 ) ;
  assign n4980 = ( ~n1605 & n4978 ) | ( ~n1605 & n4979 ) | ( n4978 & n4979 ) ;
  assign n4981 = ( ~x1147 & n1602 ) | ( ~x1147 & n1605 ) | ( n1602 & n1605 ) ;
  assign n4982 = ( ~n4977 & n4980 ) | ( ~n4977 & n4981 ) | ( n4980 & n4981 ) ;
  assign n4983 = ~x300 & x301 ;
  assign n4984 = ( x311 & n4942 ) | ( x311 & ~n4983 ) | ( n4942 & ~n4983 ) ;
  assign n4985 = ( x55 & n4942 ) | ( x55 & ~n4984 ) | ( n4942 & ~n4984 ) ;
  assign n4986 = n4983 & n4984 ;
  assign n4987 = ( x311 & n4985 ) | ( x311 & ~n4986 ) | ( n4985 & ~n4986 ) ;
  assign n4988 = ( x55 & ~n3143 ) | ( x55 & n4941 ) | ( ~n3143 & n4941 ) ;
  assign n4989 = ( x312 & n4942 ) | ( x312 & ~n4988 ) | ( n4942 & ~n4988 ) ;
  assign n4990 = x313 & x954 ;
  assign n4991 = x110 | x111 ;
  assign n4992 = ( ~n1960 & n3332 ) | ( ~n1960 & n4991 ) | ( n3332 & n4991 ) ;
  assign n4993 = n2823 & n4992 ;
  assign n4994 = ~x313 & x954 ;
  assign n4995 = ( ~n4990 & n4993 ) | ( ~n4990 & n4994 ) | ( n4993 & n4994 ) ;
  assign n4996 = n2760 | n3496 ;
  assign n4997 = n3543 | n4996 ;
  assign n4998 = ~x340 & n4880 ;
  assign n4999 = ~x1080 & n4998 ;
  assign n5000 = x315 & ~n4998 ;
  assign n5001 = ( n4998 & ~n4999 ) | ( n4998 & n5000 ) | ( ~n4999 & n5000 ) ;
  assign n5002 = x316 & ~n4998 ;
  assign n5003 = x1047 & n4998 ;
  assign n5004 = n5002 | n5003 ;
  assign n5005 = ~x330 & n4880 ;
  assign n5006 = ~x1078 & n5005 ;
  assign n5007 = x317 & ~n5005 ;
  assign n5008 = ( n5005 & ~n5006 ) | ( n5005 & n5007 ) | ( ~n5006 & n5007 ) ;
  assign n5009 = ~x341 & n4880 ;
  assign n5010 = ~x1074 & n5009 ;
  assign n5011 = x318 & ~n5009 ;
  assign n5012 = ( n5009 & ~n5010 ) | ( n5009 & n5011 ) | ( ~n5010 & n5011 ) ;
  assign n5013 = x319 & ~n5009 ;
  assign n5014 = x1072 & n5009 ;
  assign n5015 = n5013 | n5014 ;
  assign n5016 = x320 & ~n4998 ;
  assign n5017 = x1048 & n4998 ;
  assign n5018 = n5016 | n5017 ;
  assign n5019 = x321 & ~n4998 ;
  assign n5020 = x1058 & n4998 ;
  assign n5021 = n5019 | n5020 ;
  assign n5022 = x322 & ~n4998 ;
  assign n5023 = x1051 & n4998 ;
  assign n5024 = n5022 | n5023 ;
  assign n5025 = x323 & ~n4998 ;
  assign n5026 = x1065 & n4998 ;
  assign n5027 = n5025 | n5026 ;
  assign n5028 = x324 & ~n5009 ;
  assign n5029 = x1086 & n5009 ;
  assign n5030 = n5028 | n5029 ;
  assign n5031 = x325 & ~n5009 ;
  assign n5032 = x1063 & n5009 ;
  assign n5033 = n5031 | n5032 ;
  assign n5034 = x326 & ~n5009 ;
  assign n5035 = x1057 & n5009 ;
  assign n5036 = n5034 | n5035 ;
  assign n5037 = x327 & ~n4998 ;
  assign n5038 = x1040 & n4998 ;
  assign n5039 = n5037 | n5038 ;
  assign n5040 = x328 & ~n5009 ;
  assign n5041 = x1058 & n5009 ;
  assign n5042 = n5040 | n5041 ;
  assign n5043 = x329 & ~n5009 ;
  assign n5044 = x1043 & n5009 ;
  assign n5045 = n5043 | n5044 ;
  assign n5046 = x330 | n4880 ;
  assign n5047 = x1092 & ~n4308 ;
  assign n5048 = ( n4998 & ~n5046 ) | ( n4998 & n5047 ) | ( ~n5046 & n5047 ) ;
  assign n5049 = x331 | n4880 ;
  assign n5050 = ( n5009 & n5047 ) | ( n5009 & ~n5049 ) | ( n5047 & ~n5049 ) ;
  assign n5051 = n1483 | n2824 ;
  assign n5052 = n2823 & n5051 ;
  assign n5053 = n1309 & ~n2128 ;
  assign n5054 = ( ~n4285 & n5052 ) | ( ~n4285 & n5053 ) | ( n5052 & n5053 ) ;
  assign n5055 = n4285 | n5054 ;
  assign n5056 = ( n2618 & n5052 ) | ( n2618 & n5055 ) | ( n5052 & n5055 ) ;
  assign n5057 = x333 & ~n5009 ;
  assign n5058 = x1040 & n5009 ;
  assign n5059 = n5057 | n5058 ;
  assign n5060 = x334 & ~n5009 ;
  assign n5061 = x1065 & n5009 ;
  assign n5062 = n5060 | n5061 ;
  assign n5063 = x335 & ~n5009 ;
  assign n5064 = x1069 & n5009 ;
  assign n5065 = n5063 | n5064 ;
  assign n5066 = x336 & ~n5005 ;
  assign n5067 = x1070 & n5005 ;
  assign n5068 = n5066 | n5067 ;
  assign n5069 = x337 & ~n5005 ;
  assign n5070 = x1044 & n5005 ;
  assign n5071 = n5069 | n5070 ;
  assign n5072 = x338 & ~n5005 ;
  assign n5073 = x1072 & n5005 ;
  assign n5074 = n5072 | n5073 ;
  assign n5075 = x339 & ~n5005 ;
  assign n5076 = x1086 & n5005 ;
  assign n5077 = n5075 | n5076 ;
  assign n5078 = x340 & ~n4880 ;
  assign n5079 = x331 & n4880 ;
  assign n5080 = ( n5047 & n5078 ) | ( n5047 & n5079 ) | ( n5078 & n5079 ) ;
  assign n5081 = x341 | n4880 ;
  assign n5082 = ( n5005 & n5047 ) | ( n5005 & ~n5081 ) | ( n5047 & ~n5081 ) ;
  assign n5083 = x342 & ~n4998 ;
  assign n5084 = x1049 & n4998 ;
  assign n5085 = n5083 | n5084 ;
  assign n5086 = x343 & ~n4998 ;
  assign n5087 = x1062 & n4998 ;
  assign n5088 = n5086 | n5087 ;
  assign n5089 = x344 & ~n4998 ;
  assign n5090 = x1069 & n4998 ;
  assign n5091 = n5089 | n5090 ;
  assign n5092 = x345 & ~n4998 ;
  assign n5093 = x1039 & n4998 ;
  assign n5094 = n5092 | n5093 ;
  assign n5095 = x346 & ~n4998 ;
  assign n5096 = x1067 & n4998 ;
  assign n5097 = n5095 | n5096 ;
  assign n5098 = x347 & ~n4998 ;
  assign n5099 = x1055 & n4998 ;
  assign n5100 = n5098 | n5099 ;
  assign n5101 = x348 & ~n4998 ;
  assign n5102 = x1087 & n4998 ;
  assign n5103 = n5101 | n5102 ;
  assign n5104 = x349 & ~n4998 ;
  assign n5105 = x1043 & n4998 ;
  assign n5106 = n5104 | n5105 ;
  assign n5107 = x350 & ~n4998 ;
  assign n5108 = x1035 & n4998 ;
  assign n5109 = n5107 | n5108 ;
  assign n5110 = x351 & ~n4998 ;
  assign n5111 = x1079 & n4998 ;
  assign n5112 = n5110 | n5111 ;
  assign n5113 = x352 & ~n4998 ;
  assign n5114 = x1078 & n4998 ;
  assign n5115 = n5113 | n5114 ;
  assign n5116 = x353 & ~n4998 ;
  assign n5117 = x1063 & n4998 ;
  assign n5118 = n5116 | n5117 ;
  assign n5119 = x354 & ~n4998 ;
  assign n5120 = x1045 & n4998 ;
  assign n5121 = n5119 | n5120 ;
  assign n5122 = x355 & ~n4998 ;
  assign n5123 = x1084 & n4998 ;
  assign n5124 = n5122 | n5123 ;
  assign n5125 = x356 & ~n4998 ;
  assign n5126 = x1081 & n4998 ;
  assign n5127 = n5125 | n5126 ;
  assign n5128 = x357 & ~n4998 ;
  assign n5129 = x1076 & n4998 ;
  assign n5130 = n5128 | n5129 ;
  assign n5131 = x358 & ~n4998 ;
  assign n5132 = x1071 & n4998 ;
  assign n5133 = n5131 | n5132 ;
  assign n5134 = x359 & ~n4998 ;
  assign n5135 = x1068 & n4998 ;
  assign n5136 = n5134 | n5135 ;
  assign n5137 = x360 & ~n4998 ;
  assign n5138 = x1042 & n4998 ;
  assign n5139 = n5137 | n5138 ;
  assign n5140 = x361 & ~n4998 ;
  assign n5141 = x1059 & n4998 ;
  assign n5142 = n5140 | n5141 ;
  assign n5143 = x362 & ~n4998 ;
  assign n5144 = x1070 & n4998 ;
  assign n5145 = n5143 | n5144 ;
  assign n5146 = x363 & ~n5005 ;
  assign n5147 = x1049 & n5005 ;
  assign n5148 = n5146 | n5147 ;
  assign n5149 = x364 & ~n5005 ;
  assign n5150 = x1062 & n5005 ;
  assign n5151 = n5149 | n5150 ;
  assign n5152 = x365 & ~n5005 ;
  assign n5153 = x1065 & n5005 ;
  assign n5154 = n5152 | n5153 ;
  assign n5155 = x366 & ~n5005 ;
  assign n5156 = x1069 & n5005 ;
  assign n5157 = n5155 | n5156 ;
  assign n5158 = x367 & ~n5005 ;
  assign n5159 = x1039 & n5005 ;
  assign n5160 = n5158 | n5159 ;
  assign n5161 = x368 & ~n5005 ;
  assign n5162 = x1067 & n5005 ;
  assign n5163 = n5161 | n5162 ;
  assign n5164 = x369 & ~n5005 ;
  assign n5165 = x1080 & n5005 ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = x370 & ~n5005 ;
  assign n5168 = x1055 & n5005 ;
  assign n5169 = n5167 | n5168 ;
  assign n5170 = x371 & ~n5005 ;
  assign n5171 = x1051 & n5005 ;
  assign n5172 = n5170 | n5171 ;
  assign n5173 = x372 & ~n5005 ;
  assign n5174 = x1048 & n5005 ;
  assign n5175 = n5173 | n5174 ;
  assign n5176 = x373 & ~n5005 ;
  assign n5177 = x1087 & n5005 ;
  assign n5178 = n5176 | n5177 ;
  assign n5179 = x374 & ~n5005 ;
  assign n5180 = x1035 & n5005 ;
  assign n5181 = n5179 | n5180 ;
  assign n5182 = x375 & ~n5005 ;
  assign n5183 = x1047 & n5005 ;
  assign n5184 = n5182 | n5183 ;
  assign n5185 = x376 & ~n5005 ;
  assign n5186 = x1079 & n5005 ;
  assign n5187 = n5185 | n5186 ;
  assign n5188 = x377 & ~n5005 ;
  assign n5189 = x1074 & n5005 ;
  assign n5190 = n5188 | n5189 ;
  assign n5191 = x378 & ~n5005 ;
  assign n5192 = x1063 & n5005 ;
  assign n5193 = n5191 | n5192 ;
  assign n5194 = x379 & ~n5005 ;
  assign n5195 = x1045 & n5005 ;
  assign n5196 = n5194 | n5195 ;
  assign n5197 = x380 & ~n5005 ;
  assign n5198 = x1084 & n5005 ;
  assign n5199 = n5197 | n5198 ;
  assign n5200 = x381 & ~n5005 ;
  assign n5201 = x1081 & n5005 ;
  assign n5202 = n5200 | n5201 ;
  assign n5203 = x382 & ~n5005 ;
  assign n5204 = x1076 & n5005 ;
  assign n5205 = n5203 | n5204 ;
  assign n5206 = x383 & ~n5005 ;
  assign n5207 = x1071 & n5005 ;
  assign n5208 = n5206 | n5207 ;
  assign n5209 = x384 & ~n5005 ;
  assign n5210 = x1068 & n5005 ;
  assign n5211 = n5209 | n5210 ;
  assign n5212 = x385 & ~n5005 ;
  assign n5213 = x1042 & n5005 ;
  assign n5214 = n5212 | n5213 ;
  assign n5215 = x386 & ~n5005 ;
  assign n5216 = x1059 & n5005 ;
  assign n5217 = n5215 | n5216 ;
  assign n5218 = x387 & ~n5005 ;
  assign n5219 = x1053 & n5005 ;
  assign n5220 = n5218 | n5219 ;
  assign n5221 = x388 & ~n5005 ;
  assign n5222 = x1037 & n5005 ;
  assign n5223 = n5221 | n5222 ;
  assign n5224 = x389 & ~n5005 ;
  assign n5225 = x1036 & n5005 ;
  assign n5226 = n5224 | n5225 ;
  assign n5227 = x390 & ~n5009 ;
  assign n5228 = x1049 & n5009 ;
  assign n5229 = n5227 | n5228 ;
  assign n5230 = x391 & ~n5009 ;
  assign n5231 = x1062 & n5009 ;
  assign n5232 = n5230 | n5231 ;
  assign n5233 = x392 & ~n5009 ;
  assign n5234 = x1039 & n5009 ;
  assign n5235 = n5233 | n5234 ;
  assign n5236 = x393 & ~n5009 ;
  assign n5237 = x1067 & n5009 ;
  assign n5238 = n5236 | n5237 ;
  assign n5239 = x394 & ~n5009 ;
  assign n5240 = x1080 & n5009 ;
  assign n5241 = n5239 | n5240 ;
  assign n5242 = x395 & ~n5009 ;
  assign n5243 = x1055 & n5009 ;
  assign n5244 = n5242 | n5243 ;
  assign n5245 = x396 & ~n5009 ;
  assign n5246 = x1051 & n5009 ;
  assign n5247 = n5245 | n5246 ;
  assign n5248 = x397 & ~n5009 ;
  assign n5249 = x1048 & n5009 ;
  assign n5250 = n5248 | n5249 ;
  assign n5251 = x398 & ~n5009 ;
  assign n5252 = x1087 & n5009 ;
  assign n5253 = n5251 | n5252 ;
  assign n5254 = x399 & ~n5009 ;
  assign n5255 = x1047 & n5009 ;
  assign n5256 = n5254 | n5255 ;
  assign n5257 = x400 & ~n5009 ;
  assign n5258 = x1035 & n5009 ;
  assign n5259 = n5257 | n5258 ;
  assign n5260 = x401 & ~n5009 ;
  assign n5261 = x1079 & n5009 ;
  assign n5262 = n5260 | n5261 ;
  assign n5263 = x402 & ~n5009 ;
  assign n5264 = x1078 & n5009 ;
  assign n5265 = n5263 | n5264 ;
  assign n5266 = x403 & ~n5009 ;
  assign n5267 = x1045 & n5009 ;
  assign n5268 = n5266 | n5267 ;
  assign n5269 = x404 & ~n5009 ;
  assign n5270 = x1084 & n5009 ;
  assign n5271 = n5269 | n5270 ;
  assign n5272 = x405 & ~n5009 ;
  assign n5273 = x1081 & n5009 ;
  assign n5274 = n5272 | n5273 ;
  assign n5275 = x406 & ~n5009 ;
  assign n5276 = x1076 & n5009 ;
  assign n5277 = n5275 | n5276 ;
  assign n5278 = x407 & ~n5009 ;
  assign n5279 = x1071 & n5009 ;
  assign n5280 = n5278 | n5279 ;
  assign n5281 = x408 & ~n5009 ;
  assign n5282 = x1068 & n5009 ;
  assign n5283 = n5281 | n5282 ;
  assign n5284 = x409 & ~n5009 ;
  assign n5285 = x1042 & n5009 ;
  assign n5286 = n5284 | n5285 ;
  assign n5287 = x410 & ~n5009 ;
  assign n5288 = x1059 & n5009 ;
  assign n5289 = n5287 | n5288 ;
  assign n5290 = x411 & ~n5009 ;
  assign n5291 = x1053 & n5009 ;
  assign n5292 = n5290 | n5291 ;
  assign n5293 = x412 & ~n5009 ;
  assign n5294 = x1037 & n5009 ;
  assign n5295 = n5293 | n5294 ;
  assign n5296 = x413 & ~n5009 ;
  assign n5297 = x1036 & n5009 ;
  assign n5298 = n5296 | n5297 ;
  assign n5299 = ~x331 & n4880 ;
  assign n5300 = x414 & ~n5299 ;
  assign n5301 = ~x1049 & n5299 ;
  assign n5302 = ( n5299 & n5300 ) | ( n5299 & ~n5301 ) | ( n5300 & ~n5301 ) ;
  assign n5303 = x415 & ~n5299 ;
  assign n5304 = x1062 & n5299 ;
  assign n5305 = n5303 | n5304 ;
  assign n5306 = x416 & ~n5299 ;
  assign n5307 = x1069 & n5299 ;
  assign n5308 = n5306 | n5307 ;
  assign n5309 = x417 & ~n5299 ;
  assign n5310 = x1039 & n5299 ;
  assign n5311 = n5309 | n5310 ;
  assign n5312 = x418 & ~n5299 ;
  assign n5313 = x1067 & n5299 ;
  assign n5314 = n5312 | n5313 ;
  assign n5315 = x419 & ~n5299 ;
  assign n5316 = x1080 & n5299 ;
  assign n5317 = n5315 | n5316 ;
  assign n5318 = x420 & ~n5299 ;
  assign n5319 = x1055 & n5299 ;
  assign n5320 = n5318 | n5319 ;
  assign n5321 = x421 & ~n5299 ;
  assign n5322 = x1051 & n5299 ;
  assign n5323 = n5321 | n5322 ;
  assign n5324 = x422 & ~n5299 ;
  assign n5325 = x1048 & n5299 ;
  assign n5326 = n5324 | n5325 ;
  assign n5327 = x423 & ~n5299 ;
  assign n5328 = x1087 & n5299 ;
  assign n5329 = n5327 | n5328 ;
  assign n5330 = x424 & ~n5299 ;
  assign n5331 = x1047 & n5299 ;
  assign n5332 = n5330 | n5331 ;
  assign n5333 = x425 & ~n5299 ;
  assign n5334 = x1035 & n5299 ;
  assign n5335 = n5333 | n5334 ;
  assign n5336 = x426 & ~n5299 ;
  assign n5337 = x1079 & n5299 ;
  assign n5338 = n5336 | n5337 ;
  assign n5339 = x427 & ~n5299 ;
  assign n5340 = x1078 & n5299 ;
  assign n5341 = n5339 | n5340 ;
  assign n5342 = x428 & ~n5299 ;
  assign n5343 = x1045 & n5299 ;
  assign n5344 = n5342 | n5343 ;
  assign n5345 = x429 & ~n5299 ;
  assign n5346 = x1084 & n5299 ;
  assign n5347 = n5345 | n5346 ;
  assign n5348 = x430 & ~n5299 ;
  assign n5349 = x1076 & n5299 ;
  assign n5350 = n5348 | n5349 ;
  assign n5351 = x431 & ~n5299 ;
  assign n5352 = x1071 & n5299 ;
  assign n5353 = n5351 | n5352 ;
  assign n5354 = x432 & ~n5299 ;
  assign n5355 = x1068 & n5299 ;
  assign n5356 = n5354 | n5355 ;
  assign n5357 = x433 & ~n5299 ;
  assign n5358 = x1042 & n5299 ;
  assign n5359 = n5357 | n5358 ;
  assign n5360 = x434 & ~n5299 ;
  assign n5361 = x1059 & n5299 ;
  assign n5362 = n5360 | n5361 ;
  assign n5363 = x435 & ~n5299 ;
  assign n5364 = x1053 & n5299 ;
  assign n5365 = n5363 | n5364 ;
  assign n5366 = x436 & ~n5299 ;
  assign n5367 = x1037 & n5299 ;
  assign n5368 = n5366 | n5367 ;
  assign n5369 = x437 & ~n5299 ;
  assign n5370 = x1070 & n5299 ;
  assign n5371 = n5369 | n5370 ;
  assign n5372 = x438 & ~n5299 ;
  assign n5373 = x1036 & n5299 ;
  assign n5374 = n5372 | n5373 ;
  assign n5375 = x439 & ~n5005 ;
  assign n5376 = x1057 & n5005 ;
  assign n5377 = n5375 | n5376 ;
  assign n5378 = x440 & ~n5005 ;
  assign n5379 = x1043 & n5005 ;
  assign n5380 = n5378 | n5379 ;
  assign n5381 = x441 & ~n4998 ;
  assign n5382 = x1044 & n4998 ;
  assign n5383 = n5381 | n5382 ;
  assign n5384 = x442 & ~n5005 ;
  assign n5385 = x1058 & n5005 ;
  assign n5386 = n5384 | n5385 ;
  assign n5387 = x443 & ~n5299 ;
  assign n5388 = x1044 & n5299 ;
  assign n5389 = n5387 | n5388 ;
  assign n5390 = x444 & ~n5299 ;
  assign n5391 = x1072 & n5299 ;
  assign n5392 = n5390 | n5391 ;
  assign n5393 = x445 & ~n5299 ;
  assign n5394 = x1081 & n5299 ;
  assign n5395 = n5393 | n5394 ;
  assign n5396 = x446 & ~n5299 ;
  assign n5397 = x1086 & n5299 ;
  assign n5398 = n5396 | n5397 ;
  assign n5399 = x447 & ~n5005 ;
  assign n5400 = x1040 & n5005 ;
  assign n5401 = n5399 | n5400 ;
  assign n5402 = x448 & ~n5299 ;
  assign n5403 = x1074 & n5299 ;
  assign n5404 = n5402 | n5403 ;
  assign n5405 = x449 & ~n5299 ;
  assign n5406 = x1057 & n5299 ;
  assign n5407 = n5405 | n5406 ;
  assign n5408 = x450 & ~n4998 ;
  assign n5409 = x1036 & n4998 ;
  assign n5410 = n5408 | n5409 ;
  assign n5411 = x451 & ~n5299 ;
  assign n5412 = x1063 & n5299 ;
  assign n5413 = n5411 | n5412 ;
  assign n5414 = x452 & ~n4998 ;
  assign n5415 = x1053 & n4998 ;
  assign n5416 = n5414 | n5415 ;
  assign n5417 = x453 & ~n5299 ;
  assign n5418 = x1040 & n5299 ;
  assign n5419 = n5417 | n5418 ;
  assign n5420 = x454 & ~n5299 ;
  assign n5421 = x1043 & n5299 ;
  assign n5422 = n5420 | n5421 ;
  assign n5423 = x455 & ~n4998 ;
  assign n5424 = x1037 & n4998 ;
  assign n5425 = n5423 | n5424 ;
  assign n5426 = x456 & ~n5009 ;
  assign n5427 = x1044 & n5009 ;
  assign n5428 = n5426 | n5427 ;
  assign n5429 = ~x600 & x804 ;
  assign n5430 = ( ~x601 & x804 ) | ( ~x601 & x810 ) | ( x804 & x810 ) ;
  assign n5431 = n5429 | n5430 ;
  assign n5432 = x605 & ~x815 ;
  assign n5433 = ( x821 & n5431 ) | ( x821 & ~n5432 ) | ( n5431 & ~n5432 ) ;
  assign n5434 = x594 & x600 ;
  assign n5435 = x821 & n5434 ;
  assign n5436 = x804 & x990 ;
  assign n5437 = x810 & ~x815 ;
  assign n5438 = ( n5435 & ~n5436 ) | ( n5435 & n5437 ) | ( ~n5436 & n5437 ) ;
  assign n5439 = n5436 & n5438 ;
  assign n5440 = x597 & x601 ;
  assign n5441 = x605 & n5440 ;
  assign n5442 = x595 & x596 ;
  assign n5443 = ( ~x599 & x810 ) | ( ~x599 & n5437 ) | ( x810 & n5437 ) ;
  assign n5444 = n5442 & ~n5443 ;
  assign n5445 = ~x595 & x810 ;
  assign n5446 = ( x804 & ~n5444 ) | ( x804 & n5445 ) | ( ~n5444 & n5445 ) ;
  assign n5447 = n5441 & ~n5446 ;
  assign n5448 = ( n5435 & n5439 ) | ( n5435 & n5447 ) | ( n5439 & n5447 ) ;
  assign n5449 = ( x821 & ~n5433 ) | ( x821 & n5448 ) | ( ~n5433 & n5448 ) ;
  assign n5450 = x458 & ~n4998 ;
  assign n5451 = x1072 & n4998 ;
  assign n5452 = n5450 | n5451 ;
  assign n5453 = x459 & ~n5299 ;
  assign n5454 = x1058 & n5299 ;
  assign n5455 = n5453 | n5454 ;
  assign n5456 = x460 & ~n4998 ;
  assign n5457 = x1086 & n4998 ;
  assign n5458 = n5456 | n5457 ;
  assign n5459 = x461 & ~n4998 ;
  assign n5460 = x1057 & n4998 ;
  assign n5461 = n5459 | n5460 ;
  assign n5462 = x462 & ~n4998 ;
  assign n5463 = x1074 & n4998 ;
  assign n5464 = n5462 | n5463 ;
  assign n5465 = x463 & ~n5009 ;
  assign n5466 = x1070 & n5009 ;
  assign n5467 = n5465 | n5466 ;
  assign n5468 = x464 & ~n5299 ;
  assign n5469 = x1065 & n5299 ;
  assign n5470 = n5468 | n5469 ;
  assign n5471 = ( x926 & n1599 ) | ( x926 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5472 = ( ~x243 & n1607 ) | ( ~x243 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5473 = x1157 | n5472 ;
  assign n5474 = ( n1606 & n5472 ) | ( n1606 & n5473 ) | ( n5472 & n5473 ) ;
  assign n5475 = n5471 | n5474 ;
  assign n5476 = ( x275 & n1607 ) | ( x275 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5477 = ( x943 & n1599 ) | ( x943 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5478 = ( x1151 & n1602 ) | ( x1151 & ~n1605 ) | ( n1602 & ~n1605 ) ;
  assign n5479 = ( x1151 & n5477 ) | ( x1151 & ~n5478 ) | ( n5477 & ~n5478 ) ;
  assign n5480 = n5476 | n5479 ;
  assign n5481 = n3205 & n4316 ;
  assign n5482 = x40 & ~x287 ;
  assign n5483 = ( ~x1001 & n1990 ) | ( ~x1001 & n5482 ) | ( n1990 & n5482 ) ;
  assign n5484 = n5482 & ~n5483 ;
  assign n5485 = n1995 & n5484 ;
  assign n5486 = ( n5481 & n5484 ) | ( n5481 & ~n5485 ) | ( n5484 & ~n5485 ) ;
  assign n5487 = x468 & ~n2797 ;
  assign n5488 = ( x468 & ~n2618 ) | ( x468 & n5487 ) | ( ~n2618 & n5487 ) ;
  assign n5489 = n3039 | n5488 ;
  assign n5490 = ( ~x263 & n1607 ) | ( ~x263 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5491 = ( x942 & n1599 ) | ( x942 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5492 = ( x1156 & n1602 ) | ( x1156 & ~n1605 ) | ( n1602 & ~n1605 ) ;
  assign n5493 = ( x1156 & n5491 ) | ( x1156 & ~n5492 ) | ( n5491 & ~n5492 ) ;
  assign n5494 = n5490 | n5493 ;
  assign n5495 = ( x267 & n1607 ) | ( x267 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5496 = ( x925 & n1599 ) | ( x925 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5497 = ( x1155 & n1602 ) | ( x1155 & ~n1605 ) | ( n1602 & ~n1605 ) ;
  assign n5498 = ( x1155 & n5496 ) | ( x1155 & ~n5497 ) | ( n5496 & ~n5497 ) ;
  assign n5499 = n5495 | n5498 ;
  assign n5500 = ( x253 & n1607 ) | ( x253 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5501 = ( x941 & n1599 ) | ( x941 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5502 = x1153 | n5501 ;
  assign n5503 = ( n1606 & n5501 ) | ( n1606 & n5502 ) | ( n5501 & n5502 ) ;
  assign n5504 = n5500 | n5503 ;
  assign n5505 = ( x254 & n1607 ) | ( x254 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5506 = ( x923 & n1599 ) | ( x923 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5507 = ( x1154 & n1602 ) | ( x1154 & ~n1605 ) | ( n1602 & ~n1605 ) ;
  assign n5508 = ( x1154 & n5506 ) | ( x1154 & ~n5507 ) | ( n5506 & ~n5507 ) ;
  assign n5509 = n5505 | n5508 ;
  assign n5510 = ( x268 & n1607 ) | ( x268 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5511 = ( x922 & n1599 ) | ( x922 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5512 = ( x1152 & n1602 ) | ( x1152 & ~n1605 ) | ( n1602 & ~n1605 ) ;
  assign n5513 = ( x1152 & n5511 ) | ( x1152 & ~n5512 ) | ( n5511 & ~n5512 ) ;
  assign n5514 = n5510 | n5513 ;
  assign n5515 = ( x931 & n1599 ) | ( x931 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5516 = ( x272 & n1607 ) | ( x272 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5517 = x1150 | n5516 ;
  assign n5518 = ( n1606 & n5516 ) | ( n1606 & n5517 ) | ( n5516 & n5517 ) ;
  assign n5519 = n5515 | n5518 ;
  assign n5520 = ( x936 & n1599 ) | ( x936 & n1600 ) | ( n1599 & n1600 ) ;
  assign n5521 = ( x283 & n1607 ) | ( x283 & n1608 ) | ( n1607 & n1608 ) ;
  assign n5522 = x1149 | n5521 ;
  assign n5523 = ( n1606 & n5521 ) | ( n1606 & n5522 ) | ( n5521 & n5522 ) ;
  assign n5524 = n5520 | n5523 ;
  assign n5525 = x71 & n3092 ;
  assign n5526 = x84 | n5525 ;
  assign n5527 = ( n2982 & n5525 ) | ( n2982 & n5526 ) | ( n5525 & n5526 ) ;
  assign n5528 = x71 & ~n3214 ;
  assign n5529 = x248 & n4136 ;
  assign n5530 = x481 & ~n4136 ;
  assign n5531 = n5529 | n5530 ;
  assign n5532 = x249 & n4160 ;
  assign n5533 = x482 & ~n4160 ;
  assign n5534 = n5532 | n5533 ;
  assign n5535 = x242 & n4179 ;
  assign n5536 = x483 & ~n4179 ;
  assign n5537 = n5535 | n5536 ;
  assign n5538 = x249 & n4179 ;
  assign n5539 = x484 & ~n4179 ;
  assign n5540 = n5538 | n5539 ;
  assign n5541 = x234 & n4241 ;
  assign n5542 = x485 & ~n4241 ;
  assign n5543 = n5541 | n5542 ;
  assign n5544 = x244 & n4241 ;
  assign n5545 = x486 & ~n4241 ;
  assign n5546 = n5544 | n5545 ;
  assign n5547 = x246 & n4136 ;
  assign n5548 = x487 & ~n4136 ;
  assign n5549 = n5547 | n5548 ;
  assign n5550 = ~x239 & n4136 ;
  assign n5551 = x488 & ~n4136 ;
  assign n5552 = n5550 | n5551 ;
  assign n5553 = x242 & n4241 ;
  assign n5554 = x489 & ~n4241 ;
  assign n5555 = n5553 | n5554 ;
  assign n5556 = x241 & n4179 ;
  assign n5557 = x490 & ~n4179 ;
  assign n5558 = n5556 | n5557 ;
  assign n5559 = x238 & n4179 ;
  assign n5560 = x491 & ~n4179 ;
  assign n5561 = n5559 | n5560 ;
  assign n5562 = x240 & n4179 ;
  assign n5563 = x492 & ~n4179 ;
  assign n5564 = n5562 | n5563 ;
  assign n5565 = x244 & n4179 ;
  assign n5566 = x493 & ~n4179 ;
  assign n5567 = n5565 | n5566 ;
  assign n5568 = ~x239 & n4179 ;
  assign n5569 = x494 & ~n4179 ;
  assign n5570 = n5568 | n5569 ;
  assign n5571 = x235 & n4179 ;
  assign n5572 = x495 & ~n4179 ;
  assign n5573 = n5571 | n5572 ;
  assign n5574 = x249 & n4172 ;
  assign n5575 = x496 & ~n4172 ;
  assign n5576 = n5574 | n5575 ;
  assign n5577 = ~x239 & n4172 ;
  assign n5578 = x497 & ~n4172 ;
  assign n5579 = n5577 | n5578 ;
  assign n5580 = x238 & n4160 ;
  assign n5581 = x498 & ~n4160 ;
  assign n5582 = n5580 | n5581 ;
  assign n5583 = x246 & n4172 ;
  assign n5584 = x499 & ~n4172 ;
  assign n5585 = n5583 | n5584 ;
  assign n5586 = x241 & n4172 ;
  assign n5587 = x500 & ~n4172 ;
  assign n5588 = n5586 | n5587 ;
  assign n5589 = x248 & n4172 ;
  assign n5590 = x501 & ~n4172 ;
  assign n5591 = n5589 | n5590 ;
  assign n5592 = x247 & n4172 ;
  assign n5593 = x502 & ~n4172 ;
  assign n5594 = n5592 | n5593 ;
  assign n5595 = x245 & n4172 ;
  assign n5596 = x503 & ~n4172 ;
  assign n5597 = n5595 | n5596 ;
  assign n5598 = x242 & n4167 ;
  assign n5599 = x504 & ~n4167 ;
  assign n5600 = n5598 | n5599 ;
  assign n5601 = x234 & n4172 ;
  assign n5602 = x505 & ~n4172 ;
  assign n5603 = n5601 | n5602 ;
  assign n5604 = x241 & n4167 ;
  assign n5605 = x506 & ~n4167 ;
  assign n5606 = n5604 | n5605 ;
  assign n5607 = x238 & n4167 ;
  assign n5608 = x507 & ~n4167 ;
  assign n5609 = n5607 | n5608 ;
  assign n5610 = x247 & n4167 ;
  assign n5611 = x508 & ~n4167 ;
  assign n5612 = n5610 | n5611 ;
  assign n5613 = x245 & n4167 ;
  assign n5614 = x509 & ~n4167 ;
  assign n5615 = n5613 | n5614 ;
  assign n5616 = x242 & n4136 ;
  assign n5617 = x510 & ~n4136 ;
  assign n5618 = n5616 | n5617 ;
  assign n5619 = x234 & n4136 ;
  assign n5620 = x511 & ~n4136 ;
  assign n5621 = n5619 | n5620 ;
  assign n5622 = x235 & n4136 ;
  assign n5623 = x512 & ~n4136 ;
  assign n5624 = n5622 | n5623 ;
  assign n5625 = x244 & n4136 ;
  assign n5626 = x513 & ~n4136 ;
  assign n5627 = n5625 | n5626 ;
  assign n5628 = x245 & n4136 ;
  assign n5629 = x514 & ~n4136 ;
  assign n5630 = n5628 | n5629 ;
  assign n5631 = x240 & n4136 ;
  assign n5632 = x515 & ~n4136 ;
  assign n5633 = n5631 | n5632 ;
  assign n5634 = x247 & n4136 ;
  assign n5635 = x516 & ~n4136 ;
  assign n5636 = n5634 | n5635 ;
  assign n5637 = x238 & n4136 ;
  assign n5638 = x517 & ~n4136 ;
  assign n5639 = n5637 | n5638 ;
  assign n5640 = x234 & n4151 ;
  assign n5641 = x518 & ~n4151 ;
  assign n5642 = n5640 | n5641 ;
  assign n5643 = ~x239 & n4151 ;
  assign n5644 = x519 & ~n4151 ;
  assign n5645 = n5643 | n5644 ;
  assign n5646 = x246 & n4151 ;
  assign n5647 = x520 & ~n4151 ;
  assign n5648 = n5646 | n5647 ;
  assign n5649 = x248 & n4151 ;
  assign n5650 = x521 & ~n4151 ;
  assign n5651 = n5649 | n5650 ;
  assign n5652 = x238 & n4151 ;
  assign n5653 = x522 & ~n4151 ;
  assign n5654 = n5652 | n5653 ;
  assign n5655 = x234 & n4251 ;
  assign n5656 = x523 & ~n4251 ;
  assign n5657 = n5655 | n5656 ;
  assign n5658 = ~x239 & n4251 ;
  assign n5659 = x524 & ~n4251 ;
  assign n5660 = n5658 | n5659 ;
  assign n5661 = x245 & n4251 ;
  assign n5662 = x525 & ~n4251 ;
  assign n5663 = n5661 | n5662 ;
  assign n5664 = x246 & n4251 ;
  assign n5665 = x526 & ~n4251 ;
  assign n5666 = n5664 | n5665 ;
  assign n5667 = x247 & n4251 ;
  assign n5668 = x527 & ~n4251 ;
  assign n5669 = n5667 | n5668 ;
  assign n5670 = x249 & n4251 ;
  assign n5671 = x528 & ~n4251 ;
  assign n5672 = n5670 | n5671 ;
  assign n5673 = x238 & n4251 ;
  assign n5674 = x529 & ~n4251 ;
  assign n5675 = n5673 | n5674 ;
  assign n5676 = x240 & n4251 ;
  assign n5677 = x530 & ~n4251 ;
  assign n5678 = n5676 | n5677 ;
  assign n5679 = x235 & n4160 ;
  assign n5680 = x531 & ~n4160 ;
  assign n5681 = n5679 | n5680 ;
  assign n5682 = x247 & n4160 ;
  assign n5683 = x532 & ~n4160 ;
  assign n5684 = n5682 | n5683 ;
  assign n5685 = x235 & n4167 ;
  assign n5686 = x533 & ~n4167 ;
  assign n5687 = n5685 | n5686 ;
  assign n5688 = ~x239 & n4167 ;
  assign n5689 = x534 & ~n4167 ;
  assign n5690 = n5688 | n5689 ;
  assign n5691 = x240 & n4167 ;
  assign n5692 = x535 & ~n4167 ;
  assign n5693 = n5691 | n5692 ;
  assign n5694 = x246 & n4167 ;
  assign n5695 = x536 & ~n4167 ;
  assign n5696 = n5694 | n5695 ;
  assign n5697 = x248 & n4167 ;
  assign n5698 = x537 & ~n4167 ;
  assign n5699 = n5697 | n5698 ;
  assign n5700 = x249 & n4167 ;
  assign n5701 = x538 & ~n4167 ;
  assign n5702 = n5700 | n5701 ;
  assign n5703 = x242 & n4172 ;
  assign n5704 = x539 & ~n4172 ;
  assign n5705 = n5703 | n5704 ;
  assign n5706 = x235 & n4172 ;
  assign n5707 = x540 & ~n4172 ;
  assign n5708 = n5706 | n5707 ;
  assign n5709 = x244 & n4172 ;
  assign n5710 = x541 & ~n4172 ;
  assign n5711 = n5709 | n5710 ;
  assign n5712 = x240 & n4172 ;
  assign n5713 = x542 & ~n4172 ;
  assign n5714 = n5712 | n5713 ;
  assign n5715 = x238 & n4172 ;
  assign n5716 = x543 & ~n4172 ;
  assign n5717 = n5715 | n5716 ;
  assign n5718 = x234 & n4179 ;
  assign n5719 = x544 & ~n4179 ;
  assign n5720 = n5718 | n5719 ;
  assign n5721 = x245 & n4179 ;
  assign n5722 = x545 & ~n4179 ;
  assign n5723 = n5721 | n5722 ;
  assign n5724 = x246 & n4179 ;
  assign n5725 = x546 & ~n4179 ;
  assign n5726 = n5724 | n5725 ;
  assign n5727 = x247 & n4179 ;
  assign n5728 = x547 & ~n4179 ;
  assign n5729 = n5727 | n5728 ;
  assign n5730 = x248 & n4179 ;
  assign n5731 = x548 & ~n4179 ;
  assign n5732 = n5730 | n5731 ;
  assign n5733 = x235 & n4241 ;
  assign n5734 = x549 & ~n4241 ;
  assign n5735 = n5733 | n5734 ;
  assign n5736 = ~x239 & n4241 ;
  assign n5737 = x550 & ~n4241 ;
  assign n5738 = n5736 | n5737 ;
  assign n5739 = x240 & n4241 ;
  assign n5740 = x551 & ~n4241 ;
  assign n5741 = n5739 | n5740 ;
  assign n5742 = x247 & n4241 ;
  assign n5743 = x552 & ~n4241 ;
  assign n5744 = n5742 | n5743 ;
  assign n5745 = x241 & n4241 ;
  assign n5746 = x553 & ~n4241 ;
  assign n5747 = n5745 | n5746 ;
  assign n5748 = x248 & n4241 ;
  assign n5749 = x554 & ~n4241 ;
  assign n5750 = n5748 | n5749 ;
  assign n5751 = x249 & n4241 ;
  assign n5752 = x555 & ~n4241 ;
  assign n5753 = n5751 | n5752 ;
  assign n5754 = x242 & n4160 ;
  assign n5755 = x556 & ~n4160 ;
  assign n5756 = n5754 | n5755 ;
  assign n5757 = x234 & n4167 ;
  assign n5758 = x557 & ~n4167 ;
  assign n5759 = n5757 | n5758 ;
  assign n5760 = x244 & n4167 ;
  assign n5761 = x558 & ~n4167 ;
  assign n5762 = n5760 | n5761 ;
  assign n5763 = x241 & n4136 ;
  assign n5764 = x559 & ~n4136 ;
  assign n5765 = n5763 | n5764 ;
  assign n5766 = x240 & n4160 ;
  assign n5767 = x560 & ~n4160 ;
  assign n5768 = n5766 | n5767 ;
  assign n5769 = x247 & n4151 ;
  assign n5770 = x561 & ~n4151 ;
  assign n5771 = n5769 | n5770 ;
  assign n5772 = x241 & n4160 ;
  assign n5773 = x562 & ~n4160 ;
  assign n5774 = n5772 | n5773 ;
  assign n5775 = x246 & n4241 ;
  assign n5776 = x563 & ~n4241 ;
  assign n5777 = n5775 | n5776 ;
  assign n5778 = x246 & n4160 ;
  assign n5779 = x564 & ~n4160 ;
  assign n5780 = n5778 | n5779 ;
  assign n5781 = x248 & n4160 ;
  assign n5782 = x565 & ~n4160 ;
  assign n5783 = n5781 | n5782 ;
  assign n5784 = x244 & n4160 ;
  assign n5785 = x566 & ~n4160 ;
  assign n5786 = n5784 | n5785 ;
  assign n5787 = x230 & n1430 ;
  assign n5788 = n3823 & n3824 ;
  assign n5789 = ( n3773 & ~n3775 ) | ( n3773 & n5788 ) | ( ~n3775 & n5788 ) ;
  assign n5790 = n5787 & n5789 ;
  assign n5791 = x567 | n5787 ;
  assign n5792 = ( x1092 & n5790 ) | ( x1092 & ~n5791 ) | ( n5790 & ~n5791 ) ;
  assign n5793 = x245 & n4160 ;
  assign n5794 = x568 & ~n4160 ;
  assign n5795 = n5793 | n5794 ;
  assign n5796 = ~x239 & n4160 ;
  assign n5797 = x569 & ~n4160 ;
  assign n5798 = n5796 | n5797 ;
  assign n5799 = x234 & n4160 ;
  assign n5800 = x570 & ~n4160 ;
  assign n5801 = n5799 | n5800 ;
  assign n5802 = x241 & n4251 ;
  assign n5803 = x571 & ~n4251 ;
  assign n5804 = n5802 | n5803 ;
  assign n5805 = x244 & n4251 ;
  assign n5806 = x572 & ~n4251 ;
  assign n5807 = n5805 | n5806 ;
  assign n5808 = x242 & n4251 ;
  assign n5809 = x573 & ~n4251 ;
  assign n5810 = n5808 | n5809 ;
  assign n5811 = x241 & n4151 ;
  assign n5812 = x574 & ~n4151 ;
  assign n5813 = n5811 | n5812 ;
  assign n5814 = x235 & n4251 ;
  assign n5815 = x575 & ~n4251 ;
  assign n5816 = n5814 | n5815 ;
  assign n5817 = x248 & n4251 ;
  assign n5818 = x576 & ~n4251 ;
  assign n5819 = n5817 | n5818 ;
  assign n5820 = x238 & n4241 ;
  assign n5821 = x577 & ~n4241 ;
  assign n5822 = n5820 | n5821 ;
  assign n5823 = x249 & n4151 ;
  assign n5824 = x578 & ~n4151 ;
  assign n5825 = n5823 | n5824 ;
  assign n5826 = x249 & n4136 ;
  assign n5827 = x579 & ~n4136 ;
  assign n5828 = n5826 | n5827 ;
  assign n5829 = x245 & n4241 ;
  assign n5830 = x580 & ~n4241 ;
  assign n5831 = n5829 | n5830 ;
  assign n5832 = x235 & n4151 ;
  assign n5833 = x581 & ~n4151 ;
  assign n5834 = n5832 | n5833 ;
  assign n5835 = x240 & n4151 ;
  assign n5836 = x582 & ~n4151 ;
  assign n5837 = n5835 | n5836 ;
  assign n5838 = x245 & n4151 ;
  assign n5839 = x584 & ~n4151 ;
  assign n5840 = n5838 | n5839 ;
  assign n5841 = x244 & n4151 ;
  assign n5842 = x585 & ~n4151 ;
  assign n5843 = n5841 | n5842 ;
  assign n5844 = x242 & n4151 ;
  assign n5845 = x586 & ~n4151 ;
  assign n5846 = n5844 | n5845 ;
  assign n5847 = ~x230 & x587 ;
  assign n5848 = x230 | x587 ;
  assign n5849 = ( n3775 & n5847 ) | ( n3775 & n5848 ) | ( n5847 & n5848 ) ;
  assign n5850 = ~x123 & x824 ;
  assign n5851 = x950 & n5850 ;
  assign n5852 = x588 & ~n5851 ;
  assign n5853 = x591 & n5851 ;
  assign n5854 = ( n5047 & n5852 ) | ( n5047 & n5853 ) | ( n5852 & n5853 ) ;
  assign n5855 = x201 & x233 ;
  assign n5856 = x202 & ~x233 ;
  assign n5857 = ( x237 & n5855 ) | ( x237 & n5856 ) | ( n5855 & n5856 ) ;
  assign n5858 = x203 & ~x233 ;
  assign n5859 = x220 & x233 ;
  assign n5860 = ( ~x237 & n5858 ) | ( ~x237 & n5859 ) | ( n5858 & n5859 ) ;
  assign n5861 = n5857 | n5860 ;
  assign n5862 = n2105 & ~n5861 ;
  assign n5863 = x218 & ~x237 ;
  assign n5864 = x205 & x237 ;
  assign n5865 = ( ~x233 & n5863 ) | ( ~x233 & n5864 ) | ( n5863 & n5864 ) ;
  assign n5866 = x206 & ~x237 ;
  assign n5867 = x204 & x237 ;
  assign n5868 = ( x233 & n5866 ) | ( x233 & n5867 ) | ( n5866 & n5867 ) ;
  assign n5869 = n5865 | n5868 ;
  assign n5870 = n2037 | n5869 ;
  assign n5871 = ( n5862 & ~n5869 ) | ( n5862 & n5870 ) | ( ~n5869 & n5870 ) ;
  assign n5872 = ~x588 & n5851 ;
  assign n5873 = x590 | n5851 ;
  assign n5874 = ( n5047 & n5872 ) | ( n5047 & ~n5873 ) | ( n5872 & ~n5873 ) ;
  assign n5875 = x591 & ~n5851 ;
  assign n5876 = x592 & n5851 ;
  assign n5877 = ( n5047 & n5875 ) | ( n5047 & n5876 ) | ( n5875 & n5876 ) ;
  assign n5878 = x592 & ~n5851 ;
  assign n5879 = x590 & n5851 ;
  assign n5880 = ( n5047 & n5878 ) | ( n5047 & n5879 ) | ( n5878 & n5879 ) ;
  assign n5881 = x235 & ~x549 ;
  assign n5882 = ( x242 & ~x489 ) | ( x242 & n5881 ) | ( ~x489 & n5881 ) ;
  assign n5883 = ~x238 & x577 ;
  assign n5884 = ( ~x242 & x489 ) | ( ~x242 & n5883 ) | ( x489 & n5883 ) ;
  assign n5885 = n5882 | n5884 ;
  assign n5886 = ( x245 & ~x580 ) | ( x245 & n5885 ) | ( ~x580 & n5885 ) ;
  assign n5887 = ~x246 & x563 ;
  assign n5888 = ( ~x245 & x580 ) | ( ~x245 & n5887 ) | ( x580 & n5887 ) ;
  assign n5889 = n5886 | n5888 ;
  assign n5890 = x241 & ~x553 ;
  assign n5891 = ~x247 & x552 ;
  assign n5892 = x248 & ~x554 ;
  assign n5893 = ( ~n4158 & n5891 ) | ( ~n4158 & n5892 ) | ( n5891 & n5892 ) ;
  assign n5894 = ( ~n4158 & n5890 ) | ( ~n4158 & n5893 ) | ( n5890 & n5893 ) ;
  assign n5895 = n4158 | n5894 ;
  assign n5896 = x244 & ~x486 ;
  assign n5897 = x239 & x550 ;
  assign n5898 = x246 & ~x563 ;
  assign n5899 = ( ~n5896 & n5897 ) | ( ~n5896 & n5898 ) | ( n5897 & n5898 ) ;
  assign n5900 = x238 & ~x577 ;
  assign n5901 = ( ~n5896 & n5899 ) | ( ~n5896 & n5900 ) | ( n5899 & n5900 ) ;
  assign n5902 = n5896 | n5901 ;
  assign n5903 = x240 & ~x551 ;
  assign n5904 = ~x235 & x549 ;
  assign n5905 = ~x241 & x553 ;
  assign n5906 = x247 & ~x552 ;
  assign n5907 = ( ~n5903 & n5905 ) | ( ~n5903 & n5906 ) | ( n5905 & n5906 ) ;
  assign n5908 = ( ~n5903 & n5904 ) | ( ~n5903 & n5907 ) | ( n5904 & n5907 ) ;
  assign n5909 = n5903 | n5908 ;
  assign n5910 = ~x240 & x551 ;
  assign n5911 = ~x248 & x554 ;
  assign n5912 = x239 | x550 ;
  assign n5913 = ~x244 & x486 ;
  assign n5914 = ( n5910 & n5912 ) | ( n5910 & ~n5913 ) | ( n5912 & ~n5913 ) ;
  assign n5915 = ( n5910 & ~n5911 ) | ( n5910 & n5914 ) | ( ~n5911 & n5914 ) ;
  assign n5916 = ~n5910 & n5915 ;
  assign n5917 = ( n5895 & ~n5909 ) | ( n5895 & n5916 ) | ( ~n5909 & n5916 ) ;
  assign n5918 = ( n5895 & ~n5902 ) | ( n5895 & n5917 ) | ( ~n5902 & n5917 ) ;
  assign n5919 = ~n5895 & n5918 ;
  assign n5920 = ~x249 & x555 ;
  assign n5921 = ( ~x234 & x485 ) | ( ~x234 & n5920 ) | ( x485 & n5920 ) ;
  assign n5922 = x249 & ~x555 ;
  assign n5923 = ( x234 & ~x485 ) | ( x234 & n5922 ) | ( ~x485 & n5922 ) ;
  assign n5924 = n5921 | n5923 ;
  assign n5925 = ( n2037 & ~n5919 ) | ( n2037 & n5924 ) | ( ~n5919 & n5924 ) ;
  assign n5926 = ( n2037 & n5889 ) | ( n2037 & n5925 ) | ( n5889 & n5925 ) ;
  assign n5927 = n2037 & ~n5926 ;
  assign n5928 = ( x247 & ~x508 ) | ( x247 & n4132 ) | ( ~x508 & n4132 ) ;
  assign n5929 = ~x244 & x558 ;
  assign n5930 = ( x247 & ~x508 ) | ( x247 & n5929 ) | ( ~x508 & n5929 ) ;
  assign n5931 = n5928 & ~n5930 ;
  assign n5932 = x241 & ~x506 ;
  assign n5933 = ( x248 & ~x537 ) | ( x248 & n5932 ) | ( ~x537 & n5932 ) ;
  assign n5934 = ~x242 & x504 ;
  assign n5935 = ( ~x248 & x537 ) | ( ~x248 & n5934 ) | ( x537 & n5934 ) ;
  assign n5936 = n5933 | n5935 ;
  assign n5937 = n5931 & ~n5936 ;
  assign n5938 = x239 & x534 ;
  assign n5939 = ( x249 & ~x538 ) | ( x249 & n5938 ) | ( ~x538 & n5938 ) ;
  assign n5940 = n5937 & ~n5939 ;
  assign n5941 = x235 & ~x533 ;
  assign n5942 = ( x238 & ~x507 ) | ( x238 & n5941 ) | ( ~x507 & n5941 ) ;
  assign n5943 = ~x234 & x557 ;
  assign n5944 = ( ~x238 & x507 ) | ( ~x238 & n5943 ) | ( x507 & n5943 ) ;
  assign n5945 = n5942 | n5944 ;
  assign n5946 = x234 & ~x557 ;
  assign n5947 = ~x235 & x533 ;
  assign n5948 = x245 & ~x509 ;
  assign n5949 = x242 & ~x504 ;
  assign n5950 = ( ~n5946 & n5948 ) | ( ~n5946 & n5949 ) | ( n5948 & n5949 ) ;
  assign n5951 = ( ~n5946 & n5947 ) | ( ~n5946 & n5950 ) | ( n5947 & n5950 ) ;
  assign n5952 = n5946 | n5951 ;
  assign n5953 = ( n5937 & n5945 ) | ( n5937 & n5952 ) | ( n5945 & n5952 ) ;
  assign n5954 = x244 & ~x558 ;
  assign n5955 = ( x240 & ~x535 ) | ( x240 & n5954 ) | ( ~x535 & n5954 ) ;
  assign n5956 = ~x245 & x509 ;
  assign n5957 = ( ~x240 & x535 ) | ( ~x240 & n5956 ) | ( x535 & n5956 ) ;
  assign n5958 = n5955 | n5957 ;
  assign n5959 = ~x241 & x506 ;
  assign n5960 = ( ~x246 & x536 ) | ( ~x246 & n5959 ) | ( x536 & n5959 ) ;
  assign n5961 = x239 | x534 ;
  assign n5962 = ( ~x246 & x536 ) | ( ~x246 & n5961 ) | ( x536 & n5961 ) ;
  assign n5963 = ~n5960 & n5962 ;
  assign n5964 = ~n5958 & n5963 ;
  assign n5965 = ( x249 & ~x538 ) | ( x249 & n5964 ) | ( ~x538 & n5964 ) ;
  assign n5966 = ( n5940 & n5953 ) | ( n5940 & ~n5965 ) | ( n5953 & ~n5965 ) ;
  assign n5967 = n5940 & ~n5966 ;
  assign n5968 = ~x246 & x499 ;
  assign n5969 = ( x241 & ~x500 ) | ( x241 & n5968 ) | ( ~x500 & n5968 ) ;
  assign n5970 = x245 & ~x503 ;
  assign n5971 = x234 & ~x505 ;
  assign n5972 = ~x244 & x541 ;
  assign n5973 = x246 & ~x499 ;
  assign n5974 = ( ~n5970 & n5972 ) | ( ~n5970 & n5973 ) | ( n5972 & n5973 ) ;
  assign n5975 = ( ~n5970 & n5971 ) | ( ~n5970 & n5974 ) | ( n5971 & n5974 ) ;
  assign n5976 = n5970 | n5975 ;
  assign n5977 = ~n5969 & n5976 ;
  assign n5978 = ~x234 & x505 ;
  assign n5979 = ( x249 & ~x496 ) | ( x249 & n5978 ) | ( ~x496 & n5978 ) ;
  assign n5980 = x244 & ~x541 ;
  assign n5981 = ( ~x249 & x496 ) | ( ~x249 & n5980 ) | ( x496 & n5980 ) ;
  assign n5982 = n5979 | n5981 ;
  assign n5983 = ( x248 & ~x501 ) | ( x248 & n4149 ) | ( ~x501 & n4149 ) ;
  assign n5984 = x239 & x497 ;
  assign n5985 = ( x248 & ~x501 ) | ( x248 & n5984 ) | ( ~x501 & n5984 ) ;
  assign n5986 = n5983 & ~n5985 ;
  assign n5987 = ~x245 & x503 ;
  assign n5988 = ( x238 & ~x543 ) | ( x238 & n5987 ) | ( ~x543 & n5987 ) ;
  assign n5989 = x235 & ~x540 ;
  assign n5990 = ( ~x238 & x543 ) | ( ~x238 & n5989 ) | ( x543 & n5989 ) ;
  assign n5991 = n5988 | n5990 ;
  assign n5992 = n5986 & ~n5991 ;
  assign n5993 = ~n5982 & n5992 ;
  assign n5994 = ( n5969 & ~n5977 ) | ( n5969 & n5993 ) | ( ~n5977 & n5993 ) ;
  assign n5995 = x239 | x497 ;
  assign n5996 = ( x240 & ~x542 ) | ( x240 & n5995 ) | ( ~x542 & n5995 ) ;
  assign n5997 = ~x235 & x540 ;
  assign n5998 = ( x240 & ~x542 ) | ( x240 & n5997 ) | ( ~x542 & n5997 ) ;
  assign n5999 = n5996 & ~n5998 ;
  assign n6000 = ~x247 & x502 ;
  assign n6001 = ( ~x242 & x539 ) | ( ~x242 & n6000 ) | ( x539 & n6000 ) ;
  assign n6002 = x247 & ~x502 ;
  assign n6003 = ( x242 & ~x539 ) | ( x242 & n6002 ) | ( ~x539 & n6002 ) ;
  assign n6004 = n6001 | n6003 ;
  assign n6005 = n5999 & ~n6004 ;
  assign n6006 = ( x241 & ~x500 ) | ( x241 & n6005 ) | ( ~x500 & n6005 ) ;
  assign n6007 = ( n5969 & n5994 ) | ( n5969 & ~n6006 ) | ( n5994 & ~n6006 ) ;
  assign n6008 = ( n5967 & n5994 ) | ( n5967 & ~n6007 ) | ( n5994 & ~n6007 ) ;
  assign n6009 = x249 & ~x484 ;
  assign n6010 = ( x245 & ~x545 ) | ( x245 & n6009 ) | ( ~x545 & n6009 ) ;
  assign n6011 = ~x248 & x548 ;
  assign n6012 = ( ~x245 & x545 ) | ( ~x245 & n6011 ) | ( x545 & n6011 ) ;
  assign n6013 = n6010 | n6012 ;
  assign n6014 = ~x238 & x491 ;
  assign n6015 = ( x244 & ~x493 ) | ( x244 & n6014 ) | ( ~x493 & n6014 ) ;
  assign n6016 = x248 & ~x548 ;
  assign n6017 = ( ~x244 & x493 ) | ( ~x244 & n6016 ) | ( x493 & n6016 ) ;
  assign n6018 = n6015 | n6017 ;
  assign n6019 = n6013 | n6018 ;
  assign n6020 = ( ~x246 & x546 ) | ( ~x246 & n6019 ) | ( x546 & n6019 ) ;
  assign n6021 = ~x249 & x484 ;
  assign n6022 = ( x246 & ~x546 ) | ( x246 & n6021 ) | ( ~x546 & n6021 ) ;
  assign n6023 = n6020 | n6022 ;
  assign n6024 = ~x235 & x495 ;
  assign n6025 = ( x241 & ~x490 ) | ( x241 & n6024 ) | ( ~x490 & n6024 ) ;
  assign n6026 = x239 & x494 ;
  assign n6027 = ( ~x241 & x490 ) | ( ~x241 & n6026 ) | ( x490 & n6026 ) ;
  assign n6028 = n6025 | n6027 ;
  assign n6029 = x240 & ~x492 ;
  assign n6030 = ( x234 & ~x544 ) | ( x234 & n6029 ) | ( ~x544 & n6029 ) ;
  assign n6031 = x247 & ~x547 ;
  assign n6032 = ( ~x234 & x544 ) | ( ~x234 & n6031 ) | ( x544 & n6031 ) ;
  assign n6033 = n6030 | n6032 ;
  assign n6034 = n6028 | n6033 ;
  assign n6035 = ~x242 & x483 ;
  assign n6036 = x235 & ~x495 ;
  assign n6037 = ( n4177 & n6035 ) | ( n4177 & n6036 ) | ( n6035 & n6036 ) ;
  assign n6038 = x238 & ~x491 ;
  assign n6039 = ( n4177 & n6037 ) | ( n4177 & n6038 ) | ( n6037 & n6038 ) ;
  assign n6040 = n4177 & ~n6039 ;
  assign n6041 = ~x247 & x547 ;
  assign n6042 = x239 | x494 ;
  assign n6043 = ~x240 & x492 ;
  assign n6044 = x242 & ~x483 ;
  assign n6045 = ( ~n6041 & n6043 ) | ( ~n6041 & n6044 ) | ( n6043 & n6044 ) ;
  assign n6046 = ( n6041 & n6042 ) | ( n6041 & ~n6045 ) | ( n6042 & ~n6045 ) ;
  assign n6047 = ~n6041 & n6046 ;
  assign n6048 = ( n6034 & n6040 ) | ( n6034 & n6047 ) | ( n6040 & n6047 ) ;
  assign n6049 = ~n6034 & n6048 ;
  assign n6050 = ~n6023 & n6049 ;
  assign n6051 = n6008 | n6050 ;
  assign n6052 = ( n2037 & n5927 ) | ( n2037 & n6051 ) | ( n5927 & n6051 ) ;
  assign n6053 = ( x234 & ~x518 ) | ( x234 & n4149 ) | ( ~x518 & n4149 ) ;
  assign n6054 = x244 & ~x585 ;
  assign n6055 = ( x234 & ~x518 ) | ( x234 & n6054 ) | ( ~x518 & n6054 ) ;
  assign n6056 = n6053 & ~n6055 ;
  assign n6057 = x240 & ~x582 ;
  assign n6058 = ( ~x248 & x521 ) | ( ~x248 & n6057 ) | ( x521 & n6057 ) ;
  assign n6059 = x239 | x519 ;
  assign n6060 = ( ~x248 & x521 ) | ( ~x248 & n6059 ) | ( x521 & n6059 ) ;
  assign n6061 = ~n6058 & n6060 ;
  assign n6062 = n6056 & n6061 ;
  assign n6063 = x239 & x519 ;
  assign n6064 = ( x235 & ~x581 ) | ( x235 & n6063 ) | ( ~x581 & n6063 ) ;
  assign n6065 = n6062 & ~n6064 ;
  assign n6066 = ~x249 & x578 ;
  assign n6067 = ( ~x245 & x584 ) | ( ~x245 & n6066 ) | ( x584 & n6066 ) ;
  assign n6068 = x249 & ~x578 ;
  assign n6069 = ( x245 & ~x584 ) | ( x245 & n6068 ) | ( ~x584 & n6068 ) ;
  assign n6070 = n6067 | n6069 ;
  assign n6071 = x247 & ~x561 ;
  assign n6072 = ~x238 & x522 ;
  assign n6073 = ~x246 & x520 ;
  assign n6074 = ( ~n6071 & n6072 ) | ( ~n6071 & n6073 ) | ( n6072 & n6073 ) ;
  assign n6075 = ~x240 & x582 ;
  assign n6076 = ( ~n6071 & n6074 ) | ( ~n6071 & n6075 ) | ( n6074 & n6075 ) ;
  assign n6077 = n6071 | n6076 ;
  assign n6078 = ( n6062 & n6070 ) | ( n6062 & n6077 ) | ( n6070 & n6077 ) ;
  assign n6079 = ~x244 & x585 ;
  assign n6080 = ( x242 & ~x586 ) | ( x242 & n6079 ) | ( ~x586 & n6079 ) ;
  assign n6081 = x238 & ~x522 ;
  assign n6082 = ( ~x242 & x586 ) | ( ~x242 & n6081 ) | ( x586 & n6081 ) ;
  assign n6083 = n6080 | n6082 ;
  assign n6084 = x246 & ~x520 ;
  assign n6085 = ( x241 & ~x574 ) | ( x241 & n6084 ) | ( ~x574 & n6084 ) ;
  assign n6086 = ~x247 & x561 ;
  assign n6087 = ( ~x241 & x574 ) | ( ~x241 & n6086 ) | ( x574 & n6086 ) ;
  assign n6088 = n6085 | n6087 ;
  assign n6089 = n6083 | n6088 ;
  assign n6090 = ( ~x235 & x581 ) | ( ~x235 & n6089 ) | ( x581 & n6089 ) ;
  assign n6091 = ( n6065 & n6078 ) | ( n6065 & n6090 ) | ( n6078 & n6090 ) ;
  assign n6092 = n6065 & ~n6091 ;
  assign n6093 = ( x242 & ~x573 ) | ( x242 & n4177 ) | ( ~x573 & n4177 ) ;
  assign n6094 = x235 & ~x575 ;
  assign n6095 = ( x242 & ~x573 ) | ( x242 & n6094 ) | ( ~x573 & n6094 ) ;
  assign n6096 = n6093 & ~n6095 ;
  assign n6097 = x239 | x524 ;
  assign n6098 = ( x248 & ~x576 ) | ( x248 & n6097 ) | ( ~x576 & n6097 ) ;
  assign n6099 = ~x246 & x526 ;
  assign n6100 = ( x248 & ~x576 ) | ( x248 & n6099 ) | ( ~x576 & n6099 ) ;
  assign n6101 = n6098 & ~n6100 ;
  assign n6102 = ~x244 & x572 ;
  assign n6103 = ( x245 & ~x525 ) | ( x245 & n6102 ) | ( ~x525 & n6102 ) ;
  assign n6104 = x239 & x524 ;
  assign n6105 = ( ~x245 & x525 ) | ( ~x245 & n6104 ) | ( x525 & n6104 ) ;
  assign n6106 = n6103 | n6105 ;
  assign n6107 = ( n6096 & ~n6101 ) | ( n6096 & n6106 ) | ( ~n6101 & n6106 ) ;
  assign n6108 = ~x235 & x575 ;
  assign n6109 = ( x247 & ~x527 ) | ( x247 & n6108 ) | ( ~x527 & n6108 ) ;
  assign n6110 = ~x238 & x529 ;
  assign n6111 = ( ~x247 & x527 ) | ( ~x247 & n6110 ) | ( x527 & n6110 ) ;
  assign n6112 = n6109 | n6111 ;
  assign n6113 = ( n6096 & n6107 ) | ( n6096 & n6112 ) | ( n6107 & n6112 ) ;
  assign n6114 = n6096 & ~n6113 ;
  assign n6115 = ~x234 & x523 ;
  assign n6116 = ( x240 & ~x530 ) | ( x240 & n6115 ) | ( ~x530 & n6115 ) ;
  assign n6117 = n6114 | n6116 ;
  assign n6118 = ~x241 & x571 ;
  assign n6119 = x238 & ~x529 ;
  assign n6120 = x244 & ~x572 ;
  assign n6121 = x246 & ~x526 ;
  assign n6122 = ( ~n6118 & n6120 ) | ( ~n6118 & n6121 ) | ( n6120 & n6121 ) ;
  assign n6123 = ( ~n6118 & n6119 ) | ( ~n6118 & n6122 ) | ( n6119 & n6122 ) ;
  assign n6124 = n6118 | n6123 ;
  assign n6125 = x241 & ~x571 ;
  assign n6126 = ( x249 & ~x528 ) | ( x249 & n6125 ) | ( ~x528 & n6125 ) ;
  assign n6127 = x234 & ~x523 ;
  assign n6128 = ( ~x249 & x528 ) | ( ~x249 & n6127 ) | ( x528 & n6127 ) ;
  assign n6129 = n6126 | n6128 ;
  assign n6130 = n6124 | n6129 ;
  assign n6131 = ( ~x240 & x530 ) | ( ~x240 & n6130 ) | ( x530 & n6130 ) ;
  assign n6132 = ( n6116 & n6117 ) | ( n6116 & n6131 ) | ( n6117 & n6131 ) ;
  assign n6133 = ( n6092 & n6117 ) | ( n6092 & ~n6132 ) | ( n6117 & ~n6132 ) ;
  assign n6134 = ~x235 & x531 ;
  assign n6135 = ( x242 & ~x556 ) | ( x242 & n6134 ) | ( ~x556 & n6134 ) ;
  assign n6136 = x247 & ~x532 ;
  assign n6137 = ( ~x242 & x556 ) | ( ~x242 & n6136 ) | ( x556 & n6136 ) ;
  assign n6138 = n6135 | n6137 ;
  assign n6139 = ~x238 & x498 ;
  assign n6140 = ( x246 & ~x564 ) | ( x246 & n6139 ) | ( ~x564 & n6139 ) ;
  assign n6141 = x244 & ~x566 ;
  assign n6142 = ( ~x246 & x564 ) | ( ~x246 & n6141 ) | ( x564 & n6141 ) ;
  assign n6143 = n6140 | n6142 ;
  assign n6144 = ~x244 & x566 ;
  assign n6145 = ( x245 & ~x568 ) | ( x245 & n6144 ) | ( ~x568 & n6144 ) ;
  assign n6146 = x248 & ~x565 ;
  assign n6147 = ( ~x245 & x568 ) | ( ~x245 & n6146 ) | ( x568 & n6146 ) ;
  assign n6148 = n6145 | n6147 ;
  assign n6149 = ( ~n6138 & n6143 ) | ( ~n6138 & n6148 ) | ( n6143 & n6148 ) ;
  assign n6150 = ( x241 & ~x562 ) | ( x241 & n4158 ) | ( ~x562 & n4158 ) ;
  assign n6151 = x238 & ~x498 ;
  assign n6152 = ( ~x241 & x562 ) | ( ~x241 & n6151 ) | ( x562 & n6151 ) ;
  assign n6153 = n6150 | n6152 ;
  assign n6154 = ( ~n6138 & n6149 ) | ( ~n6138 & n6153 ) | ( n6149 & n6153 ) ;
  assign n6155 = n6138 | n6154 ;
  assign n6156 = ~x240 & x560 ;
  assign n6157 = ( x239 & x569 ) | ( x239 & n6156 ) | ( x569 & n6156 ) ;
  assign n6158 = x240 & ~x560 ;
  assign n6159 = ( x239 & x569 ) | ( x239 & ~n6158 ) | ( x569 & ~n6158 ) ;
  assign n6160 = ~n6157 & n6159 ;
  assign n6161 = ~x248 & x565 ;
  assign n6162 = ( x234 & ~x570 ) | ( x234 & n6161 ) | ( ~x570 & n6161 ) ;
  assign n6163 = x249 & ~x482 ;
  assign n6164 = ( ~x234 & x570 ) | ( ~x234 & n6163 ) | ( x570 & n6163 ) ;
  assign n6165 = n6162 | n6164 ;
  assign n6166 = ( n6155 & n6160 ) | ( n6155 & ~n6165 ) | ( n6160 & ~n6165 ) ;
  assign n6167 = ~x247 & x532 ;
  assign n6168 = ~x249 & x482 ;
  assign n6169 = x235 & ~x531 ;
  assign n6170 = ( ~n6167 & n6168 ) | ( ~n6167 & n6169 ) | ( n6168 & n6169 ) ;
  assign n6171 = n6167 | n6170 ;
  assign n6172 = ( n6155 & n6166 ) | ( n6155 & ~n6171 ) | ( n6166 & ~n6171 ) ;
  assign n6173 = ~n6155 & n6172 ;
  assign n6174 = x242 & ~x510 ;
  assign n6175 = ( x241 & ~x559 ) | ( x241 & n6174 ) | ( ~x559 & n6174 ) ;
  assign n6176 = n2105 & ~n6175 ;
  assign n6177 = x238 & ~x517 ;
  assign n6178 = ~x244 & x513 ;
  assign n6179 = ( n4132 & n6177 ) | ( n4132 & n6178 ) | ( n6177 & n6178 ) ;
  assign n6180 = ~x242 & x510 ;
  assign n6181 = ( n4132 & n6179 ) | ( n4132 & n6180 ) | ( n6179 & n6180 ) ;
  assign n6182 = n4132 & ~n6181 ;
  assign n6183 = x248 & ~x481 ;
  assign n6184 = ( x240 & ~x515 ) | ( x240 & n6183 ) | ( ~x515 & n6183 ) ;
  assign n6185 = ~x245 & x514 ;
  assign n6186 = ( ~x240 & x515 ) | ( ~x240 & n6185 ) | ( x515 & n6185 ) ;
  assign n6187 = n6184 | n6186 ;
  assign n6188 = x247 & ~x516 ;
  assign n6189 = x234 & ~x511 ;
  assign n6190 = x235 & ~x512 ;
  assign n6191 = ~x248 & x481 ;
  assign n6192 = ( ~n6188 & n6190 ) | ( ~n6188 & n6191 ) | ( n6190 & n6191 ) ;
  assign n6193 = ( ~n6188 & n6189 ) | ( ~n6188 & n6192 ) | ( n6189 & n6192 ) ;
  assign n6194 = n6188 | n6193 ;
  assign n6195 = ( n6182 & n6187 ) | ( n6182 & n6194 ) | ( n6187 & n6194 ) ;
  assign n6196 = ~x235 & x512 ;
  assign n6197 = x245 & ~x514 ;
  assign n6198 = x249 & ~x579 ;
  assign n6199 = x244 & ~x513 ;
  assign n6200 = ( ~n6196 & n6198 ) | ( ~n6196 & n6199 ) | ( n6198 & n6199 ) ;
  assign n6201 = ( ~n6196 & n6197 ) | ( ~n6196 & n6200 ) | ( n6197 & n6200 ) ;
  assign n6202 = n6196 | n6201 ;
  assign n6203 = ( n6182 & n6195 ) | ( n6182 & n6202 ) | ( n6195 & n6202 ) ;
  assign n6204 = n6182 & ~n6203 ;
  assign n6205 = ~x234 & x511 ;
  assign n6206 = ( x246 & ~x487 ) | ( x246 & n6205 ) | ( ~x487 & n6205 ) ;
  assign n6207 = ~x238 & x517 ;
  assign n6208 = ( ~x246 & x487 ) | ( ~x246 & n6207 ) | ( x487 & n6207 ) ;
  assign n6209 = n6206 | n6208 ;
  assign n6210 = ~x249 & x579 ;
  assign n6211 = ( x239 & x488 ) | ( x239 & ~n6210 ) | ( x488 & ~n6210 ) ;
  assign n6212 = ~x247 & x516 ;
  assign n6213 = ( x239 & x488 ) | ( x239 & n6212 ) | ( x488 & n6212 ) ;
  assign n6214 = n6211 & ~n6213 ;
  assign n6215 = ~n6209 & n6214 ;
  assign n6216 = ( x241 & ~x559 ) | ( x241 & n6215 ) | ( ~x559 & n6215 ) ;
  assign n6217 = n6204 & n6216 ;
  assign n6218 = n6176 & n6217 ;
  assign n6219 = ( n2105 & n6173 ) | ( n2105 & n6218 ) | ( n6173 & n6218 ) ;
  assign n6220 = ( n2105 & n6133 ) | ( n2105 & n6219 ) | ( n6133 & n6219 ) ;
  assign n6221 = n6052 | n6220 ;
  assign n6222 = ~x806 & x990 ;
  assign n6223 = x600 & n6222 ;
  assign n6224 = ( x332 & x594 ) | ( x332 & n6223 ) | ( x594 & n6223 ) ;
  assign n6225 = ( ~x332 & x594 ) | ( ~x332 & n6223 ) | ( x594 & n6223 ) ;
  assign n6226 = ~n6224 & n6225 ;
  assign n6227 = ~x806 & n5434 ;
  assign n6228 = ( x595 & ~n5441 ) | ( x595 & n6227 ) | ( ~n5441 & n6227 ) ;
  assign n6229 = n6227 & ~n6228 ;
  assign n6230 = ( x332 & n5441 ) | ( x332 & n6228 ) | ( n5441 & n6228 ) ;
  assign n6231 = ( x595 & n6229 ) | ( x595 & ~n6230 ) | ( n6229 & ~n6230 ) ;
  assign n6232 = n5434 & n6222 ;
  assign n6233 = x595 & x597 ;
  assign n6234 = n6232 & n6233 ;
  assign n6235 = x596 & n6234 ;
  assign n6236 = ( ~x332 & x596 ) | ( ~x332 & n6234 ) | ( x596 & n6234 ) ;
  assign n6237 = ~n6235 & n6236 ;
  assign n6238 = ( ~x332 & x597 ) | ( ~x332 & n6232 ) | ( x597 & n6232 ) ;
  assign n6239 = ( x332 & x597 ) | ( x332 & n6232 ) | ( x597 & n6232 ) ;
  assign n6240 = n6238 & ~n6239 ;
  assign n6241 = x740 & x780 ;
  assign n6242 = n1981 & n6241 ;
  assign n6243 = x598 | n6242 ;
  assign n6244 = x882 | n1208 ;
  assign n6245 = x947 & ~n6244 ;
  assign n6246 = ( n6242 & n6243 ) | ( n6242 & ~n6245 ) | ( n6243 & ~n6245 ) ;
  assign n6247 = ( x332 & x599 ) | ( x332 & n6235 ) | ( x599 & n6235 ) ;
  assign n6248 = ( ~x332 & x599 ) | ( ~x332 & n6235 ) | ( x599 & n6235 ) ;
  assign n6249 = ~n6247 & n6248 ;
  assign n6250 = ( ~x332 & x600 ) | ( ~x332 & n6222 ) | ( x600 & n6222 ) ;
  assign n6251 = ~n6223 & n6250 ;
  assign n6252 = ~x806 & x989 ;
  assign n6253 = x601 & x806 ;
  assign n6254 = ( ~x332 & n6252 ) | ( ~x332 & n6253 ) | ( n6252 & n6253 ) ;
  assign n6255 = ~x230 & x602 ;
  assign n6256 = x230 | x602 ;
  assign n6257 = ( n3825 & n6255 ) | ( n3825 & n6256 ) | ( n6255 & n6256 ) ;
  assign n6258 = ~x872 & x966 ;
  assign n6259 = ~x871 & n6258 ;
  assign n6260 = x1038 & x1060 ;
  assign n6261 = x980 | x1061 ;
  assign n6262 = n6260 & ~n6261 ;
  assign n6263 = x832 & x952 ;
  assign n6264 = n6262 & n6263 ;
  assign n6265 = x603 | n6264 ;
  assign n6266 = ~x1100 & n6264 ;
  assign n6267 = ( x966 & n6265 ) | ( x966 & ~n6266 ) | ( n6265 & ~n6266 ) ;
  assign n6268 = ~n6259 & n6267 ;
  assign n6269 = ~x681 & x823 ;
  assign n6270 = ~n1983 & n6269 ;
  assign n6271 = x779 & n6270 ;
  assign n6272 = x604 & ~x907 ;
  assign n6273 = ~x299 & x983 ;
  assign n6274 = ( x604 & n6272 ) | ( x604 & ~n6273 ) | ( n6272 & ~n6273 ) ;
  assign n6275 = ~n6270 & n6274 ;
  assign n6276 = ( n6270 & ~n6271 ) | ( n6270 & n6275 ) | ( ~n6271 & n6275 ) ;
  assign n6277 = ( x332 & ~x605 ) | ( x332 & x806 ) | ( ~x605 & x806 ) ;
  assign n6278 = ( x332 & x605 ) | ( x332 & ~x806 ) | ( x605 & ~x806 ) ;
  assign n6279 = n6277 | n6278 ;
  assign n6280 = ~x1104 & n6264 ;
  assign n6281 = x837 & x966 ;
  assign n6282 = x606 | n6264 ;
  assign n6283 = ( ~x966 & n6281 ) | ( ~x966 & n6282 ) | ( n6281 & n6282 ) ;
  assign n6284 = ( ~n6280 & n6281 ) | ( ~n6280 & n6283 ) | ( n6281 & n6283 ) ;
  assign n6285 = x1107 & n6264 ;
  assign n6286 = x607 & ~n6264 ;
  assign n6287 = ( ~x966 & n6285 ) | ( ~x966 & n6286 ) | ( n6285 & n6286 ) ;
  assign n6288 = x608 & ~n6264 ;
  assign n6289 = x1116 & n6264 ;
  assign n6290 = ( ~x966 & n6288 ) | ( ~x966 & n6289 ) | ( n6288 & n6289 ) ;
  assign n6291 = x1118 & n6264 ;
  assign n6292 = x609 & ~n6264 ;
  assign n6293 = ( ~x966 & n6291 ) | ( ~x966 & n6292 ) | ( n6291 & n6292 ) ;
  assign n6294 = x1113 & n6264 ;
  assign n6295 = x610 & ~n6264 ;
  assign n6296 = ( ~x966 & n6294 ) | ( ~x966 & n6295 ) | ( n6294 & n6295 ) ;
  assign n6297 = x611 & ~n6264 ;
  assign n6298 = x1114 & n6264 ;
  assign n6299 = ( ~x966 & n6297 ) | ( ~x966 & n6298 ) | ( n6297 & n6298 ) ;
  assign n6300 = x1111 & n6264 ;
  assign n6301 = x612 & ~n6264 ;
  assign n6302 = ( ~x966 & n6300 ) | ( ~x966 & n6301 ) | ( n6300 & n6301 ) ;
  assign n6303 = x613 & ~n6264 ;
  assign n6304 = x1115 & n6264 ;
  assign n6305 = ( ~x966 & n6303 ) | ( ~x966 & n6304 ) | ( n6303 & n6304 ) ;
  assign n6306 = x871 & x966 ;
  assign n6307 = ~x1102 & n6264 ;
  assign n6308 = x614 | n6264 ;
  assign n6309 = ( ~x966 & n6306 ) | ( ~x966 & n6308 ) | ( n6306 & n6308 ) ;
  assign n6310 = ( n6306 & ~n6307 ) | ( n6306 & n6309 ) | ( ~n6307 & n6309 ) ;
  assign n6311 = x779 & x797 ;
  assign n6312 = n1985 & n6311 ;
  assign n6313 = x615 & ~n6312 ;
  assign n6314 = x907 & ~n6244 ;
  assign n6315 = ( ~n6312 & n6313 ) | ( ~n6312 & n6314 ) | ( n6313 & n6314 ) ;
  assign n6316 = ~x1101 & n6264 ;
  assign n6317 = x872 & x966 ;
  assign n6318 = x616 & ~n6258 ;
  assign n6319 = ( ~n6258 & n6264 ) | ( ~n6258 & n6318 ) | ( n6264 & n6318 ) ;
  assign n6320 = ( ~n6316 & n6317 ) | ( ~n6316 & n6319 ) | ( n6317 & n6319 ) ;
  assign n6321 = x617 | n6264 ;
  assign n6322 = x850 & x966 ;
  assign n6323 = ~x1105 & n6264 ;
  assign n6324 = ( x966 & ~n6322 ) | ( x966 & n6323 ) | ( ~n6322 & n6323 ) ;
  assign n6325 = ( n6321 & n6322 ) | ( n6321 & ~n6324 ) | ( n6322 & ~n6324 ) ;
  assign n6326 = x618 & ~n6264 ;
  assign n6327 = x1117 & n6264 ;
  assign n6328 = ( ~x966 & n6326 ) | ( ~x966 & n6327 ) | ( n6326 & n6327 ) ;
  assign n6329 = x1122 & n6264 ;
  assign n6330 = x619 & ~n6264 ;
  assign n6331 = ( ~x966 & n6329 ) | ( ~x966 & n6330 ) | ( n6329 & n6330 ) ;
  assign n6332 = x1112 & n6264 ;
  assign n6333 = x620 & ~n6264 ;
  assign n6334 = ( ~x966 & n6332 ) | ( ~x966 & n6333 ) | ( n6332 & n6333 ) ;
  assign n6335 = x1108 & n6264 ;
  assign n6336 = x621 & ~n6264 ;
  assign n6337 = ( ~x966 & n6335 ) | ( ~x966 & n6336 ) | ( n6335 & n6336 ) ;
  assign n6338 = x622 & ~n6264 ;
  assign n6339 = x1109 & n6264 ;
  assign n6340 = ( ~x966 & n6338 ) | ( ~x966 & n6339 ) | ( n6338 & n6339 ) ;
  assign n6341 = x1106 & n6264 ;
  assign n6342 = x623 & ~n6264 ;
  assign n6343 = ( ~x966 & n6341 ) | ( ~x966 & n6342 ) | ( n6341 & n6342 ) ;
  assign n6344 = ~x642 & x831 ;
  assign n6345 = ~n1979 & n6344 ;
  assign n6346 = x780 & n6345 ;
  assign n6347 = x624 & ~x947 ;
  assign n6348 = ( x624 & ~n6273 ) | ( x624 & n6347 ) | ( ~n6273 & n6347 ) ;
  assign n6349 = ~n6345 & n6348 ;
  assign n6350 = ( n6345 & ~n6346 ) | ( n6345 & n6349 ) | ( ~n6346 & n6349 ) ;
  assign n6351 = x832 & ~x973 ;
  assign n6352 = ~x1054 & x1066 ;
  assign n6353 = ( x1088 & ~n6351 ) | ( x1088 & n6352 ) | ( ~n6351 & n6352 ) ;
  assign n6354 = n6351 & n6353 ;
  assign n6355 = ~x953 & n6354 ;
  assign n6356 = x1116 & n6355 ;
  assign n6357 = x625 & ~n6355 ;
  assign n6358 = ( ~x962 & n6356 ) | ( ~x962 & n6357 ) | ( n6356 & n6357 ) ;
  assign n6359 = x1121 & n6264 ;
  assign n6360 = x626 & ~n6264 ;
  assign n6361 = ( ~x966 & n6359 ) | ( ~x966 & n6360 ) | ( n6359 & n6360 ) ;
  assign n6362 = x1117 & n6355 ;
  assign n6363 = x627 & ~n6355 ;
  assign n6364 = ( ~x962 & n6362 ) | ( ~x962 & n6363 ) | ( n6362 & n6363 ) ;
  assign n6365 = x628 & ~n6355 ;
  assign n6366 = x1119 & n6355 ;
  assign n6367 = ( ~x962 & n6365 ) | ( ~x962 & n6366 ) | ( n6365 & n6366 ) ;
  assign n6368 = x1119 & n6264 ;
  assign n6369 = x629 & ~n6264 ;
  assign n6370 = ( ~x966 & n6368 ) | ( ~x966 & n6369 ) | ( n6368 & n6369 ) ;
  assign n6371 = x1120 & n6264 ;
  assign n6372 = x630 & ~n6264 ;
  assign n6373 = ( ~x966 & n6371 ) | ( ~x966 & n6372 ) | ( n6371 & n6372 ) ;
  assign n6374 = x631 | n6355 ;
  assign n6375 = x1113 & n6355 ;
  assign n6376 = ( x962 & n6374 ) | ( x962 & ~n6375 ) | ( n6374 & ~n6375 ) ;
  assign n6377 = x1115 & n6355 ;
  assign n6378 = x632 | n6355 ;
  assign n6379 = ( x962 & ~n6377 ) | ( x962 & n6378 ) | ( ~n6377 & n6378 ) ;
  assign n6380 = x1110 & n6264 ;
  assign n6381 = x633 & ~n6264 ;
  assign n6382 = ( ~x966 & n6380 ) | ( ~x966 & n6381 ) | ( n6380 & n6381 ) ;
  assign n6383 = x1110 & n6355 ;
  assign n6384 = x634 & ~n6355 ;
  assign n6385 = ( ~x962 & n6383 ) | ( ~x962 & n6384 ) | ( n6383 & n6384 ) ;
  assign n6386 = x635 | n6355 ;
  assign n6387 = x1112 & n6355 ;
  assign n6388 = ( x962 & n6386 ) | ( x962 & ~n6387 ) | ( n6386 & ~n6387 ) ;
  assign n6389 = x636 & ~n6264 ;
  assign n6390 = x1127 & n6264 ;
  assign n6391 = ( ~x966 & n6389 ) | ( ~x966 & n6390 ) | ( n6389 & n6390 ) ;
  assign n6392 = x1105 & n6355 ;
  assign n6393 = x637 & ~n6355 ;
  assign n6394 = ( ~x962 & n6392 ) | ( ~x962 & n6393 ) | ( n6392 & n6393 ) ;
  assign n6395 = x638 & ~n6355 ;
  assign n6396 = x1107 & n6355 ;
  assign n6397 = ( ~x962 & n6395 ) | ( ~x962 & n6396 ) | ( n6395 & n6396 ) ;
  assign n6398 = x1109 & n6355 ;
  assign n6399 = x639 & ~n6355 ;
  assign n6400 = ( ~x962 & n6398 ) | ( ~x962 & n6399 ) | ( n6398 & n6399 ) ;
  assign n6401 = x1128 & n6264 ;
  assign n6402 = x640 & ~n6264 ;
  assign n6403 = ( ~x966 & n6401 ) | ( ~x966 & n6402 ) | ( n6401 & n6402 ) ;
  assign n6404 = x641 & ~n6355 ;
  assign n6405 = x1121 & n6355 ;
  assign n6406 = ( ~x962 & n6404 ) | ( ~x962 & n6405 ) | ( n6404 & n6405 ) ;
  assign n6407 = x1103 & n6264 ;
  assign n6408 = x642 & ~n6264 ;
  assign n6409 = ( ~x966 & n6407 ) | ( ~x966 & n6408 ) | ( n6407 & n6408 ) ;
  assign n6410 = x643 & ~n6355 ;
  assign n6411 = x1104 & n6355 ;
  assign n6412 = ( ~x962 & n6410 ) | ( ~x962 & n6411 ) | ( n6410 & n6411 ) ;
  assign n6413 = x644 & ~n6264 ;
  assign n6414 = x1123 & n6264 ;
  assign n6415 = ( ~x966 & n6413 ) | ( ~x966 & n6414 ) | ( n6413 & n6414 ) ;
  assign n6416 = x1125 & n6264 ;
  assign n6417 = x645 & ~n6264 ;
  assign n6418 = ( ~x966 & n6416 ) | ( ~x966 & n6417 ) | ( n6416 & n6417 ) ;
  assign n6419 = x1114 & n6355 ;
  assign n6420 = x646 | n6355 ;
  assign n6421 = ( x962 & ~n6419 ) | ( x962 & n6420 ) | ( ~n6419 & n6420 ) ;
  assign n6422 = x1120 & n6355 ;
  assign n6423 = x647 & ~n6355 ;
  assign n6424 = ( ~x962 & n6422 ) | ( ~x962 & n6423 ) | ( n6422 & n6423 ) ;
  assign n6425 = x648 & ~n6355 ;
  assign n6426 = x1122 & n6355 ;
  assign n6427 = ( ~x962 & n6425 ) | ( ~x962 & n6426 ) | ( n6425 & n6426 ) ;
  assign n6428 = x1126 & n6355 ;
  assign n6429 = x649 | n6355 ;
  assign n6430 = ( x962 & ~n6428 ) | ( x962 & n6429 ) | ( ~n6428 & n6429 ) ;
  assign n6431 = x650 | n6355 ;
  assign n6432 = x1127 & n6355 ;
  assign n6433 = ( x962 & n6431 ) | ( x962 & ~n6432 ) | ( n6431 & ~n6432 ) ;
  assign n6434 = x1130 & n6264 ;
  assign n6435 = x651 & ~n6264 ;
  assign n6436 = ( ~x966 & n6434 ) | ( ~x966 & n6435 ) | ( n6434 & n6435 ) ;
  assign n6437 = x1131 & n6264 ;
  assign n6438 = x652 & ~n6264 ;
  assign n6439 = ( ~x966 & n6437 ) | ( ~x966 & n6438 ) | ( n6437 & n6438 ) ;
  assign n6440 = x1129 & n6264 ;
  assign n6441 = x653 & ~n6264 ;
  assign n6442 = ( ~x966 & n6440 ) | ( ~x966 & n6441 ) | ( n6440 & n6441 ) ;
  assign n6443 = x1130 & n6355 ;
  assign n6444 = x654 | n6355 ;
  assign n6445 = ( x962 & ~n6443 ) | ( x962 & n6444 ) | ( ~n6443 & n6444 ) ;
  assign n6446 = x655 | n6355 ;
  assign n6447 = x1124 & n6355 ;
  assign n6448 = ( x962 & n6446 ) | ( x962 & ~n6447 ) | ( n6446 & ~n6447 ) ;
  assign n6449 = x656 & ~n6264 ;
  assign n6450 = x1126 & n6264 ;
  assign n6451 = ( ~x966 & n6449 ) | ( ~x966 & n6450 ) | ( n6449 & n6450 ) ;
  assign n6452 = x657 | n6355 ;
  assign n6453 = x1131 & n6355 ;
  assign n6454 = ( x962 & n6452 ) | ( x962 & ~n6453 ) | ( n6452 & ~n6453 ) ;
  assign n6455 = x1124 & n6264 ;
  assign n6456 = x658 & ~n6264 ;
  assign n6457 = ( ~x966 & n6455 ) | ( ~x966 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6458 = x269 | x281 ;
  assign n6459 = ( x266 & x280 ) | ( x266 & x992 ) | ( x280 & x992 ) ;
  assign n6460 = ~x280 & n6459 ;
  assign n6461 = ~n6458 & n6460 ;
  assign n6462 = ~x282 & n6461 ;
  assign n6463 = x270 | x277 ;
  assign n6464 = n6462 & ~n6463 ;
  assign n6465 = ( ~x264 & x265 ) | ( ~x264 & n6464 ) | ( x265 & n6464 ) ;
  assign n6466 = ~x265 & n6465 ;
  assign n6467 = x274 & ~n6466 ;
  assign n6468 = ~x274 & n6466 ;
  assign n6469 = n6467 | n6468 ;
  assign n6470 = x1118 & n6355 ;
  assign n6471 = x660 & ~n6355 ;
  assign n6472 = ( ~x962 & n6470 ) | ( ~x962 & n6471 ) | ( n6470 & n6471 ) ;
  assign n6473 = x1101 & n6355 ;
  assign n6474 = x661 & ~n6355 ;
  assign n6475 = ( ~x962 & n6473 ) | ( ~x962 & n6474 ) | ( n6473 & n6474 ) ;
  assign n6476 = x662 & ~n6355 ;
  assign n6477 = x1102 & n6355 ;
  assign n6478 = ( ~x962 & n6476 ) | ( ~x962 & n6477 ) | ( n6476 & n6477 ) ;
  assign n6479 = x1137 | x1138 ;
  assign n6480 = n2180 & ~n6479 ;
  assign n6481 = x634 & ~x1134 ;
  assign n6482 = x700 & x1134 ;
  assign n6483 = ( x1135 & n6481 ) | ( x1135 & n6482 ) | ( n6481 & n6482 ) ;
  assign n6484 = x766 & x1134 ;
  assign n6485 = x633 & ~x1134 ;
  assign n6486 = ( ~x1135 & n6484 ) | ( ~x1135 & n6485 ) | ( n6484 & n6485 ) ;
  assign n6487 = ( x1136 & n6483 ) | ( x1136 & n6486 ) | ( n6483 & n6486 ) ;
  assign n6488 = x784 & x1135 ;
  assign n6489 = x815 & ~x1135 ;
  assign n6490 = ( ~x1134 & n6488 ) | ( ~x1134 & n6489 ) | ( n6488 & n6489 ) ;
  assign n6491 = x1134 & ~x1135 ;
  assign n6492 = x855 & n6491 ;
  assign n6493 = ( ~x1136 & n6490 ) | ( ~x1136 & n6492 ) | ( n6490 & n6492 ) ;
  assign n6494 = n6487 | n6493 ;
  assign n6495 = n6480 & n6494 ;
  assign n6496 = x199 & x1065 ;
  assign n6497 = x223 | x224 ;
  assign n6498 = ~n2180 & n6497 ;
  assign n6499 = ~x199 & x257 ;
  assign n6500 = ( n6496 & n6498 ) | ( n6496 & n6499 ) | ( n6498 & n6499 ) ;
  assign n6501 = n6495 | n6500 ;
  assign n6502 = n2180 | n6497 ;
  assign n6503 = x464 & n2185 ;
  assign n6504 = x334 & n2314 ;
  assign n6505 = n6503 | n6504 ;
  assign n6506 = ~x588 & n2381 ;
  assign n6507 = x323 & n6506 ;
  assign n6508 = n6505 | n6507 ;
  assign n6509 = ~n2312 & n2378 ;
  assign n6510 = x365 & n6509 ;
  assign n6511 = ( ~n6502 & n6508 ) | ( ~n6502 & n6510 ) | ( n6508 & n6510 ) ;
  assign n6512 = n6501 | n6511 ;
  assign n6513 = x1136 & n6480 ;
  assign n6514 = x614 & ~x1135 ;
  assign n6515 = x662 & x1135 ;
  assign n6516 = ( ~x1134 & n6514 ) | ( ~x1134 & n6515 ) | ( n6514 & n6515 ) ;
  assign n6517 = x772 & ~x1135 ;
  assign n6518 = x727 & x1135 ;
  assign n6519 = ( x1134 & n6517 ) | ( x1134 & n6518 ) | ( n6517 & n6518 ) ;
  assign n6520 = ( n6513 & n6516 ) | ( n6513 & n6519 ) | ( n6516 & n6519 ) ;
  assign n6521 = x429 & n2185 ;
  assign n6522 = x355 & n6506 ;
  assign n6523 = ( ~n6502 & n6521 ) | ( ~n6502 & n6522 ) | ( n6521 & n6522 ) ;
  assign n6524 = n6520 | n6523 ;
  assign n6525 = x872 & n6491 ;
  assign n6526 = ~x1136 & n6480 ;
  assign n6527 = x811 & ~x1135 ;
  assign n6528 = x785 & x1135 ;
  assign n6529 = ( ~x1134 & n6527 ) | ( ~x1134 & n6528 ) | ( n6527 & n6528 ) ;
  assign n6530 = ( n6525 & n6526 ) | ( n6525 & n6529 ) | ( n6526 & n6529 ) ;
  assign n6531 = x199 & x1084 ;
  assign n6532 = ~x199 & x292 ;
  assign n6533 = ( n6498 & n6531 ) | ( n6498 & n6532 ) | ( n6531 & n6532 ) ;
  assign n6534 = n6502 & ~n6533 ;
  assign n6535 = x404 & n2314 ;
  assign n6536 = x380 & n6509 ;
  assign n6537 = n6535 | n6536 ;
  assign n6538 = ( n6533 & ~n6534 ) | ( n6533 & n6537 ) | ( ~n6534 & n6537 ) ;
  assign n6539 = ( ~n6524 & n6530 ) | ( ~n6524 & n6538 ) | ( n6530 & n6538 ) ;
  assign n6540 = n6524 | n6539 ;
  assign n6541 = x665 & ~n6355 ;
  assign n6542 = x1108 & n6355 ;
  assign n6543 = ( ~x962 & n6541 ) | ( ~x962 & n6542 ) | ( n6541 & n6542 ) ;
  assign n6544 = x790 & ~x1136 ;
  assign n6545 = x638 & x1136 ;
  assign n6546 = ( x1135 & n6544 ) | ( x1135 & n6545 ) | ( n6544 & n6545 ) ;
  assign n6547 = x799 | x1136 ;
  assign n6548 = x607 & x1136 ;
  assign n6549 = ( x1135 & n6547 ) | ( x1135 & ~n6548 ) | ( n6547 & ~n6548 ) ;
  assign n6550 = ( x1134 & ~n6546 ) | ( x1134 & n6549 ) | ( ~n6546 & n6549 ) ;
  assign n6551 = x1135 & x1136 ;
  assign n6552 = x691 & n6551 ;
  assign n6553 = x764 & x1136 ;
  assign n6554 = x873 & ~x1136 ;
  assign n6555 = ( ~x1135 & n6553 ) | ( ~x1135 & n6554 ) | ( n6553 & n6554 ) ;
  assign n6556 = ( x1134 & n6552 ) | ( x1134 & n6555 ) | ( n6552 & n6555 ) ;
  assign n6557 = n6550 & ~n6556 ;
  assign n6558 = n6480 & ~n6557 ;
  assign n6559 = ~x199 & x297 ;
  assign n6560 = x199 & x1044 ;
  assign n6561 = ( n6498 & n6559 ) | ( n6498 & n6560 ) | ( n6559 & n6560 ) ;
  assign n6562 = n6558 | n6561 ;
  assign n6563 = x456 & n2314 ;
  assign n6564 = x443 & n2185 ;
  assign n6565 = x337 & n6509 ;
  assign n6566 = ( ~n2314 & n6564 ) | ( ~n2314 & n6565 ) | ( n6564 & n6565 ) ;
  assign n6567 = ( ~n6502 & n6563 ) | ( ~n6502 & n6566 ) | ( n6563 & n6566 ) ;
  assign n6568 = ~n6502 & n6506 ;
  assign n6569 = x441 & ~n6568 ;
  assign n6570 = ( x441 & n6567 ) | ( x441 & ~n6569 ) | ( n6567 & ~n6569 ) ;
  assign n6571 = n6562 | n6570 ;
  assign n6572 = ~x199 & x294 ;
  assign n6573 = x199 & x1072 ;
  assign n6574 = ( n6498 & n6572 ) | ( n6498 & n6573 ) | ( n6572 & n6573 ) ;
  assign n6575 = x1134 | x1136 ;
  assign n6576 = x809 & ~n6575 ;
  assign n6577 = x1134 & x1136 ;
  assign n6578 = ~x763 & n6577 ;
  assign n6579 = ( ~x1135 & n6576 ) | ( ~x1135 & n6578 ) | ( n6576 & n6578 ) ;
  assign n6580 = n6480 & n6579 ;
  assign n6581 = x1134 & x1135 ;
  assign n6582 = x681 & x1136 ;
  assign n6583 = ( x1135 & n6581 ) | ( x1135 & ~n6582 ) | ( n6581 & ~n6582 ) ;
  assign n6584 = ~x642 & x1136 ;
  assign n6585 = ( ~x1135 & n6491 ) | ( ~x1135 & n6584 ) | ( n6491 & n6584 ) ;
  assign n6586 = ( x871 & x1134 ) | ( x871 & n6577 ) | ( x1134 & n6577 ) ;
  assign n6587 = n6585 & ~n6586 ;
  assign n6588 = x792 & ~n6575 ;
  assign n6589 = x699 & n6577 ;
  assign n6590 = n6588 | n6589 ;
  assign n6591 = ( n6583 & n6587 ) | ( n6583 & ~n6590 ) | ( n6587 & ~n6590 ) ;
  assign n6592 = ( n6480 & n6580 ) | ( n6480 & n6591 ) | ( n6580 & n6591 ) ;
  assign n6593 = ( n6480 & n6574 ) | ( n6480 & ~n6592 ) | ( n6574 & ~n6592 ) ;
  assign n6594 = ~n6502 & n6509 ;
  assign n6595 = x338 & n6594 ;
  assign n6596 = x458 & n2381 ;
  assign n6597 = x319 & n2314 ;
  assign n6598 = ( ~x588 & n6596 ) | ( ~x588 & n6597 ) | ( n6596 & n6597 ) ;
  assign n6599 = x444 & n2185 ;
  assign n6600 = ( ~n6502 & n6598 ) | ( ~n6502 & n6599 ) | ( n6598 & n6599 ) ;
  assign n6601 = ( ~n6502 & n6595 ) | ( ~n6502 & n6600 ) | ( n6595 & n6600 ) ;
  assign n6602 = n6593 | n6601 ;
  assign n6603 = x414 & n2185 ;
  assign n6604 = x342 & n6506 ;
  assign n6605 = n6603 | n6604 ;
  assign n6606 = x363 & n6509 ;
  assign n6607 = x390 & n2314 ;
  assign n6608 = n6606 | n6607 ;
  assign n6609 = ( ~n6502 & n6605 ) | ( ~n6502 & n6608 ) | ( n6605 & n6608 ) ;
  assign n6610 = x837 & n6491 ;
  assign n6611 = x981 & ~x1135 ;
  assign n6612 = x778 & x1135 ;
  assign n6613 = ( ~x1134 & n6611 ) | ( ~x1134 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6614 = ( n6526 & n6610 ) | ( n6526 & n6613 ) | ( n6610 & n6613 ) ;
  assign n6615 = x759 & ~x1135 ;
  assign n6616 = x696 & x1135 ;
  assign n6617 = ( x1134 & n6615 ) | ( x1134 & n6616 ) | ( n6615 & n6616 ) ;
  assign n6618 = x603 & ~x1135 ;
  assign n6619 = x680 & x1135 ;
  assign n6620 = ( ~x1134 & n6618 ) | ( ~x1134 & n6619 ) | ( n6618 & n6619 ) ;
  assign n6621 = ( n6513 & n6617 ) | ( n6513 & n6620 ) | ( n6617 & n6620 ) ;
  assign n6622 = ~x199 & x291 ;
  assign n6623 = x199 & x1049 ;
  assign n6624 = ( n6498 & n6622 ) | ( n6498 & n6623 ) | ( n6622 & n6623 ) ;
  assign n6625 = n6621 | n6624 ;
  assign n6626 = ( ~n6609 & n6614 ) | ( ~n6609 & n6625 ) | ( n6614 & n6625 ) ;
  assign n6627 = n6609 | n6626 ;
  assign n6628 = x1125 & n6355 ;
  assign n6629 = x669 | n6355 ;
  assign n6630 = ( x962 & ~n6628 ) | ( x962 & n6629 ) | ( ~n6628 & n6629 ) ;
  assign n6631 = n6491 & n6526 ;
  assign n6632 = x852 & n6631 ;
  assign n6633 = ~x723 & n6581 ;
  assign n6634 = ~x745 & n6491 ;
  assign n6635 = x612 & ~x1135 ;
  assign n6636 = ~x695 & x1135 ;
  assign n6637 = ( ~x1134 & n6635 ) | ( ~x1134 & n6636 ) | ( n6635 & n6636 ) ;
  assign n6638 = n6634 | n6637 ;
  assign n6639 = ( n6513 & n6633 ) | ( n6513 & n6638 ) | ( n6633 & n6638 ) ;
  assign n6640 = x415 & n2185 ;
  assign n6641 = x343 & n6506 ;
  assign n6642 = ( ~n6502 & n6640 ) | ( ~n6502 & n6641 ) | ( n6640 & n6641 ) ;
  assign n6643 = x391 & n2314 ;
  assign n6644 = x364 & n6509 ;
  assign n6645 = ( ~n6502 & n6643 ) | ( ~n6502 & n6644 ) | ( n6643 & n6644 ) ;
  assign n6646 = x199 & x1062 ;
  assign n6647 = ~x199 & x258 ;
  assign n6648 = ( n6498 & n6646 ) | ( n6498 & n6647 ) | ( n6646 & n6647 ) ;
  assign n6649 = n6645 | n6648 ;
  assign n6650 = ( ~n6632 & n6642 ) | ( ~n6632 & n6649 ) | ( n6642 & n6649 ) ;
  assign n6651 = ( ~n6632 & n6639 ) | ( ~n6632 & n6650 ) | ( n6639 & n6650 ) ;
  assign n6652 = n6632 | n6651 ;
  assign n6653 = x865 & x1134 ;
  assign n6654 = ~x1136 & n6653 ;
  assign n6655 = ~x741 & x1134 ;
  assign n6656 = x611 & ~x1134 ;
  assign n6657 = ( x1136 & n6655 ) | ( x1136 & n6656 ) | ( n6655 & n6656 ) ;
  assign n6658 = ( ~x1135 & n6654 ) | ( ~x1135 & n6657 ) | ( n6654 & n6657 ) ;
  assign n6659 = ~x724 & x1134 ;
  assign n6660 = x646 | x1134 ;
  assign n6661 = ( n6551 & n6659 ) | ( n6551 & ~n6660 ) | ( n6659 & ~n6660 ) ;
  assign n6662 = ( n6480 & n6658 ) | ( n6480 & n6661 ) | ( n6658 & n6661 ) ;
  assign n6663 = x199 & x1040 ;
  assign n6664 = ~x199 & x261 ;
  assign n6665 = ( n6498 & n6663 ) | ( n6498 & n6664 ) | ( n6663 & n6664 ) ;
  assign n6666 = n6662 | n6665 ;
  assign n6667 = x453 & n2185 ;
  assign n6668 = x447 & n6509 ;
  assign n6669 = x333 & n2314 ;
  assign n6670 = ( ~n6667 & n6668 ) | ( ~n6667 & n6669 ) | ( n6668 & n6669 ) ;
  assign n6671 = n6667 | n6670 ;
  assign n6672 = x327 & n6568 ;
  assign n6673 = ( ~n6502 & n6671 ) | ( ~n6502 & n6672 ) | ( n6671 & n6672 ) ;
  assign n6674 = n6666 | n6673 ;
  assign n6675 = x736 & n6551 ;
  assign n6676 = x758 & x1136 ;
  assign n6677 = x850 & ~x1136 ;
  assign n6678 = ( ~x1135 & n6676 ) | ( ~x1135 & n6677 ) | ( n6676 & n6677 ) ;
  assign n6679 = ( x1134 & n6675 ) | ( x1134 & n6678 ) | ( n6675 & n6678 ) ;
  assign n6680 = ~x1135 & x1136 ;
  assign n6681 = x616 & n6680 ;
  assign n6682 = x781 & x1135 ;
  assign n6683 = x808 & ~x1135 ;
  assign n6684 = ( ~x1136 & n6682 ) | ( ~x1136 & n6683 ) | ( n6682 & n6683 ) ;
  assign n6685 = n6681 | n6684 ;
  assign n6686 = x661 & n6551 ;
  assign n6687 = ( ~x1134 & n6685 ) | ( ~x1134 & n6686 ) | ( n6685 & n6686 ) ;
  assign n6688 = ( n6480 & n6679 ) | ( n6480 & n6687 ) | ( n6679 & n6687 ) ;
  assign n6689 = x199 & x1048 ;
  assign n6690 = ~x199 & x290 ;
  assign n6691 = ( n6498 & n6689 ) | ( n6498 & n6690 ) | ( n6689 & n6690 ) ;
  assign n6692 = n6688 | n6691 ;
  assign n6693 = x397 & n2314 ;
  assign n6694 = x372 & n6509 ;
  assign n6695 = x422 & n2185 ;
  assign n6696 = ( ~n6693 & n6694 ) | ( ~n6693 & n6695 ) | ( n6694 & n6695 ) ;
  assign n6697 = n6693 | n6696 ;
  assign n6698 = x320 & n6568 ;
  assign n6699 = ( ~n6502 & n6697 ) | ( ~n6502 & n6698 ) | ( n6697 & n6698 ) ;
  assign n6700 = n6692 | n6699 ;
  assign n6701 = x1135 | x1136 ;
  assign n6702 = x814 | n6701 ;
  assign n6703 = x1134 & ~n6680 ;
  assign n6704 = ( ~x749 & x1134 ) | ( ~x749 & n6703 ) | ( x1134 & n6703 ) ;
  assign n6705 = x706 & n6551 ;
  assign n6706 = x866 & ~n6701 ;
  assign n6707 = ( n6704 & n6705 ) | ( n6704 & n6706 ) | ( n6705 & n6706 ) ;
  assign n6708 = n6704 & ~n6707 ;
  assign n6709 = ( x788 & x1136 ) | ( x788 & n6701 ) | ( x1136 & n6701 ) ;
  assign n6710 = x617 & n6680 ;
  assign n6711 = ( ~x1136 & n6709 ) | ( ~x1136 & n6710 ) | ( n6709 & n6710 ) ;
  assign n6712 = x637 | x1134 ;
  assign n6713 = ( x1134 & n6551 ) | ( x1134 & n6712 ) | ( n6551 & n6712 ) ;
  assign n6714 = ( n6702 & n6711 ) | ( n6702 & n6713 ) | ( n6711 & n6713 ) ;
  assign n6715 = ( n6702 & n6708 ) | ( n6702 & ~n6714 ) | ( n6708 & ~n6714 ) ;
  assign n6716 = n6480 & ~n6715 ;
  assign n6717 = x387 & n6594 ;
  assign n6718 = x435 & n2185 ;
  assign n6719 = x411 & n2314 ;
  assign n6720 = n6718 | n6719 ;
  assign n6721 = x452 & n6568 ;
  assign n6722 = ( ~n6502 & n6720 ) | ( ~n6502 & n6721 ) | ( n6720 & n6721 ) ;
  assign n6723 = ~x199 & x295 ;
  assign n6724 = x199 & x1053 ;
  assign n6725 = ( n6498 & n6723 ) | ( n6498 & n6724 ) | ( n6723 & n6724 ) ;
  assign n6726 = ( ~n6716 & n6722 ) | ( ~n6716 & n6725 ) | ( n6722 & n6725 ) ;
  assign n6727 = ( ~n6716 & n6717 ) | ( ~n6716 & n6726 ) | ( n6717 & n6726 ) ;
  assign n6728 = n6716 | n6727 ;
  assign n6729 = x639 & x1136 ;
  assign n6730 = x783 & ~x1136 ;
  assign n6731 = ( x1135 & n6729 ) | ( x1135 & n6730 ) | ( n6729 & n6730 ) ;
  assign n6732 = x622 & x1136 ;
  assign n6733 = x804 & ~x1136 ;
  assign n6734 = ( ~x1135 & n6732 ) | ( ~x1135 & n6733 ) | ( n6732 & n6733 ) ;
  assign n6735 = ( ~x1134 & n6731 ) | ( ~x1134 & n6734 ) | ( n6731 & n6734 ) ;
  assign n6736 = ~x743 & n6680 ;
  assign n6737 = ( x859 & x1134 ) | ( x859 & n6577 ) | ( x1134 & n6577 ) ;
  assign n6738 = x735 & x1136 ;
  assign n6739 = x1135 & ~n6738 ;
  assign n6740 = ( n6736 & n6737 ) | ( n6736 & ~n6739 ) | ( n6737 & ~n6739 ) ;
  assign n6741 = ~n6736 & n6740 ;
  assign n6742 = ( n6480 & n6735 ) | ( n6480 & n6741 ) | ( n6735 & n6741 ) ;
  assign n6743 = x199 & x1070 ;
  assign n6744 = ~x199 & x256 ;
  assign n6745 = ( n6498 & n6743 ) | ( n6498 & n6744 ) | ( n6743 & n6744 ) ;
  assign n6746 = n6742 | n6745 ;
  assign n6747 = x336 & n6594 ;
  assign n6748 = x463 & n2314 ;
  assign n6749 = x437 & n2185 ;
  assign n6750 = n6748 | n6749 ;
  assign n6751 = x362 & n6506 ;
  assign n6752 = n6750 | n6751 ;
  assign n6753 = ( ~n6502 & n6747 ) | ( ~n6502 & n6752 ) | ( n6747 & n6752 ) ;
  assign n6754 = n6746 | n6753 ;
  assign n6755 = x436 & n2185 ;
  assign n6756 = x388 & n6509 ;
  assign n6757 = ( x455 & x588 ) | ( x455 & n2381 ) | ( x588 & n2381 ) ;
  assign n6758 = x412 & n2314 ;
  assign n6759 = ( ~x588 & n6757 ) | ( ~x588 & n6758 ) | ( n6757 & n6758 ) ;
  assign n6760 = ( ~n6755 & n6756 ) | ( ~n6755 & n6759 ) | ( n6756 & n6759 ) ;
  assign n6761 = ( ~n6502 & n6755 ) | ( ~n6502 & n6760 ) | ( n6755 & n6760 ) ;
  assign n6762 = x199 & x1037 ;
  assign n6763 = ~x199 & x296 ;
  assign n6764 = ( n6498 & n6762 ) | ( n6498 & n6763 ) | ( n6762 & n6763 ) ;
  assign n6765 = x623 & n6680 ;
  assign n6766 = x803 | x1135 ;
  assign n6767 = x789 & x1135 ;
  assign n6768 = ( x1136 & n6766 ) | ( x1136 & ~n6767 ) | ( n6766 & ~n6767 ) ;
  assign n6769 = ~n6765 & n6768 ;
  assign n6770 = x710 | x1134 ;
  assign n6771 = ( x1134 & n6551 ) | ( x1134 & n6770 ) | ( n6551 & n6770 ) ;
  assign n6772 = n6769 & ~n6771 ;
  assign n6773 = ( ~x748 & x1134 ) | ( ~x748 & n6703 ) | ( x1134 & n6703 ) ;
  assign n6774 = x876 & ~n6701 ;
  assign n6775 = x730 & n6551 ;
  assign n6776 = ( n6773 & n6774 ) | ( n6773 & n6775 ) | ( n6774 & n6775 ) ;
  assign n6777 = ( n6772 & n6773 ) | ( n6772 & ~n6776 ) | ( n6773 & ~n6776 ) ;
  assign n6778 = n6480 & ~n6777 ;
  assign n6779 = ( ~n6761 & n6764 ) | ( ~n6761 & n6778 ) | ( n6764 & n6778 ) ;
  assign n6780 = n6761 | n6779 ;
  assign n6781 = x881 & n6491 ;
  assign n6782 = x787 & x1135 ;
  assign n6783 = x812 | x1135 ;
  assign n6784 = ( x1134 & ~n6782 ) | ( x1134 & n6783 ) | ( ~n6782 & n6783 ) ;
  assign n6785 = ( n6526 & n6781 ) | ( n6526 & ~n6784 ) | ( n6781 & ~n6784 ) ;
  assign n6786 = x643 & x1135 ;
  assign n6787 = x606 & ~x1135 ;
  assign n6788 = ( ~x1134 & n6786 ) | ( ~x1134 & n6787 ) | ( n6786 & n6787 ) ;
  assign n6789 = x746 & ~x1135 ;
  assign n6790 = x729 & x1135 ;
  assign n6791 = ( x1134 & n6789 ) | ( x1134 & n6790 ) | ( n6789 & n6790 ) ;
  assign n6792 = ( n6513 & n6788 ) | ( n6513 & n6791 ) | ( n6788 & n6791 ) ;
  assign n6793 = n6785 | n6792 ;
  assign n6794 = x434 & n2185 ;
  assign n6795 = x361 & n6506 ;
  assign n6796 = x410 & n2314 ;
  assign n6797 = x386 & n6509 ;
  assign n6798 = n6796 | n6797 ;
  assign n6799 = n6795 | n6798 ;
  assign n6800 = ( ~n6502 & n6794 ) | ( ~n6502 & n6799 ) | ( n6794 & n6799 ) ;
  assign n6801 = n6793 | n6800 ;
  assign n6802 = x199 & x1059 ;
  assign n6803 = ~x199 & x293 ;
  assign n6804 = ( n6498 & n6802 ) | ( n6498 & n6803 ) | ( n6802 & n6803 ) ;
  assign n6805 = n6801 | n6804 ;
  assign n6806 = x870 & ~x1136 ;
  assign n6807 = n6491 & n6806 ;
  assign n6808 = x635 | x1134 ;
  assign n6809 = ~x704 & x1134 ;
  assign n6810 = ( x1135 & ~n6808 ) | ( x1135 & n6809 ) | ( ~n6808 & n6809 ) ;
  assign n6811 = x620 & ~x1134 ;
  assign n6812 = ~x742 & x1134 ;
  assign n6813 = ( ~x1135 & n6811 ) | ( ~x1135 & n6812 ) | ( n6811 & n6812 ) ;
  assign n6814 = ( x1136 & n6810 ) | ( x1136 & n6813 ) | ( n6810 & n6813 ) ;
  assign n6815 = ( n6480 & n6807 ) | ( n6480 & n6814 ) | ( n6807 & n6814 ) ;
  assign n6816 = x199 & x1069 ;
  assign n6817 = ~x199 & x259 ;
  assign n6818 = ( n6498 & n6816 ) | ( n6498 & n6817 ) | ( n6816 & n6817 ) ;
  assign n6819 = n6815 | n6818 ;
  assign n6820 = x366 & n6509 ;
  assign n6821 = x335 & n2314 ;
  assign n6822 = n6820 | n6821 ;
  assign n6823 = x416 & n2185 ;
  assign n6824 = x344 & n6506 ;
  assign n6825 = n6823 | n6824 ;
  assign n6826 = ( ~n6502 & n6822 ) | ( ~n6502 & n6825 ) | ( n6822 & n6825 ) ;
  assign n6827 = n6819 | n6826 ;
  assign n6828 = x856 & n6631 ;
  assign n6829 = x346 & n6568 ;
  assign n6830 = n6828 | n6829 ;
  assign n6831 = ~x688 & n6581 ;
  assign n6832 = ~x1134 & x1135 ;
  assign n6833 = ~x632 & n6832 ;
  assign n6834 = ~x760 & x1134 ;
  assign n6835 = x613 & ~x1134 ;
  assign n6836 = ( ~x1135 & n6834 ) | ( ~x1135 & n6835 ) | ( n6834 & n6835 ) ;
  assign n6837 = ( ~n6831 & n6833 ) | ( ~n6831 & n6836 ) | ( n6833 & n6836 ) ;
  assign n6838 = ( n6513 & n6831 ) | ( n6513 & n6837 ) | ( n6831 & n6837 ) ;
  assign n6839 = ~x199 & x260 ;
  assign n6840 = x199 & x1067 ;
  assign n6841 = ( n6498 & n6839 ) | ( n6498 & n6840 ) | ( n6839 & n6840 ) ;
  assign n6842 = x418 & n2185 ;
  assign n6843 = x368 & n6509 ;
  assign n6844 = x393 & n2314 ;
  assign n6845 = n6843 | n6844 ;
  assign n6846 = ( ~n6502 & n6842 ) | ( ~n6502 & n6845 ) | ( n6842 & n6845 ) ;
  assign n6847 = ( ~n6830 & n6841 ) | ( ~n6830 & n6846 ) | ( n6841 & n6846 ) ;
  assign n6848 = ( ~n6830 & n6838 ) | ( ~n6830 & n6847 ) | ( n6838 & n6847 ) ;
  assign n6849 = n6830 | n6848 ;
  assign n6850 = x665 & ~x1134 ;
  assign n6851 = x690 & x1134 ;
  assign n6852 = ( x1135 & n6850 ) | ( x1135 & n6851 ) | ( n6850 & n6851 ) ;
  assign n6853 = x621 & ~x1134 ;
  assign n6854 = x739 & x1134 ;
  assign n6855 = ( ~x1135 & n6853 ) | ( ~x1135 & n6854 ) | ( n6853 & n6854 ) ;
  assign n6856 = ( x1136 & n6852 ) | ( x1136 & n6855 ) | ( n6852 & n6855 ) ;
  assign n6857 = x810 & ~x1135 ;
  assign n6858 = x791 & x1135 ;
  assign n6859 = ( ~n6575 & n6857 ) | ( ~n6575 & n6858 ) | ( n6857 & n6858 ) ;
  assign n6860 = n6856 | n6859 ;
  assign n6861 = x874 & ~x1136 ;
  assign n6862 = n6491 & n6861 ;
  assign n6863 = ( n6480 & n6860 ) | ( n6480 & n6862 ) | ( n6860 & n6862 ) ;
  assign n6864 = ~x199 & x255 ;
  assign n6865 = x199 & x1036 ;
  assign n6866 = ( n6498 & n6864 ) | ( n6498 & n6865 ) | ( n6864 & n6865 ) ;
  assign n6867 = n6863 | n6866 ;
  assign n6868 = x450 & n6568 ;
  assign n6869 = x413 & n2314 ;
  assign n6870 = x438 & n2185 ;
  assign n6871 = x389 & n6509 ;
  assign n6872 = ( ~n6869 & n6870 ) | ( ~n6869 & n6871 ) | ( n6870 & n6871 ) ;
  assign n6873 = n6869 | n6872 ;
  assign n6874 = ( ~n6502 & n6868 ) | ( ~n6502 & n6873 ) | ( n6868 & n6873 ) ;
  assign n6875 = n6867 | n6874 ;
  assign n6876 = x680 & ~n6355 ;
  assign n6877 = x1100 & n6355 ;
  assign n6878 = ( ~x962 & n6876 ) | ( ~x962 & n6877 ) | ( n6876 & n6877 ) ;
  assign n6879 = x1103 & n6355 ;
  assign n6880 = x681 & ~n6355 ;
  assign n6881 = ( ~x962 & n6879 ) | ( ~x962 & n6880 ) | ( n6879 & n6880 ) ;
  assign n6882 = x848 & ~x1136 ;
  assign n6883 = n6491 & n6882 ;
  assign n6884 = ~x757 & x1134 ;
  assign n6885 = x610 & ~x1134 ;
  assign n6886 = ( ~x1135 & n6884 ) | ( ~x1135 & n6885 ) | ( n6884 & n6885 ) ;
  assign n6887 = ~x686 & x1134 ;
  assign n6888 = x631 | x1134 ;
  assign n6889 = ( x1135 & n6887 ) | ( x1135 & ~n6888 ) | ( n6887 & ~n6888 ) ;
  assign n6890 = ( x1136 & n6886 ) | ( x1136 & n6889 ) | ( n6886 & n6889 ) ;
  assign n6891 = ( n6480 & n6883 ) | ( n6480 & n6890 ) | ( n6883 & n6890 ) ;
  assign n6892 = x199 & x1039 ;
  assign n6893 = ~x199 & x251 ;
  assign n6894 = ( n6498 & n6892 ) | ( n6498 & n6893 ) | ( n6892 & n6893 ) ;
  assign n6895 = n6891 | n6894 ;
  assign n6896 = x417 & n2185 ;
  assign n6897 = x345 & n6506 ;
  assign n6898 = x392 & n2314 ;
  assign n6899 = x367 & n6509 ;
  assign n6900 = n6898 | n6899 ;
  assign n6901 = n6897 | n6900 ;
  assign n6902 = ( ~n6502 & n6896 ) | ( ~n6502 & n6901 ) | ( n6896 & n6901 ) ;
  assign n6903 = n6895 | n6902 ;
  assign n6904 = x953 & n6354 ;
  assign n6905 = x684 | n6904 ;
  assign n6906 = x1130 & n6904 ;
  assign n6907 = ( x962 & n6905 ) | ( x962 & ~n6906 ) | ( n6905 & ~n6906 ) ;
  assign n6908 = x382 & n6509 ;
  assign n6909 = x406 & n2314 ;
  assign n6910 = n6908 | n6909 ;
  assign n6911 = x430 & n2185 ;
  assign n6912 = x357 & n6506 ;
  assign n6913 = n6911 | n6912 ;
  assign n6914 = ( ~n6502 & n6910 ) | ( ~n6502 & n6913 ) | ( n6910 & n6913 ) ;
  assign n6915 = x199 & x1076 ;
  assign n6916 = ( n4681 & n6498 ) | ( n4681 & n6915 ) | ( n6498 & n6915 ) ;
  assign n6917 = x860 & x1134 ;
  assign n6918 = x813 & ~x1134 ;
  assign n6919 = ( ~n6701 & n6917 ) | ( ~n6701 & n6918 ) | ( n6917 & n6918 ) ;
  assign n6920 = x657 | x1134 ;
  assign n6921 = ~x728 & x1134 ;
  assign n6922 = ( x1135 & ~n6920 ) | ( x1135 & n6921 ) | ( ~n6920 & n6921 ) ;
  assign n6923 = x652 & ~x1134 ;
  assign n6924 = ~x744 & x1134 ;
  assign n6925 = ( ~x1135 & n6923 ) | ( ~x1135 & n6924 ) | ( n6923 & n6924 ) ;
  assign n6926 = ( x1136 & n6922 ) | ( x1136 & n6925 ) | ( n6922 & n6925 ) ;
  assign n6927 = n6919 | n6926 ;
  assign n6928 = n6480 & n6927 ;
  assign n6929 = ( ~n6914 & n6916 ) | ( ~n6914 & n6928 ) | ( n6916 & n6928 ) ;
  assign n6930 = n6914 | n6929 ;
  assign n6931 = x686 | n6904 ;
  assign n6932 = x1113 & n6904 ;
  assign n6933 = ( x962 & n6931 ) | ( x962 & ~n6932 ) | ( n6931 & ~n6932 ) ;
  assign n6934 = x1127 & n6904 ;
  assign n6935 = x687 & ~n6904 ;
  assign n6936 = ( ~x962 & n6934 ) | ( ~x962 & n6935 ) | ( n6934 & n6935 ) ;
  assign n6937 = x1115 & n6904 ;
  assign n6938 = x688 | n6904 ;
  assign n6939 = ( x962 & ~n6937 ) | ( x962 & n6938 ) | ( ~n6937 & n6938 ) ;
  assign n6940 = x351 & n6506 ;
  assign n6941 = x426 & n2185 ;
  assign n6942 = x401 & n2314 ;
  assign n6943 = n6941 | n6942 ;
  assign n6944 = n6940 | n6943 ;
  assign n6945 = x376 & n6594 ;
  assign n6946 = ( ~n6502 & n6944 ) | ( ~n6502 & n6945 ) | ( n6944 & n6945 ) ;
  assign n6947 = ( x655 & x1135 ) | ( x655 & n6581 ) | ( x1135 & n6581 ) ;
  assign n6948 = ( ~x703 & x1135 ) | ( ~x703 & n6832 ) | ( x1135 & n6832 ) ;
  assign n6949 = ( ~x1136 & n6947 ) | ( ~x1136 & n6948 ) | ( n6947 & n6948 ) ;
  assign n6950 = n6480 & ~n6949 ;
  assign n6951 = x199 & x1079 ;
  assign n6952 = ( n4651 & n6498 ) | ( n4651 & n6951 ) | ( n6498 & n6951 ) ;
  assign n6953 = n6950 | n6952 ;
  assign n6954 = ~x1135 & n6480 ;
  assign n6955 = x658 & ~x1134 ;
  assign n6956 = ~x752 & x1134 ;
  assign n6957 = ( x1136 & n6955 ) | ( x1136 & n6956 ) | ( n6955 & n6956 ) ;
  assign n6958 = x798 & ~x1134 ;
  assign n6959 = x843 & x1134 ;
  assign n6960 = ( ~x1136 & n6958 ) | ( ~x1136 & n6959 ) | ( n6958 & n6959 ) ;
  assign n6961 = n6957 | n6960 ;
  assign n6962 = n6954 & ~n6961 ;
  assign n6963 = ( n6946 & n6953 ) | ( n6946 & ~n6962 ) | ( n6953 & ~n6962 ) ;
  assign n6964 = x690 & ~n6904 ;
  assign n6965 = x1108 & n6904 ;
  assign n6966 = ( ~x962 & n6964 ) | ( ~x962 & n6965 ) | ( n6964 & n6965 ) ;
  assign n6967 = x1107 & n6904 ;
  assign n6968 = x691 & ~n6904 ;
  assign n6969 = ( ~x962 & n6967 ) | ( ~x962 & n6968 ) | ( n6967 & n6968 ) ;
  assign n6970 = x317 & n6509 ;
  assign n6971 = x402 & n2314 ;
  assign n6972 = n6970 | n6971 ;
  assign n6973 = x427 & n2185 ;
  assign n6974 = x352 & n6506 ;
  assign n6975 = n6973 | n6974 ;
  assign n6976 = ( ~n6502 & n6972 ) | ( ~n6502 & n6975 ) | ( n6972 & n6975 ) ;
  assign n6977 = x199 & x1078 ;
  assign n6978 = ( n4663 & n6498 ) | ( n4663 & n6977 ) | ( n6498 & n6977 ) ;
  assign n6979 = n6976 | n6978 ;
  assign n6980 = x656 & ~x1135 ;
  assign n6981 = ~x649 & x1135 ;
  assign n6982 = ( ~x1134 & n6980 ) | ( ~x1134 & n6981 ) | ( n6980 & n6981 ) ;
  assign n6983 = ( x844 & n6480 ) | ( x844 & ~n6491 ) | ( n6480 & ~n6491 ) ;
  assign n6984 = ( x801 & n6491 ) | ( x801 & n6954 ) | ( n6491 & n6954 ) ;
  assign n6985 = ( n6513 & n6983 ) | ( n6513 & n6984 ) | ( n6983 & n6984 ) ;
  assign n6986 = x726 & n6581 ;
  assign n6987 = x770 & x1136 ;
  assign n6988 = ( x1136 & ~n6491 ) | ( x1136 & n6987 ) | ( ~n6491 & n6987 ) ;
  assign n6989 = ( n6982 & ~n6986 ) | ( n6982 & n6988 ) | ( ~n6986 & n6988 ) ;
  assign n6990 = ( n6982 & n6985 ) | ( n6982 & ~n6989 ) | ( n6985 & ~n6989 ) ;
  assign n6991 = n6979 | n6990 ;
  assign n6992 = x693 | n6355 ;
  assign n6993 = x1129 & n6355 ;
  assign n6994 = ( x962 & n6992 ) | ( x962 & ~n6993 ) | ( n6992 & ~n6993 ) ;
  assign n6995 = x694 | n6904 ;
  assign n6996 = x1128 & n6904 ;
  assign n6997 = ( x962 & n6995 ) | ( x962 & ~n6996 ) | ( n6995 & ~n6996 ) ;
  assign n6998 = x1111 & n6355 ;
  assign n6999 = x695 | n6355 ;
  assign n7000 = ( x962 & ~n6998 ) | ( x962 & n6999 ) | ( ~n6998 & n6999 ) ;
  assign n7001 = x1100 & n6904 ;
  assign n7002 = x696 & ~n6904 ;
  assign n7003 = ( ~x962 & n7001 ) | ( ~x962 & n7002 ) | ( n7001 & n7002 ) ;
  assign n7004 = x697 | n6904 ;
  assign n7005 = x1129 & n6904 ;
  assign n7006 = ( x962 & n7004 ) | ( x962 & ~n7005 ) | ( n7004 & ~n7005 ) ;
  assign n7007 = x698 | n6904 ;
  assign n7008 = x1116 & n6904 ;
  assign n7009 = ( x962 & n7007 ) | ( x962 & ~n7008 ) | ( n7007 & ~n7008 ) ;
  assign n7010 = x699 & ~n6904 ;
  assign n7011 = x1103 & n6904 ;
  assign n7012 = ( ~x962 & n7010 ) | ( ~x962 & n7011 ) | ( n7010 & n7011 ) ;
  assign n7013 = x700 & ~n6904 ;
  assign n7014 = x1110 & n6904 ;
  assign n7015 = ( ~x962 & n7013 ) | ( ~x962 & n7014 ) | ( n7013 & n7014 ) ;
  assign n7016 = x701 | n6904 ;
  assign n7017 = x1123 & n6904 ;
  assign n7018 = ( x962 & n7016 ) | ( x962 & ~n7017 ) | ( n7016 & ~n7017 ) ;
  assign n7019 = x1117 & n6904 ;
  assign n7020 = x702 | n6904 ;
  assign n7021 = ( x962 & ~n7019 ) | ( x962 & n7020 ) | ( ~n7019 & n7020 ) ;
  assign n7022 = x1124 & n6904 ;
  assign n7023 = x703 & ~n6904 ;
  assign n7024 = ( ~x962 & n7022 ) | ( ~x962 & n7023 ) | ( n7022 & n7023 ) ;
  assign n7025 = x704 | n6904 ;
  assign n7026 = x1112 & n6904 ;
  assign n7027 = ( x962 & n7025 ) | ( x962 & ~n7026 ) | ( n7025 & ~n7026 ) ;
  assign n7028 = x1125 & n6904 ;
  assign n7029 = x705 & ~n6904 ;
  assign n7030 = ( ~x962 & n7028 ) | ( ~x962 & n7029 ) | ( n7028 & n7029 ) ;
  assign n7031 = x1105 & n6904 ;
  assign n7032 = x706 & ~n6904 ;
  assign n7033 = ( ~x962 & n7031 ) | ( ~x962 & n7032 ) | ( n7031 & n7032 ) ;
  assign n7034 = x395 & n2314 ;
  assign n7035 = x370 & n6509 ;
  assign n7036 = ( ~n6502 & n7034 ) | ( ~n6502 & n7035 ) | ( n7034 & n7035 ) ;
  assign n7037 = x347 & n6506 ;
  assign n7038 = x420 & n2185 ;
  assign n7039 = ( ~n6502 & n7037 ) | ( ~n6502 & n7038 ) | ( n7037 & n7038 ) ;
  assign n7040 = n7036 | n7039 ;
  assign n7041 = ~x702 & n6581 ;
  assign n7042 = x627 & n6832 ;
  assign n7043 = ~x753 & x1134 ;
  assign n7044 = x618 & ~x1134 ;
  assign n7045 = ( ~x1135 & n7043 ) | ( ~x1135 & n7044 ) | ( n7043 & n7044 ) ;
  assign n7046 = ( ~n6581 & n7042 ) | ( ~n6581 & n7045 ) | ( n7042 & n7045 ) ;
  assign n7047 = ( n6513 & n7041 ) | ( n6513 & n7046 ) | ( n7041 & n7046 ) ;
  assign n7048 = x304 | n2904 ;
  assign n7049 = ~n6498 & n7048 ;
  assign n7050 = x199 & ~x1055 ;
  assign n7051 = ~x1048 & n4339 ;
  assign n7052 = ( n2904 & n7050 ) | ( n2904 & n7051 ) | ( n7050 & n7051 ) ;
  assign n7053 = ( n7048 & n7049 ) | ( n7048 & ~n7052 ) | ( n7049 & ~n7052 ) ;
  assign n7054 = ( n7047 & ~n7049 ) | ( n7047 & n7053 ) | ( ~n7049 & n7053 ) ;
  assign n7055 = x847 & n6631 ;
  assign n7056 = ( ~n7040 & n7054 ) | ( ~n7040 & n7055 ) | ( n7054 & n7055 ) ;
  assign n7057 = n7040 | n7056 ;
  assign n7058 = x754 | x1135 ;
  assign n7059 = ~x709 & x1135 ;
  assign n7060 = ( x1134 & ~n7058 ) | ( x1134 & n7059 ) | ( ~n7058 & n7059 ) ;
  assign n7061 = x660 & n6832 ;
  assign n7062 = x1134 | x1135 ;
  assign n7063 = x609 & ~n7062 ;
  assign n7064 = ( ~n7060 & n7061 ) | ( ~n7060 & n7063 ) | ( n7061 & n7063 ) ;
  assign n7065 = ( n6513 & n7060 ) | ( n6513 & n7064 ) | ( n7060 & n7064 ) ;
  assign n7066 = x305 | n2904 ;
  assign n7067 = x199 & ~x1058 ;
  assign n7068 = ~x1084 & n4339 ;
  assign n7069 = ( n6498 & n7067 ) | ( n6498 & n7068 ) | ( n7067 & n7068 ) ;
  assign n7070 = ( ~n6498 & n7066 ) | ( ~n6498 & n7069 ) | ( n7066 & n7069 ) ;
  assign n7071 = ( n7065 & n7066 ) | ( n7065 & ~n7070 ) | ( n7066 & ~n7070 ) ;
  assign n7072 = x321 & n6568 ;
  assign n7073 = ~x459 & n2185 ;
  assign n7074 = x328 & n2314 ;
  assign n7075 = x442 & n6509 ;
  assign n7076 = n2185 | n7075 ;
  assign n7077 = ( ~n7073 & n7074 ) | ( ~n7073 & n7076 ) | ( n7074 & n7076 ) ;
  assign n7078 = ( ~n6502 & n7072 ) | ( ~n6502 & n7077 ) | ( n7072 & n7077 ) ;
  assign n7079 = x857 & n6631 ;
  assign n7080 = ( ~n7071 & n7078 ) | ( ~n7071 & n7079 ) | ( n7078 & n7079 ) ;
  assign n7081 = n7071 | n7080 ;
  assign n7082 = x709 | n6904 ;
  assign n7083 = x1118 & n6904 ;
  assign n7084 = ( x962 & n7082 ) | ( x962 & ~n7083 ) | ( n7082 & ~n7083 ) ;
  assign n7085 = x710 & ~n6355 ;
  assign n7086 = x1106 & n6355 ;
  assign n7087 = ( ~x962 & n7085 ) | ( ~x962 & n7086 ) | ( n7085 & n7086 ) ;
  assign n7088 = x398 & n2314 ;
  assign n7089 = x348 & n6506 ;
  assign n7090 = x373 & n6509 ;
  assign n7091 = x423 & n2185 ;
  assign n7092 = n7090 | n7091 ;
  assign n7093 = n7089 | n7092 ;
  assign n7094 = ( ~n6502 & n7088 ) | ( ~n6502 & n7093 ) | ( n7088 & n7093 ) ;
  assign n7095 = x306 | n2904 ;
  assign n7096 = ~x1059 & n4339 ;
  assign n7097 = x199 & ~x1087 ;
  assign n7098 = ( n7095 & n7096 ) | ( n7095 & n7097 ) | ( n7096 & n7097 ) ;
  assign n7099 = n7095 & ~n7098 ;
  assign n7100 = n6498 & n7099 ;
  assign n7101 = x858 & n6631 ;
  assign n7102 = x630 & ~n7062 ;
  assign n7103 = x647 & n6832 ;
  assign n7104 = ~x725 & x1135 ;
  assign n7105 = x755 | x1135 ;
  assign n7106 = ( x1134 & n7104 ) | ( x1134 & ~n7105 ) | ( n7104 & ~n7105 ) ;
  assign n7107 = ( ~n7102 & n7103 ) | ( ~n7102 & n7106 ) | ( n7103 & n7106 ) ;
  assign n7108 = ( n6513 & n7102 ) | ( n6513 & n7107 ) | ( n7102 & n7107 ) ;
  assign n7109 = ( ~n7094 & n7101 ) | ( ~n7094 & n7108 ) | ( n7101 & n7108 ) ;
  assign n7110 = ( ~n7094 & n7100 ) | ( ~n7094 & n7109 ) | ( n7100 & n7109 ) ;
  assign n7111 = n7094 | n7110 ;
  assign n7112 = x842 & n6631 ;
  assign n7113 = x751 | x1135 ;
  assign n7114 = ~x701 & x1135 ;
  assign n7115 = ( x1134 & ~n7113 ) | ( x1134 & n7114 ) | ( ~n7113 & n7114 ) ;
  assign n7116 = x644 & ~x1135 ;
  assign n7117 = x715 & x1135 ;
  assign n7118 = ( ~x1134 & n7116 ) | ( ~x1134 & n7117 ) | ( n7116 & n7117 ) ;
  assign n7119 = ( n6513 & n7115 ) | ( n6513 & n7118 ) | ( n7115 & n7118 ) ;
  assign n7120 = n7112 | n7119 ;
  assign n7121 = x400 & n2314 ;
  assign n7122 = x374 & n6509 ;
  assign n7123 = n7121 | n7122 ;
  assign n7124 = x350 & n6506 ;
  assign n7125 = n7123 | n7124 ;
  assign n7126 = ( x425 & ~n2185 ) | ( x425 & n6502 ) | ( ~n2185 & n6502 ) ;
  assign n7127 = x425 & ~n7126 ;
  assign n7128 = ( ~n6502 & n7125 ) | ( ~n6502 & n7127 ) | ( n7125 & n7127 ) ;
  assign n7129 = x298 | n2904 ;
  assign n7130 = ~x1044 & n4339 ;
  assign n7131 = x199 & ~x1035 ;
  assign n7132 = n7130 | n7131 ;
  assign n7133 = ( n6498 & ~n7129 ) | ( n6498 & n7132 ) | ( ~n7129 & n7132 ) ;
  assign n7134 = ( n6498 & n7128 ) | ( n6498 & ~n7133 ) | ( n7128 & ~n7133 ) ;
  assign n7135 = n7120 | n7134 ;
  assign n7136 = x396 & n2314 ;
  assign n7137 = x371 & n6509 ;
  assign n7138 = ( ~n6502 & n7136 ) | ( ~n6502 & n7137 ) | ( n7136 & n7137 ) ;
  assign n7139 = x421 & n2185 ;
  assign n7140 = x322 & n6506 ;
  assign n7141 = n7139 | n7140 ;
  assign n7142 = ( ~n6502 & n7138 ) | ( ~n6502 & n7141 ) | ( n7138 & n7141 ) ;
  assign n7143 = ~x734 & n6581 ;
  assign n7144 = ~x756 & n6491 ;
  assign n7145 = x629 & ~x1135 ;
  assign n7146 = x628 & x1135 ;
  assign n7147 = ( ~x1134 & n7145 ) | ( ~x1134 & n7146 ) | ( n7145 & n7146 ) ;
  assign n7148 = ( ~n7143 & n7144 ) | ( ~n7143 & n7147 ) | ( n7144 & n7147 ) ;
  assign n7149 = ( n6513 & n7143 ) | ( n6513 & n7148 ) | ( n7143 & n7148 ) ;
  assign n7150 = n7142 | n7149 ;
  assign n7151 = x854 & n6631 ;
  assign n7152 = ~x1072 & n4339 ;
  assign n7153 = x309 | n2904 ;
  assign n7154 = x199 & ~x1051 ;
  assign n7155 = ( n7152 & n7153 ) | ( n7152 & ~n7154 ) | ( n7153 & ~n7154 ) ;
  assign n7156 = ( n6498 & n7152 ) | ( n6498 & ~n7155 ) | ( n7152 & ~n7155 ) ;
  assign n7157 = ( n6498 & n7151 ) | ( n6498 & ~n7156 ) | ( n7151 & ~n7156 ) ;
  assign n7158 = n7150 | n7157 ;
  assign n7159 = x199 & x1057 ;
  assign n7160 = ( n4623 & n6498 ) | ( n4623 & n7159 ) | ( n6498 & n7159 ) ;
  assign n7161 = x326 & n2314 ;
  assign n7162 = x439 & n6509 ;
  assign n7163 = x449 & n2185 ;
  assign n7164 = ( ~n7161 & n7162 ) | ( ~n7161 & n7163 ) | ( n7162 & n7163 ) ;
  assign n7165 = n7161 | n7164 ;
  assign n7166 = x461 & n6568 ;
  assign n7167 = ( ~n6502 & n7165 ) | ( ~n6502 & n7166 ) | ( n7165 & n7166 ) ;
  assign n7168 = ( ~x697 & x1134 ) | ( ~x697 & n6491 ) | ( x1134 & n6491 ) ;
  assign n7169 = x762 & n6680 ;
  assign n7170 = x867 | n6577 ;
  assign n7171 = ( n7168 & n7169 ) | ( n7168 & ~n7170 ) | ( n7169 & ~n7170 ) ;
  assign n7172 = n7168 & ~n7171 ;
  assign n7173 = ( x653 & x1136 ) | ( x653 & n6551 ) | ( x1136 & n6551 ) ;
  assign n7174 = x816 & ~x1136 ;
  assign n7175 = ( ~x1134 & n7173 ) | ( ~x1134 & n7174 ) | ( n7173 & n7174 ) ;
  assign n7176 = ( n6480 & n7172 ) | ( n6480 & n7175 ) | ( n7172 & n7175 ) ;
  assign n7177 = ( x693 & x1135 ) | ( x693 & n6581 ) | ( x1135 & n6581 ) ;
  assign n7178 = ( ~x1136 & n6832 ) | ( ~x1136 & n7177 ) | ( n6832 & n7177 ) ;
  assign n7179 = n7176 & ~n7178 ;
  assign n7180 = ( ~n7160 & n7167 ) | ( ~n7160 & n7179 ) | ( n7167 & n7179 ) ;
  assign n7181 = n7160 | n7180 ;
  assign n7182 = x715 & ~n6355 ;
  assign n7183 = x1123 & n6355 ;
  assign n7184 = ( ~x962 & n7182 ) | ( ~x962 & n7183 ) | ( n7182 & n7183 ) ;
  assign n7185 = x199 & ~x1043 ;
  assign n7186 = x200 | x307 ;
  assign n7187 = x200 & ~x1053 ;
  assign n7188 = ( x199 & n7186 ) | ( x199 & ~n7187 ) | ( n7186 & ~n7187 ) ;
  assign n7189 = ( n6498 & n7185 ) | ( n6498 & n7188 ) | ( n7185 & n7188 ) ;
  assign n7190 = x626 & ~n7062 ;
  assign n7191 = x641 & n6832 ;
  assign n7192 = x738 & n6581 ;
  assign n7193 = x761 & ~x1135 ;
  assign n7194 = x1134 & ~n7193 ;
  assign n7195 = ( n7191 & ~n7192 ) | ( n7191 & n7194 ) | ( ~n7192 & n7194 ) ;
  assign n7196 = ( n6513 & n7190 ) | ( n6513 & n7195 ) | ( n7190 & n7195 ) ;
  assign n7197 = ( ~n7185 & n7189 ) | ( ~n7185 & n7196 ) | ( n7189 & n7196 ) ;
  assign n7198 = x329 & n2314 ;
  assign n7199 = x440 & n6509 ;
  assign n7200 = ( ~n6502 & n7198 ) | ( ~n6502 & n7199 ) | ( n7198 & n7199 ) ;
  assign n7201 = x349 & n6506 ;
  assign n7202 = x454 & n2185 ;
  assign n7203 = ( ~n6502 & n7201 ) | ( ~n6502 & n7202 ) | ( n7201 & n7202 ) ;
  assign n7204 = n7200 | n7203 ;
  assign n7205 = x845 & n6631 ;
  assign n7206 = ( ~n7197 & n7204 ) | ( ~n7197 & n7205 ) | ( n7204 & n7205 ) ;
  assign n7207 = n7197 | n7206 ;
  assign n7208 = x839 & x1134 ;
  assign n7209 = x800 & ~x1134 ;
  assign n7210 = ( ~x1135 & n7208 ) | ( ~x1135 & n7209 ) | ( n7208 & n7209 ) ;
  assign n7211 = n6526 & n7210 ;
  assign n7212 = x462 & n6506 ;
  assign n7213 = x318 & n2314 ;
  assign n7214 = x377 & n6509 ;
  assign n7215 = n7213 | n7214 ;
  assign n7216 = n7212 | n7215 ;
  assign n7217 = ( x448 & ~n2185 ) | ( x448 & n6502 ) | ( ~n2185 & n6502 ) ;
  assign n7218 = x448 & ~n7217 ;
  assign n7219 = ( ~n6502 & n7216 ) | ( ~n6502 & n7218 ) | ( n7216 & n7218 ) ;
  assign n7220 = x199 & x1074 ;
  assign n7221 = ( n4656 & n6498 ) | ( n4656 & n7220 ) | ( n6498 & n7220 ) ;
  assign n7222 = x645 & ~x1135 ;
  assign n7223 = ~x669 & x1135 ;
  assign n7224 = ( ~x1134 & n7222 ) | ( ~x1134 & n7223 ) | ( n7222 & n7223 ) ;
  assign n7225 = x768 | x1135 ;
  assign n7226 = x705 & x1135 ;
  assign n7227 = ( x1134 & ~n7225 ) | ( x1134 & n7226 ) | ( ~n7225 & n7226 ) ;
  assign n7228 = ( n6513 & n7224 ) | ( n6513 & n7227 ) | ( n7224 & n7227 ) ;
  assign n7229 = n7221 | n7228 ;
  assign n7230 = ( ~n7211 & n7219 ) | ( ~n7211 & n7229 ) | ( n7219 & n7229 ) ;
  assign n7231 = n7211 | n7230 ;
  assign n7232 = ~x1049 & n4339 ;
  assign n7233 = x199 & ~x1080 ;
  assign n7234 = x303 | n2904 ;
  assign n7235 = ( n4339 & ~n7233 ) | ( n4339 & n7234 ) | ( ~n7233 & n7234 ) ;
  assign n7236 = ( n6498 & n7232 ) | ( n6498 & ~n7235 ) | ( n7232 & ~n7235 ) ;
  assign n7237 = n6498 & ~n7236 ;
  assign n7238 = ~x698 & x1135 ;
  assign n7239 = x767 | x1135 ;
  assign n7240 = ( x1134 & n7238 ) | ( x1134 & ~n7239 ) | ( n7238 & ~n7239 ) ;
  assign n7241 = x625 & x1135 ;
  assign n7242 = x608 & ~x1135 ;
  assign n7243 = ( ~x1134 & n7241 ) | ( ~x1134 & n7242 ) | ( n7241 & n7242 ) ;
  assign n7244 = ( n6513 & n7240 ) | ( n6513 & n7243 ) | ( n7240 & n7243 ) ;
  assign n7245 = n7237 | n7244 ;
  assign n7246 = x853 & n6631 ;
  assign n7247 = x369 & n6509 ;
  assign n7248 = ( x315 & x588 ) | ( x315 & n2381 ) | ( x588 & n2381 ) ;
  assign n7249 = ( ~x588 & n7247 ) | ( ~x588 & n7248 ) | ( n7247 & n7248 ) ;
  assign n7250 = x394 & n2314 ;
  assign n7251 = x419 & n2185 ;
  assign n7252 = ( ~n6502 & n7250 ) | ( ~n6502 & n7251 ) | ( n7250 & n7251 ) ;
  assign n7253 = ( ~n6502 & n7249 ) | ( ~n6502 & n7252 ) | ( n7249 & n7252 ) ;
  assign n7254 = ( ~n7245 & n7246 ) | ( ~n7245 & n7253 ) | ( n7246 & n7253 ) ;
  assign n7255 = n7245 | n7254 ;
  assign n7256 = x199 & x1063 ;
  assign n7257 = ( n4669 & n6498 ) | ( n4669 & n7256 ) | ( n6498 & n7256 ) ;
  assign n7258 = x807 & ~x1134 ;
  assign n7259 = x868 & x1134 ;
  assign n7260 = ( ~x1135 & n7258 ) | ( ~x1135 & n7259 ) | ( n7258 & n7259 ) ;
  assign n7261 = ~x1136 & n7260 ;
  assign n7262 = x687 & n6581 ;
  assign n7263 = ~x650 & x1135 ;
  assign n7264 = x636 & ~x1135 ;
  assign n7265 = ( ~x1134 & n7263 ) | ( ~x1134 & n7264 ) | ( n7263 & n7264 ) ;
  assign n7266 = n7262 | n7265 ;
  assign n7267 = ~x774 & n6491 ;
  assign n7268 = ( x1136 & n7266 ) | ( x1136 & n7267 ) | ( n7266 & n7267 ) ;
  assign n7269 = ( n6480 & n7261 ) | ( n6480 & n7268 ) | ( n7261 & n7268 ) ;
  assign n7270 = n7257 | n7269 ;
  assign n7271 = x325 & n2314 ;
  assign n7272 = x451 & n2185 ;
  assign n7273 = n7271 | n7272 ;
  assign n7274 = x353 & n6506 ;
  assign n7275 = n7273 | n7274 ;
  assign n7276 = x378 & n6594 ;
  assign n7277 = ( ~n6502 & n7275 ) | ( ~n6502 & n7276 ) | ( n7275 & n7276 ) ;
  assign n7278 = n7270 | n7277 ;
  assign n7279 = x651 | x1134 ;
  assign n7280 = x750 & x1134 ;
  assign n7281 = ( n6680 & ~n7279 ) | ( n6680 & n7280 ) | ( ~n7279 & n7280 ) ;
  assign n7282 = n6480 & ~n7281 ;
  assign n7283 = x684 & x1134 ;
  assign n7284 = x654 & ~x1134 ;
  assign n7285 = ( x1135 & n7283 ) | ( x1135 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7286 = x794 & ~x1134 ;
  assign n7287 = x880 & x1134 ;
  assign n7288 = ( ~x1135 & n7286 ) | ( ~x1135 & n7287 ) | ( n7286 & n7287 ) ;
  assign n7289 = ( x1136 & ~n7285 ) | ( x1136 & n7288 ) | ( ~n7285 & n7288 ) ;
  assign n7290 = n7282 & n7289 ;
  assign n7291 = x199 & x1081 ;
  assign n7292 = ( n4687 & n6498 ) | ( n4687 & n7291 ) | ( n6498 & n7291 ) ;
  assign n7293 = n7290 | n7292 ;
  assign n7294 = x356 & n6568 ;
  assign n7295 = x445 & n2185 ;
  assign n7296 = x405 & n2314 ;
  assign n7297 = x381 & n6509 ;
  assign n7298 = ( ~n7295 & n7296 ) | ( ~n7295 & n7297 ) | ( n7296 & n7297 ) ;
  assign n7299 = n7295 | n7298 ;
  assign n7300 = ( ~n6502 & n7294 ) | ( ~n6502 & n7299 ) | ( n7294 & n7299 ) ;
  assign n7301 = n7293 | n7300 ;
  assign n7302 = ~x945 & x988 ;
  assign n7303 = x773 & n7302 ;
  assign n7304 = x747 & n7303 ;
  assign n7305 = x731 & x775 ;
  assign n7306 = n7304 & n7305 ;
  assign n7307 = x769 & n7306 ;
  assign n7308 = ~x721 & n7307 ;
  assign n7309 = ~x769 & x794 ;
  assign n7310 = ( x731 & ~x795 ) | ( x731 & n7309 ) | ( ~x795 & n7309 ) ;
  assign n7311 = x771 & ~x800 ;
  assign n7312 = ( ~x731 & x795 ) | ( ~x731 & n7311 ) | ( x795 & n7311 ) ;
  assign n7313 = n7310 | n7312 ;
  assign n7314 = ~x775 & x816 ;
  assign n7315 = ( ~x721 & x813 ) | ( ~x721 & n7314 ) | ( x813 & n7314 ) ;
  assign n7316 = x775 & ~x816 ;
  assign n7317 = ( x721 & ~x813 ) | ( x721 & n7316 ) | ( ~x813 & n7316 ) ;
  assign n7318 = n7315 | n7317 ;
  assign n7319 = n7313 | n7318 ;
  assign n7320 = ~x773 & x801 ;
  assign n7321 = ~x747 & x807 ;
  assign n7322 = ~x765 & x798 ;
  assign n7323 = x769 & ~x794 ;
  assign n7324 = ( ~n7320 & n7322 ) | ( ~n7320 & n7323 ) | ( n7322 & n7323 ) ;
  assign n7325 = ( ~n7320 & n7321 ) | ( ~n7320 & n7324 ) | ( n7321 & n7324 ) ;
  assign n7326 = n7320 | n7325 ;
  assign n7327 = x765 & ~x798 ;
  assign n7328 = ~x771 & x800 ;
  assign n7329 = x773 & ~x801 ;
  assign n7330 = ( ~n7327 & n7328 ) | ( ~n7327 & n7329 ) | ( n7328 & n7329 ) ;
  assign n7331 = x747 & ~x807 ;
  assign n7332 = ( ~n7327 & n7330 ) | ( ~n7327 & n7331 ) | ( n7330 & n7331 ) ;
  assign n7333 = n7327 | n7332 ;
  assign n7334 = ( ~n7319 & n7326 ) | ( ~n7319 & n7333 ) | ( n7326 & n7333 ) ;
  assign n7335 = n7319 | n7334 ;
  assign n7336 = x721 & ~n7307 ;
  assign n7337 = ( n7308 & n7335 ) | ( n7308 & n7336 ) | ( n7335 & n7336 ) ;
  assign n7338 = x640 & x1136 ;
  assign n7339 = x795 & ~x1136 ;
  assign n7340 = ( ~n7062 & n7338 ) | ( ~n7062 & n7339 ) | ( n7338 & n7339 ) ;
  assign n7341 = ~x776 & x1136 ;
  assign n7342 = x851 & ~x1136 ;
  assign n7343 = ( n6491 & n7341 ) | ( n6491 & n7342 ) | ( n7341 & n7342 ) ;
  assign n7344 = n7340 | n7343 ;
  assign n7345 = ~x694 & x1134 ;
  assign n7346 = x732 | x1134 ;
  assign n7347 = ( n6551 & n7345 ) | ( n6551 & ~n7346 ) | ( n7345 & ~n7346 ) ;
  assign n7348 = n7344 | n7347 ;
  assign n7349 = n6480 & n7348 ;
  assign n7350 = x199 & x1045 ;
  assign n7351 = ( n4675 & n6498 ) | ( n4675 & n7350 ) | ( n6498 & n7350 ) ;
  assign n7352 = x379 & n6594 ;
  assign n7355 = x354 & n6506 ;
  assign n7353 = x403 & n2314 ;
  assign n7354 = x428 & n2185 ;
  assign n7356 = ( n7353 & n7354 ) | ( n7353 & ~n7355 ) | ( n7354 & ~n7355 ) ;
  assign n7357 = ( ~n6502 & n7355 ) | ( ~n6502 & n7356 ) | ( n7355 & n7356 ) ;
  assign n7358 = ( ~n7349 & n7352 ) | ( ~n7349 & n7357 ) | ( n7352 & n7357 ) ;
  assign n7359 = ( ~n7349 & n7351 ) | ( ~n7349 & n7358 ) | ( n7351 & n7358 ) ;
  assign n7360 = n7349 | n7359 ;
  assign n7361 = x1111 & n6904 ;
  assign n7362 = x723 | n6904 ;
  assign n7363 = ( x962 & ~n7361 ) | ( x962 & n7362 ) | ( ~n7361 & n7362 ) ;
  assign n7364 = x724 | n6904 ;
  assign n7365 = x1114 & n6904 ;
  assign n7366 = ( x962 & n7364 ) | ( x962 & ~n7365 ) | ( n7364 & ~n7365 ) ;
  assign n7367 = x1120 & n6904 ;
  assign n7368 = x725 | n6904 ;
  assign n7369 = ( x962 & ~n7367 ) | ( x962 & n7368 ) | ( ~n7367 & n7368 ) ;
  assign n7370 = x1126 & n6904 ;
  assign n7371 = x726 & ~n6904 ;
  assign n7372 = ( ~x962 & n7370 ) | ( ~x962 & n7371 ) | ( n7370 & n7371 ) ;
  assign n7373 = x727 & ~n6904 ;
  assign n7374 = x1102 & n6904 ;
  assign n7375 = ( ~x962 & n7373 ) | ( ~x962 & n7374 ) | ( n7373 & n7374 ) ;
  assign n7376 = x728 | n6904 ;
  assign n7377 = x1131 & n6904 ;
  assign n7378 = ( x962 & n7376 ) | ( x962 & ~n7377 ) | ( n7376 & ~n7377 ) ;
  assign n7379 = x729 & ~n6904 ;
  assign n7380 = x1104 & n6904 ;
  assign n7381 = ( ~x962 & n7379 ) | ( ~x962 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7382 = x730 & ~n6904 ;
  assign n7383 = x1106 & n6904 ;
  assign n7384 = ( ~x962 & n7382 ) | ( ~x962 & n7383 ) | ( n7382 & n7383 ) ;
  assign n7385 = ~x731 & n7304 ;
  assign n7386 = x731 & ~n7304 ;
  assign n7387 = ( n7335 & n7385 ) | ( n7335 & n7386 ) | ( n7385 & n7386 ) ;
  assign n7388 = x732 | n6355 ;
  assign n7389 = x1128 & n6355 ;
  assign n7390 = ( x962 & n7388 ) | ( x962 & ~n7389 ) | ( n7388 & ~n7389 ) ;
  assign n7391 = ~x1037 & n4339 ;
  assign n7392 = x199 & ~x1047 ;
  assign n7393 = x308 | n2904 ;
  assign n7394 = ( n7391 & ~n7392 ) | ( n7391 & n7393 ) | ( ~n7392 & n7393 ) ;
  assign n7395 = ~n7391 & n7394 ;
  assign n7396 = n6498 & n7395 ;
  assign n7397 = x777 | x1135 ;
  assign n7398 = ~x737 & x1135 ;
  assign n7399 = ( x1134 & ~n7397 ) | ( x1134 & n7398 ) | ( ~n7397 & n7398 ) ;
  assign n7400 = x648 & x1135 ;
  assign n7401 = x619 & ~x1135 ;
  assign n7402 = ( ~x1134 & n7400 ) | ( ~x1134 & n7401 ) | ( n7400 & n7401 ) ;
  assign n7403 = ( n6513 & n7399 ) | ( n6513 & n7402 ) | ( n7399 & n7402 ) ;
  assign n7404 = n7396 | n7403 ;
  assign n7405 = x424 & n2185 ;
  assign n7406 = x375 & n6509 ;
  assign n7407 = x399 & n2314 ;
  assign n7408 = ( x316 & x588 ) | ( x316 & n2381 ) | ( x588 & n2381 ) ;
  assign n7409 = ( ~x588 & n7407 ) | ( ~x588 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7410 = ( ~n7405 & n7406 ) | ( ~n7405 & n7409 ) | ( n7406 & n7409 ) ;
  assign n7411 = ( ~n6502 & n7405 ) | ( ~n6502 & n7410 ) | ( n7405 & n7410 ) ;
  assign n7412 = x838 & n6631 ;
  assign n7413 = ( ~n7404 & n7411 ) | ( ~n7404 & n7412 ) | ( n7411 & n7412 ) ;
  assign n7414 = n7404 | n7413 ;
  assign n7415 = x1119 & n6904 ;
  assign n7416 = x734 | n6904 ;
  assign n7417 = ( x962 & ~n7415 ) | ( x962 & n7416 ) | ( ~n7415 & n7416 ) ;
  assign n7418 = x1109 & n6904 ;
  assign n7419 = x735 & ~n6904 ;
  assign n7420 = ( ~x962 & n7418 ) | ( ~x962 & n7419 ) | ( n7418 & n7419 ) ;
  assign n7421 = x736 & ~n6904 ;
  assign n7422 = x1101 & n6904 ;
  assign n7423 = ( ~x962 & n7421 ) | ( ~x962 & n7422 ) | ( n7421 & n7422 ) ;
  assign n7424 = x737 | n6904 ;
  assign n7425 = x1122 & n6904 ;
  assign n7426 = ( x962 & n7424 ) | ( x962 & ~n7425 ) | ( n7424 & ~n7425 ) ;
  assign n7427 = x738 | n6904 ;
  assign n7428 = x1121 & n6904 ;
  assign n7429 = ( x962 & n7427 ) | ( x962 & ~n7428 ) | ( n7427 & ~n7428 ) ;
  assign n7430 = x832 & ~x952 ;
  assign n7431 = n6262 & n7430 ;
  assign n7432 = ~x1108 & n7431 ;
  assign n7433 = x739 | n7431 ;
  assign n7434 = ( x966 & ~n7432 ) | ( x966 & n7433 ) | ( ~n7432 & n7433 ) ;
  assign n7435 = ~x1114 & n7431 ;
  assign n7436 = x741 & ~n7431 ;
  assign n7437 = ( ~x966 & n7435 ) | ( ~x966 & n7436 ) | ( n7435 & n7436 ) ;
  assign n7438 = ~x1112 & n7431 ;
  assign n7439 = x742 & ~n7431 ;
  assign n7440 = ( ~x966 & n7438 ) | ( ~x966 & n7439 ) | ( n7438 & n7439 ) ;
  assign n7441 = ~x1109 & n7431 ;
  assign n7442 = x743 | n7431 ;
  assign n7443 = ( x966 & ~n7441 ) | ( x966 & n7442 ) | ( ~n7441 & n7442 ) ;
  assign n7444 = x744 & ~n7431 ;
  assign n7445 = ~x1131 & n7431 ;
  assign n7446 = ( ~x966 & n7444 ) | ( ~x966 & n7445 ) | ( n7444 & n7445 ) ;
  assign n7447 = x745 & ~n7431 ;
  assign n7448 = ~x1111 & n7431 ;
  assign n7449 = ( ~x966 & n7447 ) | ( ~x966 & n7448 ) | ( n7447 & n7448 ) ;
  assign n7450 = ~x1104 & n7431 ;
  assign n7451 = x746 | n7431 ;
  assign n7452 = ( x966 & ~n7450 ) | ( x966 & n7451 ) | ( ~n7450 & n7451 ) ;
  assign n7453 = ( x747 & n7303 ) | ( x747 & n7335 ) | ( n7303 & n7335 ) ;
  assign n7454 = ~n7304 & n7453 ;
  assign n7455 = ~x1106 & n7431 ;
  assign n7456 = x748 | n7431 ;
  assign n7457 = ( x966 & ~n7455 ) | ( x966 & n7456 ) | ( ~n7455 & n7456 ) ;
  assign n7458 = x749 | n7431 ;
  assign n7459 = ~x1105 & n7431 ;
  assign n7460 = ( x966 & n7458 ) | ( x966 & ~n7459 ) | ( n7458 & ~n7459 ) ;
  assign n7461 = x750 & ~n7431 ;
  assign n7462 = ~x1130 & n7431 ;
  assign n7463 = ( ~x966 & n7461 ) | ( ~x966 & n7462 ) | ( n7461 & n7462 ) ;
  assign n7464 = x751 & ~n7431 ;
  assign n7465 = ~x1123 & n7431 ;
  assign n7466 = ( ~x966 & n7464 ) | ( ~x966 & n7465 ) | ( n7464 & n7465 ) ;
  assign n7467 = ~x1124 & n7431 ;
  assign n7468 = x752 & ~n7431 ;
  assign n7469 = ( ~x966 & n7467 ) | ( ~x966 & n7468 ) | ( n7467 & n7468 ) ;
  assign n7470 = ~x1117 & n7431 ;
  assign n7471 = x753 & ~n7431 ;
  assign n7472 = ( ~x966 & n7470 ) | ( ~x966 & n7471 ) | ( n7470 & n7471 ) ;
  assign n7473 = ~x1118 & n7431 ;
  assign n7474 = x754 & ~n7431 ;
  assign n7475 = ( ~x966 & n7473 ) | ( ~x966 & n7474 ) | ( n7473 & n7474 ) ;
  assign n7476 = ~x1120 & n7431 ;
  assign n7477 = x755 & ~n7431 ;
  assign n7478 = ( ~x966 & n7476 ) | ( ~x966 & n7477 ) | ( n7476 & n7477 ) ;
  assign n7479 = ~x1119 & n7431 ;
  assign n7480 = x756 & ~n7431 ;
  assign n7481 = ( ~x966 & n7479 ) | ( ~x966 & n7480 ) | ( n7479 & n7480 ) ;
  assign n7482 = ~x1113 & n7431 ;
  assign n7483 = x757 & ~n7431 ;
  assign n7484 = ( ~x966 & n7482 ) | ( ~x966 & n7483 ) | ( n7482 & n7483 ) ;
  assign n7485 = ~x1101 & n7431 ;
  assign n7486 = x758 | n7431 ;
  assign n7487 = ( x966 & ~n7485 ) | ( x966 & n7486 ) | ( ~n7485 & n7486 ) ;
  assign n7488 = ~x1100 & n7431 ;
  assign n7489 = x759 | n7431 ;
  assign n7490 = ( x966 & ~n7488 ) | ( x966 & n7489 ) | ( ~n7488 & n7489 ) ;
  assign n7491 = x760 & ~n7431 ;
  assign n7492 = ~x1115 & n7431 ;
  assign n7493 = ( ~x966 & n7491 ) | ( ~x966 & n7492 ) | ( n7491 & n7492 ) ;
  assign n7494 = ~x1121 & n7431 ;
  assign n7495 = x761 & ~n7431 ;
  assign n7496 = ( ~x966 & n7494 ) | ( ~x966 & n7495 ) | ( n7494 & n7495 ) ;
  assign n7497 = x762 & ~n7431 ;
  assign n7498 = ~x1129 & n7431 ;
  assign n7499 = ( ~x966 & n7497 ) | ( ~x966 & n7498 ) | ( n7497 & n7498 ) ;
  assign n7500 = x763 | n7431 ;
  assign n7501 = ~x1103 & n7431 ;
  assign n7502 = ( x966 & n7500 ) | ( x966 & ~n7501 ) | ( n7500 & ~n7501 ) ;
  assign n7503 = x764 | n7431 ;
  assign n7504 = ~x1107 & n7431 ;
  assign n7505 = ( x966 & n7503 ) | ( x966 & ~n7504 ) | ( n7503 & ~n7504 ) ;
  assign n7506 = x773 | x775 ;
  assign n7507 = x747 | x765 ;
  assign n7508 = x721 | x731 ;
  assign n7509 = ( ~n7506 & n7507 ) | ( ~n7506 & n7508 ) | ( n7507 & n7508 ) ;
  assign n7510 = x794 | x800 ;
  assign n7511 = ( ~n7506 & n7509 ) | ( ~n7506 & n7510 ) | ( n7509 & n7510 ) ;
  assign n7512 = n7506 | n7511 ;
  assign n7513 = x765 & ~x945 ;
  assign n7514 = ( ~n7335 & n7512 ) | ( ~n7335 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7515 = x765 & x945 ;
  assign n7516 = ( x945 & n7514 ) | ( x945 & ~n7515 ) | ( n7514 & ~n7515 ) ;
  assign n7517 = ~x1110 & n7431 ;
  assign n7518 = x766 | n7431 ;
  assign n7519 = ( x966 & ~n7517 ) | ( x966 & n7518 ) | ( ~n7517 & n7518 ) ;
  assign n7520 = x767 & ~n7431 ;
  assign n7521 = ~x1116 & n7431 ;
  assign n7522 = ( ~x966 & n7520 ) | ( ~x966 & n7521 ) | ( n7520 & n7521 ) ;
  assign n7523 = ~x1125 & n7431 ;
  assign n7524 = x768 & ~n7431 ;
  assign n7525 = ( ~x966 & n7523 ) | ( ~x966 & n7524 ) | ( n7523 & n7524 ) ;
  assign n7526 = ( x769 & n7306 ) | ( x769 & n7335 ) | ( n7306 & n7335 ) ;
  assign n7527 = ~n7307 & n7526 ;
  assign n7528 = x770 & ~n7431 ;
  assign n7529 = ~x1126 & n7431 ;
  assign n7530 = ( ~x966 & n7528 ) | ( ~x966 & n7529 ) | ( n7528 & n7529 ) ;
  assign n7531 = ~n7335 & n7512 ;
  assign n7532 = x771 & x945 ;
  assign n7533 = ~x945 & x987 ;
  assign n7534 = ( ~n7531 & n7532 ) | ( ~n7531 & n7533 ) | ( n7532 & n7533 ) ;
  assign n7535 = x772 | n7431 ;
  assign n7536 = ~x1102 & n7431 ;
  assign n7537 = ( x966 & n7535 ) | ( x966 & ~n7536 ) | ( n7535 & ~n7536 ) ;
  assign n7538 = ( x773 & n7302 ) | ( x773 & ~n7531 ) | ( n7302 & ~n7531 ) ;
  assign n7539 = ~n7303 & n7538 ;
  assign n7540 = ~x1127 & n7431 ;
  assign n7541 = x774 & ~n7431 ;
  assign n7542 = ( ~x966 & n7540 ) | ( ~x966 & n7541 ) | ( n7540 & n7541 ) ;
  assign n7543 = x771 & x773 ;
  assign n7544 = x731 & x747 ;
  assign n7545 = ( n7513 & ~n7543 ) | ( n7513 & n7544 ) | ( ~n7543 & n7544 ) ;
  assign n7546 = n7543 & n7545 ;
  assign n7547 = ~x775 & n7546 ;
  assign n7548 = x775 & ~n7546 ;
  assign n7549 = ( n7335 & n7547 ) | ( n7335 & n7548 ) | ( n7547 & n7548 ) ;
  assign n7550 = x776 & ~n7431 ;
  assign n7551 = ~x1128 & n7431 ;
  assign n7552 = ( ~x966 & n7550 ) | ( ~x966 & n7551 ) | ( n7550 & n7551 ) ;
  assign n7553 = x777 & ~n7431 ;
  assign n7554 = ~x1122 & n7431 ;
  assign n7555 = ( ~x966 & n7553 ) | ( ~x966 & n7554 ) | ( n7553 & n7554 ) ;
  assign n7556 = x1046 | x1083 ;
  assign n7557 = x832 & x956 ;
  assign n7558 = ~n7556 & n7557 ;
  assign n7559 = ~x968 & x1085 ;
  assign n7560 = n7558 & n7559 ;
  assign n7561 = ~x1100 & n7560 ;
  assign n7562 = x778 & ~n7560 ;
  assign n7563 = ( n7560 & ~n7561 ) | ( n7560 & n7562 ) | ( ~n7561 & n7562 ) ;
  assign n7564 = x779 & ~n6314 ;
  assign n7565 = x780 & ~n6245 ;
  assign n7566 = x781 & ~n7560 ;
  assign n7567 = x1101 & n7560 ;
  assign n7568 = n7566 | n7567 ;
  assign n7569 = n1990 & ~n6273 ;
  assign n7570 = n6244 & n7569 ;
  assign n7571 = x783 & ~n7560 ;
  assign n7572 = x1109 & n7560 ;
  assign n7573 = n7571 | n7572 ;
  assign n7574 = x784 & ~n7560 ;
  assign n7575 = x1110 & n7560 ;
  assign n7576 = n7574 | n7575 ;
  assign n7577 = x785 & ~n7560 ;
  assign n7578 = x1102 & n7560 ;
  assign n7579 = n7577 | n7578 ;
  assign n7580 = ~x786 & x954 ;
  assign n7581 = ( x24 & n2127 ) | ( x24 & ~n7580 ) | ( n2127 & ~n7580 ) ;
  assign n7582 = x787 & ~n7560 ;
  assign n7583 = x1104 & n7560 ;
  assign n7584 = n7582 | n7583 ;
  assign n7585 = x788 & ~n7560 ;
  assign n7586 = x1105 & n7560 ;
  assign n7587 = n7585 | n7586 ;
  assign n7588 = x789 & ~n7560 ;
  assign n7589 = x1106 & n7560 ;
  assign n7590 = n7588 | n7589 ;
  assign n7591 = x790 & ~n7560 ;
  assign n7592 = x1107 & n7560 ;
  assign n7593 = n7591 | n7592 ;
  assign n7594 = x791 & ~n7560 ;
  assign n7595 = x1108 & n7560 ;
  assign n7596 = n7594 | n7595 ;
  assign n7597 = x792 & ~n7560 ;
  assign n7598 = x1103 & n7560 ;
  assign n7599 = n7597 | n7598 ;
  assign n7600 = x968 & x1085 ;
  assign n7601 = n7558 & n7600 ;
  assign n7602 = ~x1130 & n7601 ;
  assign n7603 = x794 & ~n7601 ;
  assign n7604 = ( n7601 & ~n7602 ) | ( n7601 & n7603 ) | ( ~n7602 & n7603 ) ;
  assign n7605 = x795 & ~n7601 ;
  assign n7606 = x1128 & n7601 ;
  assign n7607 = n7605 | n7606 ;
  assign n7608 = x281 | x282 ;
  assign n7609 = ~x264 & n7608 ;
  assign n7610 = x278 & x279 ;
  assign n7611 = ( x266 & x269 ) | ( x266 & x280 ) | ( x269 & x280 ) ;
  assign n7612 = ( x266 & ~n7610 ) | ( x266 & n7611 ) | ( ~n7610 & n7611 ) ;
  assign n7613 = x266 & ~n7612 ;
  assign n7614 = ~n6463 & n7613 ;
  assign n7615 = ( ~x264 & n7608 ) | ( ~x264 & n7614 ) | ( n7608 & n7614 ) ;
  assign n7616 = x264 & ~n7614 ;
  assign n7617 = ( ~n7609 & n7615 ) | ( ~n7609 & n7616 ) | ( n7615 & n7616 ) ;
  assign n7618 = x798 & ~n7601 ;
  assign n7619 = x1124 & n7601 ;
  assign n7620 = n7618 | n7619 ;
  assign n7621 = x799 | n7601 ;
  assign n7622 = x1107 & n7601 ;
  assign n7623 = n7621 & ~n7622 ;
  assign n7624 = x800 & ~n7601 ;
  assign n7625 = x1125 & n7601 ;
  assign n7626 = n7624 | n7625 ;
  assign n7627 = x801 & ~n7601 ;
  assign n7628 = x1126 & n7601 ;
  assign n7629 = n7627 | n7628 ;
  assign n7630 = x803 | n7601 ;
  assign n7631 = x1106 & n7601 ;
  assign n7632 = n7630 & ~n7631 ;
  assign n7633 = x804 & ~n7601 ;
  assign n7634 = x1109 & n7601 ;
  assign n7635 = n7633 | n7634 ;
  assign n7636 = x270 & ~n6462 ;
  assign n7637 = ~x270 & n6462 ;
  assign n7638 = n7636 | n7637 ;
  assign n7639 = x807 & ~n7601 ;
  assign n7640 = x1127 & n7601 ;
  assign n7641 = n7639 | n7640 ;
  assign n7642 = x808 & ~n7601 ;
  assign n7643 = x1101 & n7601 ;
  assign n7644 = n7642 | n7643 ;
  assign n7645 = x809 | n7601 ;
  assign n7646 = x1103 & n7601 ;
  assign n7647 = n7645 & ~n7646 ;
  assign n7648 = x810 & ~n7601 ;
  assign n7649 = x1108 & n7601 ;
  assign n7650 = n7648 | n7649 ;
  assign n7651 = x811 & ~n7601 ;
  assign n7652 = x1102 & n7601 ;
  assign n7653 = n7651 | n7652 ;
  assign n7654 = x812 | n7601 ;
  assign n7655 = x1104 & n7601 ;
  assign n7656 = n7654 & ~n7655 ;
  assign n7657 = x813 & ~n7601 ;
  assign n7658 = x1131 & n7601 ;
  assign n7659 = n7657 | n7658 ;
  assign n7660 = x814 | n7601 ;
  assign n7661 = x1105 & n7601 ;
  assign n7662 = n7660 & ~n7661 ;
  assign n7663 = x815 & ~n7601 ;
  assign n7664 = x1110 & n7601 ;
  assign n7665 = n7663 | n7664 ;
  assign n7666 = x816 & ~n7601 ;
  assign n7667 = x1129 & n7601 ;
  assign n7668 = n7666 | n7667 ;
  assign n7669 = x269 & n6460 ;
  assign n7670 = x269 | n6460 ;
  assign n7671 = ~n7669 & n7670 ;
  assign n7672 = n3446 | n3448 ;
  assign n7673 = x264 & x265 ;
  assign n7674 = x265 & n6464 ;
  assign n7675 = ( n6465 & n7673 ) | ( n6465 & ~n7674 ) | ( n7673 & ~n7674 ) ;
  assign n7676 = x277 & n7637 ;
  assign n7677 = x277 | n7637 ;
  assign n7678 = ~n7676 & n7677 ;
  assign n7679 = x811 | x893 ;
  assign n7680 = n1426 & ~n2180 ;
  assign n7681 = ( x982 & n1433 ) | ( x982 & ~n7680 ) | ( n1433 & ~n7680 ) ;
  assign n7682 = n1957 & ~n7681 ;
  assign n7683 = ( ~x1127 & x1128 ) | ( ~x1127 & x1129 ) | ( x1128 & x1129 ) ;
  assign n7684 = ( x1127 & x1128 ) | ( x1127 & x1129 ) | ( x1128 & x1129 ) ;
  assign n7685 = ( x1127 & n7683 ) | ( x1127 & ~n7684 ) | ( n7683 & ~n7684 ) ;
  assign n7686 = ( ~x1130 & x1131 ) | ( ~x1130 & n7685 ) | ( x1131 & n7685 ) ;
  assign n7687 = ( x1130 & x1131 ) | ( x1130 & n7685 ) | ( x1131 & n7685 ) ;
  assign n7688 = ( x1130 & n7686 ) | ( x1130 & ~n7687 ) | ( n7686 & ~n7687 ) ;
  assign n7689 = ( ~x1124 & x1125 ) | ( ~x1124 & x1126 ) | ( x1125 & x1126 ) ;
  assign n7690 = ( x1124 & x1125 ) | ( x1124 & x1126 ) | ( x1125 & x1126 ) ;
  assign n7691 = ( x1124 & n7689 ) | ( x1124 & ~n7690 ) | ( n7689 & ~n7690 ) ;
  assign n7692 = n7688 & ~n7691 ;
  assign n7693 = x123 & ~n1467 ;
  assign n7694 = ( ~n7688 & n7691 ) | ( ~n7688 & n7693 ) | ( n7691 & n7693 ) ;
  assign n7695 = x825 & n7693 ;
  assign n7696 = ( n7692 & n7694 ) | ( n7692 & ~n7695 ) | ( n7694 & ~n7695 ) ;
  assign n7697 = ( ~x1116 & x1117 ) | ( ~x1116 & x1120 ) | ( x1117 & x1120 ) ;
  assign n7698 = ( x1116 & x1117 ) | ( x1116 & x1120 ) | ( x1117 & x1120 ) ;
  assign n7699 = ( x1116 & n7697 ) | ( x1116 & ~n7698 ) | ( n7697 & ~n7698 ) ;
  assign n7700 = x1122 & x1123 ;
  assign n7701 = x1122 | x1123 ;
  assign n7702 = ~n7700 & n7701 ;
  assign n7703 = x1118 & x1119 ;
  assign n7704 = x1118 | x1119 ;
  assign n7705 = ~n7703 & n7704 ;
  assign n7706 = ( x1121 & n7702 ) | ( x1121 & n7705 ) | ( n7702 & n7705 ) ;
  assign n7707 = ( ~x1121 & n7702 ) | ( ~x1121 & n7705 ) | ( n7702 & n7705 ) ;
  assign n7708 = ( x1121 & ~n7706 ) | ( x1121 & n7707 ) | ( ~n7706 & n7707 ) ;
  assign n7709 = ( n7693 & ~n7699 ) | ( n7693 & n7708 ) | ( ~n7699 & n7708 ) ;
  assign n7710 = n7699 & ~n7708 ;
  assign n7711 = x826 & n7693 ;
  assign n7712 = ( n7709 & n7710 ) | ( n7709 & ~n7711 ) | ( n7710 & ~n7711 ) ;
  assign n7713 = x827 & n7693 ;
  assign n7714 = ( x1102 & x1104 ) | ( x1102 & x1105 ) | ( x1104 & x1105 ) ;
  assign n7715 = ( ~x1102 & x1104 ) | ( ~x1102 & x1105 ) | ( x1104 & x1105 ) ;
  assign n7716 = ( x1102 & ~n7714 ) | ( x1102 & n7715 ) | ( ~n7714 & n7715 ) ;
  assign n7717 = ( ~x1106 & x1107 ) | ( ~x1106 & n7716 ) | ( x1107 & n7716 ) ;
  assign n7718 = ( x1106 & x1107 ) | ( x1106 & n7716 ) | ( x1107 & n7716 ) ;
  assign n7719 = ( x1106 & n7717 ) | ( x1106 & ~n7718 ) | ( n7717 & ~n7718 ) ;
  assign n7720 = ( x1100 & x1101 ) | ( x1100 & x1103 ) | ( x1101 & x1103 ) ;
  assign n7721 = ( ~x1100 & x1101 ) | ( ~x1100 & x1103 ) | ( x1101 & x1103 ) ;
  assign n7722 = ( x1100 & ~n7720 ) | ( x1100 & n7721 ) | ( ~n7720 & n7721 ) ;
  assign n7723 = n7719 & ~n7722 ;
  assign n7724 = ( n7693 & ~n7719 ) | ( n7693 & n7722 ) | ( ~n7719 & n7722 ) ;
  assign n7725 = ( ~n7713 & n7723 ) | ( ~n7713 & n7724 ) | ( n7723 & n7724 ) ;
  assign n7726 = ( ~x1110 & x1114 ) | ( ~x1110 & x1115 ) | ( x1114 & x1115 ) ;
  assign n7727 = ( x1110 & x1114 ) | ( x1110 & x1115 ) | ( x1114 & x1115 ) ;
  assign n7728 = ( x1110 & n7726 ) | ( x1110 & ~n7727 ) | ( n7726 & ~n7727 ) ;
  assign n7729 = ( ~x1108 & x1112 ) | ( ~x1108 & x1113 ) | ( x1112 & x1113 ) ;
  assign n7730 = ( x1108 & x1112 ) | ( x1108 & x1113 ) | ( x1112 & x1113 ) ;
  assign n7731 = ( x1108 & n7729 ) | ( x1108 & ~n7730 ) | ( n7729 & ~n7730 ) ;
  assign n7732 = ( ~x1109 & x1111 ) | ( ~x1109 & n7731 ) | ( x1111 & n7731 ) ;
  assign n7733 = ( x1109 & x1111 ) | ( x1109 & n7731 ) | ( x1111 & n7731 ) ;
  assign n7734 = ( x1109 & n7732 ) | ( x1109 & ~n7733 ) | ( n7732 & ~n7733 ) ;
  assign n7735 = n7728 & ~n7734 ;
  assign n7736 = ( n7693 & ~n7728 ) | ( n7693 & n7734 ) | ( ~n7728 & n7734 ) ;
  assign n7737 = x828 & n7693 ;
  assign n7738 = ( n7735 & n7736 ) | ( n7735 & ~n7737 ) | ( n7736 & ~n7737 ) ;
  assign n7739 = ~x951 & x1092 ;
  assign n7740 = ~n2180 & n4308 ;
  assign n7741 = ( x1092 & n7739 ) | ( x1092 & n7740 ) | ( n7739 & n7740 ) ;
  assign n7742 = x281 & n7613 ;
  assign n7743 = x281 | n7613 ;
  assign n7744 = ~n7742 & n7743 ;
  assign n7745 = ~x832 & n1431 ;
  assign n7746 = n2532 & n7745 ;
  assign n7747 = x833 & ~n1430 ;
  assign n7748 = n1431 | n7747 ;
  assign n7749 = x946 & n1430 ;
  assign n7750 = x282 & ~n6461 ;
  assign n7751 = n6462 | n7750 ;
  assign n7752 = x837 & x955 ;
  assign n7753 = ~x955 & x1049 ;
  assign n7754 = n7752 | n7753 ;
  assign n7755 = x838 & x955 ;
  assign n7756 = ~x955 & x1047 ;
  assign n7757 = n7755 | n7756 ;
  assign n7758 = x839 & x955 ;
  assign n7759 = ~x955 & x1074 ;
  assign n7760 = n7758 | n7759 ;
  assign n7761 = x840 & ~n1430 ;
  assign n7762 = x1196 & n1430 ;
  assign n7763 = n7761 | n7762 ;
  assign n7764 = x842 & x955 ;
  assign n7765 = ~x955 & x1035 ;
  assign n7766 = n7764 | n7765 ;
  assign n7767 = x843 & x955 ;
  assign n7768 = ~x955 & x1079 ;
  assign n7769 = n7767 | n7768 ;
  assign n7770 = x844 & x955 ;
  assign n7771 = ~x955 & x1078 ;
  assign n7772 = n7770 | n7771 ;
  assign n7773 = x845 & x955 ;
  assign n7774 = ~x955 & x1043 ;
  assign n7775 = n7773 | n7774 ;
  assign n7776 = ( x846 & ~n4690 ) | ( x846 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n7777 = ( x846 & n4690 ) | ( x846 & ~n4691 ) | ( n4690 & ~n4691 ) ;
  assign n7778 = ( x1134 & n7776 ) | ( x1134 & n7777 ) | ( n7776 & n7777 ) ;
  assign n7779 = x847 & x955 ;
  assign n7780 = ~x955 & x1055 ;
  assign n7781 = n7779 | n7780 ;
  assign n7782 = x848 & x955 ;
  assign n7783 = ~x955 & x1039 ;
  assign n7784 = n7782 | n7783 ;
  assign n7785 = x849 & ~n1430 ;
  assign n7786 = x1198 & n1430 ;
  assign n7787 = n7785 | n7786 ;
  assign n7788 = x850 & x955 ;
  assign n7789 = ~x955 & x1048 ;
  assign n7790 = n7788 | n7789 ;
  assign n7791 = x851 & x955 ;
  assign n7792 = ~x955 & x1045 ;
  assign n7793 = n7791 | n7792 ;
  assign n7794 = x852 & x955 ;
  assign n7795 = ~x955 & x1062 ;
  assign n7796 = n7794 | n7795 ;
  assign n7797 = x853 & x955 ;
  assign n7798 = ~x955 & x1080 ;
  assign n7799 = n7797 | n7798 ;
  assign n7800 = x854 & x955 ;
  assign n7801 = ~x955 & x1051 ;
  assign n7802 = n7800 | n7801 ;
  assign n7803 = x855 & x955 ;
  assign n7804 = ~x955 & x1065 ;
  assign n7805 = n7803 | n7804 ;
  assign n7806 = x856 & x955 ;
  assign n7807 = ~x955 & x1067 ;
  assign n7808 = n7806 | n7807 ;
  assign n7809 = x857 & x955 ;
  assign n7810 = ~x955 & x1058 ;
  assign n7811 = n7809 | n7810 ;
  assign n7812 = x858 & x955 ;
  assign n7813 = ~x955 & x1087 ;
  assign n7814 = n7812 | n7813 ;
  assign n7815 = x859 & x955 ;
  assign n7816 = ~x955 & x1070 ;
  assign n7817 = n7815 | n7816 ;
  assign n7818 = x860 & x955 ;
  assign n7819 = ~x955 & x1076 ;
  assign n7820 = n7818 | n7819 ;
  assign n7821 = ( x861 & n4690 ) | ( x861 & ~n4691 ) | ( n4690 & ~n4691 ) ;
  assign n7822 = ( x861 & ~n4690 ) | ( x861 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n7823 = ( x1141 & n7821 ) | ( x1141 & n7822 ) | ( n7821 & n7822 ) ;
  assign n7824 = ( x862 & n4690 ) | ( x862 & ~n4691 ) | ( n4690 & ~n4691 ) ;
  assign n7825 = ( x862 & ~n4690 ) | ( x862 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n7826 = ( x1139 & n7824 ) | ( x1139 & n7825 ) | ( n7824 & n7825 ) ;
  assign n7827 = x863 & ~n1430 ;
  assign n7828 = x1199 & n1430 ;
  assign n7829 = n7827 | n7828 ;
  assign n7830 = x864 & ~n1430 ;
  assign n7831 = x1197 & n1430 ;
  assign n7832 = n7830 | n7831 ;
  assign n7833 = x865 & x955 ;
  assign n7834 = ~x955 & x1040 ;
  assign n7835 = n7833 | n7834 ;
  assign n7836 = x866 & x955 ;
  assign n7837 = ~x955 & x1053 ;
  assign n7838 = n7836 | n7837 ;
  assign n7839 = x867 & x955 ;
  assign n7840 = ~x955 & x1057 ;
  assign n7841 = n7839 | n7840 ;
  assign n7842 = x868 & x955 ;
  assign n7843 = ~x955 & x1063 ;
  assign n7844 = n7842 | n7843 ;
  assign n7845 = ( x869 & ~n4690 ) | ( x869 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n7846 = ( x869 & n4690 ) | ( x869 & ~n4691 ) | ( n4690 & ~n4691 ) ;
  assign n7847 = ( x1140 & n7845 ) | ( x1140 & n7846 ) | ( n7845 & n7846 ) ;
  assign n7848 = x870 & x955 ;
  assign n7849 = ~x955 & x1069 ;
  assign n7850 = n7848 | n7849 ;
  assign n7851 = x871 & x955 ;
  assign n7852 = ~x955 & x1072 ;
  assign n7853 = n7851 | n7852 ;
  assign n7854 = x872 & x955 ;
  assign n7855 = ~x955 & x1084 ;
  assign n7856 = n7854 | n7855 ;
  assign n7857 = x873 & x955 ;
  assign n7858 = ~x955 & x1044 ;
  assign n7859 = n7857 | n7858 ;
  assign n7860 = x874 & x955 ;
  assign n7861 = ~x955 & x1036 ;
  assign n7862 = n7860 | n7861 ;
  assign n7863 = ( x875 & n4690 ) | ( x875 & ~n4691 ) | ( n4690 & ~n4691 ) ;
  assign n7864 = ( x875 & ~n4690 ) | ( x875 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n7865 = ( x1136 & n7863 ) | ( x1136 & n7864 ) | ( n7863 & n7864 ) ;
  assign n7866 = x876 & x955 ;
  assign n7867 = ~x955 & x1037 ;
  assign n7868 = n7866 | n7867 ;
  assign n7869 = ( x877 & n4690 ) | ( x877 & ~n4691 ) | ( n4690 & ~n4691 ) ;
  assign n7870 = ( x877 & ~n4690 ) | ( x877 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n7871 = ( x1138 & n7869 ) | ( x1138 & n7870 ) | ( n7869 & n7870 ) ;
  assign n7872 = ( x878 & n4690 ) | ( x878 & ~n4691 ) | ( n4690 & ~n4691 ) ;
  assign n7873 = ( x878 & ~n4690 ) | ( x878 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n7874 = ( x1137 & n7872 ) | ( x1137 & n7873 ) | ( n7872 & n7873 ) ;
  assign n7875 = ( x879 & ~n4690 ) | ( x879 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n7876 = ( x879 & n4690 ) | ( x879 & ~n4691 ) | ( n4690 & ~n4691 ) ;
  assign n7877 = ( x1135 & n7875 ) | ( x1135 & n7876 ) | ( n7875 & n7876 ) ;
  assign n7878 = x880 & x955 ;
  assign n7879 = ~x955 & x1081 ;
  assign n7880 = n7878 | n7879 ;
  assign n7881 = x881 & x955 ;
  assign n7882 = ~x955 & x1059 ;
  assign n7883 = n7881 | n7882 ;
  assign n7884 = ~x883 & n7693 ;
  assign n7885 = x1107 & ~n7693 ;
  assign n7886 = n7884 | n7885 ;
  assign n7887 = ~x884 & n7693 ;
  assign n7888 = x1124 & ~n7693 ;
  assign n7889 = n7887 | n7888 ;
  assign n7890 = ~x885 & n7693 ;
  assign n7891 = x1125 & ~n7693 ;
  assign n7892 = n7890 | n7891 ;
  assign n7893 = ~x886 & n7693 ;
  assign n7894 = x1109 & ~n7693 ;
  assign n7895 = n7893 | n7894 ;
  assign n7896 = ~x887 & n7693 ;
  assign n7897 = x1100 & ~n7693 ;
  assign n7898 = n7896 | n7897 ;
  assign n7899 = ~x888 & n7693 ;
  assign n7900 = x1120 & ~n7693 ;
  assign n7901 = n7899 | n7900 ;
  assign n7902 = ~x889 & n7693 ;
  assign n7903 = x1103 & ~n7693 ;
  assign n7904 = n7902 | n7903 ;
  assign n7905 = ~x890 & n7693 ;
  assign n7906 = x1126 & ~n7693 ;
  assign n7907 = n7905 | n7906 ;
  assign n7908 = ~x891 & n7693 ;
  assign n7909 = x1116 & ~n7693 ;
  assign n7910 = n7908 | n7909 ;
  assign n7911 = ~x892 & n7693 ;
  assign n7912 = x1101 & ~n7693 ;
  assign n7913 = n7911 | n7912 ;
  assign n7914 = x107 | n1242 ;
  assign n7915 = ~x894 & n7693 ;
  assign n7916 = x1119 & ~n7693 ;
  assign n7917 = n7915 | n7916 ;
  assign n7918 = ~x895 & n7693 ;
  assign n7919 = x1113 & ~n7693 ;
  assign n7920 = n7918 | n7919 ;
  assign n7921 = ~x896 & n7693 ;
  assign n7922 = x1118 & ~n7693 ;
  assign n7923 = n7921 | n7922 ;
  assign n7924 = ~x898 & n7693 ;
  assign n7925 = x1129 & ~n7693 ;
  assign n7926 = n7924 | n7925 ;
  assign n7927 = ~x899 & n7693 ;
  assign n7928 = x1115 & ~n7693 ;
  assign n7929 = n7927 | n7928 ;
  assign n7930 = ~x900 & n7693 ;
  assign n7931 = x1110 & ~n7693 ;
  assign n7932 = n7930 | n7931 ;
  assign n7933 = ~x902 & n7693 ;
  assign n7934 = x1111 & ~n7693 ;
  assign n7935 = n7933 | n7934 ;
  assign n7936 = ~x903 & n7693 ;
  assign n7937 = x1121 & ~n7693 ;
  assign n7938 = n7936 | n7937 ;
  assign n7939 = ~x904 & n7693 ;
  assign n7940 = x1127 & ~n7693 ;
  assign n7941 = n7939 | n7940 ;
  assign n7942 = ~x905 & n7693 ;
  assign n7943 = x1131 & ~n7693 ;
  assign n7944 = n7942 | n7943 ;
  assign n7945 = ~x906 & n7693 ;
  assign n7946 = x1128 & ~n7693 ;
  assign n7947 = n7945 | n7946 ;
  assign n7948 = ~x782 & x907 ;
  assign n7949 = x604 | x624 ;
  assign n7950 = ( ~x624 & x979 ) | ( ~x624 & n7949 ) | ( x979 & n7949 ) ;
  assign n7951 = ~x598 & x615 ;
  assign n7952 = ( x598 & x979 ) | ( x598 & n7951 ) | ( x979 & n7951 ) ;
  assign n7953 = ( x782 & n7948 ) | ( x782 & ~n7952 ) | ( n7948 & ~n7952 ) ;
  assign n7954 = ( n7948 & n7950 ) | ( n7948 & n7953 ) | ( n7950 & n7953 ) ;
  assign n7955 = ~x908 & n7693 ;
  assign n7956 = x1122 & ~n7693 ;
  assign n7957 = n7955 | n7956 ;
  assign n7958 = ~x909 & n7693 ;
  assign n7959 = x1105 & ~n7693 ;
  assign n7960 = n7958 | n7959 ;
  assign n7961 = ~x910 & n7693 ;
  assign n7962 = x1117 & ~n7693 ;
  assign n7963 = n7961 | n7962 ;
  assign n7964 = ~x911 & n7693 ;
  assign n7965 = x1130 & ~n7693 ;
  assign n7966 = n7964 | n7965 ;
  assign n7967 = ~x912 & n7693 ;
  assign n7968 = x1114 & ~n7693 ;
  assign n7969 = n7967 | n7968 ;
  assign n7970 = ~x913 & n7693 ;
  assign n7971 = x1106 & ~n7693 ;
  assign n7972 = n7970 | n7971 ;
  assign n7973 = ~x266 & x280 ;
  assign n7974 = x280 & x992 ;
  assign n7975 = ( n6459 & n7973 ) | ( n6459 & ~n7974 ) | ( n7973 & ~n7974 ) ;
  assign n7976 = ~x915 & n7693 ;
  assign n7977 = x1108 & ~n7693 ;
  assign n7978 = n7976 | n7977 ;
  assign n7979 = ~x916 & n7693 ;
  assign n7980 = x1123 & ~n7693 ;
  assign n7981 = n7979 | n7980 ;
  assign n7982 = ~x917 & n7693 ;
  assign n7983 = x1112 & ~n7693 ;
  assign n7984 = n7982 | n7983 ;
  assign n7985 = ~x918 & n7693 ;
  assign n7986 = x1104 & ~n7693 ;
  assign n7987 = n7985 | n7986 ;
  assign n7988 = ~x919 & n7693 ;
  assign n7989 = x1102 & ~n7693 ;
  assign n7990 = n7988 | n7989 ;
  assign n7991 = x920 & ~x1093 ;
  assign n7992 = x1093 & x1139 ;
  assign n7993 = n7991 | n7992 ;
  assign n7994 = x921 & ~x1093 ;
  assign n7995 = x1093 & x1140 ;
  assign n7996 = n7994 | n7995 ;
  assign n7997 = x922 & ~x1093 ;
  assign n7998 = x1093 & x1152 ;
  assign n7999 = n7997 | n7998 ;
  assign n8000 = x923 & ~x1093 ;
  assign n8001 = x1093 & x1154 ;
  assign n8002 = n8000 | n8001 ;
  assign n8003 = x311 & ~x312 ;
  assign n8004 = n4983 & n8003 ;
  assign n8005 = x925 & ~x1093 ;
  assign n8006 = x1093 & x1155 ;
  assign n8007 = n8005 | n8006 ;
  assign n8008 = x926 & ~x1093 ;
  assign n8009 = x1093 & x1157 ;
  assign n8010 = n8008 | n8009 ;
  assign n8011 = x927 & ~x1093 ;
  assign n8012 = x1093 & x1145 ;
  assign n8013 = n8011 | n8012 ;
  assign n8014 = x928 & ~x1093 ;
  assign n8015 = x1093 & x1136 ;
  assign n8016 = n8014 | n8015 ;
  assign n8017 = x929 & ~x1093 ;
  assign n8018 = x1093 & x1144 ;
  assign n8019 = n8017 | n8018 ;
  assign n8020 = x930 & ~x1093 ;
  assign n8021 = x1093 & x1134 ;
  assign n8022 = n8020 | n8021 ;
  assign n8023 = x931 & ~x1093 ;
  assign n8024 = x1093 & x1150 ;
  assign n8025 = n8023 | n8024 ;
  assign n8026 = x932 & ~x1093 ;
  assign n8027 = x1093 & x1142 ;
  assign n8028 = n8026 | n8027 ;
  assign n8029 = x933 & ~x1093 ;
  assign n8030 = x1093 & x1137 ;
  assign n8031 = n8029 | n8030 ;
  assign n8032 = x934 & ~x1093 ;
  assign n8033 = x1093 & x1147 ;
  assign n8034 = n8032 | n8033 ;
  assign n8035 = x935 & ~x1093 ;
  assign n8036 = x1093 & x1141 ;
  assign n8037 = n8035 | n8036 ;
  assign n8038 = x936 & ~x1093 ;
  assign n8039 = x1093 & x1149 ;
  assign n8040 = n8038 | n8039 ;
  assign n8041 = x937 & ~x1093 ;
  assign n8042 = x1093 & x1148 ;
  assign n8043 = n8041 | n8042 ;
  assign n8044 = x938 & ~x1093 ;
  assign n8045 = x1093 & x1135 ;
  assign n8046 = n8044 | n8045 ;
  assign n8047 = x939 & ~x1093 ;
  assign n8048 = x1093 & x1146 ;
  assign n8049 = n8047 | n8048 ;
  assign n8050 = x940 & ~x1093 ;
  assign n8051 = x1093 & x1138 ;
  assign n8052 = n8050 | n8051 ;
  assign n8053 = x941 & ~x1093 ;
  assign n8054 = x1093 & x1153 ;
  assign n8055 = n8053 | n8054 ;
  assign n8056 = x942 & ~x1093 ;
  assign n8057 = x1093 & x1156 ;
  assign n8058 = n8056 | n8057 ;
  assign n8059 = x943 & ~x1093 ;
  assign n8060 = x1093 & x1151 ;
  assign n8061 = n8059 | n8060 ;
  assign n8062 = x944 & ~x1093 ;
  assign n8063 = x1093 & x1143 ;
  assign n8064 = n8062 | n8063 ;
  assign n8065 = n1981 | n1985 ;
  assign n8066 = ~x782 & x947 ;
  assign n8067 = x624 | x979 ;
  assign n8068 = ( x782 & n8066 ) | ( x782 & n8067 ) | ( n8066 & n8067 ) ;
  assign n8069 = ~x598 & x979 ;
  assign n8070 = ( n8066 & n8068 ) | ( n8066 & ~n8069 ) | ( n8068 & ~n8069 ) ;
  assign n8071 = x266 & x992 ;
  assign n8072 = x266 | x992 ;
  assign n8073 = ~n8071 & n8072 ;
  assign n8074 = ~x949 & x954 ;
  assign n8075 = ( x313 & ~n4990 ) | ( x313 & n8074 ) | ( ~n4990 & n8074 ) ;
  assign n8076 = x957 & x1092 ;
  assign n8077 = x31 | n8076 ;
  assign n8078 = ~x782 & x960 ;
  assign n8079 = ~x230 & x961 ;
  assign n8080 = ~x782 & x963 ;
  assign n8081 = ~x230 & x967 ;
  assign n8082 = ~x230 & x969 ;
  assign n8083 = ~x782 & x970 ;
  assign n8084 = ~x230 & x971 ;
  assign n8085 = ~x782 & x972 ;
  assign n8086 = ~x230 & x974 ;
  assign n8087 = ~x782 & x975 ;
  assign n8088 = ~x230 & x977 ;
  assign n8089 = ~x782 & x978 ;
  assign n8090 = x824 & x1092 ;
  assign y0 = x668 ;
  assign y1 = x672 ;
  assign y2 = x664 ;
  assign y3 = x667 ;
  assign y4 = x676 ;
  assign y5 = x673 ;
  assign y6 = x675 ;
  assign y7 = x666 ;
  assign y8 = x679 ;
  assign y9 = x674 ;
  assign y10 = x663 ;
  assign y11 = x670 ;
  assign y12 = x677 ;
  assign y13 = x682 ;
  assign y14 = x671 ;
  assign y15 = x678 ;
  assign y16 = x718 ;
  assign y17 = x707 ;
  assign y18 = x708 ;
  assign y19 = x713 ;
  assign y20 = x711 ;
  assign y21 = x716 ;
  assign y22 = x733 ;
  assign y23 = x712 ;
  assign y24 = x689 ;
  assign y25 = x717 ;
  assign y26 = x692 ;
  assign y27 = x719 ;
  assign y28 = x722 ;
  assign y29 = x714 ;
  assign y30 = x720 ;
  assign y31 = x685 ;
  assign y32 = x837 ;
  assign y33 = x850 ;
  assign y34 = x872 ;
  assign y35 = x871 ;
  assign y36 = x881 ;
  assign y37 = x866 ;
  assign y38 = x876 ;
  assign y39 = x873 ;
  assign y40 = x874 ;
  assign y41 = x859 ;
  assign y42 = x855 ;
  assign y43 = x852 ;
  assign y44 = x870 ;
  assign y45 = x848 ;
  assign y46 = x865 ;
  assign y47 = x856 ;
  assign y48 = x853 ;
  assign y49 = x847 ;
  assign y50 = x857 ;
  assign y51 = x854 ;
  assign y52 = x858 ;
  assign y53 = x845 ;
  assign y54 = x838 ;
  assign y55 = x842 ;
  assign y56 = x843 ;
  assign y57 = x839 ;
  assign y58 = x844 ;
  assign y59 = x868 ;
  assign y60 = x851 ;
  assign y61 = x867 ;
  assign y62 = x880 ;
  assign y63 = x860 ;
  assign y64 = x1030 ;
  assign y65 = x1034 ;
  assign y66 = x1015 ;
  assign y67 = x1020 ;
  assign y68 = x1025 ;
  assign y69 = x1005 ;
  assign y70 = x996 ;
  assign y71 = x1012 ;
  assign y72 = x993 ;
  assign y73 = x1016 ;
  assign y74 = x1021 ;
  assign y75 = x1010 ;
  assign y76 = x1027 ;
  assign y77 = x1018 ;
  assign y78 = x1017 ;
  assign y79 = x1024 ;
  assign y80 = x1009 ;
  assign y81 = x1032 ;
  assign y82 = x1003 ;
  assign y83 = x997 ;
  assign y84 = x1013 ;
  assign y85 = x1011 ;
  assign y86 = x1008 ;
  assign y87 = x1019 ;
  assign y88 = x1031 ;
  assign y89 = x1022 ;
  assign y90 = x1000 ;
  assign y91 = x1023 ;
  assign y92 = x1002 ;
  assign y93 = x1026 ;
  assign y94 = x1006 ;
  assign y95 = x998 ;
  assign y96 = x31 ;
  assign y97 = x80 ;
  assign y98 = x893 ;
  assign y99 = x467 ;
  assign y100 = x78 ;
  assign y101 = x112 ;
  assign y102 = x13 ;
  assign y103 = x25 ;
  assign y104 = x226 ;
  assign y105 = x127 ;
  assign y106 = x822 ;
  assign y107 = x808 ;
  assign y108 = x227 ;
  assign y109 = x477 ;
  assign y110 = x834 ;
  assign y111 = x229 ;
  assign y112 = x12 ;
  assign y113 = x11 ;
  assign y114 = x10 ;
  assign y115 = x9 ;
  assign y116 = x8 ;
  assign y117 = x7 ;
  assign y118 = x6 ;
  assign y119 = x5 ;
  assign y120 = x4 ;
  assign y121 = x3 ;
  assign y122 = x0 ;
  assign y123 = x2 ;
  assign y124 = x1 ;
  assign y125 = x310 ;
  assign y126 = x302 ;
  assign y127 = x475 ;
  assign y128 = x474 ;
  assign y129 = x466 ;
  assign y130 = x473 ;
  assign y131 = x471 ;
  assign y132 = x472 ;
  assign y133 = x470 ;
  assign y134 = x469 ;
  assign y135 = x465 ;
  assign y136 = x1028 ;
  assign y137 = x1033 ;
  assign y138 = x995 ;
  assign y139 = x994 ;
  assign y140 = x28 ;
  assign y141 = x27 ;
  assign y142 = x26 ;
  assign y143 = x29 ;
  assign y144 = x15 ;
  assign y145 = x14 ;
  assign y146 = x21 ;
  assign y147 = x20 ;
  assign y148 = x19 ;
  assign y149 = x18 ;
  assign y150 = x17 ;
  assign y151 = x16 ;
  assign y152 = x1096 ;
  assign y153 = n1552 ;
  assign y154 = n1596 ;
  assign y155 = n1620 ;
  assign y156 = ~n1659 ;
  assign y157 = ~n1682 ;
  assign y158 = n1715 ;
  assign y159 = n1730 ;
  assign y160 = n1750 ;
  assign y161 = n1801 ;
  assign y162 = n1838 ;
  assign y163 = n1858 ;
  assign y164 = n1908 ;
  assign y165 = n1939 ;
  assign y166 = ~1'b0 ;
  assign y167 = n2033 ;
  assign y168 = x228 ;
  assign y169 = x22 ;
  assign y170 = ~x1090 ;
  assign y171 = ~n2099 ;
  assign y172 = ~n2106 ;
  assign y173 = ~n2110 ;
  assign y174 = ~n2113 ;
  assign y175 = ~n2116 ;
  assign y176 = ~n2119 ;
  assign y177 = ~n2122 ;
  assign y178 = ~n2125 ;
  assign y179 = x1089 ;
  assign y180 = x23 ;
  assign y181 = n2033 ;
  assign y182 = n2140 ;
  assign y183 = n2168 ;
  assign y184 = ~n2171 ;
  assign y185 = ~n2173 ;
  assign y186 = ~n2175 ;
  assign y187 = ~n2177 ;
  assign y188 = x37 ;
  assign y189 = n2534 ;
  assign y190 = n2574 ;
  assign y191 = n2711 ;
  assign y192 = n2790 ;
  assign y193 = n2818 ;
  assign y194 = n2822 ;
  assign y195 = n2139 ;
  assign y196 = n2834 ;
  assign y197 = n2849 ;
  assign y198 = n2852 ;
  assign y199 = n2894 ;
  assign y200 = n2915 ;
  assign y201 = n2935 ;
  assign y202 = n2946 ;
  assign y203 = n2948 ;
  assign y204 = n2952 ;
  assign y205 = n2957 ;
  assign y206 = n2959 ;
  assign y207 = n2965 ;
  assign y208 = n2981 ;
  assign y209 = n2983 ;
  assign y210 = n2993 ;
  assign y211 = n3000 ;
  assign y212 = n3005 ;
  assign y213 = n3013 ;
  assign y214 = n3017 ;
  assign y215 = n3025 ;
  assign y216 = n3027 ;
  assign y217 = n3037 ;
  assign y218 = n3042 ;
  assign y219 = n3044 ;
  assign y220 = n3047 ;
  assign y221 = n3052 ;
  assign y222 = n3055 ;
  assign y223 = n3056 ;
  assign y224 = n3064 ;
  assign y225 = n3068 ;
  assign y226 = n3071 ;
  assign y227 = n3074 ;
  assign y228 = n3087 ;
  assign y229 = n3095 ;
  assign y230 = n3103 ;
  assign y231 = n3106 ;
  assign y232 = n3119 ;
  assign y233 = n3122 ;
  assign y234 = n3127 ;
  assign y235 = n3129 ;
  assign y236 = n3131 ;
  assign y237 = n3202 ;
  assign y238 = n3204 ;
  assign y239 = n3208 ;
  assign y240 = n3210 ;
  assign y241 = n3213 ;
  assign y242 = n3216 ;
  assign y243 = n3219 ;
  assign y244 = n3221 ;
  assign y245 = n3222 ;
  assign y246 = n3226 ;
  assign y247 = n3231 ;
  assign y248 = n3234 ;
  assign y249 = n3244 ;
  assign y250 = n3248 ;
  assign y251 = n3251 ;
  assign y252 = n3255 ;
  assign y253 = n3265 ;
  assign y254 = n3270 ;
  assign y255 = n3275 ;
  assign y256 = n3279 ;
  assign y257 = n3289 ;
  assign y258 = n3293 ;
  assign y259 = n3307 ;
  assign y260 = n3308 ;
  assign y261 = n3311 ;
  assign y262 = n3317 ;
  assign y263 = x117 ;
  assign y264 = n3320 ;
  assign y265 = n3322 ;
  assign y266 = n3329 ;
  assign y267 = n3331 ;
  assign y268 = n3334 ;
  assign y269 = n3337 ;
  assign y270 = ~n3338 ;
  assign y271 = n3343 ;
  assign y272 = n3346 ;
  assign y273 = n3349 ;
  assign y274 = n3354 ;
  assign y275 = n2167 ;
  assign y276 = n3426 ;
  assign y277 = n3443 ;
  assign y278 = n3451 ;
  assign y279 = n3500 ;
  assign y280 = n2529 ;
  assign y281 = ~n3521 ;
  assign y282 = n3555 ;
  assign y283 = n3592 ;
  assign y284 = n3603 ;
  assign y285 = x131 ;
  assign y286 = n3610 ;
  assign y287 = n3629 ;
  assign y288 = n3442 ;
  assign y289 = n3659 ;
  assign y290 = n3672 ;
  assign y291 = n3692 ;
  assign y292 = n3713 ;
  assign y293 = n3726 ;
  assign y294 = n3734 ;
  assign y295 = n3741 ;
  assign y296 = n3746 ;
  assign y297 = ~n3829 ;
  assign y298 = ~n3834 ;
  assign y299 = n3839 ;
  assign y300 = ~n3844 ;
  assign y301 = n3849 ;
  assign y302 = ~n3854 ;
  assign y303 = n3859 ;
  assign y304 = ~n3864 ;
  assign y305 = ~n3869 ;
  assign y306 = ~n3874 ;
  assign y307 = ~n3879 ;
  assign y308 = ~n3884 ;
  assign y309 = n3889 ;
  assign y310 = ~n3894 ;
  assign y311 = ~n3899 ;
  assign y312 = ~n3904 ;
  assign y313 = ~n3909 ;
  assign y314 = ~n3914 ;
  assign y315 = ~n3919 ;
  assign y316 = ~n3924 ;
  assign y317 = ~n3929 ;
  assign y318 = n3934 ;
  assign y319 = ~n3939 ;
  assign y320 = ~n3944 ;
  assign y321 = ~n3949 ;
  assign y322 = ~n3954 ;
  assign y323 = n3959 ;
  assign y324 = ~n3964 ;
  assign y325 = ~n3969 ;
  assign y326 = ~n3974 ;
  assign y327 = ~n3979 ;
  assign y328 = ~n3984 ;
  assign y329 = ~n3989 ;
  assign y330 = ~n3994 ;
  assign y331 = n3999 ;
  assign y332 = ~n4004 ;
  assign y333 = ~n4009 ;
  assign y334 = ~n4014 ;
  assign y335 = ~n4019 ;
  assign y336 = ~n4024 ;
  assign y337 = ~n4029 ;
  assign y338 = ~n4034 ;
  assign y339 = ~n4039 ;
  assign y340 = ~n4044 ;
  assign y341 = ~n4049 ;
  assign y342 = ~n4054 ;
  assign y343 = ~n4059 ;
  assign y344 = ~n4064 ;
  assign y345 = ~n4069 ;
  assign y346 = n4074 ;
  assign y347 = ~n4079 ;
  assign y348 = ~n4084 ;
  assign y349 = ~n4089 ;
  assign y350 = ~n4094 ;
  assign y351 = ~n4099 ;
  assign y352 = n4105 ;
  assign y353 = n4111 ;
  assign y354 = ~n4116 ;
  assign y355 = n4121 ;
  assign y356 = n4126 ;
  assign y357 = n4131 ;
  assign y358 = ~n4148 ;
  assign y359 = ~n4157 ;
  assign y360 = ~n4166 ;
  assign y361 = ~n4171 ;
  assign y362 = ~n4176 ;
  assign y363 = ~n4185 ;
  assign y364 = ~n4190 ;
  assign y365 = ~n4195 ;
  assign y366 = ~n4200 ;
  assign y367 = n4205 ;
  assign y368 = n4210 ;
  assign y369 = ~n4215 ;
  assign y370 = ~n4220 ;
  assign y371 = ~n4225 ;
  assign y372 = n4230 ;
  assign y373 = n4235 ;
  assign y374 = ~n4240 ;
  assign y375 = ~n4245 ;
  assign y376 = n4250 ;
  assign y377 = ~n4255 ;
  assign y378 = n4260 ;
  assign y379 = n4265 ;
  assign y380 = n4270 ;
  assign y381 = n4275 ;
  assign y382 = n4291 ;
  assign y383 = n4298 ;
  assign y384 = ~n4305 ;
  assign y385 = n4315 ;
  assign y386 = x232 ;
  assign y387 = n3793 ;
  assign y388 = x236 ;
  assign y389 = n4319 ;
  assign y390 = ~n4391 ;
  assign y391 = n4414 ;
  assign y392 = n4435 ;
  assign y393 = n4295 ;
  assign y394 = ~n4465 ;
  assign y395 = n4487 ;
  assign y396 = n4499 ;
  assign y397 = n4514 ;
  assign y398 = n4525 ;
  assign y399 = n4538 ;
  assign y400 = ~n4566 ;
  assign y401 = n4572 ;
  assign y402 = n4582 ;
  assign y403 = n4592 ;
  assign y404 = n4597 ;
  assign y405 = n4607 ;
  assign y406 = n4612 ;
  assign y407 = n4616 ;
  assign y408 = n4625 ;
  assign y409 = n4630 ;
  assign y410 = n4637 ;
  assign y411 = n4647 ;
  assign y412 = n4653 ;
  assign y413 = n4659 ;
  assign y414 = n4665 ;
  assign y415 = n4671 ;
  assign y416 = n4677 ;
  assign y417 = n4683 ;
  assign y418 = n4689 ;
  assign y419 = ~n4697 ;
  assign y420 = ~n4707 ;
  assign y421 = ~n4716 ;
  assign y422 = ~n4725 ;
  assign y423 = n4734 ;
  assign y424 = n4745 ;
  assign y425 = n4752 ;
  assign y426 = ~n4761 ;
  assign y427 = ~n4770 ;
  assign y428 = n4777 ;
  assign y429 = n4784 ;
  assign y430 = n4792 ;
  assign y431 = ~n4801 ;
  assign y432 = n4807 ;
  assign y433 = n4813 ;
  assign y434 = ~n4822 ;
  assign y435 = n4831 ;
  assign y436 = n4840 ;
  assign y437 = ~n4849 ;
  assign y438 = ~n4857 ;
  assign y439 = ~n4866 ;
  assign y440 = n4875 ;
  assign y441 = ~n4879 ;
  assign y442 = n4891 ;
  assign y443 = n4896 ;
  assign y444 = ~n4898 ;
  assign y445 = n4904 ;
  assign y446 = n4908 ;
  assign y447 = n4911 ;
  assign y448 = n4914 ;
  assign y449 = n4917 ;
  assign y450 = n4920 ;
  assign y451 = n4923 ;
  assign y452 = n4926 ;
  assign y453 = n4929 ;
  assign y454 = n4932 ;
  assign y455 = n4935 ;
  assign y456 = n4939 ;
  assign y457 = n4945 ;
  assign y458 = ~n4948 ;
  assign y459 = ~n4955 ;
  assign y460 = n4958 ;
  assign y461 = n4961 ;
  assign y462 = n4964 ;
  assign y463 = n4967 ;
  assign y464 = n4970 ;
  assign y465 = n4973 ;
  assign y466 = n4976 ;
  assign y467 = ~n4982 ;
  assign y468 = ~n4987 ;
  assign y469 = n4989 ;
  assign y470 = n4995 ;
  assign y471 = ~n4997 ;
  assign y472 = n5001 ;
  assign y473 = n5004 ;
  assign y474 = n5008 ;
  assign y475 = n5012 ;
  assign y476 = n5015 ;
  assign y477 = n5018 ;
  assign y478 = n5021 ;
  assign y479 = n5024 ;
  assign y480 = n5027 ;
  assign y481 = n5030 ;
  assign y482 = n5033 ;
  assign y483 = n5036 ;
  assign y484 = n5039 ;
  assign y485 = n5042 ;
  assign y486 = n5045 ;
  assign y487 = n5048 ;
  assign y488 = n5050 ;
  assign y489 = n5056 ;
  assign y490 = n5059 ;
  assign y491 = n5062 ;
  assign y492 = n5065 ;
  assign y493 = n5068 ;
  assign y494 = n5071 ;
  assign y495 = n5074 ;
  assign y496 = n5077 ;
  assign y497 = ~n5080 ;
  assign y498 = n5082 ;
  assign y499 = n5085 ;
  assign y500 = n5088 ;
  assign y501 = n5091 ;
  assign y502 = n5094 ;
  assign y503 = n5097 ;
  assign y504 = n5100 ;
  assign y505 = n5103 ;
  assign y506 = n5106 ;
  assign y507 = n5109 ;
  assign y508 = n5112 ;
  assign y509 = n5115 ;
  assign y510 = n5118 ;
  assign y511 = n5121 ;
  assign y512 = n5124 ;
  assign y513 = n5127 ;
  assign y514 = n5130 ;
  assign y515 = n5133 ;
  assign y516 = n5136 ;
  assign y517 = n5139 ;
  assign y518 = n5142 ;
  assign y519 = n5145 ;
  assign y520 = n5148 ;
  assign y521 = n5151 ;
  assign y522 = n5154 ;
  assign y523 = n5157 ;
  assign y524 = n5160 ;
  assign y525 = n5163 ;
  assign y526 = n5166 ;
  assign y527 = n5169 ;
  assign y528 = n5172 ;
  assign y529 = n5175 ;
  assign y530 = n5178 ;
  assign y531 = n5181 ;
  assign y532 = n5184 ;
  assign y533 = n5187 ;
  assign y534 = n5190 ;
  assign y535 = n5193 ;
  assign y536 = n5196 ;
  assign y537 = n5199 ;
  assign y538 = n5202 ;
  assign y539 = n5205 ;
  assign y540 = n5208 ;
  assign y541 = n5211 ;
  assign y542 = n5214 ;
  assign y543 = n5217 ;
  assign y544 = n5220 ;
  assign y545 = n5223 ;
  assign y546 = n5226 ;
  assign y547 = n5229 ;
  assign y548 = n5232 ;
  assign y549 = n5235 ;
  assign y550 = n5238 ;
  assign y551 = n5241 ;
  assign y552 = n5244 ;
  assign y553 = n5247 ;
  assign y554 = n5250 ;
  assign y555 = n5253 ;
  assign y556 = n5256 ;
  assign y557 = n5259 ;
  assign y558 = n5262 ;
  assign y559 = n5265 ;
  assign y560 = n5268 ;
  assign y561 = n5271 ;
  assign y562 = n5274 ;
  assign y563 = n5277 ;
  assign y564 = n5280 ;
  assign y565 = n5283 ;
  assign y566 = n5286 ;
  assign y567 = n5289 ;
  assign y568 = n5292 ;
  assign y569 = n5295 ;
  assign y570 = n5298 ;
  assign y571 = n5302 ;
  assign y572 = n5305 ;
  assign y573 = n5308 ;
  assign y574 = n5311 ;
  assign y575 = n5314 ;
  assign y576 = n5317 ;
  assign y577 = n5320 ;
  assign y578 = n5323 ;
  assign y579 = n5326 ;
  assign y580 = n5329 ;
  assign y581 = n5332 ;
  assign y582 = n5335 ;
  assign y583 = n5338 ;
  assign y584 = n5341 ;
  assign y585 = n5344 ;
  assign y586 = n5347 ;
  assign y587 = n5350 ;
  assign y588 = n5353 ;
  assign y589 = n5356 ;
  assign y590 = n5359 ;
  assign y591 = n5362 ;
  assign y592 = n5365 ;
  assign y593 = n5368 ;
  assign y594 = n5371 ;
  assign y595 = n5374 ;
  assign y596 = n5377 ;
  assign y597 = n5380 ;
  assign y598 = n5383 ;
  assign y599 = n5386 ;
  assign y600 = n5389 ;
  assign y601 = n5392 ;
  assign y602 = n5395 ;
  assign y603 = n5398 ;
  assign y604 = n5401 ;
  assign y605 = n5404 ;
  assign y606 = n5407 ;
  assign y607 = n5410 ;
  assign y608 = n5413 ;
  assign y609 = n5416 ;
  assign y610 = n5419 ;
  assign y611 = n5422 ;
  assign y612 = n5425 ;
  assign y613 = n5428 ;
  assign y614 = n5449 ;
  assign y615 = n5452 ;
  assign y616 = n5455 ;
  assign y617 = n5458 ;
  assign y618 = n5461 ;
  assign y619 = n5464 ;
  assign y620 = n5467 ;
  assign y621 = n5470 ;
  assign y622 = n5475 ;
  assign y623 = n5480 ;
  assign y624 = n5486 ;
  assign y625 = n5489 ;
  assign y626 = n5494 ;
  assign y627 = n5499 ;
  assign y628 = n5504 ;
  assign y629 = n5509 ;
  assign y630 = n5514 ;
  assign y631 = n5519 ;
  assign y632 = n5524 ;
  assign y633 = n5527 ;
  assign y634 = ~n4993 ;
  assign y635 = n5528 ;
  assign y636 = x583 ;
  assign y637 = n4880 ;
  assign y638 = n5531 ;
  assign y639 = n5534 ;
  assign y640 = n5537 ;
  assign y641 = n5540 ;
  assign y642 = n5543 ;
  assign y643 = n5546 ;
  assign y644 = n5549 ;
  assign y645 = ~n5552 ;
  assign y646 = n5555 ;
  assign y647 = n5558 ;
  assign y648 = n5561 ;
  assign y649 = n5564 ;
  assign y650 = n5567 ;
  assign y651 = ~n5570 ;
  assign y652 = n5573 ;
  assign y653 = n5576 ;
  assign y654 = ~n5579 ;
  assign y655 = n5582 ;
  assign y656 = n5585 ;
  assign y657 = n5588 ;
  assign y658 = n5591 ;
  assign y659 = n5594 ;
  assign y660 = n5597 ;
  assign y661 = n5600 ;
  assign y662 = n5603 ;
  assign y663 = n5606 ;
  assign y664 = n5609 ;
  assign y665 = n5612 ;
  assign y666 = n5615 ;
  assign y667 = n5618 ;
  assign y668 = n5621 ;
  assign y669 = n5624 ;
  assign y670 = n5627 ;
  assign y671 = n5630 ;
  assign y672 = n5633 ;
  assign y673 = n5636 ;
  assign y674 = n5639 ;
  assign y675 = n5642 ;
  assign y676 = ~n5645 ;
  assign y677 = n5648 ;
  assign y678 = n5651 ;
  assign y679 = n5654 ;
  assign y680 = n5657 ;
  assign y681 = ~n5660 ;
  assign y682 = n5663 ;
  assign y683 = n5666 ;
  assign y684 = n5669 ;
  assign y685 = n5672 ;
  assign y686 = n5675 ;
  assign y687 = n5678 ;
  assign y688 = n5681 ;
  assign y689 = n5684 ;
  assign y690 = n5687 ;
  assign y691 = ~n5690 ;
  assign y692 = n5693 ;
  assign y693 = n5696 ;
  assign y694 = n5699 ;
  assign y695 = n5702 ;
  assign y696 = n5705 ;
  assign y697 = n5708 ;
  assign y698 = n5711 ;
  assign y699 = n5714 ;
  assign y700 = n5717 ;
  assign y701 = n5720 ;
  assign y702 = n5723 ;
  assign y703 = n5726 ;
  assign y704 = n5729 ;
  assign y705 = n5732 ;
  assign y706 = n5735 ;
  assign y707 = ~n5738 ;
  assign y708 = n5741 ;
  assign y709 = n5744 ;
  assign y710 = n5747 ;
  assign y711 = n5750 ;
  assign y712 = n5753 ;
  assign y713 = n5756 ;
  assign y714 = n5759 ;
  assign y715 = n5762 ;
  assign y716 = n5765 ;
  assign y717 = n5768 ;
  assign y718 = n5771 ;
  assign y719 = n5774 ;
  assign y720 = n5777 ;
  assign y721 = n5780 ;
  assign y722 = n5783 ;
  assign y723 = n5786 ;
  assign y724 = n5792 ;
  assign y725 = n5795 ;
  assign y726 = ~n5798 ;
  assign y727 = n5801 ;
  assign y728 = n5804 ;
  assign y729 = n5807 ;
  assign y730 = n5810 ;
  assign y731 = n5813 ;
  assign y732 = n5816 ;
  assign y733 = n5819 ;
  assign y734 = n5822 ;
  assign y735 = n5825 ;
  assign y736 = n5828 ;
  assign y737 = n5831 ;
  assign y738 = n5834 ;
  assign y739 = n5837 ;
  assign y740 = n1960 ;
  assign y741 = n5840 ;
  assign y742 = n5843 ;
  assign y743 = n5846 ;
  assign y744 = n5849 ;
  assign y745 = n5854 ;
  assign y746 = n5871 ;
  assign y747 = ~n5874 ;
  assign y748 = n5877 ;
  assign y749 = n5880 ;
  assign y750 = n6221 ;
  assign y751 = n6226 ;
  assign y752 = n6231 ;
  assign y753 = n6237 ;
  assign y754 = n6240 ;
  assign y755 = n6246 ;
  assign y756 = n6249 ;
  assign y757 = n6251 ;
  assign y758 = n6254 ;
  assign y759 = n6257 ;
  assign y760 = n6268 ;
  assign y761 = n6276 ;
  assign y762 = ~n6279 ;
  assign y763 = n6284 ;
  assign y764 = n6287 ;
  assign y765 = n6290 ;
  assign y766 = n6293 ;
  assign y767 = n6296 ;
  assign y768 = n6299 ;
  assign y769 = n6302 ;
  assign y770 = n6305 ;
  assign y771 = n6310 ;
  assign y772 = ~n6315 ;
  assign y773 = n6320 ;
  assign y774 = n6325 ;
  assign y775 = n6328 ;
  assign y776 = n6331 ;
  assign y777 = n6334 ;
  assign y778 = n6337 ;
  assign y779 = n6340 ;
  assign y780 = n6343 ;
  assign y781 = n6350 ;
  assign y782 = n6358 ;
  assign y783 = n6361 ;
  assign y784 = n6364 ;
  assign y785 = n6367 ;
  assign y786 = n6370 ;
  assign y787 = n6373 ;
  assign y788 = ~n6376 ;
  assign y789 = ~n6379 ;
  assign y790 = n6382 ;
  assign y791 = n6385 ;
  assign y792 = ~n6388 ;
  assign y793 = n6391 ;
  assign y794 = n6394 ;
  assign y795 = n6397 ;
  assign y796 = n6400 ;
  assign y797 = n6403 ;
  assign y798 = n6406 ;
  assign y799 = n6409 ;
  assign y800 = n6412 ;
  assign y801 = n6415 ;
  assign y802 = n6418 ;
  assign y803 = ~n6421 ;
  assign y804 = n6424 ;
  assign y805 = n6427 ;
  assign y806 = ~n6430 ;
  assign y807 = ~n6433 ;
  assign y808 = n6436 ;
  assign y809 = n6439 ;
  assign y810 = n6442 ;
  assign y811 = ~n6445 ;
  assign y812 = ~n6448 ;
  assign y813 = n6451 ;
  assign y814 = ~n6454 ;
  assign y815 = n6457 ;
  assign y816 = ~n6469 ;
  assign y817 = n6472 ;
  assign y818 = n6475 ;
  assign y819 = n6478 ;
  assign y820 = n6512 ;
  assign y821 = n6540 ;
  assign y822 = n6543 ;
  assign y823 = n6571 ;
  assign y824 = n6602 ;
  assign y825 = n6627 ;
  assign y826 = ~n6630 ;
  assign y827 = n6652 ;
  assign y828 = n6674 ;
  assign y829 = n6700 ;
  assign y830 = n6728 ;
  assign y831 = n6754 ;
  assign y832 = n6780 ;
  assign y833 = n6805 ;
  assign y834 = n6827 ;
  assign y835 = n6849 ;
  assign y836 = n6875 ;
  assign y837 = n6878 ;
  assign y838 = n6881 ;
  assign y839 = n6903 ;
  assign y840 = n1434 ;
  assign y841 = ~n6907 ;
  assign y842 = n6930 ;
  assign y843 = ~n6933 ;
  assign y844 = n6936 ;
  assign y845 = ~n6939 ;
  assign y846 = n6963 ;
  assign y847 = n6966 ;
  assign y848 = n6969 ;
  assign y849 = n6991 ;
  assign y850 = ~n6994 ;
  assign y851 = ~n6997 ;
  assign y852 = ~n7000 ;
  assign y853 = n7003 ;
  assign y854 = ~n7006 ;
  assign y855 = ~n7009 ;
  assign y856 = n7012 ;
  assign y857 = n7015 ;
  assign y858 = ~n7018 ;
  assign y859 = ~n7021 ;
  assign y860 = n7024 ;
  assign y861 = ~n7027 ;
  assign y862 = n7030 ;
  assign y863 = n7033 ;
  assign y864 = n7057 ;
  assign y865 = n7081 ;
  assign y866 = ~n7084 ;
  assign y867 = n7087 ;
  assign y868 = n7111 ;
  assign y869 = n7135 ;
  assign y870 = n7158 ;
  assign y871 = n7181 ;
  assign y872 = n7184 ;
  assign y873 = n7207 ;
  assign y874 = n7231 ;
  assign y875 = n7255 ;
  assign y876 = n7278 ;
  assign y877 = n7301 ;
  assign y878 = n7337 ;
  assign y879 = n7360 ;
  assign y880 = ~n7363 ;
  assign y881 = ~n7366 ;
  assign y882 = ~n7369 ;
  assign y883 = n7372 ;
  assign y884 = n7375 ;
  assign y885 = ~n7378 ;
  assign y886 = n7381 ;
  assign y887 = n7384 ;
  assign y888 = n7387 ;
  assign y889 = ~n7390 ;
  assign y890 = n7414 ;
  assign y891 = ~n7417 ;
  assign y892 = n7420 ;
  assign y893 = n7423 ;
  assign y894 = ~n7426 ;
  assign y895 = ~n7429 ;
  assign y896 = n7434 ;
  assign y897 = n6264 ;
  assign y898 = ~n7437 ;
  assign y899 = ~n7440 ;
  assign y900 = n7443 ;
  assign y901 = ~n7446 ;
  assign y902 = ~n7449 ;
  assign y903 = n7452 ;
  assign y904 = n7454 ;
  assign y905 = n7457 ;
  assign y906 = n7460 ;
  assign y907 = ~n7463 ;
  assign y908 = ~n7466 ;
  assign y909 = ~n7469 ;
  assign y910 = ~n7472 ;
  assign y911 = ~n7475 ;
  assign y912 = ~n7478 ;
  assign y913 = ~n7481 ;
  assign y914 = ~n7484 ;
  assign y915 = n7487 ;
  assign y916 = n7490 ;
  assign y917 = ~n7493 ;
  assign y918 = ~n7496 ;
  assign y919 = ~n7499 ;
  assign y920 = n7502 ;
  assign y921 = n7505 ;
  assign y922 = ~n7516 ;
  assign y923 = n7519 ;
  assign y924 = ~n7522 ;
  assign y925 = ~n7525 ;
  assign y926 = n7527 ;
  assign y927 = ~n7530 ;
  assign y928 = n7534 ;
  assign y929 = n7537 ;
  assign y930 = n7539 ;
  assign y931 = ~n7542 ;
  assign y932 = n7549 ;
  assign y933 = ~n7552 ;
  assign y934 = ~n7555 ;
  assign y935 = n7563 ;
  assign y936 = ~n7564 ;
  assign y937 = ~n7565 ;
  assign y938 = n7568 ;
  assign y939 = ~n7570 ;
  assign y940 = n7573 ;
  assign y941 = n7576 ;
  assign y942 = n7579 ;
  assign y943 = ~n7581 ;
  assign y944 = n7584 ;
  assign y945 = n7587 ;
  assign y946 = n7590 ;
  assign y947 = n7593 ;
  assign y948 = n7596 ;
  assign y949 = n7599 ;
  assign y950 = ~n1995 ;
  assign y951 = n7604 ;
  assign y952 = n7607 ;
  assign y953 = ~n7617 ;
  assign y954 = n6355 ;
  assign y955 = n7620 ;
  assign y956 = ~n7623 ;
  assign y957 = n7626 ;
  assign y958 = n7629 ;
  assign y959 = n6468 ;
  assign y960 = ~n7632 ;
  assign y961 = n7635 ;
  assign y962 = ~n7638 ;
  assign y963 = n7531 ;
  assign y964 = n7641 ;
  assign y965 = n7644 ;
  assign y966 = ~n7647 ;
  assign y967 = n7650 ;
  assign y968 = n7653 ;
  assign y969 = ~n7656 ;
  assign y970 = n7659 ;
  assign y971 = ~n7662 ;
  assign y972 = n7665 ;
  assign y973 = n7668 ;
  assign y974 = ~n7671 ;
  assign y975 = n7672 ;
  assign y976 = ~n7675 ;
  assign y977 = ~n7678 ;
  assign y978 = ~n7335 ;
  assign y979 = ~n7679 ;
  assign y980 = n6904 ;
  assign y981 = n7682 ;
  assign y982 = n7696 ;
  assign y983 = n7712 ;
  assign y984 = n7725 ;
  assign y985 = n7738 ;
  assign y986 = n7741 ;
  assign y987 = ~n7744 ;
  assign y988 = n7431 ;
  assign y989 = n7746 ;
  assign y990 = n7748 ;
  assign y991 = n7749 ;
  assign y992 = ~n7751 ;
  assign y993 = n7754 ;
  assign y994 = n7757 ;
  assign y995 = n7760 ;
  assign y996 = n7763 ;
  assign y997 = ~n2628 ;
  assign y998 = n7766 ;
  assign y999 = n7769 ;
  assign y1000 = n7772 ;
  assign y1001 = n7775 ;
  assign y1002 = n7778 ;
  assign y1003 = n7781 ;
  assign y1004 = n7784 ;
  assign y1005 = n7787 ;
  assign y1006 = n7790 ;
  assign y1007 = n7793 ;
  assign y1008 = n7796 ;
  assign y1009 = n7799 ;
  assign y1010 = n7802 ;
  assign y1011 = n7805 ;
  assign y1012 = n7808 ;
  assign y1013 = n7811 ;
  assign y1014 = n7814 ;
  assign y1015 = n7817 ;
  assign y1016 = n7820 ;
  assign y1017 = n7823 ;
  assign y1018 = n7826 ;
  assign y1019 = n7829 ;
  assign y1020 = n7832 ;
  assign y1021 = n7835 ;
  assign y1022 = n7838 ;
  assign y1023 = n7841 ;
  assign y1024 = n7844 ;
  assign y1025 = n7847 ;
  assign y1026 = n7850 ;
  assign y1027 = n7853 ;
  assign y1028 = n7856 ;
  assign y1029 = n7859 ;
  assign y1030 = n7862 ;
  assign y1031 = n7865 ;
  assign y1032 = n7868 ;
  assign y1033 = n7871 ;
  assign y1034 = n7874 ;
  assign y1035 = n7877 ;
  assign y1036 = n7880 ;
  assign y1037 = n7883 ;
  assign y1038 = n1208 ;
  assign y1039 = n7886 ;
  assign y1040 = n7889 ;
  assign y1041 = n7892 ;
  assign y1042 = n7895 ;
  assign y1043 = n7898 ;
  assign y1044 = n7901 ;
  assign y1045 = n7904 ;
  assign y1046 = n7907 ;
  assign y1047 = n7910 ;
  assign y1048 = n7913 ;
  assign y1049 = n7914 ;
  assign y1050 = n7917 ;
  assign y1051 = n7920 ;
  assign y1052 = n7923 ;
  assign y1053 = x67 ;
  assign y1054 = n7926 ;
  assign y1055 = n7929 ;
  assign y1056 = n7932 ;
  assign y1057 = n1950 ;
  assign y1058 = n7935 ;
  assign y1059 = n7938 ;
  assign y1060 = n7941 ;
  assign y1061 = n7944 ;
  assign y1062 = n7947 ;
  assign y1063 = n7954 ;
  assign y1064 = n7957 ;
  assign y1065 = n7960 ;
  assign y1066 = n7963 ;
  assign y1067 = n7966 ;
  assign y1068 = n7969 ;
  assign y1069 = n7972 ;
  assign y1070 = ~n7975 ;
  assign y1071 = n7978 ;
  assign y1072 = n7981 ;
  assign y1073 = n7984 ;
  assign y1074 = n7987 ;
  assign y1075 = n7990 ;
  assign y1076 = n7993 ;
  assign y1077 = n7996 ;
  assign y1078 = n7999 ;
  assign y1079 = n8002 ;
  assign y1080 = n8004 ;
  assign y1081 = n8007 ;
  assign y1082 = n8010 ;
  assign y1083 = n8013 ;
  assign y1084 = n8016 ;
  assign y1085 = n8019 ;
  assign y1086 = n8022 ;
  assign y1087 = n8025 ;
  assign y1088 = n8028 ;
  assign y1089 = n8031 ;
  assign y1090 = n8034 ;
  assign y1091 = n8037 ;
  assign y1092 = n8040 ;
  assign y1093 = n8043 ;
  assign y1094 = n8046 ;
  assign y1095 = n8049 ;
  assign y1096 = n8052 ;
  assign y1097 = n8055 ;
  assign y1098 = n8058 ;
  assign y1099 = n8061 ;
  assign y1100 = n8064 ;
  assign y1101 = n8065 ;
  assign y1102 = n5787 ;
  assign y1103 = n8070 ;
  assign y1104 = n8073 ;
  assign y1105 = ~n8075 ;
  assign y1106 = n1433 ;
  assign y1107 = n1428 ;
  assign y1108 = x1134 ;
  assign y1109 = x964 ;
  assign y1110 = ~x954 ;
  assign y1111 = x965 ;
  assign y1112 = n8077 ;
  assign y1113 = x991 ;
  assign y1114 = x985 ;
  assign y1115 = n8078 ;
  assign y1116 = n8079 ;
  assign y1117 = x1014 ;
  assign y1118 = n8080 ;
  assign y1119 = x1029 ;
  assign y1120 = x1004 ;
  assign y1121 = x1007 ;
  assign y1122 = n8081 ;
  assign y1123 = x1135 ;
  assign y1124 = n8082 ;
  assign y1125 = n8083 ;
  assign y1126 = n8084 ;
  assign y1127 = n8085 ;
  assign y1128 = n8086 ;
  assign y1129 = n8087 ;
  assign y1130 = ~x278 ;
  assign y1131 = n8088 ;
  assign y1132 = n8089 ;
  assign y1133 = ~n7951 ;
  assign y1134 = x1064 ;
  assign y1135 = n8090 ;
  assign y1136 = x299 ;
  assign y1137 = n7949 ;
  assign y1138 = x1075 ;
  assign y1139 = x1052 ;
  assign y1140 = x771 ;
  assign y1141 = x765 ;
  assign y1142 = x605 ;
  assign y1143 = x601 ;
  assign y1144 = x278 ;
  assign y1145 = x279 ;
  assign y1146 = ~x915 ;
  assign y1147 = ~x825 ;
  assign y1148 = ~x826 ;
  assign y1149 = ~x913 ;
  assign y1150 = ~x894 ;
  assign y1151 = ~x905 ;
  assign y1152 = x1095 ;
  assign y1153 = ~x890 ;
  assign y1154 = x1094 ;
  assign y1155 = ~x906 ;
  assign y1156 = ~x896 ;
  assign y1157 = ~x909 ;
  assign y1158 = ~x911 ;
  assign y1159 = ~x908 ;
  assign y1160 = ~x891 ;
  assign y1161 = ~x902 ;
  assign y1162 = ~x903 ;
  assign y1163 = ~x883 ;
  assign y1164 = ~x888 ;
  assign y1165 = ~x919 ;
  assign y1166 = ~x886 ;
  assign y1167 = ~x912 ;
  assign y1168 = ~x895 ;
  assign y1169 = ~x916 ;
  assign y1170 = ~x889 ;
  assign y1171 = ~x900 ;
  assign y1172 = ~x885 ;
  assign y1173 = ~x904 ;
  assign y1174 = ~x899 ;
  assign y1175 = ~x918 ;
  assign y1176 = ~x898 ;
  assign y1177 = ~x917 ;
  assign y1178 = ~x827 ;
  assign y1179 = ~x887 ;
  assign y1180 = ~x884 ;
  assign y1181 = ~x910 ;
  assign y1182 = ~x828 ;
  assign y1183 = ~x892 ;
  assign y1184 = x1187 ;
  assign y1185 = x1172 ;
  assign y1186 = x1170 ;
  assign y1187 = x1138 ;
  assign y1188 = x1177 ;
  assign y1189 = x1178 ;
  assign y1190 = x863 ;
  assign y1191 = x1203 ;
  assign y1192 = x1185 ;
  assign y1193 = x1171 ;
  assign y1194 = x1192 ;
  assign y1195 = x1137 ;
  assign y1196 = x1186 ;
  assign y1197 = x1165 ;
  assign y1198 = x1164 ;
  assign y1199 = x1098 ;
  assign y1200 = x1183 ;
  assign y1201 = x230 ;
  assign y1202 = x1169 ;
  assign y1203 = x1136 ;
  assign y1204 = x1181 ;
  assign y1205 = x849 ;
  assign y1206 = x1193 ;
  assign y1207 = x1182 ;
  assign y1208 = x1168 ;
  assign y1209 = x1175 ;
  assign y1210 = x1191 ;
  assign y1211 = x1099 ;
  assign y1212 = x1174 ;
  assign y1213 = x1179 ;
  assign y1214 = x1202 ;
  assign y1215 = x1176 ;
  assign y1216 = x1173 ;
  assign y1217 = x1201 ;
  assign y1218 = x1167 ;
  assign y1219 = x840 ;
  assign y1220 = x1189 ;
  assign y1221 = x1195 ;
  assign y1222 = x864 ;
  assign y1223 = x1190 ;
  assign y1224 = x1188 ;
  assign y1225 = x1180 ;
  assign y1226 = x1194 ;
  assign y1227 = x1097 ;
  assign y1228 = x1166 ;
  assign y1229 = x1200 ;
  assign y1230 = x1184 ;
endmodule
