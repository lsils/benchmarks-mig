module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 ;
  assign n129 = x0 & x64 ;
  assign n130 = x2 & n129 ;
  assign n131 = ~x64 & x65 ;
  assign n132 = x64 & x65 ;
  assign n133 = ( x64 & n131 ) | ( x64 & ~n132 ) | ( n131 & ~n132 ) ;
  assign n134 = ~x1 & x2 ;
  assign n135 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n136 = ( ~x2 & n134 ) | ( ~x2 & n135 ) | ( n134 & n135 ) ;
  assign n137 = n133 & n136 ;
  assign n138 = ~x0 & x1 ;
  assign n139 = x64 & n138 ;
  assign n140 = x65 | n139 ;
  assign n141 = x0 & ~n136 ;
  assign n142 = ( n139 & n140 ) | ( n139 & n141 ) | ( n140 & n141 ) ;
  assign n143 = ( n130 & n137 ) | ( n130 & n142 ) | ( n137 & n142 ) ;
  assign n144 = n137 | n142 ;
  assign n145 = ~n130 & n144 ;
  assign n146 = ( n130 & ~n143 ) | ( n130 & n145 ) | ( ~n143 & n145 ) ;
  assign n147 = ( x2 & n130 ) | ( x2 & n144 ) | ( n130 & n144 ) ;
  assign n148 = x65 & n138 ;
  assign n149 = x66 | n148 ;
  assign n150 = ( n141 & n148 ) | ( n141 & n149 ) | ( n148 & n149 ) ;
  assign n151 = ~x66 & n131 ;
  assign n152 = x66 & ~n131 ;
  assign n153 = ( n136 & n151 ) | ( n136 & n152 ) | ( n151 & n152 ) ;
  assign n154 = x2 & ~n135 ;
  assign n155 = ( x64 & n153 ) | ( x64 & n154 ) | ( n153 & n154 ) ;
  assign n156 = ( ~n150 & n153 ) | ( ~n150 & n155 ) | ( n153 & n155 ) ;
  assign n157 = n150 | n156 ;
  assign n158 = n147 | n157 ;
  assign n159 = ( n147 & n157 ) | ( n147 & ~n158 ) | ( n157 & ~n158 ) ;
  assign n160 = n158 & ~n159 ;
  assign n161 = ( x65 & x66 ) | ( x65 & n132 ) | ( x66 & n132 ) ;
  assign n162 = ( x66 & x67 ) | ( x66 & n161 ) | ( x67 & n161 ) ;
  assign n163 = ( x66 & ~x67 ) | ( x66 & n161 ) | ( ~x67 & n161 ) ;
  assign n164 = ( x67 & ~n162 ) | ( x67 & n163 ) | ( ~n162 & n163 ) ;
  assign n165 = n136 & n164 ;
  assign n166 = x66 & n138 ;
  assign n167 = x67 | n166 ;
  assign n168 = ( n141 & n166 ) | ( n141 & n167 ) | ( n166 & n167 ) ;
  assign n169 = x65 & n154 ;
  assign n170 = n168 | n169 ;
  assign n171 = ( ~x2 & n165 ) | ( ~x2 & n170 ) | ( n165 & n170 ) ;
  assign n172 = ( n165 & n170 ) | ( n165 & ~n171 ) | ( n170 & ~n171 ) ;
  assign n173 = ( x2 & n171 ) | ( x2 & ~n172 ) | ( n171 & ~n172 ) ;
  assign n174 = x2 & x3 ;
  assign n175 = x2 | x3 ;
  assign n176 = ~n174 & n175 ;
  assign n177 = x64 & n176 ;
  assign n178 = x2 & ~n158 ;
  assign n179 = ( n173 & n177 ) | ( n173 & n178 ) | ( n177 & n178 ) ;
  assign n180 = ( ~n173 & n177 ) | ( ~n173 & n178 ) | ( n177 & n178 ) ;
  assign n181 = ( n173 & ~n179 ) | ( n173 & n180 ) | ( ~n179 & n180 ) ;
  assign n182 = x5 & n177 ;
  assign n183 = x4 | x5 ;
  assign n184 = ( x4 & x5 ) | ( x4 & ~n183 ) | ( x5 & ~n183 ) ;
  assign n185 = n183 & ~n184 ;
  assign n186 = n176 & n185 ;
  assign n187 = n133 & n186 ;
  assign n188 = ~x2 & x4 ;
  assign n189 = x3 & x4 ;
  assign n190 = ( n174 & n188 ) | ( n174 & ~n189 ) | ( n188 & ~n189 ) ;
  assign n191 = x64 & n190 ;
  assign n192 = ( n176 & ~n183 ) | ( n176 & n184 ) | ( ~n183 & n184 ) ;
  assign n193 = x65 | n191 ;
  assign n194 = ( n191 & n192 ) | ( n191 & n193 ) | ( n192 & n193 ) ;
  assign n195 = ( n182 & n187 ) | ( n182 & n194 ) | ( n187 & n194 ) ;
  assign n196 = n187 | n194 ;
  assign n197 = ~n182 & n196 ;
  assign n198 = ( n182 & ~n195 ) | ( n182 & n197 ) | ( ~n195 & n197 ) ;
  assign n199 = ( x67 & x68 ) | ( x67 & n162 ) | ( x68 & n162 ) ;
  assign n200 = ( x67 & ~x68 ) | ( x67 & n162 ) | ( ~x68 & n162 ) ;
  assign n201 = ( x68 & ~n199 ) | ( x68 & n200 ) | ( ~n199 & n200 ) ;
  assign n202 = n136 & n201 ;
  assign n203 = x67 & n138 ;
  assign n204 = x68 | n203 ;
  assign n205 = ( n141 & n203 ) | ( n141 & n204 ) | ( n203 & n204 ) ;
  assign n206 = x66 & n154 ;
  assign n207 = n205 | n206 ;
  assign n208 = ( x2 & n202 ) | ( x2 & ~n207 ) | ( n202 & ~n207 ) ;
  assign n209 = ( ~x2 & n207 ) | ( ~x2 & n208 ) | ( n207 & n208 ) ;
  assign n210 = ( ~n202 & n208 ) | ( ~n202 & n209 ) | ( n208 & n209 ) ;
  assign n211 = ( n179 & n198 ) | ( n179 & n210 ) | ( n198 & n210 ) ;
  assign n212 = ( ~n179 & n198 ) | ( ~n179 & n210 ) | ( n198 & n210 ) ;
  assign n213 = ( n179 & ~n211 ) | ( n179 & n212 ) | ( ~n211 & n212 ) ;
  assign n214 = ( x5 & n182 ) | ( x5 & n196 ) | ( n182 & n196 ) ;
  assign n215 = n151 | n152 ;
  assign n216 = x66 & n192 ;
  assign n217 = ( n176 & ~n192 ) | ( n176 & n216 ) | ( ~n192 & n216 ) ;
  assign n218 = ( n215 & n216 ) | ( n215 & n217 ) | ( n216 & n217 ) ;
  assign n219 = ( x2 & ~x4 ) | ( x2 & n185 ) | ( ~x4 & n185 ) ;
  assign n220 = ( ~n175 & n189 ) | ( ~n175 & n219 ) | ( n189 & n219 ) ;
  assign n221 = x64 & n220 ;
  assign n222 = x65 & n190 ;
  assign n223 = ( ~n218 & n221 ) | ( ~n218 & n222 ) | ( n221 & n222 ) ;
  assign n224 = n218 | n223 ;
  assign n225 = n214 | n224 ;
  assign n226 = ( n214 & n224 ) | ( n214 & ~n225 ) | ( n224 & ~n225 ) ;
  assign n227 = n225 & ~n226 ;
  assign n228 = ( x68 & x69 ) | ( x68 & n199 ) | ( x69 & n199 ) ;
  assign n229 = ( x68 & ~x69 ) | ( x68 & n199 ) | ( ~x69 & n199 ) ;
  assign n230 = ( x69 & ~n228 ) | ( x69 & n229 ) | ( ~n228 & n229 ) ;
  assign n231 = n136 & n230 ;
  assign n232 = x68 & n138 ;
  assign n233 = x69 | n232 ;
  assign n234 = ( n141 & n232 ) | ( n141 & n233 ) | ( n232 & n233 ) ;
  assign n235 = x67 & n154 ;
  assign n236 = n234 | n235 ;
  assign n237 = ( x2 & n231 ) | ( x2 & ~n236 ) | ( n231 & ~n236 ) ;
  assign n238 = ( ~x2 & n236 ) | ( ~x2 & n237 ) | ( n236 & n237 ) ;
  assign n239 = ( ~n231 & n237 ) | ( ~n231 & n238 ) | ( n237 & n238 ) ;
  assign n240 = ( n211 & n227 ) | ( n211 & n239 ) | ( n227 & n239 ) ;
  assign n241 = ( n211 & ~n227 ) | ( n211 & n239 ) | ( ~n227 & n239 ) ;
  assign n242 = ( n227 & ~n240 ) | ( n227 & n241 ) | ( ~n240 & n241 ) ;
  assign n243 = ( x69 & x70 ) | ( x69 & n228 ) | ( x70 & n228 ) ;
  assign n244 = ( x69 & ~x70 ) | ( x69 & n228 ) | ( ~x70 & n228 ) ;
  assign n245 = ( x70 & ~n243 ) | ( x70 & n244 ) | ( ~n243 & n244 ) ;
  assign n246 = n136 & n245 ;
  assign n247 = x69 & n138 ;
  assign n248 = x70 | n247 ;
  assign n249 = ( n141 & n247 ) | ( n141 & n248 ) | ( n247 & n248 ) ;
  assign n250 = x68 & n154 ;
  assign n251 = n249 | n250 ;
  assign n252 = ( x2 & n246 ) | ( x2 & ~n251 ) | ( n246 & ~n251 ) ;
  assign n253 = ( ~x2 & n251 ) | ( ~x2 & n252 ) | ( n251 & n252 ) ;
  assign n254 = ( ~n246 & n252 ) | ( ~n246 & n253 ) | ( n252 & n253 ) ;
  assign n255 = x66 & n190 ;
  assign n256 = x67 | n255 ;
  assign n257 = ( n192 & n255 ) | ( n192 & n256 ) | ( n255 & n256 ) ;
  assign n258 = x65 & n220 ;
  assign n259 = n257 | n258 ;
  assign n260 = n164 & n186 ;
  assign n261 = ( x5 & n259 ) | ( x5 & ~n260 ) | ( n259 & ~n260 ) ;
  assign n262 = ( ~x5 & n260 ) | ( ~x5 & n261 ) | ( n260 & n261 ) ;
  assign n263 = ( ~n259 & n261 ) | ( ~n259 & n262 ) | ( n261 & n262 ) ;
  assign n264 = x5 & x6 ;
  assign n265 = x5 | x6 ;
  assign n266 = ~n264 & n265 ;
  assign n267 = x64 & n266 ;
  assign n268 = x5 & ~n225 ;
  assign n269 = ( n263 & n267 ) | ( n263 & n268 ) | ( n267 & n268 ) ;
  assign n270 = ( ~n263 & n267 ) | ( ~n263 & n268 ) | ( n267 & n268 ) ;
  assign n271 = ( n263 & ~n269 ) | ( n263 & n270 ) | ( ~n269 & n270 ) ;
  assign n272 = ( n240 & n254 ) | ( n240 & n271 ) | ( n254 & n271 ) ;
  assign n273 = ( ~n240 & n254 ) | ( ~n240 & n271 ) | ( n254 & n271 ) ;
  assign n274 = ( n240 & ~n272 ) | ( n240 & n273 ) | ( ~n272 & n273 ) ;
  assign n275 = ( x70 & x71 ) | ( x70 & n243 ) | ( x71 & n243 ) ;
  assign n276 = ( x70 & ~x71 ) | ( x70 & n243 ) | ( ~x71 & n243 ) ;
  assign n277 = ( x71 & ~n275 ) | ( x71 & n276 ) | ( ~n275 & n276 ) ;
  assign n278 = n136 & n277 ;
  assign n279 = x70 & n138 ;
  assign n280 = x71 | n279 ;
  assign n281 = ( n141 & n279 ) | ( n141 & n280 ) | ( n279 & n280 ) ;
  assign n282 = x69 & n154 ;
  assign n283 = n281 | n282 ;
  assign n284 = ( x2 & n278 ) | ( x2 & ~n283 ) | ( n278 & ~n283 ) ;
  assign n285 = ( ~x2 & n283 ) | ( ~x2 & n284 ) | ( n283 & n284 ) ;
  assign n286 = ( ~n278 & n284 ) | ( ~n278 & n285 ) | ( n284 & n285 ) ;
  assign n287 = x8 & n267 ;
  assign n288 = x7 | x8 ;
  assign n289 = ( x7 & x8 ) | ( x7 & ~n288 ) | ( x8 & ~n288 ) ;
  assign n290 = n288 & ~n289 ;
  assign n291 = n266 & n290 ;
  assign n292 = n133 & n291 ;
  assign n293 = ~x5 & x7 ;
  assign n294 = x6 & x7 ;
  assign n295 = ( n264 & n293 ) | ( n264 & ~n294 ) | ( n293 & ~n294 ) ;
  assign n296 = x64 & n295 ;
  assign n297 = ( n266 & ~n288 ) | ( n266 & n289 ) | ( ~n288 & n289 ) ;
  assign n298 = x65 | n296 ;
  assign n299 = ( n296 & n297 ) | ( n296 & n298 ) | ( n297 & n298 ) ;
  assign n300 = ( n287 & n292 ) | ( n287 & n299 ) | ( n292 & n299 ) ;
  assign n301 = n292 | n299 ;
  assign n302 = ~n287 & n301 ;
  assign n303 = ( n287 & ~n300 ) | ( n287 & n302 ) | ( ~n300 & n302 ) ;
  assign n304 = x67 & n190 ;
  assign n305 = x68 | n304 ;
  assign n306 = ( n192 & n304 ) | ( n192 & n305 ) | ( n304 & n305 ) ;
  assign n307 = x66 & n220 ;
  assign n308 = n306 | n307 ;
  assign n309 = n186 & n201 ;
  assign n310 = ( x5 & n308 ) | ( x5 & ~n309 ) | ( n308 & ~n309 ) ;
  assign n311 = ( ~x5 & n309 ) | ( ~x5 & n310 ) | ( n309 & n310 ) ;
  assign n312 = ( ~n308 & n310 ) | ( ~n308 & n311 ) | ( n310 & n311 ) ;
  assign n313 = ( n269 & n303 ) | ( n269 & n312 ) | ( n303 & n312 ) ;
  assign n314 = ( ~n269 & n303 ) | ( ~n269 & n312 ) | ( n303 & n312 ) ;
  assign n315 = ( n269 & ~n313 ) | ( n269 & n314 ) | ( ~n313 & n314 ) ;
  assign n316 = ( n272 & n286 ) | ( n272 & n315 ) | ( n286 & n315 ) ;
  assign n317 = ( ~n272 & n286 ) | ( ~n272 & n315 ) | ( n286 & n315 ) ;
  assign n318 = ( n272 & ~n316 ) | ( n272 & n317 ) | ( ~n316 & n317 ) ;
  assign n319 = n186 & n230 ;
  assign n320 = x68 & n190 ;
  assign n321 = x69 | n320 ;
  assign n322 = ( n192 & n320 ) | ( n192 & n321 ) | ( n320 & n321 ) ;
  assign n323 = x67 & n220 ;
  assign n324 = n322 | n323 ;
  assign n325 = ( ~x5 & n319 ) | ( ~x5 & n324 ) | ( n319 & n324 ) ;
  assign n326 = ( n319 & n324 ) | ( n319 & ~n325 ) | ( n324 & ~n325 ) ;
  assign n327 = ( x5 & n325 ) | ( x5 & ~n326 ) | ( n325 & ~n326 ) ;
  assign n328 = ( x8 & n287 ) | ( x8 & n301 ) | ( n287 & n301 ) ;
  assign n329 = ( x5 & ~x7 ) | ( x5 & n290 ) | ( ~x7 & n290 ) ;
  assign n330 = ( ~n265 & n294 ) | ( ~n265 & n329 ) | ( n294 & n329 ) ;
  assign n331 = x64 & n330 ;
  assign n332 = x65 & n295 ;
  assign n333 = x66 | n332 ;
  assign n334 = ( n297 & n332 ) | ( n297 & n333 ) | ( n332 & n333 ) ;
  assign n335 = ( n151 & n152 ) | ( n151 & n291 ) | ( n152 & n291 ) ;
  assign n336 = ( ~n331 & n334 ) | ( ~n331 & n335 ) | ( n334 & n335 ) ;
  assign n337 = n331 | n336 ;
  assign n338 = n328 | n337 ;
  assign n339 = ( n328 & n337 ) | ( n328 & ~n338 ) | ( n337 & ~n338 ) ;
  assign n340 = n338 & ~n339 ;
  assign n341 = ( n313 & n327 ) | ( n313 & n340 ) | ( n327 & n340 ) ;
  assign n342 = ( ~n313 & n327 ) | ( ~n313 & n340 ) | ( n327 & n340 ) ;
  assign n343 = ( n313 & ~n341 ) | ( n313 & n342 ) | ( ~n341 & n342 ) ;
  assign n344 = ( x71 & x72 ) | ( x71 & n275 ) | ( x72 & n275 ) ;
  assign n345 = ( x71 & ~x72 ) | ( x71 & n275 ) | ( ~x72 & n275 ) ;
  assign n346 = ( x72 & ~n344 ) | ( x72 & n345 ) | ( ~n344 & n345 ) ;
  assign n347 = n136 & n346 ;
  assign n348 = x71 & n138 ;
  assign n349 = x72 | n348 ;
  assign n350 = ( n141 & n348 ) | ( n141 & n349 ) | ( n348 & n349 ) ;
  assign n351 = x70 & n154 ;
  assign n352 = n350 | n351 ;
  assign n353 = ( x2 & n347 ) | ( x2 & ~n352 ) | ( n347 & ~n352 ) ;
  assign n354 = ( ~x2 & n352 ) | ( ~x2 & n353 ) | ( n352 & n353 ) ;
  assign n355 = ( ~n347 & n353 ) | ( ~n347 & n354 ) | ( n353 & n354 ) ;
  assign n356 = ( n316 & n343 ) | ( n316 & n355 ) | ( n343 & n355 ) ;
  assign n357 = ( ~n316 & n343 ) | ( ~n316 & n355 ) | ( n343 & n355 ) ;
  assign n358 = ( n316 & ~n356 ) | ( n316 & n357 ) | ( ~n356 & n357 ) ;
  assign n359 = x66 & n295 ;
  assign n360 = x67 | n359 ;
  assign n361 = ( n297 & n359 ) | ( n297 & n360 ) | ( n359 & n360 ) ;
  assign n362 = x65 & n330 ;
  assign n363 = n361 | n362 ;
  assign n364 = n164 & n291 ;
  assign n365 = ( x8 & n363 ) | ( x8 & ~n364 ) | ( n363 & ~n364 ) ;
  assign n366 = ( ~x8 & n364 ) | ( ~x8 & n365 ) | ( n364 & n365 ) ;
  assign n367 = ( ~n363 & n365 ) | ( ~n363 & n366 ) | ( n365 & n366 ) ;
  assign n368 = x8 & x9 ;
  assign n369 = x8 | x9 ;
  assign n370 = ~n368 & n369 ;
  assign n371 = x64 & n370 ;
  assign n372 = x8 & ~n338 ;
  assign n373 = ( n367 & n371 ) | ( n367 & n372 ) | ( n371 & n372 ) ;
  assign n374 = ( ~n367 & n371 ) | ( ~n367 & n372 ) | ( n371 & n372 ) ;
  assign n375 = ( n367 & ~n373 ) | ( n367 & n374 ) | ( ~n373 & n374 ) ;
  assign n376 = n186 & n245 ;
  assign n377 = x69 & n190 ;
  assign n378 = x70 | n377 ;
  assign n379 = ( n192 & n377 ) | ( n192 & n378 ) | ( n377 & n378 ) ;
  assign n380 = x68 & n220 ;
  assign n381 = n379 | n380 ;
  assign n382 = ( x5 & n376 ) | ( x5 & ~n381 ) | ( n376 & ~n381 ) ;
  assign n383 = ( ~x5 & n381 ) | ( ~x5 & n382 ) | ( n381 & n382 ) ;
  assign n384 = ( ~n376 & n382 ) | ( ~n376 & n383 ) | ( n382 & n383 ) ;
  assign n385 = ( n341 & n375 ) | ( n341 & n384 ) | ( n375 & n384 ) ;
  assign n386 = ( ~n341 & n375 ) | ( ~n341 & n384 ) | ( n375 & n384 ) ;
  assign n387 = ( n341 & ~n385 ) | ( n341 & n386 ) | ( ~n385 & n386 ) ;
  assign n388 = ( x72 & x73 ) | ( x72 & n344 ) | ( x73 & n344 ) ;
  assign n389 = ( x72 & ~x73 ) | ( x72 & n344 ) | ( ~x73 & n344 ) ;
  assign n390 = ( x73 & ~n388 ) | ( x73 & n389 ) | ( ~n388 & n389 ) ;
  assign n391 = n136 & n390 ;
  assign n392 = x72 & n138 ;
  assign n393 = x73 | n392 ;
  assign n394 = ( n141 & n392 ) | ( n141 & n393 ) | ( n392 & n393 ) ;
  assign n395 = x71 & n154 ;
  assign n396 = n394 | n395 ;
  assign n397 = ( x2 & n391 ) | ( x2 & ~n396 ) | ( n391 & ~n396 ) ;
  assign n398 = ( ~x2 & n396 ) | ( ~x2 & n397 ) | ( n396 & n397 ) ;
  assign n399 = ( ~n391 & n397 ) | ( ~n391 & n398 ) | ( n397 & n398 ) ;
  assign n400 = ( n356 & n387 ) | ( n356 & n399 ) | ( n387 & n399 ) ;
  assign n401 = ( ~n356 & n387 ) | ( ~n356 & n399 ) | ( n387 & n399 ) ;
  assign n402 = ( n356 & ~n400 ) | ( n356 & n401 ) | ( ~n400 & n401 ) ;
  assign n403 = x11 & n371 ;
  assign n404 = x10 | x11 ;
  assign n405 = ( x10 & x11 ) | ( x10 & ~n404 ) | ( x11 & ~n404 ) ;
  assign n406 = n404 & ~n405 ;
  assign n407 = n370 & n406 ;
  assign n408 = n133 & n407 ;
  assign n409 = ~x8 & x10 ;
  assign n410 = x9 & x10 ;
  assign n411 = ( n368 & n409 ) | ( n368 & ~n410 ) | ( n409 & ~n410 ) ;
  assign n412 = x64 & n411 ;
  assign n413 = ( n370 & ~n404 ) | ( n370 & n405 ) | ( ~n404 & n405 ) ;
  assign n414 = x65 | n412 ;
  assign n415 = ( n412 & n413 ) | ( n412 & n414 ) | ( n413 & n414 ) ;
  assign n416 = ( n403 & n408 ) | ( n403 & n415 ) | ( n408 & n415 ) ;
  assign n417 = n408 | n415 ;
  assign n418 = ~n403 & n417 ;
  assign n419 = ( n403 & ~n416 ) | ( n403 & n418 ) | ( ~n416 & n418 ) ;
  assign n420 = x67 & n295 ;
  assign n421 = x68 | n420 ;
  assign n422 = ( n297 & n420 ) | ( n297 & n421 ) | ( n420 & n421 ) ;
  assign n423 = x66 & n330 ;
  assign n424 = n422 | n423 ;
  assign n425 = n201 & n291 ;
  assign n426 = ( x8 & n424 ) | ( x8 & ~n425 ) | ( n424 & ~n425 ) ;
  assign n427 = ( ~x8 & n425 ) | ( ~x8 & n426 ) | ( n425 & n426 ) ;
  assign n428 = ( ~n424 & n426 ) | ( ~n424 & n427 ) | ( n426 & n427 ) ;
  assign n429 = ( n373 & n419 ) | ( n373 & n428 ) | ( n419 & n428 ) ;
  assign n430 = ( ~n373 & n419 ) | ( ~n373 & n428 ) | ( n419 & n428 ) ;
  assign n431 = ( n373 & ~n429 ) | ( n373 & n430 ) | ( ~n429 & n430 ) ;
  assign n432 = n186 & n277 ;
  assign n433 = x70 & n190 ;
  assign n434 = x71 | n433 ;
  assign n435 = ( n192 & n433 ) | ( n192 & n434 ) | ( n433 & n434 ) ;
  assign n436 = x69 & n220 ;
  assign n437 = n435 | n436 ;
  assign n438 = ( x5 & n432 ) | ( x5 & ~n437 ) | ( n432 & ~n437 ) ;
  assign n439 = ( ~x5 & n437 ) | ( ~x5 & n438 ) | ( n437 & n438 ) ;
  assign n440 = ( ~n432 & n438 ) | ( ~n432 & n439 ) | ( n438 & n439 ) ;
  assign n441 = ( n385 & n431 ) | ( n385 & n440 ) | ( n431 & n440 ) ;
  assign n442 = ( ~n385 & n431 ) | ( ~n385 & n440 ) | ( n431 & n440 ) ;
  assign n443 = ( n385 & ~n441 ) | ( n385 & n442 ) | ( ~n441 & n442 ) ;
  assign n444 = ( x73 & x74 ) | ( x73 & n388 ) | ( x74 & n388 ) ;
  assign n445 = ( x73 & ~x74 ) | ( x73 & n388 ) | ( ~x74 & n388 ) ;
  assign n446 = ( x74 & ~n444 ) | ( x74 & n445 ) | ( ~n444 & n445 ) ;
  assign n447 = n136 & n446 ;
  assign n448 = x73 & n138 ;
  assign n449 = x74 | n448 ;
  assign n450 = ( n141 & n448 ) | ( n141 & n449 ) | ( n448 & n449 ) ;
  assign n451 = x72 & n154 ;
  assign n452 = n450 | n451 ;
  assign n453 = ( x2 & n447 ) | ( x2 & ~n452 ) | ( n447 & ~n452 ) ;
  assign n454 = ( ~x2 & n452 ) | ( ~x2 & n453 ) | ( n452 & n453 ) ;
  assign n455 = ( ~n447 & n453 ) | ( ~n447 & n454 ) | ( n453 & n454 ) ;
  assign n456 = ( n400 & n443 ) | ( n400 & n455 ) | ( n443 & n455 ) ;
  assign n457 = ( ~n400 & n443 ) | ( ~n400 & n455 ) | ( n443 & n455 ) ;
  assign n458 = ( n400 & ~n456 ) | ( n400 & n457 ) | ( ~n456 & n457 ) ;
  assign n459 = ( x74 & x75 ) | ( x74 & n444 ) | ( x75 & n444 ) ;
  assign n460 = ( x74 & ~x75 ) | ( x74 & n444 ) | ( ~x75 & n444 ) ;
  assign n461 = ( x75 & ~n459 ) | ( x75 & n460 ) | ( ~n459 & n460 ) ;
  assign n462 = n136 & n461 ;
  assign n463 = x74 & n138 ;
  assign n464 = x75 | n463 ;
  assign n465 = ( n141 & n463 ) | ( n141 & n464 ) | ( n463 & n464 ) ;
  assign n466 = x73 & n154 ;
  assign n467 = n465 | n466 ;
  assign n468 = ( x2 & n462 ) | ( x2 & ~n467 ) | ( n462 & ~n467 ) ;
  assign n469 = ( ~x2 & n467 ) | ( ~x2 & n468 ) | ( n467 & n468 ) ;
  assign n470 = ( ~n462 & n468 ) | ( ~n462 & n469 ) | ( n468 & n469 ) ;
  assign n471 = n186 & n346 ;
  assign n472 = x71 & n190 ;
  assign n473 = x72 | n472 ;
  assign n474 = ( n192 & n472 ) | ( n192 & n473 ) | ( n472 & n473 ) ;
  assign n475 = x70 & n220 ;
  assign n476 = n474 | n475 ;
  assign n477 = ( x5 & n471 ) | ( x5 & ~n476 ) | ( n471 & ~n476 ) ;
  assign n478 = ( ~x5 & n476 ) | ( ~x5 & n477 ) | ( n476 & n477 ) ;
  assign n479 = ( ~n471 & n477 ) | ( ~n471 & n478 ) | ( n477 & n478 ) ;
  assign n480 = n230 & n291 ;
  assign n481 = x68 & n295 ;
  assign n482 = x69 | n481 ;
  assign n483 = ( n297 & n481 ) | ( n297 & n482 ) | ( n481 & n482 ) ;
  assign n484 = x67 & n330 ;
  assign n485 = n483 | n484 ;
  assign n486 = ( ~x8 & n480 ) | ( ~x8 & n485 ) | ( n480 & n485 ) ;
  assign n487 = ( n480 & n485 ) | ( n480 & ~n486 ) | ( n485 & ~n486 ) ;
  assign n488 = ( x8 & n486 ) | ( x8 & ~n487 ) | ( n486 & ~n487 ) ;
  assign n489 = ( x11 & n403 ) | ( x11 & n417 ) | ( n403 & n417 ) ;
  assign n490 = ( x8 & ~x10 ) | ( x8 & n406 ) | ( ~x10 & n406 ) ;
  assign n491 = ( ~n369 & n410 ) | ( ~n369 & n490 ) | ( n410 & n490 ) ;
  assign n492 = x64 & n491 ;
  assign n493 = x65 & n411 ;
  assign n494 = x66 | n493 ;
  assign n495 = ( n413 & n493 ) | ( n413 & n494 ) | ( n493 & n494 ) ;
  assign n496 = ( n151 & n152 ) | ( n151 & n407 ) | ( n152 & n407 ) ;
  assign n497 = ( ~n492 & n495 ) | ( ~n492 & n496 ) | ( n495 & n496 ) ;
  assign n498 = n492 | n497 ;
  assign n499 = n489 | n498 ;
  assign n500 = ( n489 & n498 ) | ( n489 & ~n499 ) | ( n498 & ~n499 ) ;
  assign n501 = n499 & ~n500 ;
  assign n502 = ( n429 & n488 ) | ( n429 & n501 ) | ( n488 & n501 ) ;
  assign n503 = ( ~n429 & n488 ) | ( ~n429 & n501 ) | ( n488 & n501 ) ;
  assign n504 = ( n429 & ~n502 ) | ( n429 & n503 ) | ( ~n502 & n503 ) ;
  assign n505 = ( n441 & n479 ) | ( n441 & n504 ) | ( n479 & n504 ) ;
  assign n506 = ( ~n441 & n479 ) | ( ~n441 & n504 ) | ( n479 & n504 ) ;
  assign n507 = ( n441 & ~n505 ) | ( n441 & n506 ) | ( ~n505 & n506 ) ;
  assign n508 = ( n456 & n470 ) | ( n456 & n507 ) | ( n470 & n507 ) ;
  assign n509 = ( ~n456 & n470 ) | ( ~n456 & n507 ) | ( n470 & n507 ) ;
  assign n510 = ( n456 & ~n508 ) | ( n456 & n509 ) | ( ~n508 & n509 ) ;
  assign n511 = x66 & n411 ;
  assign n512 = x67 | n511 ;
  assign n513 = ( n413 & n511 ) | ( n413 & n512 ) | ( n511 & n512 ) ;
  assign n514 = x65 & n491 ;
  assign n515 = n513 | n514 ;
  assign n516 = n164 & n407 ;
  assign n517 = ( x11 & n515 ) | ( x11 & ~n516 ) | ( n515 & ~n516 ) ;
  assign n518 = ( ~x11 & n516 ) | ( ~x11 & n517 ) | ( n516 & n517 ) ;
  assign n519 = ( ~n515 & n517 ) | ( ~n515 & n518 ) | ( n517 & n518 ) ;
  assign n520 = x11 & x12 ;
  assign n521 = x11 | x12 ;
  assign n522 = ~n520 & n521 ;
  assign n523 = x64 & n522 ;
  assign n524 = x11 & ~n499 ;
  assign n525 = ( n519 & n523 ) | ( n519 & n524 ) | ( n523 & n524 ) ;
  assign n526 = ( ~n519 & n523 ) | ( ~n519 & n524 ) | ( n523 & n524 ) ;
  assign n527 = ( n519 & ~n525 ) | ( n519 & n526 ) | ( ~n525 & n526 ) ;
  assign n528 = n245 & n291 ;
  assign n529 = x69 & n295 ;
  assign n530 = x70 | n529 ;
  assign n531 = ( n297 & n529 ) | ( n297 & n530 ) | ( n529 & n530 ) ;
  assign n532 = x68 & n330 ;
  assign n533 = n531 | n532 ;
  assign n534 = ( x8 & n528 ) | ( x8 & ~n533 ) | ( n528 & ~n533 ) ;
  assign n535 = ( ~x8 & n533 ) | ( ~x8 & n534 ) | ( n533 & n534 ) ;
  assign n536 = ( ~n528 & n534 ) | ( ~n528 & n535 ) | ( n534 & n535 ) ;
  assign n537 = ( n502 & n527 ) | ( n502 & n536 ) | ( n527 & n536 ) ;
  assign n538 = ( ~n502 & n527 ) | ( ~n502 & n536 ) | ( n527 & n536 ) ;
  assign n539 = ( n502 & ~n537 ) | ( n502 & n538 ) | ( ~n537 & n538 ) ;
  assign n540 = n186 & n390 ;
  assign n541 = x72 & n190 ;
  assign n542 = x73 | n541 ;
  assign n543 = ( n192 & n541 ) | ( n192 & n542 ) | ( n541 & n542 ) ;
  assign n544 = x71 & n220 ;
  assign n545 = n543 | n544 ;
  assign n546 = ( x5 & n540 ) | ( x5 & ~n545 ) | ( n540 & ~n545 ) ;
  assign n547 = ( ~x5 & n545 ) | ( ~x5 & n546 ) | ( n545 & n546 ) ;
  assign n548 = ( ~n540 & n546 ) | ( ~n540 & n547 ) | ( n546 & n547 ) ;
  assign n549 = ( n505 & n539 ) | ( n505 & n548 ) | ( n539 & n548 ) ;
  assign n550 = ( n505 & ~n539 ) | ( n505 & n548 ) | ( ~n539 & n548 ) ;
  assign n551 = ( n539 & ~n549 ) | ( n539 & n550 ) | ( ~n549 & n550 ) ;
  assign n552 = ( x75 & x76 ) | ( x75 & n459 ) | ( x76 & n459 ) ;
  assign n553 = ( x75 & ~x76 ) | ( x75 & n459 ) | ( ~x76 & n459 ) ;
  assign n554 = ( x76 & ~n552 ) | ( x76 & n553 ) | ( ~n552 & n553 ) ;
  assign n555 = n136 & n554 ;
  assign n556 = x75 & n138 ;
  assign n557 = x76 | n556 ;
  assign n558 = ( n141 & n556 ) | ( n141 & n557 ) | ( n556 & n557 ) ;
  assign n559 = x74 & n154 ;
  assign n560 = n558 | n559 ;
  assign n561 = ( x2 & n555 ) | ( x2 & ~n560 ) | ( n555 & ~n560 ) ;
  assign n562 = ( ~x2 & n560 ) | ( ~x2 & n561 ) | ( n560 & n561 ) ;
  assign n563 = ( ~n555 & n561 ) | ( ~n555 & n562 ) | ( n561 & n562 ) ;
  assign n564 = ( n508 & n551 ) | ( n508 & n563 ) | ( n551 & n563 ) ;
  assign n565 = ( ~n508 & n551 ) | ( ~n508 & n563 ) | ( n551 & n563 ) ;
  assign n566 = ( n508 & ~n564 ) | ( n508 & n565 ) | ( ~n564 & n565 ) ;
  assign n567 = ( x76 & x77 ) | ( x76 & n552 ) | ( x77 & n552 ) ;
  assign n568 = ( x76 & ~x77 ) | ( x76 & n552 ) | ( ~x77 & n552 ) ;
  assign n569 = ( x77 & ~n567 ) | ( x77 & n568 ) | ( ~n567 & n568 ) ;
  assign n570 = n136 & n569 ;
  assign n571 = x76 & n138 ;
  assign n572 = x77 | n571 ;
  assign n573 = ( n141 & n571 ) | ( n141 & n572 ) | ( n571 & n572 ) ;
  assign n574 = x75 & n154 ;
  assign n575 = n573 | n574 ;
  assign n576 = ( x2 & n570 ) | ( x2 & ~n575 ) | ( n570 & ~n575 ) ;
  assign n577 = ( ~x2 & n575 ) | ( ~x2 & n576 ) | ( n575 & n576 ) ;
  assign n578 = ( ~n570 & n576 ) | ( ~n570 & n577 ) | ( n576 & n577 ) ;
  assign n579 = x14 & n523 ;
  assign n580 = x13 | x14 ;
  assign n581 = ( x13 & x14 ) | ( x13 & ~n580 ) | ( x14 & ~n580 ) ;
  assign n582 = n580 & ~n581 ;
  assign n583 = n522 & n582 ;
  assign n584 = n133 & n583 ;
  assign n585 = ~x11 & x13 ;
  assign n586 = x12 & x13 ;
  assign n587 = ( n520 & n585 ) | ( n520 & ~n586 ) | ( n585 & ~n586 ) ;
  assign n588 = x64 & n587 ;
  assign n589 = ( n522 & ~n580 ) | ( n522 & n581 ) | ( ~n580 & n581 ) ;
  assign n590 = x65 | n588 ;
  assign n591 = ( n588 & n589 ) | ( n588 & n590 ) | ( n589 & n590 ) ;
  assign n592 = ( n579 & n584 ) | ( n579 & n591 ) | ( n584 & n591 ) ;
  assign n593 = n584 | n591 ;
  assign n594 = ~n579 & n593 ;
  assign n595 = ( n579 & ~n592 ) | ( n579 & n594 ) | ( ~n592 & n594 ) ;
  assign n596 = x67 & n411 ;
  assign n597 = x68 | n596 ;
  assign n598 = ( n413 & n596 ) | ( n413 & n597 ) | ( n596 & n597 ) ;
  assign n599 = x66 & n491 ;
  assign n600 = n598 | n599 ;
  assign n601 = n201 & n407 ;
  assign n602 = ( x11 & n600 ) | ( x11 & ~n601 ) | ( n600 & ~n601 ) ;
  assign n603 = ( ~x11 & n601 ) | ( ~x11 & n602 ) | ( n601 & n602 ) ;
  assign n604 = ( ~n600 & n602 ) | ( ~n600 & n603 ) | ( n602 & n603 ) ;
  assign n605 = ( n525 & n595 ) | ( n525 & n604 ) | ( n595 & n604 ) ;
  assign n606 = ( ~n525 & n595 ) | ( ~n525 & n604 ) | ( n595 & n604 ) ;
  assign n607 = ( n525 & ~n605 ) | ( n525 & n606 ) | ( ~n605 & n606 ) ;
  assign n608 = n277 & n291 ;
  assign n609 = x70 & n295 ;
  assign n610 = x71 | n609 ;
  assign n611 = ( n297 & n609 ) | ( n297 & n610 ) | ( n609 & n610 ) ;
  assign n612 = x69 & n330 ;
  assign n613 = n611 | n612 ;
  assign n614 = ( x8 & n608 ) | ( x8 & ~n613 ) | ( n608 & ~n613 ) ;
  assign n615 = ( ~x8 & n613 ) | ( ~x8 & n614 ) | ( n613 & n614 ) ;
  assign n616 = ( ~n608 & n614 ) | ( ~n608 & n615 ) | ( n614 & n615 ) ;
  assign n617 = ( n537 & n607 ) | ( n537 & n616 ) | ( n607 & n616 ) ;
  assign n618 = ( ~n537 & n607 ) | ( ~n537 & n616 ) | ( n607 & n616 ) ;
  assign n619 = ( n537 & ~n617 ) | ( n537 & n618 ) | ( ~n617 & n618 ) ;
  assign n620 = n186 & n446 ;
  assign n621 = x73 & n190 ;
  assign n622 = x74 | n621 ;
  assign n623 = ( n192 & n621 ) | ( n192 & n622 ) | ( n621 & n622 ) ;
  assign n624 = x72 & n220 ;
  assign n625 = n623 | n624 ;
  assign n626 = ( x5 & n620 ) | ( x5 & ~n625 ) | ( n620 & ~n625 ) ;
  assign n627 = ( ~x5 & n625 ) | ( ~x5 & n626 ) | ( n625 & n626 ) ;
  assign n628 = ( ~n620 & n626 ) | ( ~n620 & n627 ) | ( n626 & n627 ) ;
  assign n629 = ( n549 & n619 ) | ( n549 & n628 ) | ( n619 & n628 ) ;
  assign n630 = ( ~n549 & n619 ) | ( ~n549 & n628 ) | ( n619 & n628 ) ;
  assign n631 = ( n549 & ~n629 ) | ( n549 & n630 ) | ( ~n629 & n630 ) ;
  assign n632 = ( n564 & n578 ) | ( n564 & n631 ) | ( n578 & n631 ) ;
  assign n633 = ( ~n564 & n578 ) | ( ~n564 & n631 ) | ( n578 & n631 ) ;
  assign n634 = ( n564 & ~n632 ) | ( n564 & n633 ) | ( ~n632 & n633 ) ;
  assign n635 = ( x77 & x78 ) | ( x77 & n567 ) | ( x78 & n567 ) ;
  assign n636 = ( x77 & ~x78 ) | ( x77 & n567 ) | ( ~x78 & n567 ) ;
  assign n637 = ( x78 & ~n635 ) | ( x78 & n636 ) | ( ~n635 & n636 ) ;
  assign n638 = n136 & n637 ;
  assign n639 = x77 & n138 ;
  assign n640 = x78 | n639 ;
  assign n641 = ( n141 & n639 ) | ( n141 & n640 ) | ( n639 & n640 ) ;
  assign n642 = x76 & n154 ;
  assign n643 = n641 | n642 ;
  assign n644 = ( x2 & n638 ) | ( x2 & ~n643 ) | ( n638 & ~n643 ) ;
  assign n645 = ( ~x2 & n643 ) | ( ~x2 & n644 ) | ( n643 & n644 ) ;
  assign n646 = ( ~n638 & n644 ) | ( ~n638 & n645 ) | ( n644 & n645 ) ;
  assign n647 = n186 & n461 ;
  assign n648 = x74 & n190 ;
  assign n649 = x75 | n648 ;
  assign n650 = ( n192 & n648 ) | ( n192 & n649 ) | ( n648 & n649 ) ;
  assign n651 = x73 & n220 ;
  assign n652 = n650 | n651 ;
  assign n653 = ( x5 & n647 ) | ( x5 & ~n652 ) | ( n647 & ~n652 ) ;
  assign n654 = ( ~x5 & n652 ) | ( ~x5 & n653 ) | ( n652 & n653 ) ;
  assign n655 = ( ~n647 & n653 ) | ( ~n647 & n654 ) | ( n653 & n654 ) ;
  assign n656 = n291 & n346 ;
  assign n657 = x71 & n295 ;
  assign n658 = x72 | n657 ;
  assign n659 = ( n297 & n657 ) | ( n297 & n658 ) | ( n657 & n658 ) ;
  assign n660 = x70 & n330 ;
  assign n661 = n659 | n660 ;
  assign n662 = ( x8 & n656 ) | ( x8 & ~n661 ) | ( n656 & ~n661 ) ;
  assign n663 = ( ~x8 & n661 ) | ( ~x8 & n662 ) | ( n661 & n662 ) ;
  assign n664 = ( ~n656 & n662 ) | ( ~n656 & n663 ) | ( n662 & n663 ) ;
  assign n665 = n230 & n407 ;
  assign n666 = x68 & n411 ;
  assign n667 = x69 | n666 ;
  assign n668 = ( n413 & n666 ) | ( n413 & n667 ) | ( n666 & n667 ) ;
  assign n669 = x67 & n491 ;
  assign n670 = n668 | n669 ;
  assign n671 = ( ~x11 & n665 ) | ( ~x11 & n670 ) | ( n665 & n670 ) ;
  assign n672 = ( n665 & n670 ) | ( n665 & ~n671 ) | ( n670 & ~n671 ) ;
  assign n673 = ( x11 & n671 ) | ( x11 & ~n672 ) | ( n671 & ~n672 ) ;
  assign n674 = ( x14 & n579 ) | ( x14 & n593 ) | ( n579 & n593 ) ;
  assign n675 = ( x11 & ~x13 ) | ( x11 & n582 ) | ( ~x13 & n582 ) ;
  assign n676 = ( ~n521 & n586 ) | ( ~n521 & n675 ) | ( n586 & n675 ) ;
  assign n677 = x64 & n676 ;
  assign n678 = x65 & n587 ;
  assign n679 = x66 | n678 ;
  assign n680 = ( n589 & n678 ) | ( n589 & n679 ) | ( n678 & n679 ) ;
  assign n681 = ( n151 & n152 ) | ( n151 & n583 ) | ( n152 & n583 ) ;
  assign n682 = ( ~n677 & n680 ) | ( ~n677 & n681 ) | ( n680 & n681 ) ;
  assign n683 = n677 | n682 ;
  assign n684 = n674 | n683 ;
  assign n685 = ( n674 & n683 ) | ( n674 & ~n684 ) | ( n683 & ~n684 ) ;
  assign n686 = n684 & ~n685 ;
  assign n687 = ( n605 & n673 ) | ( n605 & n686 ) | ( n673 & n686 ) ;
  assign n688 = ( ~n605 & n673 ) | ( ~n605 & n686 ) | ( n673 & n686 ) ;
  assign n689 = ( n605 & ~n687 ) | ( n605 & n688 ) | ( ~n687 & n688 ) ;
  assign n690 = ( n617 & n664 ) | ( n617 & n689 ) | ( n664 & n689 ) ;
  assign n691 = ( ~n617 & n664 ) | ( ~n617 & n689 ) | ( n664 & n689 ) ;
  assign n692 = ( n617 & ~n690 ) | ( n617 & n691 ) | ( ~n690 & n691 ) ;
  assign n693 = ( n629 & n655 ) | ( n629 & n692 ) | ( n655 & n692 ) ;
  assign n694 = ( ~n629 & n655 ) | ( ~n629 & n692 ) | ( n655 & n692 ) ;
  assign n695 = ( n629 & ~n693 ) | ( n629 & n694 ) | ( ~n693 & n694 ) ;
  assign n696 = ( n632 & n646 ) | ( n632 & n695 ) | ( n646 & n695 ) ;
  assign n697 = ( ~n632 & n646 ) | ( ~n632 & n695 ) | ( n646 & n695 ) ;
  assign n698 = ( n632 & ~n696 ) | ( n632 & n697 ) | ( ~n696 & n697 ) ;
  assign n699 = ( x78 & x79 ) | ( x78 & n635 ) | ( x79 & n635 ) ;
  assign n700 = ( x78 & ~x79 ) | ( x78 & n635 ) | ( ~x79 & n635 ) ;
  assign n701 = ( x79 & ~n699 ) | ( x79 & n700 ) | ( ~n699 & n700 ) ;
  assign n702 = n136 & n701 ;
  assign n703 = x78 & n138 ;
  assign n704 = x79 | n703 ;
  assign n705 = ( n141 & n703 ) | ( n141 & n704 ) | ( n703 & n704 ) ;
  assign n706 = x77 & n154 ;
  assign n707 = n705 | n706 ;
  assign n708 = ( x2 & n702 ) | ( x2 & ~n707 ) | ( n702 & ~n707 ) ;
  assign n709 = ( ~x2 & n707 ) | ( ~x2 & n708 ) | ( n707 & n708 ) ;
  assign n710 = ( ~n702 & n708 ) | ( ~n702 & n709 ) | ( n708 & n709 ) ;
  assign n711 = n186 & n554 ;
  assign n712 = x75 & n190 ;
  assign n713 = x76 | n712 ;
  assign n714 = ( n192 & n712 ) | ( n192 & n713 ) | ( n712 & n713 ) ;
  assign n715 = x74 & n220 ;
  assign n716 = n714 | n715 ;
  assign n717 = ( x5 & n711 ) | ( x5 & ~n716 ) | ( n711 & ~n716 ) ;
  assign n718 = ( ~x5 & n716 ) | ( ~x5 & n717 ) | ( n716 & n717 ) ;
  assign n719 = ( ~n711 & n717 ) | ( ~n711 & n718 ) | ( n717 & n718 ) ;
  assign n720 = n291 & n390 ;
  assign n721 = x72 & n295 ;
  assign n722 = x73 | n721 ;
  assign n723 = ( n297 & n721 ) | ( n297 & n722 ) | ( n721 & n722 ) ;
  assign n724 = x71 & n330 ;
  assign n725 = n723 | n724 ;
  assign n726 = ( x8 & n720 ) | ( x8 & ~n725 ) | ( n720 & ~n725 ) ;
  assign n727 = ( ~x8 & n725 ) | ( ~x8 & n726 ) | ( n725 & n726 ) ;
  assign n728 = ( ~n720 & n726 ) | ( ~n720 & n727 ) | ( n726 & n727 ) ;
  assign n729 = x66 & n587 ;
  assign n730 = x67 | n729 ;
  assign n731 = ( n589 & n729 ) | ( n589 & n730 ) | ( n729 & n730 ) ;
  assign n732 = x65 & n676 ;
  assign n733 = n731 | n732 ;
  assign n734 = n164 & n583 ;
  assign n735 = ( x14 & n733 ) | ( x14 & ~n734 ) | ( n733 & ~n734 ) ;
  assign n736 = ( ~x14 & n734 ) | ( ~x14 & n735 ) | ( n734 & n735 ) ;
  assign n737 = ( ~n733 & n735 ) | ( ~n733 & n736 ) | ( n735 & n736 ) ;
  assign n738 = x14 & x15 ;
  assign n739 = x14 | x15 ;
  assign n740 = ~n738 & n739 ;
  assign n741 = x64 & n740 ;
  assign n742 = x14 & ~n684 ;
  assign n743 = ( n737 & n741 ) | ( n737 & n742 ) | ( n741 & n742 ) ;
  assign n744 = ( ~n737 & n741 ) | ( ~n737 & n742 ) | ( n741 & n742 ) ;
  assign n745 = ( n737 & ~n743 ) | ( n737 & n744 ) | ( ~n743 & n744 ) ;
  assign n746 = n245 & n407 ;
  assign n747 = x69 & n411 ;
  assign n748 = x70 | n747 ;
  assign n749 = ( n413 & n747 ) | ( n413 & n748 ) | ( n747 & n748 ) ;
  assign n750 = x68 & n491 ;
  assign n751 = n749 | n750 ;
  assign n752 = ( x11 & n746 ) | ( x11 & ~n751 ) | ( n746 & ~n751 ) ;
  assign n753 = ( ~x11 & n751 ) | ( ~x11 & n752 ) | ( n751 & n752 ) ;
  assign n754 = ( ~n746 & n752 ) | ( ~n746 & n753 ) | ( n752 & n753 ) ;
  assign n755 = ( n687 & n745 ) | ( n687 & n754 ) | ( n745 & n754 ) ;
  assign n756 = ( ~n687 & n745 ) | ( ~n687 & n754 ) | ( n745 & n754 ) ;
  assign n757 = ( n687 & ~n755 ) | ( n687 & n756 ) | ( ~n755 & n756 ) ;
  assign n758 = ( n690 & n728 ) | ( n690 & n757 ) | ( n728 & n757 ) ;
  assign n759 = ( ~n690 & n728 ) | ( ~n690 & n757 ) | ( n728 & n757 ) ;
  assign n760 = ( n690 & ~n758 ) | ( n690 & n759 ) | ( ~n758 & n759 ) ;
  assign n761 = ( n693 & n719 ) | ( n693 & n760 ) | ( n719 & n760 ) ;
  assign n762 = ( ~n693 & n719 ) | ( ~n693 & n760 ) | ( n719 & n760 ) ;
  assign n763 = ( n693 & ~n761 ) | ( n693 & n762 ) | ( ~n761 & n762 ) ;
  assign n764 = ( n696 & n710 ) | ( n696 & n763 ) | ( n710 & n763 ) ;
  assign n765 = ( ~n696 & n710 ) | ( ~n696 & n763 ) | ( n710 & n763 ) ;
  assign n766 = ( n696 & ~n764 ) | ( n696 & n765 ) | ( ~n764 & n765 ) ;
  assign n767 = ( x79 & x80 ) | ( x79 & n699 ) | ( x80 & n699 ) ;
  assign n768 = ( x79 & ~x80 ) | ( x79 & n699 ) | ( ~x80 & n699 ) ;
  assign n769 = ( x80 & ~n767 ) | ( x80 & n768 ) | ( ~n767 & n768 ) ;
  assign n770 = n136 & n769 ;
  assign n771 = x79 & n138 ;
  assign n772 = x80 | n771 ;
  assign n773 = ( n141 & n771 ) | ( n141 & n772 ) | ( n771 & n772 ) ;
  assign n774 = x78 & n154 ;
  assign n775 = n773 | n774 ;
  assign n776 = ( x2 & n770 ) | ( x2 & ~n775 ) | ( n770 & ~n775 ) ;
  assign n777 = ( ~x2 & n775 ) | ( ~x2 & n776 ) | ( n775 & n776 ) ;
  assign n778 = ( ~n770 & n776 ) | ( ~n770 & n777 ) | ( n776 & n777 ) ;
  assign n779 = n186 & n569 ;
  assign n780 = x76 & n190 ;
  assign n781 = x77 | n780 ;
  assign n782 = ( n192 & n780 ) | ( n192 & n781 ) | ( n780 & n781 ) ;
  assign n783 = x75 & n220 ;
  assign n784 = n782 | n783 ;
  assign n785 = ( x5 & n779 ) | ( x5 & ~n784 ) | ( n779 & ~n784 ) ;
  assign n786 = ( ~x5 & n784 ) | ( ~x5 & n785 ) | ( n784 & n785 ) ;
  assign n787 = ( ~n779 & n785 ) | ( ~n779 & n786 ) | ( n785 & n786 ) ;
  assign n788 = n291 & n446 ;
  assign n789 = x73 & n295 ;
  assign n790 = x74 | n789 ;
  assign n791 = ( n297 & n789 ) | ( n297 & n790 ) | ( n789 & n790 ) ;
  assign n792 = x72 & n330 ;
  assign n793 = n791 | n792 ;
  assign n794 = ( x8 & n788 ) | ( x8 & ~n793 ) | ( n788 & ~n793 ) ;
  assign n795 = ( ~x8 & n793 ) | ( ~x8 & n794 ) | ( n793 & n794 ) ;
  assign n796 = ( ~n788 & n794 ) | ( ~n788 & n795 ) | ( n794 & n795 ) ;
  assign n797 = n277 & n407 ;
  assign n798 = x70 & n411 ;
  assign n799 = x71 | n798 ;
  assign n800 = ( n413 & n798 ) | ( n413 & n799 ) | ( n798 & n799 ) ;
  assign n801 = x69 & n491 ;
  assign n802 = n800 | n801 ;
  assign n803 = ( x11 & n797 ) | ( x11 & ~n802 ) | ( n797 & ~n802 ) ;
  assign n804 = ( ~x11 & n802 ) | ( ~x11 & n803 ) | ( n802 & n803 ) ;
  assign n805 = ( ~n797 & n803 ) | ( ~n797 & n804 ) | ( n803 & n804 ) ;
  assign n806 = x17 & n741 ;
  assign n807 = x16 | x17 ;
  assign n808 = ( x16 & x17 ) | ( x16 & ~n807 ) | ( x17 & ~n807 ) ;
  assign n809 = n807 & ~n808 ;
  assign n810 = n740 & n809 ;
  assign n811 = n133 & n810 ;
  assign n812 = ~x14 & x16 ;
  assign n813 = x15 & x16 ;
  assign n814 = ( n738 & n812 ) | ( n738 & ~n813 ) | ( n812 & ~n813 ) ;
  assign n815 = x64 & n814 ;
  assign n816 = ( n740 & ~n807 ) | ( n740 & n808 ) | ( ~n807 & n808 ) ;
  assign n817 = x65 | n815 ;
  assign n818 = ( n815 & n816 ) | ( n815 & n817 ) | ( n816 & n817 ) ;
  assign n819 = ( n806 & n811 ) | ( n806 & n818 ) | ( n811 & n818 ) ;
  assign n820 = n811 | n818 ;
  assign n821 = ~n806 & n820 ;
  assign n822 = ( n806 & ~n819 ) | ( n806 & n821 ) | ( ~n819 & n821 ) ;
  assign n823 = x67 & n587 ;
  assign n824 = x68 | n823 ;
  assign n825 = ( n589 & n823 ) | ( n589 & n824 ) | ( n823 & n824 ) ;
  assign n826 = x66 & n676 ;
  assign n827 = n825 | n826 ;
  assign n828 = n201 & n583 ;
  assign n829 = ( x14 & n827 ) | ( x14 & ~n828 ) | ( n827 & ~n828 ) ;
  assign n830 = ( ~x14 & n828 ) | ( ~x14 & n829 ) | ( n828 & n829 ) ;
  assign n831 = ( ~n827 & n829 ) | ( ~n827 & n830 ) | ( n829 & n830 ) ;
  assign n832 = ( n743 & n822 ) | ( n743 & n831 ) | ( n822 & n831 ) ;
  assign n833 = ( ~n743 & n822 ) | ( ~n743 & n831 ) | ( n822 & n831 ) ;
  assign n834 = ( n743 & ~n832 ) | ( n743 & n833 ) | ( ~n832 & n833 ) ;
  assign n835 = ( n755 & n805 ) | ( n755 & n834 ) | ( n805 & n834 ) ;
  assign n836 = ( ~n755 & n805 ) | ( ~n755 & n834 ) | ( n805 & n834 ) ;
  assign n837 = ( n755 & ~n835 ) | ( n755 & n836 ) | ( ~n835 & n836 ) ;
  assign n838 = ( n758 & n796 ) | ( n758 & n837 ) | ( n796 & n837 ) ;
  assign n839 = ( ~n758 & n796 ) | ( ~n758 & n837 ) | ( n796 & n837 ) ;
  assign n840 = ( n758 & ~n838 ) | ( n758 & n839 ) | ( ~n838 & n839 ) ;
  assign n841 = ( n761 & n787 ) | ( n761 & n840 ) | ( n787 & n840 ) ;
  assign n842 = ( ~n761 & n787 ) | ( ~n761 & n840 ) | ( n787 & n840 ) ;
  assign n843 = ( n761 & ~n841 ) | ( n761 & n842 ) | ( ~n841 & n842 ) ;
  assign n844 = ( n764 & n778 ) | ( n764 & n843 ) | ( n778 & n843 ) ;
  assign n845 = ( ~n764 & n778 ) | ( ~n764 & n843 ) | ( n778 & n843 ) ;
  assign n846 = ( n764 & ~n844 ) | ( n764 & n845 ) | ( ~n844 & n845 ) ;
  assign n847 = n186 & n637 ;
  assign n848 = x77 & n190 ;
  assign n849 = x78 | n848 ;
  assign n850 = ( n192 & n848 ) | ( n192 & n849 ) | ( n848 & n849 ) ;
  assign n851 = x76 & n220 ;
  assign n852 = n850 | n851 ;
  assign n853 = ( x5 & n847 ) | ( x5 & ~n852 ) | ( n847 & ~n852 ) ;
  assign n854 = ( ~x5 & n852 ) | ( ~x5 & n853 ) | ( n852 & n853 ) ;
  assign n855 = ( ~n847 & n853 ) | ( ~n847 & n854 ) | ( n853 & n854 ) ;
  assign n856 = n291 & n461 ;
  assign n857 = x74 & n295 ;
  assign n858 = x75 | n857 ;
  assign n859 = ( n297 & n857 ) | ( n297 & n858 ) | ( n857 & n858 ) ;
  assign n860 = x73 & n330 ;
  assign n861 = n859 | n860 ;
  assign n862 = ( x8 & n856 ) | ( x8 & ~n861 ) | ( n856 & ~n861 ) ;
  assign n863 = ( ~x8 & n861 ) | ( ~x8 & n862 ) | ( n861 & n862 ) ;
  assign n864 = ( ~n856 & n862 ) | ( ~n856 & n863 ) | ( n862 & n863 ) ;
  assign n865 = n346 & n407 ;
  assign n866 = x71 & n411 ;
  assign n867 = x72 | n866 ;
  assign n868 = ( n413 & n866 ) | ( n413 & n867 ) | ( n866 & n867 ) ;
  assign n869 = x70 & n491 ;
  assign n870 = n868 | n869 ;
  assign n871 = ( x11 & n865 ) | ( x11 & ~n870 ) | ( n865 & ~n870 ) ;
  assign n872 = ( ~x11 & n870 ) | ( ~x11 & n871 ) | ( n870 & n871 ) ;
  assign n873 = ( ~n865 & n871 ) | ( ~n865 & n872 ) | ( n871 & n872 ) ;
  assign n874 = n230 & n583 ;
  assign n875 = x68 & n587 ;
  assign n876 = x69 | n875 ;
  assign n877 = ( n589 & n875 ) | ( n589 & n876 ) | ( n875 & n876 ) ;
  assign n878 = x67 & n676 ;
  assign n879 = n877 | n878 ;
  assign n880 = ( ~x14 & n874 ) | ( ~x14 & n879 ) | ( n874 & n879 ) ;
  assign n881 = ( n874 & n879 ) | ( n874 & ~n880 ) | ( n879 & ~n880 ) ;
  assign n882 = ( x14 & n880 ) | ( x14 & ~n881 ) | ( n880 & ~n881 ) ;
  assign n883 = ( x17 & n806 ) | ( x17 & n820 ) | ( n806 & n820 ) ;
  assign n884 = ( x14 & ~x16 ) | ( x14 & n809 ) | ( ~x16 & n809 ) ;
  assign n885 = ( ~n739 & n813 ) | ( ~n739 & n884 ) | ( n813 & n884 ) ;
  assign n886 = x64 & n885 ;
  assign n887 = x65 & n814 ;
  assign n888 = x66 | n887 ;
  assign n889 = ( n816 & n887 ) | ( n816 & n888 ) | ( n887 & n888 ) ;
  assign n890 = ( n151 & n152 ) | ( n151 & n810 ) | ( n152 & n810 ) ;
  assign n891 = ( ~n886 & n889 ) | ( ~n886 & n890 ) | ( n889 & n890 ) ;
  assign n892 = n886 | n891 ;
  assign n893 = n883 | n892 ;
  assign n894 = ( n883 & n892 ) | ( n883 & ~n893 ) | ( n892 & ~n893 ) ;
  assign n895 = n893 & ~n894 ;
  assign n896 = ( n832 & n882 ) | ( n832 & n895 ) | ( n882 & n895 ) ;
  assign n897 = ( ~n832 & n882 ) | ( ~n832 & n895 ) | ( n882 & n895 ) ;
  assign n898 = ( n832 & ~n896 ) | ( n832 & n897 ) | ( ~n896 & n897 ) ;
  assign n899 = ( n835 & n873 ) | ( n835 & n898 ) | ( n873 & n898 ) ;
  assign n900 = ( ~n835 & n873 ) | ( ~n835 & n898 ) | ( n873 & n898 ) ;
  assign n901 = ( n835 & ~n899 ) | ( n835 & n900 ) | ( ~n899 & n900 ) ;
  assign n902 = ( n838 & n864 ) | ( n838 & n901 ) | ( n864 & n901 ) ;
  assign n903 = ( ~n838 & n864 ) | ( ~n838 & n901 ) | ( n864 & n901 ) ;
  assign n904 = ( n838 & ~n902 ) | ( n838 & n903 ) | ( ~n902 & n903 ) ;
  assign n905 = ( n841 & n855 ) | ( n841 & n904 ) | ( n855 & n904 ) ;
  assign n906 = ( ~n841 & n855 ) | ( ~n841 & n904 ) | ( n855 & n904 ) ;
  assign n907 = ( n841 & ~n905 ) | ( n841 & n906 ) | ( ~n905 & n906 ) ;
  assign n908 = ( x80 & x81 ) | ( x80 & n767 ) | ( x81 & n767 ) ;
  assign n909 = ( x80 & ~x81 ) | ( x80 & n767 ) | ( ~x81 & n767 ) ;
  assign n910 = ( x81 & ~n908 ) | ( x81 & n909 ) | ( ~n908 & n909 ) ;
  assign n911 = n136 & n910 ;
  assign n912 = x80 & n138 ;
  assign n913 = x81 | n912 ;
  assign n914 = ( n141 & n912 ) | ( n141 & n913 ) | ( n912 & n913 ) ;
  assign n915 = x79 & n154 ;
  assign n916 = n914 | n915 ;
  assign n917 = ( x2 & n911 ) | ( x2 & ~n916 ) | ( n911 & ~n916 ) ;
  assign n918 = ( ~x2 & n916 ) | ( ~x2 & n917 ) | ( n916 & n917 ) ;
  assign n919 = ( ~n911 & n917 ) | ( ~n911 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ( n844 & n907 ) | ( n844 & n919 ) | ( n907 & n919 ) ;
  assign n921 = ( ~n844 & n907 ) | ( ~n844 & n919 ) | ( n907 & n919 ) ;
  assign n922 = ( n844 & ~n920 ) | ( n844 & n921 ) | ( ~n920 & n921 ) ;
  assign n923 = n186 & n701 ;
  assign n924 = x78 & n190 ;
  assign n925 = x79 | n924 ;
  assign n926 = ( n192 & n924 ) | ( n192 & n925 ) | ( n924 & n925 ) ;
  assign n927 = x77 & n220 ;
  assign n928 = n926 | n927 ;
  assign n929 = ( x5 & n923 ) | ( x5 & ~n928 ) | ( n923 & ~n928 ) ;
  assign n930 = ( ~x5 & n928 ) | ( ~x5 & n929 ) | ( n928 & n929 ) ;
  assign n931 = ( ~n923 & n929 ) | ( ~n923 & n930 ) | ( n929 & n930 ) ;
  assign n932 = n291 & n554 ;
  assign n933 = x75 & n295 ;
  assign n934 = x76 | n933 ;
  assign n935 = ( n297 & n933 ) | ( n297 & n934 ) | ( n933 & n934 ) ;
  assign n936 = x74 & n330 ;
  assign n937 = n935 | n936 ;
  assign n938 = ( x8 & n932 ) | ( x8 & ~n937 ) | ( n932 & ~n937 ) ;
  assign n939 = ( ~x8 & n937 ) | ( ~x8 & n938 ) | ( n937 & n938 ) ;
  assign n940 = ( ~n932 & n938 ) | ( ~n932 & n939 ) | ( n938 & n939 ) ;
  assign n941 = n390 & n407 ;
  assign n942 = x72 & n411 ;
  assign n943 = x73 | n942 ;
  assign n944 = ( n413 & n942 ) | ( n413 & n943 ) | ( n942 & n943 ) ;
  assign n945 = x71 & n491 ;
  assign n946 = n944 | n945 ;
  assign n947 = ( x11 & n941 ) | ( x11 & ~n946 ) | ( n941 & ~n946 ) ;
  assign n948 = ( ~x11 & n946 ) | ( ~x11 & n947 ) | ( n946 & n947 ) ;
  assign n949 = ( ~n941 & n947 ) | ( ~n941 & n948 ) | ( n947 & n948 ) ;
  assign n950 = x66 & n814 ;
  assign n951 = x67 | n950 ;
  assign n952 = ( n816 & n950 ) | ( n816 & n951 ) | ( n950 & n951 ) ;
  assign n953 = x65 & n885 ;
  assign n954 = n952 | n953 ;
  assign n955 = n164 & n810 ;
  assign n956 = ( x17 & n954 ) | ( x17 & ~n955 ) | ( n954 & ~n955 ) ;
  assign n957 = ( ~x17 & n955 ) | ( ~x17 & n956 ) | ( n955 & n956 ) ;
  assign n958 = ( ~n954 & n956 ) | ( ~n954 & n957 ) | ( n956 & n957 ) ;
  assign n959 = x17 & x18 ;
  assign n960 = x17 | x18 ;
  assign n961 = ~n959 & n960 ;
  assign n962 = x64 & n961 ;
  assign n963 = x17 & ~n893 ;
  assign n964 = ( n958 & n962 ) | ( n958 & n963 ) | ( n962 & n963 ) ;
  assign n965 = ( ~n958 & n962 ) | ( ~n958 & n963 ) | ( n962 & n963 ) ;
  assign n966 = ( n958 & ~n964 ) | ( n958 & n965 ) | ( ~n964 & n965 ) ;
  assign n967 = n245 & n583 ;
  assign n968 = x69 & n587 ;
  assign n969 = x70 | n968 ;
  assign n970 = ( n589 & n968 ) | ( n589 & n969 ) | ( n968 & n969 ) ;
  assign n971 = x68 & n676 ;
  assign n972 = n970 | n971 ;
  assign n973 = ( x14 & n967 ) | ( x14 & ~n972 ) | ( n967 & ~n972 ) ;
  assign n974 = ( ~x14 & n972 ) | ( ~x14 & n973 ) | ( n972 & n973 ) ;
  assign n975 = ( ~n967 & n973 ) | ( ~n967 & n974 ) | ( n973 & n974 ) ;
  assign n976 = ( n896 & n966 ) | ( n896 & n975 ) | ( n966 & n975 ) ;
  assign n977 = ( ~n896 & n966 ) | ( ~n896 & n975 ) | ( n966 & n975 ) ;
  assign n978 = ( n896 & ~n976 ) | ( n896 & n977 ) | ( ~n976 & n977 ) ;
  assign n979 = ( n899 & n949 ) | ( n899 & n978 ) | ( n949 & n978 ) ;
  assign n980 = ( ~n899 & n949 ) | ( ~n899 & n978 ) | ( n949 & n978 ) ;
  assign n981 = ( n899 & ~n979 ) | ( n899 & n980 ) | ( ~n979 & n980 ) ;
  assign n982 = ( n902 & n940 ) | ( n902 & n981 ) | ( n940 & n981 ) ;
  assign n983 = ( ~n902 & n940 ) | ( ~n902 & n981 ) | ( n940 & n981 ) ;
  assign n984 = ( n902 & ~n982 ) | ( n902 & n983 ) | ( ~n982 & n983 ) ;
  assign n985 = ( n905 & n931 ) | ( n905 & n984 ) | ( n931 & n984 ) ;
  assign n986 = ( ~n905 & n931 ) | ( ~n905 & n984 ) | ( n931 & n984 ) ;
  assign n987 = ( n905 & ~n985 ) | ( n905 & n986 ) | ( ~n985 & n986 ) ;
  assign n988 = ( x81 & x82 ) | ( x81 & n908 ) | ( x82 & n908 ) ;
  assign n989 = ( x81 & ~x82 ) | ( x81 & n908 ) | ( ~x82 & n908 ) ;
  assign n990 = ( x82 & ~n988 ) | ( x82 & n989 ) | ( ~n988 & n989 ) ;
  assign n991 = n136 & n990 ;
  assign n992 = x81 & n138 ;
  assign n993 = x82 | n992 ;
  assign n994 = ( n141 & n992 ) | ( n141 & n993 ) | ( n992 & n993 ) ;
  assign n995 = x80 & n154 ;
  assign n996 = n994 | n995 ;
  assign n997 = ( x2 & n991 ) | ( x2 & ~n996 ) | ( n991 & ~n996 ) ;
  assign n998 = ( ~x2 & n996 ) | ( ~x2 & n997 ) | ( n996 & n997 ) ;
  assign n999 = ( ~n991 & n997 ) | ( ~n991 & n998 ) | ( n997 & n998 ) ;
  assign n1000 = ( n920 & n987 ) | ( n920 & n999 ) | ( n987 & n999 ) ;
  assign n1001 = ( ~n920 & n987 ) | ( ~n920 & n999 ) | ( n987 & n999 ) ;
  assign n1002 = ( n920 & ~n1000 ) | ( n920 & n1001 ) | ( ~n1000 & n1001 ) ;
  assign n1003 = n277 & n583 ;
  assign n1004 = x70 & n587 ;
  assign n1005 = x71 | n1004 ;
  assign n1006 = ( n589 & n1004 ) | ( n589 & n1005 ) | ( n1004 & n1005 ) ;
  assign n1007 = x69 & n676 ;
  assign n1008 = n1006 | n1007 ;
  assign n1009 = ( x14 & n1003 ) | ( x14 & ~n1008 ) | ( n1003 & ~n1008 ) ;
  assign n1010 = ( ~x14 & n1008 ) | ( ~x14 & n1009 ) | ( n1008 & n1009 ) ;
  assign n1011 = ( ~n1003 & n1009 ) | ( ~n1003 & n1010 ) | ( n1009 & n1010 ) ;
  assign n1012 = x20 & n962 ;
  assign n1013 = x19 | x20 ;
  assign n1014 = ( x19 & x20 ) | ( x19 & ~n1013 ) | ( x20 & ~n1013 ) ;
  assign n1015 = n1013 & ~n1014 ;
  assign n1016 = n961 & n1015 ;
  assign n1017 = n133 & n1016 ;
  assign n1018 = ~x17 & x19 ;
  assign n1019 = x18 & x19 ;
  assign n1020 = ( n959 & n1018 ) | ( n959 & ~n1019 ) | ( n1018 & ~n1019 ) ;
  assign n1021 = x64 & n1020 ;
  assign n1022 = ( n961 & ~n1013 ) | ( n961 & n1014 ) | ( ~n1013 & n1014 ) ;
  assign n1023 = x65 | n1021 ;
  assign n1024 = ( n1021 & n1022 ) | ( n1021 & n1023 ) | ( n1022 & n1023 ) ;
  assign n1025 = ( n1012 & n1017 ) | ( n1012 & n1024 ) | ( n1017 & n1024 ) ;
  assign n1026 = n1017 | n1024 ;
  assign n1027 = ~n1012 & n1026 ;
  assign n1028 = ( n1012 & ~n1025 ) | ( n1012 & n1027 ) | ( ~n1025 & n1027 ) ;
  assign n1029 = x67 & n814 ;
  assign n1030 = x68 | n1029 ;
  assign n1031 = ( n816 & n1029 ) | ( n816 & n1030 ) | ( n1029 & n1030 ) ;
  assign n1032 = x66 & n885 ;
  assign n1033 = n1031 | n1032 ;
  assign n1034 = n201 & n810 ;
  assign n1035 = ( x17 & n1033 ) | ( x17 & ~n1034 ) | ( n1033 & ~n1034 ) ;
  assign n1036 = ( ~x17 & n1034 ) | ( ~x17 & n1035 ) | ( n1034 & n1035 ) ;
  assign n1037 = ( ~n1033 & n1035 ) | ( ~n1033 & n1036 ) | ( n1035 & n1036 ) ;
  assign n1038 = ( n964 & n1028 ) | ( n964 & n1037 ) | ( n1028 & n1037 ) ;
  assign n1039 = ( ~n964 & n1028 ) | ( ~n964 & n1037 ) | ( n1028 & n1037 ) ;
  assign n1040 = ( n964 & ~n1038 ) | ( n964 & n1039 ) | ( ~n1038 & n1039 ) ;
  assign n1041 = ( n976 & n1011 ) | ( n976 & n1040 ) | ( n1011 & n1040 ) ;
  assign n1042 = ( ~n976 & n1011 ) | ( ~n976 & n1040 ) | ( n1011 & n1040 ) ;
  assign n1043 = ( n976 & ~n1041 ) | ( n976 & n1042 ) | ( ~n1041 & n1042 ) ;
  assign n1044 = n407 & n446 ;
  assign n1045 = x73 & n411 ;
  assign n1046 = x74 | n1045 ;
  assign n1047 = ( n413 & n1045 ) | ( n413 & n1046 ) | ( n1045 & n1046 ) ;
  assign n1048 = x72 & n491 ;
  assign n1049 = n1047 | n1048 ;
  assign n1050 = ( x11 & n1044 ) | ( x11 & ~n1049 ) | ( n1044 & ~n1049 ) ;
  assign n1051 = ( ~x11 & n1049 ) | ( ~x11 & n1050 ) | ( n1049 & n1050 ) ;
  assign n1052 = ( ~n1044 & n1050 ) | ( ~n1044 & n1051 ) | ( n1050 & n1051 ) ;
  assign n1053 = ( n979 & n1043 ) | ( n979 & n1052 ) | ( n1043 & n1052 ) ;
  assign n1054 = ( ~n979 & n1043 ) | ( ~n979 & n1052 ) | ( n1043 & n1052 ) ;
  assign n1055 = ( n979 & ~n1053 ) | ( n979 & n1054 ) | ( ~n1053 & n1054 ) ;
  assign n1056 = n291 & n569 ;
  assign n1057 = x76 & n295 ;
  assign n1058 = x77 | n1057 ;
  assign n1059 = ( n297 & n1057 ) | ( n297 & n1058 ) | ( n1057 & n1058 ) ;
  assign n1060 = x75 & n330 ;
  assign n1061 = n1059 | n1060 ;
  assign n1062 = ( x8 & n1056 ) | ( x8 & ~n1061 ) | ( n1056 & ~n1061 ) ;
  assign n1063 = ( ~x8 & n1061 ) | ( ~x8 & n1062 ) | ( n1061 & n1062 ) ;
  assign n1064 = ( ~n1056 & n1062 ) | ( ~n1056 & n1063 ) | ( n1062 & n1063 ) ;
  assign n1065 = ( n982 & n1055 ) | ( n982 & n1064 ) | ( n1055 & n1064 ) ;
  assign n1066 = ( n982 & ~n1055 ) | ( n982 & n1064 ) | ( ~n1055 & n1064 ) ;
  assign n1067 = ( n1055 & ~n1065 ) | ( n1055 & n1066 ) | ( ~n1065 & n1066 ) ;
  assign n1068 = n186 & n769 ;
  assign n1069 = x79 & n190 ;
  assign n1070 = x80 | n1069 ;
  assign n1071 = ( n192 & n1069 ) | ( n192 & n1070 ) | ( n1069 & n1070 ) ;
  assign n1072 = x78 & n220 ;
  assign n1073 = n1071 | n1072 ;
  assign n1074 = ( x5 & n1068 ) | ( x5 & ~n1073 ) | ( n1068 & ~n1073 ) ;
  assign n1075 = ( ~x5 & n1073 ) | ( ~x5 & n1074 ) | ( n1073 & n1074 ) ;
  assign n1076 = ( ~n1068 & n1074 ) | ( ~n1068 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1077 = ( n985 & n1067 ) | ( n985 & n1076 ) | ( n1067 & n1076 ) ;
  assign n1078 = ( ~n985 & n1067 ) | ( ~n985 & n1076 ) | ( n1067 & n1076 ) ;
  assign n1079 = ( n985 & ~n1077 ) | ( n985 & n1078 ) | ( ~n1077 & n1078 ) ;
  assign n1080 = ( x82 & x83 ) | ( x82 & n988 ) | ( x83 & n988 ) ;
  assign n1081 = ( x82 & ~x83 ) | ( x82 & n988 ) | ( ~x83 & n988 ) ;
  assign n1082 = ( x83 & ~n1080 ) | ( x83 & n1081 ) | ( ~n1080 & n1081 ) ;
  assign n1083 = n136 & n1082 ;
  assign n1084 = x82 & n138 ;
  assign n1085 = x83 | n1084 ;
  assign n1086 = ( n141 & n1084 ) | ( n141 & n1085 ) | ( n1084 & n1085 ) ;
  assign n1087 = x81 & n154 ;
  assign n1088 = n1086 | n1087 ;
  assign n1089 = ( x2 & n1083 ) | ( x2 & ~n1088 ) | ( n1083 & ~n1088 ) ;
  assign n1090 = ( ~x2 & n1088 ) | ( ~x2 & n1089 ) | ( n1088 & n1089 ) ;
  assign n1091 = ( ~n1083 & n1089 ) | ( ~n1083 & n1090 ) | ( n1089 & n1090 ) ;
  assign n1092 = ( n1000 & n1079 ) | ( n1000 & n1091 ) | ( n1079 & n1091 ) ;
  assign n1093 = ( ~n1000 & n1079 ) | ( ~n1000 & n1091 ) | ( n1079 & n1091 ) ;
  assign n1094 = ( n1000 & ~n1092 ) | ( n1000 & n1093 ) | ( ~n1092 & n1093 ) ;
  assign n1095 = ( x83 & x84 ) | ( x83 & n1080 ) | ( x84 & n1080 ) ;
  assign n1096 = ( x83 & ~x84 ) | ( x83 & n1080 ) | ( ~x84 & n1080 ) ;
  assign n1097 = ( x84 & ~n1095 ) | ( x84 & n1096 ) | ( ~n1095 & n1096 ) ;
  assign n1098 = n136 & n1097 ;
  assign n1099 = x83 & n138 ;
  assign n1100 = x84 | n1099 ;
  assign n1101 = ( n141 & n1099 ) | ( n141 & n1100 ) | ( n1099 & n1100 ) ;
  assign n1102 = x82 & n154 ;
  assign n1103 = n1101 | n1102 ;
  assign n1104 = ( x2 & n1098 ) | ( x2 & ~n1103 ) | ( n1098 & ~n1103 ) ;
  assign n1105 = ( ~x2 & n1103 ) | ( ~x2 & n1104 ) | ( n1103 & n1104 ) ;
  assign n1106 = ( ~n1098 & n1104 ) | ( ~n1098 & n1105 ) | ( n1104 & n1105 ) ;
  assign n1107 = n186 & n910 ;
  assign n1108 = x80 & n190 ;
  assign n1109 = x81 | n1108 ;
  assign n1110 = ( n192 & n1108 ) | ( n192 & n1109 ) | ( n1108 & n1109 ) ;
  assign n1111 = x79 & n220 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = ( x5 & n1107 ) | ( x5 & ~n1112 ) | ( n1107 & ~n1112 ) ;
  assign n1114 = ( ~x5 & n1112 ) | ( ~x5 & n1113 ) | ( n1112 & n1113 ) ;
  assign n1115 = ( ~n1107 & n1113 ) | ( ~n1107 & n1114 ) | ( n1113 & n1114 ) ;
  assign n1116 = n407 & n461 ;
  assign n1117 = x74 & n411 ;
  assign n1118 = x75 | n1117 ;
  assign n1119 = ( n413 & n1117 ) | ( n413 & n1118 ) | ( n1117 & n1118 ) ;
  assign n1120 = x73 & n491 ;
  assign n1121 = n1119 | n1120 ;
  assign n1122 = ( x11 & n1116 ) | ( x11 & ~n1121 ) | ( n1116 & ~n1121 ) ;
  assign n1123 = ( ~x11 & n1121 ) | ( ~x11 & n1122 ) | ( n1121 & n1122 ) ;
  assign n1124 = ( ~n1116 & n1122 ) | ( ~n1116 & n1123 ) | ( n1122 & n1123 ) ;
  assign n1125 = n346 & n583 ;
  assign n1126 = x71 & n587 ;
  assign n1127 = x72 | n1126 ;
  assign n1128 = ( n589 & n1126 ) | ( n589 & n1127 ) | ( n1126 & n1127 ) ;
  assign n1129 = x70 & n676 ;
  assign n1130 = n1128 | n1129 ;
  assign n1131 = ( x14 & n1125 ) | ( x14 & ~n1130 ) | ( n1125 & ~n1130 ) ;
  assign n1132 = ( ~x14 & n1130 ) | ( ~x14 & n1131 ) | ( n1130 & n1131 ) ;
  assign n1133 = ( ~n1125 & n1131 ) | ( ~n1125 & n1132 ) | ( n1131 & n1132 ) ;
  assign n1134 = n230 & n810 ;
  assign n1135 = x68 & n814 ;
  assign n1136 = x69 | n1135 ;
  assign n1137 = ( n816 & n1135 ) | ( n816 & n1136 ) | ( n1135 & n1136 ) ;
  assign n1138 = x67 & n885 ;
  assign n1139 = n1137 | n1138 ;
  assign n1140 = ( ~x17 & n1134 ) | ( ~x17 & n1139 ) | ( n1134 & n1139 ) ;
  assign n1141 = ( n1134 & n1139 ) | ( n1134 & ~n1140 ) | ( n1139 & ~n1140 ) ;
  assign n1142 = ( x17 & n1140 ) | ( x17 & ~n1141 ) | ( n1140 & ~n1141 ) ;
  assign n1143 = ( x20 & n1012 ) | ( x20 & n1026 ) | ( n1012 & n1026 ) ;
  assign n1144 = ( x17 & ~x19 ) | ( x17 & n1015 ) | ( ~x19 & n1015 ) ;
  assign n1145 = ( ~n960 & n1019 ) | ( ~n960 & n1144 ) | ( n1019 & n1144 ) ;
  assign n1146 = x64 & n1145 ;
  assign n1147 = x65 & n1020 ;
  assign n1148 = x66 | n1147 ;
  assign n1149 = ( n1022 & n1147 ) | ( n1022 & n1148 ) | ( n1147 & n1148 ) ;
  assign n1150 = ( n151 & n152 ) | ( n151 & n1016 ) | ( n152 & n1016 ) ;
  assign n1151 = ( ~n1146 & n1149 ) | ( ~n1146 & n1150 ) | ( n1149 & n1150 ) ;
  assign n1152 = n1146 | n1151 ;
  assign n1153 = n1143 | n1152 ;
  assign n1154 = ( n1143 & n1152 ) | ( n1143 & ~n1153 ) | ( n1152 & ~n1153 ) ;
  assign n1155 = n1153 & ~n1154 ;
  assign n1156 = ( n1038 & n1142 ) | ( n1038 & n1155 ) | ( n1142 & n1155 ) ;
  assign n1157 = ( ~n1038 & n1142 ) | ( ~n1038 & n1155 ) | ( n1142 & n1155 ) ;
  assign n1158 = ( n1038 & ~n1156 ) | ( n1038 & n1157 ) | ( ~n1156 & n1157 ) ;
  assign n1159 = ( n1041 & n1133 ) | ( n1041 & n1158 ) | ( n1133 & n1158 ) ;
  assign n1160 = ( ~n1041 & n1133 ) | ( ~n1041 & n1158 ) | ( n1133 & n1158 ) ;
  assign n1161 = ( n1041 & ~n1159 ) | ( n1041 & n1160 ) | ( ~n1159 & n1160 ) ;
  assign n1162 = ( n1053 & n1124 ) | ( n1053 & n1161 ) | ( n1124 & n1161 ) ;
  assign n1163 = ( ~n1053 & n1124 ) | ( ~n1053 & n1161 ) | ( n1124 & n1161 ) ;
  assign n1164 = ( n1053 & ~n1162 ) | ( n1053 & n1163 ) | ( ~n1162 & n1163 ) ;
  assign n1165 = n291 & n637 ;
  assign n1166 = x77 & n295 ;
  assign n1167 = x78 | n1166 ;
  assign n1168 = ( n297 & n1166 ) | ( n297 & n1167 ) | ( n1166 & n1167 ) ;
  assign n1169 = x76 & n330 ;
  assign n1170 = n1168 | n1169 ;
  assign n1171 = ( x8 & n1165 ) | ( x8 & ~n1170 ) | ( n1165 & ~n1170 ) ;
  assign n1172 = ( ~x8 & n1170 ) | ( ~x8 & n1171 ) | ( n1170 & n1171 ) ;
  assign n1173 = ( ~n1165 & n1171 ) | ( ~n1165 & n1172 ) | ( n1171 & n1172 ) ;
  assign n1174 = ( n1065 & n1164 ) | ( n1065 & n1173 ) | ( n1164 & n1173 ) ;
  assign n1175 = ( ~n1065 & n1164 ) | ( ~n1065 & n1173 ) | ( n1164 & n1173 ) ;
  assign n1176 = ( n1065 & ~n1174 ) | ( n1065 & n1175 ) | ( ~n1174 & n1175 ) ;
  assign n1177 = ( n1077 & n1115 ) | ( n1077 & n1176 ) | ( n1115 & n1176 ) ;
  assign n1178 = ( ~n1077 & n1115 ) | ( ~n1077 & n1176 ) | ( n1115 & n1176 ) ;
  assign n1179 = ( n1077 & ~n1177 ) | ( n1077 & n1178 ) | ( ~n1177 & n1178 ) ;
  assign n1180 = ( n1092 & n1106 ) | ( n1092 & n1179 ) | ( n1106 & n1179 ) ;
  assign n1181 = ( ~n1092 & n1106 ) | ( ~n1092 & n1179 ) | ( n1106 & n1179 ) ;
  assign n1182 = ( n1092 & ~n1180 ) | ( n1092 & n1181 ) | ( ~n1180 & n1181 ) ;
  assign n1183 = n291 & n701 ;
  assign n1184 = x78 & n295 ;
  assign n1185 = x79 | n1184 ;
  assign n1186 = ( n297 & n1184 ) | ( n297 & n1185 ) | ( n1184 & n1185 ) ;
  assign n1187 = x77 & n330 ;
  assign n1188 = n1186 | n1187 ;
  assign n1189 = ( x8 & n1183 ) | ( x8 & ~n1188 ) | ( n1183 & ~n1188 ) ;
  assign n1190 = ( ~x8 & n1188 ) | ( ~x8 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1191 = ( ~n1183 & n1189 ) | ( ~n1183 & n1190 ) | ( n1189 & n1190 ) ;
  assign n1192 = n407 & n554 ;
  assign n1193 = x75 & n411 ;
  assign n1194 = x76 | n1193 ;
  assign n1195 = ( n413 & n1193 ) | ( n413 & n1194 ) | ( n1193 & n1194 ) ;
  assign n1196 = x74 & n491 ;
  assign n1197 = n1195 | n1196 ;
  assign n1198 = ( x11 & n1192 ) | ( x11 & ~n1197 ) | ( n1192 & ~n1197 ) ;
  assign n1199 = ( ~x11 & n1197 ) | ( ~x11 & n1198 ) | ( n1197 & n1198 ) ;
  assign n1200 = ( ~n1192 & n1198 ) | ( ~n1192 & n1199 ) | ( n1198 & n1199 ) ;
  assign n1201 = n390 & n583 ;
  assign n1202 = x72 & n587 ;
  assign n1203 = x73 | n1202 ;
  assign n1204 = ( n589 & n1202 ) | ( n589 & n1203 ) | ( n1202 & n1203 ) ;
  assign n1205 = x71 & n676 ;
  assign n1206 = n1204 | n1205 ;
  assign n1207 = ( x14 & n1201 ) | ( x14 & ~n1206 ) | ( n1201 & ~n1206 ) ;
  assign n1208 = ( ~x14 & n1206 ) | ( ~x14 & n1207 ) | ( n1206 & n1207 ) ;
  assign n1209 = ( ~n1201 & n1207 ) | ( ~n1201 & n1208 ) | ( n1207 & n1208 ) ;
  assign n1210 = x66 & n1020 ;
  assign n1211 = x67 | n1210 ;
  assign n1212 = ( n1022 & n1210 ) | ( n1022 & n1211 ) | ( n1210 & n1211 ) ;
  assign n1213 = x65 & n1145 ;
  assign n1214 = n1212 | n1213 ;
  assign n1215 = n164 & n1016 ;
  assign n1216 = ( x20 & n1214 ) | ( x20 & ~n1215 ) | ( n1214 & ~n1215 ) ;
  assign n1217 = ( ~x20 & n1215 ) | ( ~x20 & n1216 ) | ( n1215 & n1216 ) ;
  assign n1218 = ( ~n1214 & n1216 ) | ( ~n1214 & n1217 ) | ( n1216 & n1217 ) ;
  assign n1219 = x20 & x21 ;
  assign n1220 = x20 | x21 ;
  assign n1221 = ~n1219 & n1220 ;
  assign n1222 = x64 & n1221 ;
  assign n1223 = x20 & ~n1153 ;
  assign n1224 = ( n1218 & n1222 ) | ( n1218 & n1223 ) | ( n1222 & n1223 ) ;
  assign n1225 = ( ~n1218 & n1222 ) | ( ~n1218 & n1223 ) | ( n1222 & n1223 ) ;
  assign n1226 = ( n1218 & ~n1224 ) | ( n1218 & n1225 ) | ( ~n1224 & n1225 ) ;
  assign n1227 = n245 & n810 ;
  assign n1228 = x69 & n814 ;
  assign n1229 = x70 | n1228 ;
  assign n1230 = ( n816 & n1228 ) | ( n816 & n1229 ) | ( n1228 & n1229 ) ;
  assign n1231 = x68 & n885 ;
  assign n1232 = n1230 | n1231 ;
  assign n1233 = ( x17 & n1227 ) | ( x17 & ~n1232 ) | ( n1227 & ~n1232 ) ;
  assign n1234 = ( ~x17 & n1232 ) | ( ~x17 & n1233 ) | ( n1232 & n1233 ) ;
  assign n1235 = ( ~n1227 & n1233 ) | ( ~n1227 & n1234 ) | ( n1233 & n1234 ) ;
  assign n1236 = ( n1156 & n1226 ) | ( n1156 & n1235 ) | ( n1226 & n1235 ) ;
  assign n1237 = ( ~n1156 & n1226 ) | ( ~n1156 & n1235 ) | ( n1226 & n1235 ) ;
  assign n1238 = ( n1156 & ~n1236 ) | ( n1156 & n1237 ) | ( ~n1236 & n1237 ) ;
  assign n1239 = ( n1159 & n1209 ) | ( n1159 & n1238 ) | ( n1209 & n1238 ) ;
  assign n1240 = ( ~n1159 & n1209 ) | ( ~n1159 & n1238 ) | ( n1209 & n1238 ) ;
  assign n1241 = ( n1159 & ~n1239 ) | ( n1159 & n1240 ) | ( ~n1239 & n1240 ) ;
  assign n1242 = ( n1162 & n1200 ) | ( n1162 & n1241 ) | ( n1200 & n1241 ) ;
  assign n1243 = ( ~n1162 & n1200 ) | ( ~n1162 & n1241 ) | ( n1200 & n1241 ) ;
  assign n1244 = ( n1162 & ~n1242 ) | ( n1162 & n1243 ) | ( ~n1242 & n1243 ) ;
  assign n1245 = ( n1174 & n1191 ) | ( n1174 & n1244 ) | ( n1191 & n1244 ) ;
  assign n1246 = ( ~n1174 & n1191 ) | ( ~n1174 & n1244 ) | ( n1191 & n1244 ) ;
  assign n1247 = ( n1174 & ~n1245 ) | ( n1174 & n1246 ) | ( ~n1245 & n1246 ) ;
  assign n1248 = n186 & n990 ;
  assign n1249 = x81 & n190 ;
  assign n1250 = x82 | n1249 ;
  assign n1251 = ( n192 & n1249 ) | ( n192 & n1250 ) | ( n1249 & n1250 ) ;
  assign n1252 = x80 & n220 ;
  assign n1253 = n1251 | n1252 ;
  assign n1254 = ( x5 & n1248 ) | ( x5 & ~n1253 ) | ( n1248 & ~n1253 ) ;
  assign n1255 = ( ~x5 & n1253 ) | ( ~x5 & n1254 ) | ( n1253 & n1254 ) ;
  assign n1256 = ( ~n1248 & n1254 ) | ( ~n1248 & n1255 ) | ( n1254 & n1255 ) ;
  assign n1257 = ( n1177 & n1247 ) | ( n1177 & n1256 ) | ( n1247 & n1256 ) ;
  assign n1258 = ( ~n1177 & n1247 ) | ( ~n1177 & n1256 ) | ( n1247 & n1256 ) ;
  assign n1259 = ( n1177 & ~n1257 ) | ( n1177 & n1258 ) | ( ~n1257 & n1258 ) ;
  assign n1260 = ( x84 & x85 ) | ( x84 & n1095 ) | ( x85 & n1095 ) ;
  assign n1261 = ( x84 & ~x85 ) | ( x84 & n1095 ) | ( ~x85 & n1095 ) ;
  assign n1262 = ( x85 & ~n1260 ) | ( x85 & n1261 ) | ( ~n1260 & n1261 ) ;
  assign n1263 = n136 & n1262 ;
  assign n1264 = x84 & n138 ;
  assign n1265 = x85 | n1264 ;
  assign n1266 = ( n141 & n1264 ) | ( n141 & n1265 ) | ( n1264 & n1265 ) ;
  assign n1267 = x83 & n154 ;
  assign n1268 = n1266 | n1267 ;
  assign n1269 = ( x2 & n1263 ) | ( x2 & ~n1268 ) | ( n1263 & ~n1268 ) ;
  assign n1270 = ( ~x2 & n1268 ) | ( ~x2 & n1269 ) | ( n1268 & n1269 ) ;
  assign n1271 = ( ~n1263 & n1269 ) | ( ~n1263 & n1270 ) | ( n1269 & n1270 ) ;
  assign n1272 = ( n1180 & n1259 ) | ( n1180 & n1271 ) | ( n1259 & n1271 ) ;
  assign n1273 = ( ~n1180 & n1259 ) | ( ~n1180 & n1271 ) | ( n1259 & n1271 ) ;
  assign n1274 = ( n1180 & ~n1272 ) | ( n1180 & n1273 ) | ( ~n1272 & n1273 ) ;
  assign n1275 = n291 & n769 ;
  assign n1276 = x79 & n295 ;
  assign n1277 = x80 | n1276 ;
  assign n1278 = ( n297 & n1276 ) | ( n297 & n1277 ) | ( n1276 & n1277 ) ;
  assign n1279 = x78 & n330 ;
  assign n1280 = n1278 | n1279 ;
  assign n1281 = ( x8 & n1275 ) | ( x8 & ~n1280 ) | ( n1275 & ~n1280 ) ;
  assign n1282 = ( ~x8 & n1280 ) | ( ~x8 & n1281 ) | ( n1280 & n1281 ) ;
  assign n1283 = ( ~n1275 & n1281 ) | ( ~n1275 & n1282 ) | ( n1281 & n1282 ) ;
  assign n1284 = n277 & n810 ;
  assign n1285 = x70 & n814 ;
  assign n1286 = x71 | n1285 ;
  assign n1287 = ( n816 & n1285 ) | ( n816 & n1286 ) | ( n1285 & n1286 ) ;
  assign n1288 = x69 & n885 ;
  assign n1289 = n1287 | n1288 ;
  assign n1290 = ( x17 & n1284 ) | ( x17 & ~n1289 ) | ( n1284 & ~n1289 ) ;
  assign n1291 = ( ~x17 & n1289 ) | ( ~x17 & n1290 ) | ( n1289 & n1290 ) ;
  assign n1292 = ( ~n1284 & n1290 ) | ( ~n1284 & n1291 ) | ( n1290 & n1291 ) ;
  assign n1293 = x23 & n1222 ;
  assign n1294 = x22 | x23 ;
  assign n1295 = ( x22 & x23 ) | ( x22 & ~n1294 ) | ( x23 & ~n1294 ) ;
  assign n1296 = n1294 & ~n1295 ;
  assign n1297 = n1221 & n1296 ;
  assign n1298 = n133 & n1297 ;
  assign n1299 = ~x20 & x22 ;
  assign n1300 = x21 & x22 ;
  assign n1301 = ( n1219 & n1299 ) | ( n1219 & ~n1300 ) | ( n1299 & ~n1300 ) ;
  assign n1302 = x64 & n1301 ;
  assign n1303 = ( n1221 & ~n1294 ) | ( n1221 & n1295 ) | ( ~n1294 & n1295 ) ;
  assign n1304 = x65 | n1302 ;
  assign n1305 = ( n1302 & n1303 ) | ( n1302 & n1304 ) | ( n1303 & n1304 ) ;
  assign n1306 = ( n1293 & n1298 ) | ( n1293 & n1305 ) | ( n1298 & n1305 ) ;
  assign n1307 = n1298 | n1305 ;
  assign n1308 = ~n1293 & n1307 ;
  assign n1309 = ( n1293 & ~n1306 ) | ( n1293 & n1308 ) | ( ~n1306 & n1308 ) ;
  assign n1310 = x67 & n1020 ;
  assign n1311 = x68 | n1310 ;
  assign n1312 = ( n1022 & n1310 ) | ( n1022 & n1311 ) | ( n1310 & n1311 ) ;
  assign n1313 = x66 & n1145 ;
  assign n1314 = n1312 | n1313 ;
  assign n1315 = n201 & n1016 ;
  assign n1316 = ( x20 & n1314 ) | ( x20 & ~n1315 ) | ( n1314 & ~n1315 ) ;
  assign n1317 = ( ~x20 & n1315 ) | ( ~x20 & n1316 ) | ( n1315 & n1316 ) ;
  assign n1318 = ( ~n1314 & n1316 ) | ( ~n1314 & n1317 ) | ( n1316 & n1317 ) ;
  assign n1319 = ( n1224 & n1309 ) | ( n1224 & n1318 ) | ( n1309 & n1318 ) ;
  assign n1320 = ( ~n1224 & n1309 ) | ( ~n1224 & n1318 ) | ( n1309 & n1318 ) ;
  assign n1321 = ( n1224 & ~n1319 ) | ( n1224 & n1320 ) | ( ~n1319 & n1320 ) ;
  assign n1322 = ( n1236 & n1292 ) | ( n1236 & n1321 ) | ( n1292 & n1321 ) ;
  assign n1323 = ( ~n1236 & n1292 ) | ( ~n1236 & n1321 ) | ( n1292 & n1321 ) ;
  assign n1324 = ( n1236 & ~n1322 ) | ( n1236 & n1323 ) | ( ~n1322 & n1323 ) ;
  assign n1325 = n446 & n583 ;
  assign n1326 = x73 & n587 ;
  assign n1327 = x74 | n1326 ;
  assign n1328 = ( n589 & n1326 ) | ( n589 & n1327 ) | ( n1326 & n1327 ) ;
  assign n1329 = x72 & n676 ;
  assign n1330 = n1328 | n1329 ;
  assign n1331 = ( x14 & n1325 ) | ( x14 & ~n1330 ) | ( n1325 & ~n1330 ) ;
  assign n1332 = ( ~x14 & n1330 ) | ( ~x14 & n1331 ) | ( n1330 & n1331 ) ;
  assign n1333 = ( ~n1325 & n1331 ) | ( ~n1325 & n1332 ) | ( n1331 & n1332 ) ;
  assign n1334 = ( n1239 & n1324 ) | ( n1239 & n1333 ) | ( n1324 & n1333 ) ;
  assign n1335 = ( ~n1239 & n1324 ) | ( ~n1239 & n1333 ) | ( n1324 & n1333 ) ;
  assign n1336 = ( n1239 & ~n1334 ) | ( n1239 & n1335 ) | ( ~n1334 & n1335 ) ;
  assign n1337 = n407 & n569 ;
  assign n1338 = x76 & n411 ;
  assign n1339 = x77 | n1338 ;
  assign n1340 = ( n413 & n1338 ) | ( n413 & n1339 ) | ( n1338 & n1339 ) ;
  assign n1341 = x75 & n491 ;
  assign n1342 = n1340 | n1341 ;
  assign n1343 = ( x11 & n1337 ) | ( x11 & ~n1342 ) | ( n1337 & ~n1342 ) ;
  assign n1344 = ( ~x11 & n1342 ) | ( ~x11 & n1343 ) | ( n1342 & n1343 ) ;
  assign n1345 = ( ~n1337 & n1343 ) | ( ~n1337 & n1344 ) | ( n1343 & n1344 ) ;
  assign n1346 = ( n1242 & n1336 ) | ( n1242 & n1345 ) | ( n1336 & n1345 ) ;
  assign n1347 = ( ~n1242 & n1336 ) | ( ~n1242 & n1345 ) | ( n1336 & n1345 ) ;
  assign n1348 = ( n1242 & ~n1346 ) | ( n1242 & n1347 ) | ( ~n1346 & n1347 ) ;
  assign n1349 = ( n1245 & n1283 ) | ( n1245 & n1348 ) | ( n1283 & n1348 ) ;
  assign n1350 = ( ~n1245 & n1283 ) | ( ~n1245 & n1348 ) | ( n1283 & n1348 ) ;
  assign n1351 = ( n1245 & ~n1349 ) | ( n1245 & n1350 ) | ( ~n1349 & n1350 ) ;
  assign n1352 = n186 & n1082 ;
  assign n1353 = x82 & n190 ;
  assign n1354 = x83 | n1353 ;
  assign n1355 = ( n192 & n1353 ) | ( n192 & n1354 ) | ( n1353 & n1354 ) ;
  assign n1356 = x81 & n220 ;
  assign n1357 = n1355 | n1356 ;
  assign n1358 = ( x5 & n1352 ) | ( x5 & ~n1357 ) | ( n1352 & ~n1357 ) ;
  assign n1359 = ( ~x5 & n1357 ) | ( ~x5 & n1358 ) | ( n1357 & n1358 ) ;
  assign n1360 = ( ~n1352 & n1358 ) | ( ~n1352 & n1359 ) | ( n1358 & n1359 ) ;
  assign n1361 = ( n1257 & n1351 ) | ( n1257 & n1360 ) | ( n1351 & n1360 ) ;
  assign n1362 = ( ~n1257 & n1351 ) | ( ~n1257 & n1360 ) | ( n1351 & n1360 ) ;
  assign n1363 = ( n1257 & ~n1361 ) | ( n1257 & n1362 ) | ( ~n1361 & n1362 ) ;
  assign n1364 = ( x85 & x86 ) | ( x85 & n1260 ) | ( x86 & n1260 ) ;
  assign n1365 = ( x85 & ~x86 ) | ( x85 & n1260 ) | ( ~x86 & n1260 ) ;
  assign n1366 = ( x86 & ~n1364 ) | ( x86 & n1365 ) | ( ~n1364 & n1365 ) ;
  assign n1367 = n136 & n1366 ;
  assign n1368 = x85 & n138 ;
  assign n1369 = x86 | n1368 ;
  assign n1370 = ( n141 & n1368 ) | ( n141 & n1369 ) | ( n1368 & n1369 ) ;
  assign n1371 = x84 & n154 ;
  assign n1372 = n1370 | n1371 ;
  assign n1373 = ( x2 & n1367 ) | ( x2 & ~n1372 ) | ( n1367 & ~n1372 ) ;
  assign n1374 = ( ~x2 & n1372 ) | ( ~x2 & n1373 ) | ( n1372 & n1373 ) ;
  assign n1375 = ( ~n1367 & n1373 ) | ( ~n1367 & n1374 ) | ( n1373 & n1374 ) ;
  assign n1376 = ( n1272 & n1363 ) | ( n1272 & n1375 ) | ( n1363 & n1375 ) ;
  assign n1377 = ( ~n1272 & n1363 ) | ( ~n1272 & n1375 ) | ( n1363 & n1375 ) ;
  assign n1378 = ( n1272 & ~n1376 ) | ( n1272 & n1377 ) | ( ~n1376 & n1377 ) ;
  assign n1379 = n186 & n1097 ;
  assign n1380 = x83 & n190 ;
  assign n1381 = x84 | n1380 ;
  assign n1382 = ( n192 & n1380 ) | ( n192 & n1381 ) | ( n1380 & n1381 ) ;
  assign n1383 = x82 & n220 ;
  assign n1384 = n1382 | n1383 ;
  assign n1385 = ( x5 & n1379 ) | ( x5 & ~n1384 ) | ( n1379 & ~n1384 ) ;
  assign n1386 = ( ~x5 & n1384 ) | ( ~x5 & n1385 ) | ( n1384 & n1385 ) ;
  assign n1387 = ( ~n1379 & n1385 ) | ( ~n1379 & n1386 ) | ( n1385 & n1386 ) ;
  assign n1388 = n291 & n910 ;
  assign n1389 = x80 & n295 ;
  assign n1390 = x81 | n1389 ;
  assign n1391 = ( n297 & n1389 ) | ( n297 & n1390 ) | ( n1389 & n1390 ) ;
  assign n1392 = x79 & n330 ;
  assign n1393 = n1391 | n1392 ;
  assign n1394 = ( x8 & n1388 ) | ( x8 & ~n1393 ) | ( n1388 & ~n1393 ) ;
  assign n1395 = ( ~x8 & n1393 ) | ( ~x8 & n1394 ) | ( n1393 & n1394 ) ;
  assign n1396 = ( ~n1388 & n1394 ) | ( ~n1388 & n1395 ) | ( n1394 & n1395 ) ;
  assign n1397 = n461 & n583 ;
  assign n1398 = x74 & n587 ;
  assign n1399 = x75 | n1398 ;
  assign n1400 = ( n589 & n1398 ) | ( n589 & n1399 ) | ( n1398 & n1399 ) ;
  assign n1401 = x73 & n676 ;
  assign n1402 = n1400 | n1401 ;
  assign n1403 = ( x14 & n1397 ) | ( x14 & ~n1402 ) | ( n1397 & ~n1402 ) ;
  assign n1404 = ( ~x14 & n1402 ) | ( ~x14 & n1403 ) | ( n1402 & n1403 ) ;
  assign n1405 = ( ~n1397 & n1403 ) | ( ~n1397 & n1404 ) | ( n1403 & n1404 ) ;
  assign n1406 = n346 & n810 ;
  assign n1407 = x71 & n814 ;
  assign n1408 = x72 | n1407 ;
  assign n1409 = ( n816 & n1407 ) | ( n816 & n1408 ) | ( n1407 & n1408 ) ;
  assign n1410 = x70 & n885 ;
  assign n1411 = n1409 | n1410 ;
  assign n1412 = ( x17 & n1406 ) | ( x17 & ~n1411 ) | ( n1406 & ~n1411 ) ;
  assign n1413 = ( ~x17 & n1411 ) | ( ~x17 & n1412 ) | ( n1411 & n1412 ) ;
  assign n1414 = ( ~n1406 & n1412 ) | ( ~n1406 & n1413 ) | ( n1412 & n1413 ) ;
  assign n1415 = n230 & n1016 ;
  assign n1416 = x68 & n1020 ;
  assign n1417 = x69 | n1416 ;
  assign n1418 = ( n1022 & n1416 ) | ( n1022 & n1417 ) | ( n1416 & n1417 ) ;
  assign n1419 = x67 & n1145 ;
  assign n1420 = n1418 | n1419 ;
  assign n1421 = ( ~x20 & n1415 ) | ( ~x20 & n1420 ) | ( n1415 & n1420 ) ;
  assign n1422 = ( n1415 & n1420 ) | ( n1415 & ~n1421 ) | ( n1420 & ~n1421 ) ;
  assign n1423 = ( x20 & n1421 ) | ( x20 & ~n1422 ) | ( n1421 & ~n1422 ) ;
  assign n1424 = ( x23 & n1293 ) | ( x23 & n1307 ) | ( n1293 & n1307 ) ;
  assign n1425 = ( x20 & ~x22 ) | ( x20 & n1296 ) | ( ~x22 & n1296 ) ;
  assign n1426 = ( ~n1220 & n1300 ) | ( ~n1220 & n1425 ) | ( n1300 & n1425 ) ;
  assign n1427 = x64 & n1426 ;
  assign n1428 = x65 & n1301 ;
  assign n1429 = x66 | n1428 ;
  assign n1430 = ( n1303 & n1428 ) | ( n1303 & n1429 ) | ( n1428 & n1429 ) ;
  assign n1431 = ( n151 & n152 ) | ( n151 & n1297 ) | ( n152 & n1297 ) ;
  assign n1432 = ( ~n1427 & n1430 ) | ( ~n1427 & n1431 ) | ( n1430 & n1431 ) ;
  assign n1433 = n1427 | n1432 ;
  assign n1434 = n1424 | n1433 ;
  assign n1435 = ( n1424 & n1433 ) | ( n1424 & ~n1434 ) | ( n1433 & ~n1434 ) ;
  assign n1436 = n1434 & ~n1435 ;
  assign n1437 = ( n1319 & n1423 ) | ( n1319 & n1436 ) | ( n1423 & n1436 ) ;
  assign n1438 = ( ~n1319 & n1423 ) | ( ~n1319 & n1436 ) | ( n1423 & n1436 ) ;
  assign n1439 = ( n1319 & ~n1437 ) | ( n1319 & n1438 ) | ( ~n1437 & n1438 ) ;
  assign n1440 = ( n1322 & n1414 ) | ( n1322 & n1439 ) | ( n1414 & n1439 ) ;
  assign n1441 = ( ~n1322 & n1414 ) | ( ~n1322 & n1439 ) | ( n1414 & n1439 ) ;
  assign n1442 = ( n1322 & ~n1440 ) | ( n1322 & n1441 ) | ( ~n1440 & n1441 ) ;
  assign n1443 = ( n1334 & n1405 ) | ( n1334 & n1442 ) | ( n1405 & n1442 ) ;
  assign n1444 = ( ~n1334 & n1405 ) | ( ~n1334 & n1442 ) | ( n1405 & n1442 ) ;
  assign n1445 = ( n1334 & ~n1443 ) | ( n1334 & n1444 ) | ( ~n1443 & n1444 ) ;
  assign n1446 = n407 & n637 ;
  assign n1447 = x77 & n411 ;
  assign n1448 = x78 | n1447 ;
  assign n1449 = ( n413 & n1447 ) | ( n413 & n1448 ) | ( n1447 & n1448 ) ;
  assign n1450 = x76 & n491 ;
  assign n1451 = n1449 | n1450 ;
  assign n1452 = ( x11 & n1446 ) | ( x11 & ~n1451 ) | ( n1446 & ~n1451 ) ;
  assign n1453 = ( ~x11 & n1451 ) | ( ~x11 & n1452 ) | ( n1451 & n1452 ) ;
  assign n1454 = ( ~n1446 & n1452 ) | ( ~n1446 & n1453 ) | ( n1452 & n1453 ) ;
  assign n1455 = ( n1346 & n1445 ) | ( n1346 & n1454 ) | ( n1445 & n1454 ) ;
  assign n1456 = ( ~n1346 & n1445 ) | ( ~n1346 & n1454 ) | ( n1445 & n1454 ) ;
  assign n1457 = ( n1346 & ~n1455 ) | ( n1346 & n1456 ) | ( ~n1455 & n1456 ) ;
  assign n1458 = ( n1349 & n1396 ) | ( n1349 & n1457 ) | ( n1396 & n1457 ) ;
  assign n1459 = ( ~n1349 & n1396 ) | ( ~n1349 & n1457 ) | ( n1396 & n1457 ) ;
  assign n1460 = ( n1349 & ~n1458 ) | ( n1349 & n1459 ) | ( ~n1458 & n1459 ) ;
  assign n1461 = ( n1361 & n1387 ) | ( n1361 & n1460 ) | ( n1387 & n1460 ) ;
  assign n1462 = ( ~n1361 & n1387 ) | ( ~n1361 & n1460 ) | ( n1387 & n1460 ) ;
  assign n1463 = ( n1361 & ~n1461 ) | ( n1361 & n1462 ) | ( ~n1461 & n1462 ) ;
  assign n1464 = ( x86 & x87 ) | ( x86 & n1364 ) | ( x87 & n1364 ) ;
  assign n1465 = ( x86 & ~x87 ) | ( x86 & n1364 ) | ( ~x87 & n1364 ) ;
  assign n1466 = ( x87 & ~n1464 ) | ( x87 & n1465 ) | ( ~n1464 & n1465 ) ;
  assign n1467 = n136 & n1466 ;
  assign n1468 = x86 & n138 ;
  assign n1469 = x87 | n1468 ;
  assign n1470 = ( n141 & n1468 ) | ( n141 & n1469 ) | ( n1468 & n1469 ) ;
  assign n1471 = x85 & n154 ;
  assign n1472 = n1470 | n1471 ;
  assign n1473 = ( x2 & n1467 ) | ( x2 & ~n1472 ) | ( n1467 & ~n1472 ) ;
  assign n1474 = ( ~x2 & n1472 ) | ( ~x2 & n1473 ) | ( n1472 & n1473 ) ;
  assign n1475 = ( ~n1467 & n1473 ) | ( ~n1467 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1476 = ( n1376 & n1463 ) | ( n1376 & n1475 ) | ( n1463 & n1475 ) ;
  assign n1477 = ( ~n1376 & n1463 ) | ( ~n1376 & n1475 ) | ( n1463 & n1475 ) ;
  assign n1478 = ( n1376 & ~n1476 ) | ( n1376 & n1477 ) | ( ~n1476 & n1477 ) ;
  assign n1479 = ( x87 & x88 ) | ( x87 & n1464 ) | ( x88 & n1464 ) ;
  assign n1480 = ( x87 & ~x88 ) | ( x87 & n1464 ) | ( ~x88 & n1464 ) ;
  assign n1481 = ( x88 & ~n1479 ) | ( x88 & n1480 ) | ( ~n1479 & n1480 ) ;
  assign n1482 = n136 & n1481 ;
  assign n1483 = x87 & n138 ;
  assign n1484 = x88 | n1483 ;
  assign n1485 = ( n141 & n1483 ) | ( n141 & n1484 ) | ( n1483 & n1484 ) ;
  assign n1486 = x86 & n154 ;
  assign n1487 = n1485 | n1486 ;
  assign n1488 = ( x2 & n1482 ) | ( x2 & ~n1487 ) | ( n1482 & ~n1487 ) ;
  assign n1489 = ( ~x2 & n1487 ) | ( ~x2 & n1488 ) | ( n1487 & n1488 ) ;
  assign n1490 = ( ~n1482 & n1488 ) | ( ~n1482 & n1489 ) | ( n1488 & n1489 ) ;
  assign n1491 = n186 & n1262 ;
  assign n1492 = x84 & n190 ;
  assign n1493 = x85 | n1492 ;
  assign n1494 = ( n192 & n1492 ) | ( n192 & n1493 ) | ( n1492 & n1493 ) ;
  assign n1495 = x83 & n220 ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = ( x5 & n1491 ) | ( x5 & ~n1496 ) | ( n1491 & ~n1496 ) ;
  assign n1498 = ( ~x5 & n1496 ) | ( ~x5 & n1497 ) | ( n1496 & n1497 ) ;
  assign n1499 = ( ~n1491 & n1497 ) | ( ~n1491 & n1498 ) | ( n1497 & n1498 ) ;
  assign n1500 = n554 & n583 ;
  assign n1501 = x75 & n587 ;
  assign n1502 = x76 | n1501 ;
  assign n1503 = ( n589 & n1501 ) | ( n589 & n1502 ) | ( n1501 & n1502 ) ;
  assign n1504 = x74 & n676 ;
  assign n1505 = n1503 | n1504 ;
  assign n1506 = ( x14 & n1500 ) | ( x14 & ~n1505 ) | ( n1500 & ~n1505 ) ;
  assign n1507 = ( ~x14 & n1505 ) | ( ~x14 & n1506 ) | ( n1505 & n1506 ) ;
  assign n1508 = ( ~n1500 & n1506 ) | ( ~n1500 & n1507 ) | ( n1506 & n1507 ) ;
  assign n1509 = n390 & n810 ;
  assign n1510 = x72 & n814 ;
  assign n1511 = x73 | n1510 ;
  assign n1512 = ( n816 & n1510 ) | ( n816 & n1511 ) | ( n1510 & n1511 ) ;
  assign n1513 = x71 & n885 ;
  assign n1514 = n1512 | n1513 ;
  assign n1515 = ( x17 & n1509 ) | ( x17 & ~n1514 ) | ( n1509 & ~n1514 ) ;
  assign n1516 = ( ~x17 & n1514 ) | ( ~x17 & n1515 ) | ( n1514 & n1515 ) ;
  assign n1517 = ( ~n1509 & n1515 ) | ( ~n1509 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1518 = x66 & n1301 ;
  assign n1519 = x67 | n1518 ;
  assign n1520 = ( n1303 & n1518 ) | ( n1303 & n1519 ) | ( n1518 & n1519 ) ;
  assign n1521 = x65 & n1426 ;
  assign n1522 = n1520 | n1521 ;
  assign n1523 = n164 & n1297 ;
  assign n1524 = ( x23 & n1522 ) | ( x23 & ~n1523 ) | ( n1522 & ~n1523 ) ;
  assign n1525 = ( ~x23 & n1523 ) | ( ~x23 & n1524 ) | ( n1523 & n1524 ) ;
  assign n1526 = ( ~n1522 & n1524 ) | ( ~n1522 & n1525 ) | ( n1524 & n1525 ) ;
  assign n1527 = x23 & x24 ;
  assign n1528 = x23 | x24 ;
  assign n1529 = ~n1527 & n1528 ;
  assign n1530 = x64 & n1529 ;
  assign n1531 = x23 & ~n1434 ;
  assign n1532 = ( n1526 & n1530 ) | ( n1526 & n1531 ) | ( n1530 & n1531 ) ;
  assign n1533 = ( ~n1526 & n1530 ) | ( ~n1526 & n1531 ) | ( n1530 & n1531 ) ;
  assign n1534 = ( n1526 & ~n1532 ) | ( n1526 & n1533 ) | ( ~n1532 & n1533 ) ;
  assign n1535 = n245 & n1016 ;
  assign n1536 = x69 & n1020 ;
  assign n1537 = x70 | n1536 ;
  assign n1538 = ( n1022 & n1536 ) | ( n1022 & n1537 ) | ( n1536 & n1537 ) ;
  assign n1539 = x68 & n1145 ;
  assign n1540 = n1538 | n1539 ;
  assign n1541 = ( x20 & n1535 ) | ( x20 & ~n1540 ) | ( n1535 & ~n1540 ) ;
  assign n1542 = ( ~x20 & n1540 ) | ( ~x20 & n1541 ) | ( n1540 & n1541 ) ;
  assign n1543 = ( ~n1535 & n1541 ) | ( ~n1535 & n1542 ) | ( n1541 & n1542 ) ;
  assign n1544 = ( n1437 & n1534 ) | ( n1437 & n1543 ) | ( n1534 & n1543 ) ;
  assign n1545 = ( ~n1437 & n1534 ) | ( ~n1437 & n1543 ) | ( n1534 & n1543 ) ;
  assign n1546 = ( n1437 & ~n1544 ) | ( n1437 & n1545 ) | ( ~n1544 & n1545 ) ;
  assign n1547 = ( n1440 & n1517 ) | ( n1440 & n1546 ) | ( n1517 & n1546 ) ;
  assign n1548 = ( ~n1440 & n1517 ) | ( ~n1440 & n1546 ) | ( n1517 & n1546 ) ;
  assign n1549 = ( n1440 & ~n1547 ) | ( n1440 & n1548 ) | ( ~n1547 & n1548 ) ;
  assign n1550 = ( n1443 & n1508 ) | ( n1443 & n1549 ) | ( n1508 & n1549 ) ;
  assign n1551 = ( ~n1443 & n1508 ) | ( ~n1443 & n1549 ) | ( n1508 & n1549 ) ;
  assign n1552 = ( n1443 & ~n1550 ) | ( n1443 & n1551 ) | ( ~n1550 & n1551 ) ;
  assign n1553 = n407 & n701 ;
  assign n1554 = x78 & n411 ;
  assign n1555 = x79 | n1554 ;
  assign n1556 = ( n413 & n1554 ) | ( n413 & n1555 ) | ( n1554 & n1555 ) ;
  assign n1557 = x77 & n491 ;
  assign n1558 = n1556 | n1557 ;
  assign n1559 = ( x11 & n1553 ) | ( x11 & ~n1558 ) | ( n1553 & ~n1558 ) ;
  assign n1560 = ( ~x11 & n1558 ) | ( ~x11 & n1559 ) | ( n1558 & n1559 ) ;
  assign n1561 = ( ~n1553 & n1559 ) | ( ~n1553 & n1560 ) | ( n1559 & n1560 ) ;
  assign n1562 = ( n1455 & n1552 ) | ( n1455 & n1561 ) | ( n1552 & n1561 ) ;
  assign n1563 = ( ~n1455 & n1552 ) | ( ~n1455 & n1561 ) | ( n1552 & n1561 ) ;
  assign n1564 = ( n1455 & ~n1562 ) | ( n1455 & n1563 ) | ( ~n1562 & n1563 ) ;
  assign n1565 = n291 & n990 ;
  assign n1566 = x81 & n295 ;
  assign n1567 = x82 | n1566 ;
  assign n1568 = ( n297 & n1566 ) | ( n297 & n1567 ) | ( n1566 & n1567 ) ;
  assign n1569 = x80 & n330 ;
  assign n1570 = n1568 | n1569 ;
  assign n1571 = ( x8 & n1565 ) | ( x8 & ~n1570 ) | ( n1565 & ~n1570 ) ;
  assign n1572 = ( ~x8 & n1570 ) | ( ~x8 & n1571 ) | ( n1570 & n1571 ) ;
  assign n1573 = ( ~n1565 & n1571 ) | ( ~n1565 & n1572 ) | ( n1571 & n1572 ) ;
  assign n1574 = ( n1458 & n1564 ) | ( n1458 & n1573 ) | ( n1564 & n1573 ) ;
  assign n1575 = ( ~n1458 & n1564 ) | ( ~n1458 & n1573 ) | ( n1564 & n1573 ) ;
  assign n1576 = ( n1458 & ~n1574 ) | ( n1458 & n1575 ) | ( ~n1574 & n1575 ) ;
  assign n1577 = ( n1461 & n1499 ) | ( n1461 & n1576 ) | ( n1499 & n1576 ) ;
  assign n1578 = ( ~n1461 & n1499 ) | ( ~n1461 & n1576 ) | ( n1499 & n1576 ) ;
  assign n1579 = ( n1461 & ~n1577 ) | ( n1461 & n1578 ) | ( ~n1577 & n1578 ) ;
  assign n1580 = ( n1476 & n1490 ) | ( n1476 & n1579 ) | ( n1490 & n1579 ) ;
  assign n1581 = ( ~n1476 & n1490 ) | ( ~n1476 & n1579 ) | ( n1490 & n1579 ) ;
  assign n1582 = ( n1476 & ~n1580 ) | ( n1476 & n1581 ) | ( ~n1580 & n1581 ) ;
  assign n1583 = ( x88 & x89 ) | ( x88 & n1479 ) | ( x89 & n1479 ) ;
  assign n1584 = ( x88 & ~x89 ) | ( x88 & n1479 ) | ( ~x89 & n1479 ) ;
  assign n1585 = ( x89 & ~n1583 ) | ( x89 & n1584 ) | ( ~n1583 & n1584 ) ;
  assign n1586 = n136 & n1585 ;
  assign n1587 = x88 & n138 ;
  assign n1588 = x89 | n1587 ;
  assign n1589 = ( n141 & n1587 ) | ( n141 & n1588 ) | ( n1587 & n1588 ) ;
  assign n1590 = x87 & n154 ;
  assign n1591 = n1589 | n1590 ;
  assign n1592 = ( x2 & n1586 ) | ( x2 & ~n1591 ) | ( n1586 & ~n1591 ) ;
  assign n1593 = ( ~x2 & n1591 ) | ( ~x2 & n1592 ) | ( n1591 & n1592 ) ;
  assign n1594 = ( ~n1586 & n1592 ) | ( ~n1586 & n1593 ) | ( n1592 & n1593 ) ;
  assign n1595 = n186 & n1366 ;
  assign n1596 = x85 & n190 ;
  assign n1597 = x86 | n1596 ;
  assign n1598 = ( n192 & n1596 ) | ( n192 & n1597 ) | ( n1596 & n1597 ) ;
  assign n1599 = x84 & n220 ;
  assign n1600 = n1598 | n1599 ;
  assign n1601 = ( x5 & n1595 ) | ( x5 & ~n1600 ) | ( n1595 & ~n1600 ) ;
  assign n1602 = ( ~x5 & n1600 ) | ( ~x5 & n1601 ) | ( n1600 & n1601 ) ;
  assign n1603 = ( ~n1595 & n1601 ) | ( ~n1595 & n1602 ) | ( n1601 & n1602 ) ;
  assign n1604 = n277 & n1016 ;
  assign n1605 = x70 & n1020 ;
  assign n1606 = x71 | n1605 ;
  assign n1607 = ( n1022 & n1605 ) | ( n1022 & n1606 ) | ( n1605 & n1606 ) ;
  assign n1608 = x69 & n1145 ;
  assign n1609 = n1607 | n1608 ;
  assign n1610 = ( x20 & n1604 ) | ( x20 & ~n1609 ) | ( n1604 & ~n1609 ) ;
  assign n1611 = ( ~x20 & n1609 ) | ( ~x20 & n1610 ) | ( n1609 & n1610 ) ;
  assign n1612 = ( ~n1604 & n1610 ) | ( ~n1604 & n1611 ) | ( n1610 & n1611 ) ;
  assign n1613 = x26 & n1530 ;
  assign n1614 = x25 | x26 ;
  assign n1615 = ( x25 & x26 ) | ( x25 & ~n1614 ) | ( x26 & ~n1614 ) ;
  assign n1616 = n1614 & ~n1615 ;
  assign n1617 = n1529 & n1616 ;
  assign n1618 = n133 & n1617 ;
  assign n1619 = ~x23 & x25 ;
  assign n1620 = x24 & x25 ;
  assign n1621 = ( n1527 & n1619 ) | ( n1527 & ~n1620 ) | ( n1619 & ~n1620 ) ;
  assign n1622 = x64 & n1621 ;
  assign n1623 = ( n1529 & ~n1614 ) | ( n1529 & n1615 ) | ( ~n1614 & n1615 ) ;
  assign n1624 = x65 | n1622 ;
  assign n1625 = ( n1622 & n1623 ) | ( n1622 & n1624 ) | ( n1623 & n1624 ) ;
  assign n1626 = ( n1613 & n1618 ) | ( n1613 & n1625 ) | ( n1618 & n1625 ) ;
  assign n1627 = n1618 | n1625 ;
  assign n1628 = ~n1613 & n1627 ;
  assign n1629 = ( n1613 & ~n1626 ) | ( n1613 & n1628 ) | ( ~n1626 & n1628 ) ;
  assign n1630 = x67 & n1301 ;
  assign n1631 = x68 | n1630 ;
  assign n1632 = ( n1303 & n1630 ) | ( n1303 & n1631 ) | ( n1630 & n1631 ) ;
  assign n1633 = x66 & n1426 ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = n201 & n1297 ;
  assign n1636 = ( x23 & n1634 ) | ( x23 & ~n1635 ) | ( n1634 & ~n1635 ) ;
  assign n1637 = ( ~x23 & n1635 ) | ( ~x23 & n1636 ) | ( n1635 & n1636 ) ;
  assign n1638 = ( ~n1634 & n1636 ) | ( ~n1634 & n1637 ) | ( n1636 & n1637 ) ;
  assign n1639 = ( n1532 & n1629 ) | ( n1532 & n1638 ) | ( n1629 & n1638 ) ;
  assign n1640 = ( ~n1532 & n1629 ) | ( ~n1532 & n1638 ) | ( n1629 & n1638 ) ;
  assign n1641 = ( n1532 & ~n1639 ) | ( n1532 & n1640 ) | ( ~n1639 & n1640 ) ;
  assign n1642 = ( n1544 & n1612 ) | ( n1544 & n1641 ) | ( n1612 & n1641 ) ;
  assign n1643 = ( ~n1544 & n1612 ) | ( ~n1544 & n1641 ) | ( n1612 & n1641 ) ;
  assign n1644 = ( n1544 & ~n1642 ) | ( n1544 & n1643 ) | ( ~n1642 & n1643 ) ;
  assign n1645 = n446 & n810 ;
  assign n1646 = x73 & n814 ;
  assign n1647 = x74 | n1646 ;
  assign n1648 = ( n816 & n1646 ) | ( n816 & n1647 ) | ( n1646 & n1647 ) ;
  assign n1649 = x72 & n885 ;
  assign n1650 = n1648 | n1649 ;
  assign n1651 = ( x17 & n1645 ) | ( x17 & ~n1650 ) | ( n1645 & ~n1650 ) ;
  assign n1652 = ( ~x17 & n1650 ) | ( ~x17 & n1651 ) | ( n1650 & n1651 ) ;
  assign n1653 = ( ~n1645 & n1651 ) | ( ~n1645 & n1652 ) | ( n1651 & n1652 ) ;
  assign n1654 = ( n1547 & n1644 ) | ( n1547 & n1653 ) | ( n1644 & n1653 ) ;
  assign n1655 = ( ~n1547 & n1644 ) | ( ~n1547 & n1653 ) | ( n1644 & n1653 ) ;
  assign n1656 = ( n1547 & ~n1654 ) | ( n1547 & n1655 ) | ( ~n1654 & n1655 ) ;
  assign n1657 = n569 & n583 ;
  assign n1658 = x76 & n587 ;
  assign n1659 = x77 | n1658 ;
  assign n1660 = ( n589 & n1658 ) | ( n589 & n1659 ) | ( n1658 & n1659 ) ;
  assign n1661 = x75 & n676 ;
  assign n1662 = n1660 | n1661 ;
  assign n1663 = ( x14 & n1657 ) | ( x14 & ~n1662 ) | ( n1657 & ~n1662 ) ;
  assign n1664 = ( ~x14 & n1662 ) | ( ~x14 & n1663 ) | ( n1662 & n1663 ) ;
  assign n1665 = ( ~n1657 & n1663 ) | ( ~n1657 & n1664 ) | ( n1663 & n1664 ) ;
  assign n1666 = ( n1550 & n1656 ) | ( n1550 & n1665 ) | ( n1656 & n1665 ) ;
  assign n1667 = ( n1550 & ~n1656 ) | ( n1550 & n1665 ) | ( ~n1656 & n1665 ) ;
  assign n1668 = ( n1656 & ~n1666 ) | ( n1656 & n1667 ) | ( ~n1666 & n1667 ) ;
  assign n1669 = n407 & n769 ;
  assign n1670 = x79 & n411 ;
  assign n1671 = x80 | n1670 ;
  assign n1672 = ( n413 & n1670 ) | ( n413 & n1671 ) | ( n1670 & n1671 ) ;
  assign n1673 = x78 & n491 ;
  assign n1674 = n1672 | n1673 ;
  assign n1675 = ( x11 & n1669 ) | ( x11 & ~n1674 ) | ( n1669 & ~n1674 ) ;
  assign n1676 = ( ~x11 & n1674 ) | ( ~x11 & n1675 ) | ( n1674 & n1675 ) ;
  assign n1677 = ( ~n1669 & n1675 ) | ( ~n1669 & n1676 ) | ( n1675 & n1676 ) ;
  assign n1678 = ( n1562 & n1668 ) | ( n1562 & n1677 ) | ( n1668 & n1677 ) ;
  assign n1679 = ( ~n1562 & n1668 ) | ( ~n1562 & n1677 ) | ( n1668 & n1677 ) ;
  assign n1680 = ( n1562 & ~n1678 ) | ( n1562 & n1679 ) | ( ~n1678 & n1679 ) ;
  assign n1681 = n291 & n1082 ;
  assign n1682 = x82 & n295 ;
  assign n1683 = x83 | n1682 ;
  assign n1684 = ( n297 & n1682 ) | ( n297 & n1683 ) | ( n1682 & n1683 ) ;
  assign n1685 = x81 & n330 ;
  assign n1686 = n1684 | n1685 ;
  assign n1687 = ( x8 & n1681 ) | ( x8 & ~n1686 ) | ( n1681 & ~n1686 ) ;
  assign n1688 = ( ~x8 & n1686 ) | ( ~x8 & n1687 ) | ( n1686 & n1687 ) ;
  assign n1689 = ( ~n1681 & n1687 ) | ( ~n1681 & n1688 ) | ( n1687 & n1688 ) ;
  assign n1690 = ( n1574 & n1680 ) | ( n1574 & n1689 ) | ( n1680 & n1689 ) ;
  assign n1691 = ( ~n1574 & n1680 ) | ( ~n1574 & n1689 ) | ( n1680 & n1689 ) ;
  assign n1692 = ( n1574 & ~n1690 ) | ( n1574 & n1691 ) | ( ~n1690 & n1691 ) ;
  assign n1693 = ( n1577 & n1603 ) | ( n1577 & n1692 ) | ( n1603 & n1692 ) ;
  assign n1694 = ( ~n1577 & n1603 ) | ( ~n1577 & n1692 ) | ( n1603 & n1692 ) ;
  assign n1695 = ( n1577 & ~n1693 ) | ( n1577 & n1694 ) | ( ~n1693 & n1694 ) ;
  assign n1696 = ( n1580 & n1594 ) | ( n1580 & n1695 ) | ( n1594 & n1695 ) ;
  assign n1697 = ( ~n1580 & n1594 ) | ( ~n1580 & n1695 ) | ( n1594 & n1695 ) ;
  assign n1698 = ( n1580 & ~n1696 ) | ( n1580 & n1697 ) | ( ~n1696 & n1697 ) ;
  assign n1699 = ( x89 & x90 ) | ( x89 & n1583 ) | ( x90 & n1583 ) ;
  assign n1700 = ( x89 & ~x90 ) | ( x89 & n1583 ) | ( ~x90 & n1583 ) ;
  assign n1701 = ( x90 & ~n1699 ) | ( x90 & n1700 ) | ( ~n1699 & n1700 ) ;
  assign n1702 = n136 & n1701 ;
  assign n1703 = x89 & n138 ;
  assign n1704 = x90 | n1703 ;
  assign n1705 = ( n141 & n1703 ) | ( n141 & n1704 ) | ( n1703 & n1704 ) ;
  assign n1706 = x88 & n154 ;
  assign n1707 = n1705 | n1706 ;
  assign n1708 = ( x2 & n1702 ) | ( x2 & ~n1707 ) | ( n1702 & ~n1707 ) ;
  assign n1709 = ( ~x2 & n1707 ) | ( ~x2 & n1708 ) | ( n1707 & n1708 ) ;
  assign n1710 = ( ~n1702 & n1708 ) | ( ~n1702 & n1709 ) | ( n1708 & n1709 ) ;
  assign n1711 = n407 & n910 ;
  assign n1712 = x80 & n411 ;
  assign n1713 = x81 | n1712 ;
  assign n1714 = ( n413 & n1712 ) | ( n413 & n1713 ) | ( n1712 & n1713 ) ;
  assign n1715 = x79 & n491 ;
  assign n1716 = n1714 | n1715 ;
  assign n1717 = ( x11 & n1711 ) | ( x11 & ~n1716 ) | ( n1711 & ~n1716 ) ;
  assign n1718 = ( ~x11 & n1716 ) | ( ~x11 & n1717 ) | ( n1716 & n1717 ) ;
  assign n1719 = ( ~n1711 & n1717 ) | ( ~n1711 & n1718 ) | ( n1717 & n1718 ) ;
  assign n1720 = n461 & n810 ;
  assign n1721 = x74 & n814 ;
  assign n1722 = x75 | n1721 ;
  assign n1723 = ( n816 & n1721 ) | ( n816 & n1722 ) | ( n1721 & n1722 ) ;
  assign n1724 = x73 & n885 ;
  assign n1725 = n1723 | n1724 ;
  assign n1726 = ( x17 & n1720 ) | ( x17 & ~n1725 ) | ( n1720 & ~n1725 ) ;
  assign n1727 = ( ~x17 & n1725 ) | ( ~x17 & n1726 ) | ( n1725 & n1726 ) ;
  assign n1728 = ( ~n1720 & n1726 ) | ( ~n1720 & n1727 ) | ( n1726 & n1727 ) ;
  assign n1729 = n346 & n1016 ;
  assign n1730 = x71 & n1020 ;
  assign n1731 = x72 | n1730 ;
  assign n1732 = ( n1022 & n1730 ) | ( n1022 & n1731 ) | ( n1730 & n1731 ) ;
  assign n1733 = x70 & n1145 ;
  assign n1734 = n1732 | n1733 ;
  assign n1735 = ( x20 & n1729 ) | ( x20 & ~n1734 ) | ( n1729 & ~n1734 ) ;
  assign n1736 = ( ~x20 & n1734 ) | ( ~x20 & n1735 ) | ( n1734 & n1735 ) ;
  assign n1737 = ( ~n1729 & n1735 ) | ( ~n1729 & n1736 ) | ( n1735 & n1736 ) ;
  assign n1738 = n230 & n1297 ;
  assign n1739 = x68 & n1301 ;
  assign n1740 = x69 | n1739 ;
  assign n1741 = ( n1303 & n1739 ) | ( n1303 & n1740 ) | ( n1739 & n1740 ) ;
  assign n1742 = x67 & n1426 ;
  assign n1743 = n1741 | n1742 ;
  assign n1744 = ( ~x23 & n1738 ) | ( ~x23 & n1743 ) | ( n1738 & n1743 ) ;
  assign n1745 = ( n1738 & n1743 ) | ( n1738 & ~n1744 ) | ( n1743 & ~n1744 ) ;
  assign n1746 = ( x23 & n1744 ) | ( x23 & ~n1745 ) | ( n1744 & ~n1745 ) ;
  assign n1747 = ( x26 & n1613 ) | ( x26 & n1627 ) | ( n1613 & n1627 ) ;
  assign n1748 = ( x23 & ~x25 ) | ( x23 & n1616 ) | ( ~x25 & n1616 ) ;
  assign n1749 = ( ~n1528 & n1620 ) | ( ~n1528 & n1748 ) | ( n1620 & n1748 ) ;
  assign n1750 = x64 & n1749 ;
  assign n1751 = x65 & n1621 ;
  assign n1752 = x66 | n1751 ;
  assign n1753 = ( n1623 & n1751 ) | ( n1623 & n1752 ) | ( n1751 & n1752 ) ;
  assign n1754 = ( n151 & n152 ) | ( n151 & n1617 ) | ( n152 & n1617 ) ;
  assign n1755 = ( ~n1750 & n1753 ) | ( ~n1750 & n1754 ) | ( n1753 & n1754 ) ;
  assign n1756 = n1750 | n1755 ;
  assign n1757 = n1747 | n1756 ;
  assign n1758 = ( n1747 & n1756 ) | ( n1747 & ~n1757 ) | ( n1756 & ~n1757 ) ;
  assign n1759 = n1757 & ~n1758 ;
  assign n1760 = ( n1639 & n1746 ) | ( n1639 & n1759 ) | ( n1746 & n1759 ) ;
  assign n1761 = ( ~n1639 & n1746 ) | ( ~n1639 & n1759 ) | ( n1746 & n1759 ) ;
  assign n1762 = ( n1639 & ~n1760 ) | ( n1639 & n1761 ) | ( ~n1760 & n1761 ) ;
  assign n1763 = ( n1642 & n1737 ) | ( n1642 & n1762 ) | ( n1737 & n1762 ) ;
  assign n1764 = ( ~n1642 & n1737 ) | ( ~n1642 & n1762 ) | ( n1737 & n1762 ) ;
  assign n1765 = ( n1642 & ~n1763 ) | ( n1642 & n1764 ) | ( ~n1763 & n1764 ) ;
  assign n1766 = ( n1654 & n1728 ) | ( n1654 & n1765 ) | ( n1728 & n1765 ) ;
  assign n1767 = ( ~n1654 & n1728 ) | ( ~n1654 & n1765 ) | ( n1728 & n1765 ) ;
  assign n1768 = ( n1654 & ~n1766 ) | ( n1654 & n1767 ) | ( ~n1766 & n1767 ) ;
  assign n1769 = n583 & n637 ;
  assign n1770 = x77 & n587 ;
  assign n1771 = x78 | n1770 ;
  assign n1772 = ( n589 & n1770 ) | ( n589 & n1771 ) | ( n1770 & n1771 ) ;
  assign n1773 = x76 & n676 ;
  assign n1774 = n1772 | n1773 ;
  assign n1775 = ( x14 & n1769 ) | ( x14 & ~n1774 ) | ( n1769 & ~n1774 ) ;
  assign n1776 = ( ~x14 & n1774 ) | ( ~x14 & n1775 ) | ( n1774 & n1775 ) ;
  assign n1777 = ( ~n1769 & n1775 ) | ( ~n1769 & n1776 ) | ( n1775 & n1776 ) ;
  assign n1778 = ( n1666 & n1768 ) | ( n1666 & n1777 ) | ( n1768 & n1777 ) ;
  assign n1779 = ( ~n1666 & n1768 ) | ( ~n1666 & n1777 ) | ( n1768 & n1777 ) ;
  assign n1780 = ( n1666 & ~n1778 ) | ( n1666 & n1779 ) | ( ~n1778 & n1779 ) ;
  assign n1781 = ( n1678 & n1719 ) | ( n1678 & n1780 ) | ( n1719 & n1780 ) ;
  assign n1782 = ( ~n1678 & n1719 ) | ( ~n1678 & n1780 ) | ( n1719 & n1780 ) ;
  assign n1783 = ( n1678 & ~n1781 ) | ( n1678 & n1782 ) | ( ~n1781 & n1782 ) ;
  assign n1784 = n291 & n1097 ;
  assign n1785 = x83 & n295 ;
  assign n1786 = x84 | n1785 ;
  assign n1787 = ( n297 & n1785 ) | ( n297 & n1786 ) | ( n1785 & n1786 ) ;
  assign n1788 = x82 & n330 ;
  assign n1789 = n1787 | n1788 ;
  assign n1790 = ( x8 & n1784 ) | ( x8 & ~n1789 ) | ( n1784 & ~n1789 ) ;
  assign n1791 = ( ~x8 & n1789 ) | ( ~x8 & n1790 ) | ( n1789 & n1790 ) ;
  assign n1792 = ( ~n1784 & n1790 ) | ( ~n1784 & n1791 ) | ( n1790 & n1791 ) ;
  assign n1793 = ( n1690 & n1783 ) | ( n1690 & n1792 ) | ( n1783 & n1792 ) ;
  assign n1794 = ( ~n1690 & n1783 ) | ( ~n1690 & n1792 ) | ( n1783 & n1792 ) ;
  assign n1795 = ( n1690 & ~n1793 ) | ( n1690 & n1794 ) | ( ~n1793 & n1794 ) ;
  assign n1796 = n186 & n1466 ;
  assign n1797 = x86 & n190 ;
  assign n1798 = x87 | n1797 ;
  assign n1799 = ( n192 & n1797 ) | ( n192 & n1798 ) | ( n1797 & n1798 ) ;
  assign n1800 = x85 & n220 ;
  assign n1801 = n1799 | n1800 ;
  assign n1802 = ( x5 & n1796 ) | ( x5 & ~n1801 ) | ( n1796 & ~n1801 ) ;
  assign n1803 = ( ~x5 & n1801 ) | ( ~x5 & n1802 ) | ( n1801 & n1802 ) ;
  assign n1804 = ( ~n1796 & n1802 ) | ( ~n1796 & n1803 ) | ( n1802 & n1803 ) ;
  assign n1805 = ( n1693 & n1795 ) | ( n1693 & n1804 ) | ( n1795 & n1804 ) ;
  assign n1806 = ( ~n1693 & n1795 ) | ( ~n1693 & n1804 ) | ( n1795 & n1804 ) ;
  assign n1807 = ( n1693 & ~n1805 ) | ( n1693 & n1806 ) | ( ~n1805 & n1806 ) ;
  assign n1808 = ( n1696 & n1710 ) | ( n1696 & n1807 ) | ( n1710 & n1807 ) ;
  assign n1809 = ( ~n1696 & n1710 ) | ( ~n1696 & n1807 ) | ( n1710 & n1807 ) ;
  assign n1810 = ( n1696 & ~n1808 ) | ( n1696 & n1809 ) | ( ~n1808 & n1809 ) ;
  assign n1811 = n554 & n810 ;
  assign n1812 = x75 & n814 ;
  assign n1813 = x76 | n1812 ;
  assign n1814 = ( n816 & n1812 ) | ( n816 & n1813 ) | ( n1812 & n1813 ) ;
  assign n1815 = x74 & n885 ;
  assign n1816 = n1814 | n1815 ;
  assign n1817 = ( x17 & n1811 ) | ( x17 & ~n1816 ) | ( n1811 & ~n1816 ) ;
  assign n1818 = ( ~x17 & n1816 ) | ( ~x17 & n1817 ) | ( n1816 & n1817 ) ;
  assign n1819 = ( ~n1811 & n1817 ) | ( ~n1811 & n1818 ) | ( n1817 & n1818 ) ;
  assign n1820 = n390 & n1016 ;
  assign n1821 = x72 & n1020 ;
  assign n1822 = x73 | n1821 ;
  assign n1823 = ( n1022 & n1821 ) | ( n1022 & n1822 ) | ( n1821 & n1822 ) ;
  assign n1824 = x71 & n1145 ;
  assign n1825 = n1823 | n1824 ;
  assign n1826 = ( x20 & n1820 ) | ( x20 & ~n1825 ) | ( n1820 & ~n1825 ) ;
  assign n1827 = ( ~x20 & n1825 ) | ( ~x20 & n1826 ) | ( n1825 & n1826 ) ;
  assign n1828 = ( ~n1820 & n1826 ) | ( ~n1820 & n1827 ) | ( n1826 & n1827 ) ;
  assign n1829 = x66 & n1621 ;
  assign n1830 = x67 | n1829 ;
  assign n1831 = ( n1623 & n1829 ) | ( n1623 & n1830 ) | ( n1829 & n1830 ) ;
  assign n1832 = x65 & n1749 ;
  assign n1833 = n1831 | n1832 ;
  assign n1834 = n164 & n1617 ;
  assign n1835 = ( x26 & n1833 ) | ( x26 & ~n1834 ) | ( n1833 & ~n1834 ) ;
  assign n1836 = ( ~x26 & n1834 ) | ( ~x26 & n1835 ) | ( n1834 & n1835 ) ;
  assign n1837 = ( ~n1833 & n1835 ) | ( ~n1833 & n1836 ) | ( n1835 & n1836 ) ;
  assign n1838 = x26 & x27 ;
  assign n1839 = x26 | x27 ;
  assign n1840 = ~n1838 & n1839 ;
  assign n1841 = x64 & n1840 ;
  assign n1842 = x26 & ~n1757 ;
  assign n1843 = ( n1837 & n1841 ) | ( n1837 & n1842 ) | ( n1841 & n1842 ) ;
  assign n1844 = ( ~n1837 & n1841 ) | ( ~n1837 & n1842 ) | ( n1841 & n1842 ) ;
  assign n1845 = ( n1837 & ~n1843 ) | ( n1837 & n1844 ) | ( ~n1843 & n1844 ) ;
  assign n1846 = n245 & n1297 ;
  assign n1847 = x69 & n1301 ;
  assign n1848 = x70 | n1847 ;
  assign n1849 = ( n1303 & n1847 ) | ( n1303 & n1848 ) | ( n1847 & n1848 ) ;
  assign n1850 = x68 & n1426 ;
  assign n1851 = n1849 | n1850 ;
  assign n1852 = ( x23 & n1846 ) | ( x23 & ~n1851 ) | ( n1846 & ~n1851 ) ;
  assign n1853 = ( ~x23 & n1851 ) | ( ~x23 & n1852 ) | ( n1851 & n1852 ) ;
  assign n1854 = ( ~n1846 & n1852 ) | ( ~n1846 & n1853 ) | ( n1852 & n1853 ) ;
  assign n1855 = ( n1760 & n1845 ) | ( n1760 & n1854 ) | ( n1845 & n1854 ) ;
  assign n1856 = ( ~n1760 & n1845 ) | ( ~n1760 & n1854 ) | ( n1845 & n1854 ) ;
  assign n1857 = ( n1760 & ~n1855 ) | ( n1760 & n1856 ) | ( ~n1855 & n1856 ) ;
  assign n1858 = ( n1763 & n1828 ) | ( n1763 & n1857 ) | ( n1828 & n1857 ) ;
  assign n1859 = ( ~n1763 & n1828 ) | ( ~n1763 & n1857 ) | ( n1828 & n1857 ) ;
  assign n1860 = ( n1763 & ~n1858 ) | ( n1763 & n1859 ) | ( ~n1858 & n1859 ) ;
  assign n1861 = ( n1766 & n1819 ) | ( n1766 & n1860 ) | ( n1819 & n1860 ) ;
  assign n1862 = ( ~n1766 & n1819 ) | ( ~n1766 & n1860 ) | ( n1819 & n1860 ) ;
  assign n1863 = ( n1766 & ~n1861 ) | ( n1766 & n1862 ) | ( ~n1861 & n1862 ) ;
  assign n1864 = n583 & n701 ;
  assign n1865 = x78 & n587 ;
  assign n1866 = x79 | n1865 ;
  assign n1867 = ( n589 & n1865 ) | ( n589 & n1866 ) | ( n1865 & n1866 ) ;
  assign n1868 = x77 & n676 ;
  assign n1869 = n1867 | n1868 ;
  assign n1870 = ( x14 & n1864 ) | ( x14 & ~n1869 ) | ( n1864 & ~n1869 ) ;
  assign n1871 = ( ~x14 & n1869 ) | ( ~x14 & n1870 ) | ( n1869 & n1870 ) ;
  assign n1872 = ( ~n1864 & n1870 ) | ( ~n1864 & n1871 ) | ( n1870 & n1871 ) ;
  assign n1873 = ( n1778 & n1863 ) | ( n1778 & n1872 ) | ( n1863 & n1872 ) ;
  assign n1874 = ( ~n1778 & n1863 ) | ( ~n1778 & n1872 ) | ( n1863 & n1872 ) ;
  assign n1875 = ( n1778 & ~n1873 ) | ( n1778 & n1874 ) | ( ~n1873 & n1874 ) ;
  assign n1876 = n407 & n990 ;
  assign n1877 = x81 & n411 ;
  assign n1878 = x82 | n1877 ;
  assign n1879 = ( n413 & n1877 ) | ( n413 & n1878 ) | ( n1877 & n1878 ) ;
  assign n1880 = x80 & n491 ;
  assign n1881 = n1879 | n1880 ;
  assign n1882 = ( x11 & n1876 ) | ( x11 & ~n1881 ) | ( n1876 & ~n1881 ) ;
  assign n1883 = ( ~x11 & n1881 ) | ( ~x11 & n1882 ) | ( n1881 & n1882 ) ;
  assign n1884 = ( ~n1876 & n1882 ) | ( ~n1876 & n1883 ) | ( n1882 & n1883 ) ;
  assign n1885 = ( n1781 & n1875 ) | ( n1781 & n1884 ) | ( n1875 & n1884 ) ;
  assign n1886 = ( ~n1781 & n1875 ) | ( ~n1781 & n1884 ) | ( n1875 & n1884 ) ;
  assign n1887 = ( n1781 & ~n1885 ) | ( n1781 & n1886 ) | ( ~n1885 & n1886 ) ;
  assign n1888 = n291 & n1262 ;
  assign n1889 = x84 & n295 ;
  assign n1890 = x85 | n1889 ;
  assign n1891 = ( n297 & n1889 ) | ( n297 & n1890 ) | ( n1889 & n1890 ) ;
  assign n1892 = x83 & n330 ;
  assign n1893 = n1891 | n1892 ;
  assign n1894 = ( x8 & n1888 ) | ( x8 & ~n1893 ) | ( n1888 & ~n1893 ) ;
  assign n1895 = ( ~x8 & n1893 ) | ( ~x8 & n1894 ) | ( n1893 & n1894 ) ;
  assign n1896 = ( ~n1888 & n1894 ) | ( ~n1888 & n1895 ) | ( n1894 & n1895 ) ;
  assign n1897 = ( n1793 & n1887 ) | ( n1793 & n1896 ) | ( n1887 & n1896 ) ;
  assign n1898 = ( n1793 & ~n1887 ) | ( n1793 & n1896 ) | ( ~n1887 & n1896 ) ;
  assign n1899 = ( n1887 & ~n1897 ) | ( n1887 & n1898 ) | ( ~n1897 & n1898 ) ;
  assign n1900 = n186 & n1481 ;
  assign n1901 = x87 & n190 ;
  assign n1902 = x88 | n1901 ;
  assign n1903 = ( n192 & n1901 ) | ( n192 & n1902 ) | ( n1901 & n1902 ) ;
  assign n1904 = x86 & n220 ;
  assign n1905 = n1903 | n1904 ;
  assign n1906 = ( x5 & n1900 ) | ( x5 & ~n1905 ) | ( n1900 & ~n1905 ) ;
  assign n1907 = ( ~x5 & n1905 ) | ( ~x5 & n1906 ) | ( n1905 & n1906 ) ;
  assign n1908 = ( ~n1900 & n1906 ) | ( ~n1900 & n1907 ) | ( n1906 & n1907 ) ;
  assign n1909 = ( n1805 & n1899 ) | ( n1805 & n1908 ) | ( n1899 & n1908 ) ;
  assign n1910 = ( ~n1805 & n1899 ) | ( ~n1805 & n1908 ) | ( n1899 & n1908 ) ;
  assign n1911 = ( n1805 & ~n1909 ) | ( n1805 & n1910 ) | ( ~n1909 & n1910 ) ;
  assign n1912 = ( x90 & x91 ) | ( x90 & n1699 ) | ( x91 & n1699 ) ;
  assign n1913 = ( x90 & ~x91 ) | ( x90 & n1699 ) | ( ~x91 & n1699 ) ;
  assign n1914 = ( x91 & ~n1912 ) | ( x91 & n1913 ) | ( ~n1912 & n1913 ) ;
  assign n1915 = n136 & n1914 ;
  assign n1916 = x90 & n138 ;
  assign n1917 = x91 | n1916 ;
  assign n1918 = ( n141 & n1916 ) | ( n141 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1919 = x89 & n154 ;
  assign n1920 = n1918 | n1919 ;
  assign n1921 = ( x2 & n1915 ) | ( x2 & ~n1920 ) | ( n1915 & ~n1920 ) ;
  assign n1922 = ( ~x2 & n1920 ) | ( ~x2 & n1921 ) | ( n1920 & n1921 ) ;
  assign n1923 = ( ~n1915 & n1921 ) | ( ~n1915 & n1922 ) | ( n1921 & n1922 ) ;
  assign n1924 = ( n1808 & n1911 ) | ( n1808 & n1923 ) | ( n1911 & n1923 ) ;
  assign n1925 = ( ~n1808 & n1911 ) | ( ~n1808 & n1923 ) | ( n1911 & n1923 ) ;
  assign n1926 = ( n1808 & ~n1924 ) | ( n1808 & n1925 ) | ( ~n1924 & n1925 ) ;
  assign n1927 = n583 & n769 ;
  assign n1928 = x79 & n587 ;
  assign n1929 = x80 | n1928 ;
  assign n1930 = ( n589 & n1928 ) | ( n589 & n1929 ) | ( n1928 & n1929 ) ;
  assign n1931 = x78 & n676 ;
  assign n1932 = n1930 | n1931 ;
  assign n1933 = ( x14 & n1927 ) | ( x14 & ~n1932 ) | ( n1927 & ~n1932 ) ;
  assign n1934 = ( ~x14 & n1932 ) | ( ~x14 & n1933 ) | ( n1932 & n1933 ) ;
  assign n1935 = ( ~n1927 & n1933 ) | ( ~n1927 & n1934 ) | ( n1933 & n1934 ) ;
  assign n1936 = n277 & n1297 ;
  assign n1937 = x70 & n1301 ;
  assign n1938 = x71 | n1937 ;
  assign n1939 = ( n1303 & n1937 ) | ( n1303 & n1938 ) | ( n1937 & n1938 ) ;
  assign n1940 = x69 & n1426 ;
  assign n1941 = n1939 | n1940 ;
  assign n1942 = ( x23 & n1936 ) | ( x23 & ~n1941 ) | ( n1936 & ~n1941 ) ;
  assign n1943 = ( ~x23 & n1941 ) | ( ~x23 & n1942 ) | ( n1941 & n1942 ) ;
  assign n1944 = ( ~n1936 & n1942 ) | ( ~n1936 & n1943 ) | ( n1942 & n1943 ) ;
  assign n1945 = x29 & n1841 ;
  assign n1946 = x28 | x29 ;
  assign n1947 = ( x28 & x29 ) | ( x28 & ~n1946 ) | ( x29 & ~n1946 ) ;
  assign n1948 = n1946 & ~n1947 ;
  assign n1949 = n1840 & n1948 ;
  assign n1950 = n133 & n1949 ;
  assign n1951 = ~x26 & x28 ;
  assign n1952 = x27 & x28 ;
  assign n1953 = ( n1838 & n1951 ) | ( n1838 & ~n1952 ) | ( n1951 & ~n1952 ) ;
  assign n1954 = x64 & n1953 ;
  assign n1955 = ( n1840 & ~n1946 ) | ( n1840 & n1947 ) | ( ~n1946 & n1947 ) ;
  assign n1956 = x65 | n1954 ;
  assign n1957 = ( n1954 & n1955 ) | ( n1954 & n1956 ) | ( n1955 & n1956 ) ;
  assign n1958 = ( n1945 & n1950 ) | ( n1945 & n1957 ) | ( n1950 & n1957 ) ;
  assign n1959 = n1950 | n1957 ;
  assign n1960 = ~n1945 & n1959 ;
  assign n1961 = ( n1945 & ~n1958 ) | ( n1945 & n1960 ) | ( ~n1958 & n1960 ) ;
  assign n1962 = x67 & n1621 ;
  assign n1963 = x68 | n1962 ;
  assign n1964 = ( n1623 & n1962 ) | ( n1623 & n1963 ) | ( n1962 & n1963 ) ;
  assign n1965 = x66 & n1749 ;
  assign n1966 = n1964 | n1965 ;
  assign n1967 = n201 & n1617 ;
  assign n1968 = ( x26 & n1966 ) | ( x26 & ~n1967 ) | ( n1966 & ~n1967 ) ;
  assign n1969 = ( ~x26 & n1967 ) | ( ~x26 & n1968 ) | ( n1967 & n1968 ) ;
  assign n1970 = ( ~n1966 & n1968 ) | ( ~n1966 & n1969 ) | ( n1968 & n1969 ) ;
  assign n1971 = ( n1843 & n1961 ) | ( n1843 & n1970 ) | ( n1961 & n1970 ) ;
  assign n1972 = ( ~n1843 & n1961 ) | ( ~n1843 & n1970 ) | ( n1961 & n1970 ) ;
  assign n1973 = ( n1843 & ~n1971 ) | ( n1843 & n1972 ) | ( ~n1971 & n1972 ) ;
  assign n1974 = ( n1855 & n1944 ) | ( n1855 & n1973 ) | ( n1944 & n1973 ) ;
  assign n1975 = ( ~n1855 & n1944 ) | ( ~n1855 & n1973 ) | ( n1944 & n1973 ) ;
  assign n1976 = ( n1855 & ~n1974 ) | ( n1855 & n1975 ) | ( ~n1974 & n1975 ) ;
  assign n1977 = n446 & n1016 ;
  assign n1978 = x73 & n1020 ;
  assign n1979 = x74 | n1978 ;
  assign n1980 = ( n1022 & n1978 ) | ( n1022 & n1979 ) | ( n1978 & n1979 ) ;
  assign n1981 = x72 & n1145 ;
  assign n1982 = n1980 | n1981 ;
  assign n1983 = ( x20 & n1977 ) | ( x20 & ~n1982 ) | ( n1977 & ~n1982 ) ;
  assign n1984 = ( ~x20 & n1982 ) | ( ~x20 & n1983 ) | ( n1982 & n1983 ) ;
  assign n1985 = ( ~n1977 & n1983 ) | ( ~n1977 & n1984 ) | ( n1983 & n1984 ) ;
  assign n1986 = ( n1858 & n1976 ) | ( n1858 & n1985 ) | ( n1976 & n1985 ) ;
  assign n1987 = ( ~n1858 & n1976 ) | ( ~n1858 & n1985 ) | ( n1976 & n1985 ) ;
  assign n1988 = ( n1858 & ~n1986 ) | ( n1858 & n1987 ) | ( ~n1986 & n1987 ) ;
  assign n1989 = n569 & n810 ;
  assign n1990 = x76 & n814 ;
  assign n1991 = x77 | n1990 ;
  assign n1992 = ( n816 & n1990 ) | ( n816 & n1991 ) | ( n1990 & n1991 ) ;
  assign n1993 = x75 & n885 ;
  assign n1994 = n1992 | n1993 ;
  assign n1995 = ( x17 & n1989 ) | ( x17 & ~n1994 ) | ( n1989 & ~n1994 ) ;
  assign n1996 = ( ~x17 & n1994 ) | ( ~x17 & n1995 ) | ( n1994 & n1995 ) ;
  assign n1997 = ( ~n1989 & n1995 ) | ( ~n1989 & n1996 ) | ( n1995 & n1996 ) ;
  assign n1998 = ( n1861 & n1988 ) | ( n1861 & n1997 ) | ( n1988 & n1997 ) ;
  assign n1999 = ( ~n1861 & n1988 ) | ( ~n1861 & n1997 ) | ( n1988 & n1997 ) ;
  assign n2000 = ( n1861 & ~n1998 ) | ( n1861 & n1999 ) | ( ~n1998 & n1999 ) ;
  assign n2001 = ( n1873 & n1935 ) | ( n1873 & n2000 ) | ( n1935 & n2000 ) ;
  assign n2002 = ( ~n1873 & n1935 ) | ( ~n1873 & n2000 ) | ( n1935 & n2000 ) ;
  assign n2003 = ( n1873 & ~n2001 ) | ( n1873 & n2002 ) | ( ~n2001 & n2002 ) ;
  assign n2004 = n407 & n1082 ;
  assign n2005 = x82 & n411 ;
  assign n2006 = x83 | n2005 ;
  assign n2007 = ( n413 & n2005 ) | ( n413 & n2006 ) | ( n2005 & n2006 ) ;
  assign n2008 = x81 & n491 ;
  assign n2009 = n2007 | n2008 ;
  assign n2010 = ( x11 & n2004 ) | ( x11 & ~n2009 ) | ( n2004 & ~n2009 ) ;
  assign n2011 = ( ~x11 & n2009 ) | ( ~x11 & n2010 ) | ( n2009 & n2010 ) ;
  assign n2012 = ( ~n2004 & n2010 ) | ( ~n2004 & n2011 ) | ( n2010 & n2011 ) ;
  assign n2013 = ( n1885 & n2003 ) | ( n1885 & n2012 ) | ( n2003 & n2012 ) ;
  assign n2014 = ( ~n1885 & n2003 ) | ( ~n1885 & n2012 ) | ( n2003 & n2012 ) ;
  assign n2015 = ( n1885 & ~n2013 ) | ( n1885 & n2014 ) | ( ~n2013 & n2014 ) ;
  assign n2016 = n291 & n1366 ;
  assign n2017 = x85 & n295 ;
  assign n2018 = x86 | n2017 ;
  assign n2019 = ( n297 & n2017 ) | ( n297 & n2018 ) | ( n2017 & n2018 ) ;
  assign n2020 = x84 & n330 ;
  assign n2021 = n2019 | n2020 ;
  assign n2022 = ( x8 & n2016 ) | ( x8 & ~n2021 ) | ( n2016 & ~n2021 ) ;
  assign n2023 = ( ~x8 & n2021 ) | ( ~x8 & n2022 ) | ( n2021 & n2022 ) ;
  assign n2024 = ( ~n2016 & n2022 ) | ( ~n2016 & n2023 ) | ( n2022 & n2023 ) ;
  assign n2025 = ( n1897 & n2015 ) | ( n1897 & n2024 ) | ( n2015 & n2024 ) ;
  assign n2026 = ( n1897 & ~n2015 ) | ( n1897 & n2024 ) | ( ~n2015 & n2024 ) ;
  assign n2027 = ( n2015 & ~n2025 ) | ( n2015 & n2026 ) | ( ~n2025 & n2026 ) ;
  assign n2028 = n186 & n1585 ;
  assign n2029 = x88 & n190 ;
  assign n2030 = x89 | n2029 ;
  assign n2031 = ( n192 & n2029 ) | ( n192 & n2030 ) | ( n2029 & n2030 ) ;
  assign n2032 = x87 & n220 ;
  assign n2033 = n2031 | n2032 ;
  assign n2034 = ( x5 & n2028 ) | ( x5 & ~n2033 ) | ( n2028 & ~n2033 ) ;
  assign n2035 = ( ~x5 & n2033 ) | ( ~x5 & n2034 ) | ( n2033 & n2034 ) ;
  assign n2036 = ( ~n2028 & n2034 ) | ( ~n2028 & n2035 ) | ( n2034 & n2035 ) ;
  assign n2037 = ( n1909 & n2027 ) | ( n1909 & n2036 ) | ( n2027 & n2036 ) ;
  assign n2038 = ( ~n1909 & n2027 ) | ( ~n1909 & n2036 ) | ( n2027 & n2036 ) ;
  assign n2039 = ( n1909 & ~n2037 ) | ( n1909 & n2038 ) | ( ~n2037 & n2038 ) ;
  assign n2040 = ( x91 & x92 ) | ( x91 & n1912 ) | ( x92 & n1912 ) ;
  assign n2041 = ( x91 & ~x92 ) | ( x91 & n1912 ) | ( ~x92 & n1912 ) ;
  assign n2042 = ( x92 & ~n2040 ) | ( x92 & n2041 ) | ( ~n2040 & n2041 ) ;
  assign n2043 = n136 & n2042 ;
  assign n2044 = x91 & n138 ;
  assign n2045 = x92 | n2044 ;
  assign n2046 = ( n141 & n2044 ) | ( n141 & n2045 ) | ( n2044 & n2045 ) ;
  assign n2047 = x90 & n154 ;
  assign n2048 = n2046 | n2047 ;
  assign n2049 = ( x2 & n2043 ) | ( x2 & ~n2048 ) | ( n2043 & ~n2048 ) ;
  assign n2050 = ( ~x2 & n2048 ) | ( ~x2 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2051 = ( ~n2043 & n2049 ) | ( ~n2043 & n2050 ) | ( n2049 & n2050 ) ;
  assign n2052 = ( n1924 & n2039 ) | ( n1924 & n2051 ) | ( n2039 & n2051 ) ;
  assign n2053 = ( ~n1924 & n2039 ) | ( ~n1924 & n2051 ) | ( n2039 & n2051 ) ;
  assign n2054 = ( n1924 & ~n2052 ) | ( n1924 & n2053 ) | ( ~n2052 & n2053 ) ;
  assign n2055 = ( x92 & x93 ) | ( x92 & n2040 ) | ( x93 & n2040 ) ;
  assign n2056 = ( x92 & ~x93 ) | ( x92 & n2040 ) | ( ~x93 & n2040 ) ;
  assign n2057 = ( x93 & ~n2055 ) | ( x93 & n2056 ) | ( ~n2055 & n2056 ) ;
  assign n2058 = n136 & n2057 ;
  assign n2059 = x92 & n138 ;
  assign n2060 = x93 | n2059 ;
  assign n2061 = ( n141 & n2059 ) | ( n141 & n2060 ) | ( n2059 & n2060 ) ;
  assign n2062 = x91 & n154 ;
  assign n2063 = n2061 | n2062 ;
  assign n2064 = ( x2 & n2058 ) | ( x2 & ~n2063 ) | ( n2058 & ~n2063 ) ;
  assign n2065 = ( ~x2 & n2063 ) | ( ~x2 & n2064 ) | ( n2063 & n2064 ) ;
  assign n2066 = ( ~n2058 & n2064 ) | ( ~n2058 & n2065 ) | ( n2064 & n2065 ) ;
  assign n2067 = n186 & n1701 ;
  assign n2068 = x89 & n190 ;
  assign n2069 = x90 | n2068 ;
  assign n2070 = ( n192 & n2068 ) | ( n192 & n2069 ) | ( n2068 & n2069 ) ;
  assign n2071 = x88 & n220 ;
  assign n2072 = n2070 | n2071 ;
  assign n2073 = ( x5 & n2067 ) | ( x5 & ~n2072 ) | ( n2067 & ~n2072 ) ;
  assign n2074 = ( ~x5 & n2072 ) | ( ~x5 & n2073 ) | ( n2072 & n2073 ) ;
  assign n2075 = ( ~n2067 & n2073 ) | ( ~n2067 & n2074 ) | ( n2073 & n2074 ) ;
  assign n2076 = n291 & n1466 ;
  assign n2077 = x86 & n295 ;
  assign n2078 = x87 | n2077 ;
  assign n2079 = ( n297 & n2077 ) | ( n297 & n2078 ) | ( n2077 & n2078 ) ;
  assign n2080 = x85 & n330 ;
  assign n2081 = n2079 | n2080 ;
  assign n2082 = ( x8 & n2076 ) | ( x8 & ~n2081 ) | ( n2076 & ~n2081 ) ;
  assign n2083 = ( ~x8 & n2081 ) | ( ~x8 & n2082 ) | ( n2081 & n2082 ) ;
  assign n2084 = ( ~n2076 & n2082 ) | ( ~n2076 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2085 = n461 & n1016 ;
  assign n2086 = x74 & n1020 ;
  assign n2087 = x75 | n2086 ;
  assign n2088 = ( n1022 & n2086 ) | ( n1022 & n2087 ) | ( n2086 & n2087 ) ;
  assign n2089 = x73 & n1145 ;
  assign n2090 = n2088 | n2089 ;
  assign n2091 = ( x20 & n2085 ) | ( x20 & ~n2090 ) | ( n2085 & ~n2090 ) ;
  assign n2092 = ( ~x20 & n2090 ) | ( ~x20 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2093 = ( ~n2085 & n2091 ) | ( ~n2085 & n2092 ) | ( n2091 & n2092 ) ;
  assign n2094 = n346 & n1297 ;
  assign n2095 = x71 & n1301 ;
  assign n2096 = x72 | n2095 ;
  assign n2097 = ( n1303 & n2095 ) | ( n1303 & n2096 ) | ( n2095 & n2096 ) ;
  assign n2098 = x70 & n1426 ;
  assign n2099 = n2097 | n2098 ;
  assign n2100 = ( x23 & n2094 ) | ( x23 & ~n2099 ) | ( n2094 & ~n2099 ) ;
  assign n2101 = ( ~x23 & n2099 ) | ( ~x23 & n2100 ) | ( n2099 & n2100 ) ;
  assign n2102 = ( ~n2094 & n2100 ) | ( ~n2094 & n2101 ) | ( n2100 & n2101 ) ;
  assign n2103 = n230 & n1617 ;
  assign n2104 = x68 & n1621 ;
  assign n2105 = x69 | n2104 ;
  assign n2106 = ( n1623 & n2104 ) | ( n1623 & n2105 ) | ( n2104 & n2105 ) ;
  assign n2107 = x67 & n1749 ;
  assign n2108 = n2106 | n2107 ;
  assign n2109 = ( ~x26 & n2103 ) | ( ~x26 & n2108 ) | ( n2103 & n2108 ) ;
  assign n2110 = ( n2103 & n2108 ) | ( n2103 & ~n2109 ) | ( n2108 & ~n2109 ) ;
  assign n2111 = ( x26 & n2109 ) | ( x26 & ~n2110 ) | ( n2109 & ~n2110 ) ;
  assign n2112 = ( x29 & n1945 ) | ( x29 & n1959 ) | ( n1945 & n1959 ) ;
  assign n2113 = ( x26 & ~x28 ) | ( x26 & n1948 ) | ( ~x28 & n1948 ) ;
  assign n2114 = ( ~n1839 & n1952 ) | ( ~n1839 & n2113 ) | ( n1952 & n2113 ) ;
  assign n2115 = x64 & n2114 ;
  assign n2116 = x65 & n1953 ;
  assign n2117 = x66 | n2116 ;
  assign n2118 = ( n1955 & n2116 ) | ( n1955 & n2117 ) | ( n2116 & n2117 ) ;
  assign n2119 = ( n151 & n152 ) | ( n151 & n1949 ) | ( n152 & n1949 ) ;
  assign n2120 = ( ~n2115 & n2118 ) | ( ~n2115 & n2119 ) | ( n2118 & n2119 ) ;
  assign n2121 = n2115 | n2120 ;
  assign n2122 = n2112 | n2121 ;
  assign n2123 = ( n2112 & n2121 ) | ( n2112 & ~n2122 ) | ( n2121 & ~n2122 ) ;
  assign n2124 = n2122 & ~n2123 ;
  assign n2125 = ( n1971 & n2111 ) | ( n1971 & n2124 ) | ( n2111 & n2124 ) ;
  assign n2126 = ( ~n1971 & n2111 ) | ( ~n1971 & n2124 ) | ( n2111 & n2124 ) ;
  assign n2127 = ( n1971 & ~n2125 ) | ( n1971 & n2126 ) | ( ~n2125 & n2126 ) ;
  assign n2128 = ( n1974 & n2102 ) | ( n1974 & n2127 ) | ( n2102 & n2127 ) ;
  assign n2129 = ( ~n1974 & n2102 ) | ( ~n1974 & n2127 ) | ( n2102 & n2127 ) ;
  assign n2130 = ( n1974 & ~n2128 ) | ( n1974 & n2129 ) | ( ~n2128 & n2129 ) ;
  assign n2131 = ( n1986 & n2093 ) | ( n1986 & n2130 ) | ( n2093 & n2130 ) ;
  assign n2132 = ( ~n1986 & n2093 ) | ( ~n1986 & n2130 ) | ( n2093 & n2130 ) ;
  assign n2133 = ( n1986 & ~n2131 ) | ( n1986 & n2132 ) | ( ~n2131 & n2132 ) ;
  assign n2134 = n637 & n810 ;
  assign n2135 = x77 & n814 ;
  assign n2136 = x78 | n2135 ;
  assign n2137 = ( n816 & n2135 ) | ( n816 & n2136 ) | ( n2135 & n2136 ) ;
  assign n2138 = x76 & n885 ;
  assign n2139 = n2137 | n2138 ;
  assign n2140 = ( x17 & n2134 ) | ( x17 & ~n2139 ) | ( n2134 & ~n2139 ) ;
  assign n2141 = ( ~x17 & n2139 ) | ( ~x17 & n2140 ) | ( n2139 & n2140 ) ;
  assign n2142 = ( ~n2134 & n2140 ) | ( ~n2134 & n2141 ) | ( n2140 & n2141 ) ;
  assign n2143 = ( n1998 & n2133 ) | ( n1998 & n2142 ) | ( n2133 & n2142 ) ;
  assign n2144 = ( ~n1998 & n2133 ) | ( ~n1998 & n2142 ) | ( n2133 & n2142 ) ;
  assign n2145 = ( n1998 & ~n2143 ) | ( n1998 & n2144 ) | ( ~n2143 & n2144 ) ;
  assign n2146 = n583 & n910 ;
  assign n2147 = x80 & n587 ;
  assign n2148 = x81 | n2147 ;
  assign n2149 = ( n589 & n2147 ) | ( n589 & n2148 ) | ( n2147 & n2148 ) ;
  assign n2150 = x79 & n676 ;
  assign n2151 = n2149 | n2150 ;
  assign n2152 = ( x14 & n2146 ) | ( x14 & ~n2151 ) | ( n2146 & ~n2151 ) ;
  assign n2153 = ( ~x14 & n2151 ) | ( ~x14 & n2152 ) | ( n2151 & n2152 ) ;
  assign n2154 = ( ~n2146 & n2152 ) | ( ~n2146 & n2153 ) | ( n2152 & n2153 ) ;
  assign n2155 = ( n2001 & n2145 ) | ( n2001 & n2154 ) | ( n2145 & n2154 ) ;
  assign n2156 = ( ~n2001 & n2145 ) | ( ~n2001 & n2154 ) | ( n2145 & n2154 ) ;
  assign n2157 = ( n2001 & ~n2155 ) | ( n2001 & n2156 ) | ( ~n2155 & n2156 ) ;
  assign n2158 = n407 & n1097 ;
  assign n2159 = x83 & n411 ;
  assign n2160 = x84 | n2159 ;
  assign n2161 = ( n413 & n2159 ) | ( n413 & n2160 ) | ( n2159 & n2160 ) ;
  assign n2162 = x82 & n491 ;
  assign n2163 = n2161 | n2162 ;
  assign n2164 = ( x11 & n2158 ) | ( x11 & ~n2163 ) | ( n2158 & ~n2163 ) ;
  assign n2165 = ( ~x11 & n2163 ) | ( ~x11 & n2164 ) | ( n2163 & n2164 ) ;
  assign n2166 = ( ~n2158 & n2164 ) | ( ~n2158 & n2165 ) | ( n2164 & n2165 ) ;
  assign n2167 = ( n2013 & n2157 ) | ( n2013 & n2166 ) | ( n2157 & n2166 ) ;
  assign n2168 = ( ~n2013 & n2157 ) | ( ~n2013 & n2166 ) | ( n2157 & n2166 ) ;
  assign n2169 = ( n2013 & ~n2167 ) | ( n2013 & n2168 ) | ( ~n2167 & n2168 ) ;
  assign n2170 = ( n2025 & n2084 ) | ( n2025 & n2169 ) | ( n2084 & n2169 ) ;
  assign n2171 = ( ~n2025 & n2084 ) | ( ~n2025 & n2169 ) | ( n2084 & n2169 ) ;
  assign n2172 = ( n2025 & ~n2170 ) | ( n2025 & n2171 ) | ( ~n2170 & n2171 ) ;
  assign n2173 = ( n2037 & n2075 ) | ( n2037 & n2172 ) | ( n2075 & n2172 ) ;
  assign n2174 = ( ~n2037 & n2075 ) | ( ~n2037 & n2172 ) | ( n2075 & n2172 ) ;
  assign n2175 = ( n2037 & ~n2173 ) | ( n2037 & n2174 ) | ( ~n2173 & n2174 ) ;
  assign n2176 = ( n2052 & n2066 ) | ( n2052 & n2175 ) | ( n2066 & n2175 ) ;
  assign n2177 = ( ~n2052 & n2066 ) | ( ~n2052 & n2175 ) | ( n2066 & n2175 ) ;
  assign n2178 = ( n2052 & ~n2176 ) | ( n2052 & n2177 ) | ( ~n2176 & n2177 ) ;
  assign n2179 = n291 & n1481 ;
  assign n2180 = x87 & n295 ;
  assign n2181 = x88 | n2180 ;
  assign n2182 = ( n297 & n2180 ) | ( n297 & n2181 ) | ( n2180 & n2181 ) ;
  assign n2183 = x86 & n330 ;
  assign n2184 = n2182 | n2183 ;
  assign n2185 = ( x8 & n2179 ) | ( x8 & ~n2184 ) | ( n2179 & ~n2184 ) ;
  assign n2186 = ( ~x8 & n2184 ) | ( ~x8 & n2185 ) | ( n2184 & n2185 ) ;
  assign n2187 = ( ~n2179 & n2185 ) | ( ~n2179 & n2186 ) | ( n2185 & n2186 ) ;
  assign n2188 = n554 & n1016 ;
  assign n2189 = x75 & n1020 ;
  assign n2190 = x76 | n2189 ;
  assign n2191 = ( n1022 & n2189 ) | ( n1022 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2192 = x74 & n1145 ;
  assign n2193 = n2191 | n2192 ;
  assign n2194 = ( x20 & n2188 ) | ( x20 & ~n2193 ) | ( n2188 & ~n2193 ) ;
  assign n2195 = ( ~x20 & n2193 ) | ( ~x20 & n2194 ) | ( n2193 & n2194 ) ;
  assign n2196 = ( ~n2188 & n2194 ) | ( ~n2188 & n2195 ) | ( n2194 & n2195 ) ;
  assign n2197 = n390 & n1297 ;
  assign n2198 = x72 & n1301 ;
  assign n2199 = x73 | n2198 ;
  assign n2200 = ( n1303 & n2198 ) | ( n1303 & n2199 ) | ( n2198 & n2199 ) ;
  assign n2201 = x71 & n1426 ;
  assign n2202 = n2200 | n2201 ;
  assign n2203 = ( x23 & n2197 ) | ( x23 & ~n2202 ) | ( n2197 & ~n2202 ) ;
  assign n2204 = ( ~x23 & n2202 ) | ( ~x23 & n2203 ) | ( n2202 & n2203 ) ;
  assign n2205 = ( ~n2197 & n2203 ) | ( ~n2197 & n2204 ) | ( n2203 & n2204 ) ;
  assign n2206 = x66 & n1953 ;
  assign n2207 = x67 | n2206 ;
  assign n2208 = ( n1955 & n2206 ) | ( n1955 & n2207 ) | ( n2206 & n2207 ) ;
  assign n2209 = x65 & n2114 ;
  assign n2210 = n2208 | n2209 ;
  assign n2211 = n164 & n1949 ;
  assign n2212 = ( x29 & n2210 ) | ( x29 & ~n2211 ) | ( n2210 & ~n2211 ) ;
  assign n2213 = ( ~x29 & n2211 ) | ( ~x29 & n2212 ) | ( n2211 & n2212 ) ;
  assign n2214 = ( ~n2210 & n2212 ) | ( ~n2210 & n2213 ) | ( n2212 & n2213 ) ;
  assign n2215 = x29 & x30 ;
  assign n2216 = x29 | x30 ;
  assign n2217 = ~n2215 & n2216 ;
  assign n2218 = x64 & n2217 ;
  assign n2219 = x29 & ~n2122 ;
  assign n2220 = ( n2214 & n2218 ) | ( n2214 & n2219 ) | ( n2218 & n2219 ) ;
  assign n2221 = ( ~n2214 & n2218 ) | ( ~n2214 & n2219 ) | ( n2218 & n2219 ) ;
  assign n2222 = ( n2214 & ~n2220 ) | ( n2214 & n2221 ) | ( ~n2220 & n2221 ) ;
  assign n2223 = n245 & n1617 ;
  assign n2224 = x69 & n1621 ;
  assign n2225 = x70 | n2224 ;
  assign n2226 = ( n1623 & n2224 ) | ( n1623 & n2225 ) | ( n2224 & n2225 ) ;
  assign n2227 = x68 & n1749 ;
  assign n2228 = n2226 | n2227 ;
  assign n2229 = ( x26 & n2223 ) | ( x26 & ~n2228 ) | ( n2223 & ~n2228 ) ;
  assign n2230 = ( ~x26 & n2228 ) | ( ~x26 & n2229 ) | ( n2228 & n2229 ) ;
  assign n2231 = ( ~n2223 & n2229 ) | ( ~n2223 & n2230 ) | ( n2229 & n2230 ) ;
  assign n2232 = ( n2125 & n2222 ) | ( n2125 & n2231 ) | ( n2222 & n2231 ) ;
  assign n2233 = ( ~n2125 & n2222 ) | ( ~n2125 & n2231 ) | ( n2222 & n2231 ) ;
  assign n2234 = ( n2125 & ~n2232 ) | ( n2125 & n2233 ) | ( ~n2232 & n2233 ) ;
  assign n2235 = ( n2128 & n2205 ) | ( n2128 & n2234 ) | ( n2205 & n2234 ) ;
  assign n2236 = ( ~n2128 & n2205 ) | ( ~n2128 & n2234 ) | ( n2205 & n2234 ) ;
  assign n2237 = ( n2128 & ~n2235 ) | ( n2128 & n2236 ) | ( ~n2235 & n2236 ) ;
  assign n2238 = ( n2131 & n2196 ) | ( n2131 & n2237 ) | ( n2196 & n2237 ) ;
  assign n2239 = ( ~n2131 & n2196 ) | ( ~n2131 & n2237 ) | ( n2196 & n2237 ) ;
  assign n2240 = ( n2131 & ~n2238 ) | ( n2131 & n2239 ) | ( ~n2238 & n2239 ) ;
  assign n2241 = n701 & n810 ;
  assign n2242 = x78 & n814 ;
  assign n2243 = x79 | n2242 ;
  assign n2244 = ( n816 & n2242 ) | ( n816 & n2243 ) | ( n2242 & n2243 ) ;
  assign n2245 = x77 & n885 ;
  assign n2246 = n2244 | n2245 ;
  assign n2247 = ( x17 & n2241 ) | ( x17 & ~n2246 ) | ( n2241 & ~n2246 ) ;
  assign n2248 = ( ~x17 & n2246 ) | ( ~x17 & n2247 ) | ( n2246 & n2247 ) ;
  assign n2249 = ( ~n2241 & n2247 ) | ( ~n2241 & n2248 ) | ( n2247 & n2248 ) ;
  assign n2250 = ( n2143 & n2240 ) | ( n2143 & n2249 ) | ( n2240 & n2249 ) ;
  assign n2251 = ( ~n2143 & n2240 ) | ( ~n2143 & n2249 ) | ( n2240 & n2249 ) ;
  assign n2252 = ( n2143 & ~n2250 ) | ( n2143 & n2251 ) | ( ~n2250 & n2251 ) ;
  assign n2253 = n583 & n990 ;
  assign n2254 = x81 & n587 ;
  assign n2255 = x82 | n2254 ;
  assign n2256 = ( n589 & n2254 ) | ( n589 & n2255 ) | ( n2254 & n2255 ) ;
  assign n2257 = x80 & n676 ;
  assign n2258 = n2256 | n2257 ;
  assign n2259 = ( x14 & n2253 ) | ( x14 & ~n2258 ) | ( n2253 & ~n2258 ) ;
  assign n2260 = ( ~x14 & n2258 ) | ( ~x14 & n2259 ) | ( n2258 & n2259 ) ;
  assign n2261 = ( ~n2253 & n2259 ) | ( ~n2253 & n2260 ) | ( n2259 & n2260 ) ;
  assign n2262 = ( n2155 & n2252 ) | ( n2155 & n2261 ) | ( n2252 & n2261 ) ;
  assign n2263 = ( ~n2155 & n2252 ) | ( ~n2155 & n2261 ) | ( n2252 & n2261 ) ;
  assign n2264 = ( n2155 & ~n2262 ) | ( n2155 & n2263 ) | ( ~n2262 & n2263 ) ;
  assign n2265 = n407 & n1262 ;
  assign n2266 = x84 & n411 ;
  assign n2267 = x85 | n2266 ;
  assign n2268 = ( n413 & n2266 ) | ( n413 & n2267 ) | ( n2266 & n2267 ) ;
  assign n2269 = x83 & n491 ;
  assign n2270 = n2268 | n2269 ;
  assign n2271 = ( x11 & n2265 ) | ( x11 & ~n2270 ) | ( n2265 & ~n2270 ) ;
  assign n2272 = ( ~x11 & n2270 ) | ( ~x11 & n2271 ) | ( n2270 & n2271 ) ;
  assign n2273 = ( ~n2265 & n2271 ) | ( ~n2265 & n2272 ) | ( n2271 & n2272 ) ;
  assign n2274 = ( n2167 & n2264 ) | ( n2167 & n2273 ) | ( n2264 & n2273 ) ;
  assign n2275 = ( ~n2167 & n2264 ) | ( ~n2167 & n2273 ) | ( n2264 & n2273 ) ;
  assign n2276 = ( n2167 & ~n2274 ) | ( n2167 & n2275 ) | ( ~n2274 & n2275 ) ;
  assign n2277 = ( n2170 & n2187 ) | ( n2170 & n2276 ) | ( n2187 & n2276 ) ;
  assign n2278 = ( ~n2170 & n2187 ) | ( ~n2170 & n2276 ) | ( n2187 & n2276 ) ;
  assign n2279 = ( n2170 & ~n2277 ) | ( n2170 & n2278 ) | ( ~n2277 & n2278 ) ;
  assign n2280 = n186 & n1914 ;
  assign n2281 = x90 & n190 ;
  assign n2282 = x91 | n2281 ;
  assign n2283 = ( n192 & n2281 ) | ( n192 & n2282 ) | ( n2281 & n2282 ) ;
  assign n2284 = x89 & n220 ;
  assign n2285 = n2283 | n2284 ;
  assign n2286 = ( x5 & n2280 ) | ( x5 & ~n2285 ) | ( n2280 & ~n2285 ) ;
  assign n2287 = ( ~x5 & n2285 ) | ( ~x5 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2288 = ( ~n2280 & n2286 ) | ( ~n2280 & n2287 ) | ( n2286 & n2287 ) ;
  assign n2289 = ( n2173 & n2279 ) | ( n2173 & n2288 ) | ( n2279 & n2288 ) ;
  assign n2290 = ( ~n2173 & n2279 ) | ( ~n2173 & n2288 ) | ( n2279 & n2288 ) ;
  assign n2291 = ( n2173 & ~n2289 ) | ( n2173 & n2290 ) | ( ~n2289 & n2290 ) ;
  assign n2292 = ( x93 & x94 ) | ( x93 & n2055 ) | ( x94 & n2055 ) ;
  assign n2293 = ( x93 & ~x94 ) | ( x93 & n2055 ) | ( ~x94 & n2055 ) ;
  assign n2294 = ( x94 & ~n2292 ) | ( x94 & n2293 ) | ( ~n2292 & n2293 ) ;
  assign n2295 = n136 & n2294 ;
  assign n2296 = x93 & n138 ;
  assign n2297 = x94 | n2296 ;
  assign n2298 = ( n141 & n2296 ) | ( n141 & n2297 ) | ( n2296 & n2297 ) ;
  assign n2299 = x92 & n154 ;
  assign n2300 = n2298 | n2299 ;
  assign n2301 = ( x2 & n2295 ) | ( x2 & ~n2300 ) | ( n2295 & ~n2300 ) ;
  assign n2302 = ( ~x2 & n2300 ) | ( ~x2 & n2301 ) | ( n2300 & n2301 ) ;
  assign n2303 = ( ~n2295 & n2301 ) | ( ~n2295 & n2302 ) | ( n2301 & n2302 ) ;
  assign n2304 = ( n2176 & n2291 ) | ( n2176 & n2303 ) | ( n2291 & n2303 ) ;
  assign n2305 = ( ~n2176 & n2291 ) | ( ~n2176 & n2303 ) | ( n2291 & n2303 ) ;
  assign n2306 = ( n2176 & ~n2304 ) | ( n2176 & n2305 ) | ( ~n2304 & n2305 ) ;
  assign n2307 = n277 & n1617 ;
  assign n2308 = x70 & n1621 ;
  assign n2309 = x71 | n2308 ;
  assign n2310 = ( n1623 & n2308 ) | ( n1623 & n2309 ) | ( n2308 & n2309 ) ;
  assign n2311 = x69 & n1749 ;
  assign n2312 = n2310 | n2311 ;
  assign n2313 = ( x26 & n2307 ) | ( x26 & ~n2312 ) | ( n2307 & ~n2312 ) ;
  assign n2314 = ( ~x26 & n2312 ) | ( ~x26 & n2313 ) | ( n2312 & n2313 ) ;
  assign n2315 = ( ~n2307 & n2313 ) | ( ~n2307 & n2314 ) | ( n2313 & n2314 ) ;
  assign n2316 = x32 & n2218 ;
  assign n2317 = x31 | x32 ;
  assign n2318 = ( x31 & x32 ) | ( x31 & ~n2317 ) | ( x32 & ~n2317 ) ;
  assign n2319 = n2317 & ~n2318 ;
  assign n2320 = n2217 & n2319 ;
  assign n2321 = n133 & n2320 ;
  assign n2322 = ~x29 & x31 ;
  assign n2323 = x30 & x31 ;
  assign n2324 = ( n2215 & n2322 ) | ( n2215 & ~n2323 ) | ( n2322 & ~n2323 ) ;
  assign n2325 = x64 & n2324 ;
  assign n2326 = ( n2217 & ~n2317 ) | ( n2217 & n2318 ) | ( ~n2317 & n2318 ) ;
  assign n2327 = x65 | n2325 ;
  assign n2328 = ( n2325 & n2326 ) | ( n2325 & n2327 ) | ( n2326 & n2327 ) ;
  assign n2329 = ( n2316 & n2321 ) | ( n2316 & n2328 ) | ( n2321 & n2328 ) ;
  assign n2330 = n2321 | n2328 ;
  assign n2331 = ~n2316 & n2330 ;
  assign n2332 = ( n2316 & ~n2329 ) | ( n2316 & n2331 ) | ( ~n2329 & n2331 ) ;
  assign n2333 = x67 & n1953 ;
  assign n2334 = x68 | n2333 ;
  assign n2335 = ( n1955 & n2333 ) | ( n1955 & n2334 ) | ( n2333 & n2334 ) ;
  assign n2336 = x66 & n2114 ;
  assign n2337 = n2335 | n2336 ;
  assign n2338 = n201 & n1949 ;
  assign n2339 = ( x29 & n2337 ) | ( x29 & ~n2338 ) | ( n2337 & ~n2338 ) ;
  assign n2340 = ( ~x29 & n2338 ) | ( ~x29 & n2339 ) | ( n2338 & n2339 ) ;
  assign n2341 = ( ~n2337 & n2339 ) | ( ~n2337 & n2340 ) | ( n2339 & n2340 ) ;
  assign n2342 = ( n2220 & n2332 ) | ( n2220 & n2341 ) | ( n2332 & n2341 ) ;
  assign n2343 = ( ~n2220 & n2332 ) | ( ~n2220 & n2341 ) | ( n2332 & n2341 ) ;
  assign n2344 = ( n2220 & ~n2342 ) | ( n2220 & n2343 ) | ( ~n2342 & n2343 ) ;
  assign n2345 = ( n2232 & n2315 ) | ( n2232 & n2344 ) | ( n2315 & n2344 ) ;
  assign n2346 = ( ~n2232 & n2315 ) | ( ~n2232 & n2344 ) | ( n2315 & n2344 ) ;
  assign n2347 = ( n2232 & ~n2345 ) | ( n2232 & n2346 ) | ( ~n2345 & n2346 ) ;
  assign n2348 = n446 & n1297 ;
  assign n2349 = x73 & n1301 ;
  assign n2350 = x74 | n2349 ;
  assign n2351 = ( n1303 & n2349 ) | ( n1303 & n2350 ) | ( n2349 & n2350 ) ;
  assign n2352 = x72 & n1426 ;
  assign n2353 = n2351 | n2352 ;
  assign n2354 = ( x23 & n2348 ) | ( x23 & ~n2353 ) | ( n2348 & ~n2353 ) ;
  assign n2355 = ( ~x23 & n2353 ) | ( ~x23 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2356 = ( ~n2348 & n2354 ) | ( ~n2348 & n2355 ) | ( n2354 & n2355 ) ;
  assign n2357 = ( n2235 & n2347 ) | ( n2235 & n2356 ) | ( n2347 & n2356 ) ;
  assign n2358 = ( ~n2235 & n2347 ) | ( ~n2235 & n2356 ) | ( n2347 & n2356 ) ;
  assign n2359 = ( n2235 & ~n2357 ) | ( n2235 & n2358 ) | ( ~n2357 & n2358 ) ;
  assign n2360 = n569 & n1016 ;
  assign n2361 = x76 & n1020 ;
  assign n2362 = x77 | n2361 ;
  assign n2363 = ( n1022 & n2361 ) | ( n1022 & n2362 ) | ( n2361 & n2362 ) ;
  assign n2364 = x75 & n1145 ;
  assign n2365 = n2363 | n2364 ;
  assign n2366 = ( x20 & n2360 ) | ( x20 & ~n2365 ) | ( n2360 & ~n2365 ) ;
  assign n2367 = ( ~x20 & n2365 ) | ( ~x20 & n2366 ) | ( n2365 & n2366 ) ;
  assign n2368 = ( ~n2360 & n2366 ) | ( ~n2360 & n2367 ) | ( n2366 & n2367 ) ;
  assign n2369 = ( n2238 & n2359 ) | ( n2238 & n2368 ) | ( n2359 & n2368 ) ;
  assign n2370 = ( n2238 & ~n2359 ) | ( n2238 & n2368 ) | ( ~n2359 & n2368 ) ;
  assign n2371 = ( n2359 & ~n2369 ) | ( n2359 & n2370 ) | ( ~n2369 & n2370 ) ;
  assign n2372 = n769 & n810 ;
  assign n2373 = x79 & n814 ;
  assign n2374 = x80 | n2373 ;
  assign n2375 = ( n816 & n2373 ) | ( n816 & n2374 ) | ( n2373 & n2374 ) ;
  assign n2376 = x78 & n885 ;
  assign n2377 = n2375 | n2376 ;
  assign n2378 = ( x17 & n2372 ) | ( x17 & ~n2377 ) | ( n2372 & ~n2377 ) ;
  assign n2379 = ( ~x17 & n2377 ) | ( ~x17 & n2378 ) | ( n2377 & n2378 ) ;
  assign n2380 = ( ~n2372 & n2378 ) | ( ~n2372 & n2379 ) | ( n2378 & n2379 ) ;
  assign n2381 = ( n2250 & n2371 ) | ( n2250 & n2380 ) | ( n2371 & n2380 ) ;
  assign n2382 = ( ~n2250 & n2371 ) | ( ~n2250 & n2380 ) | ( n2371 & n2380 ) ;
  assign n2383 = ( n2250 & ~n2381 ) | ( n2250 & n2382 ) | ( ~n2381 & n2382 ) ;
  assign n2384 = n583 & n1082 ;
  assign n2385 = x82 & n587 ;
  assign n2386 = x83 | n2385 ;
  assign n2387 = ( n589 & n2385 ) | ( n589 & n2386 ) | ( n2385 & n2386 ) ;
  assign n2388 = x81 & n676 ;
  assign n2389 = n2387 | n2388 ;
  assign n2390 = ( x14 & n2384 ) | ( x14 & ~n2389 ) | ( n2384 & ~n2389 ) ;
  assign n2391 = ( ~x14 & n2389 ) | ( ~x14 & n2390 ) | ( n2389 & n2390 ) ;
  assign n2392 = ( ~n2384 & n2390 ) | ( ~n2384 & n2391 ) | ( n2390 & n2391 ) ;
  assign n2393 = ( n2262 & n2383 ) | ( n2262 & n2392 ) | ( n2383 & n2392 ) ;
  assign n2394 = ( ~n2262 & n2383 ) | ( ~n2262 & n2392 ) | ( n2383 & n2392 ) ;
  assign n2395 = ( n2262 & ~n2393 ) | ( n2262 & n2394 ) | ( ~n2393 & n2394 ) ;
  assign n2396 = n407 & n1366 ;
  assign n2397 = x85 & n411 ;
  assign n2398 = x86 | n2397 ;
  assign n2399 = ( n413 & n2397 ) | ( n413 & n2398 ) | ( n2397 & n2398 ) ;
  assign n2400 = x84 & n491 ;
  assign n2401 = n2399 | n2400 ;
  assign n2402 = ( x11 & n2396 ) | ( x11 & ~n2401 ) | ( n2396 & ~n2401 ) ;
  assign n2403 = ( ~x11 & n2401 ) | ( ~x11 & n2402 ) | ( n2401 & n2402 ) ;
  assign n2404 = ( ~n2396 & n2402 ) | ( ~n2396 & n2403 ) | ( n2402 & n2403 ) ;
  assign n2405 = ( n2274 & n2395 ) | ( n2274 & n2404 ) | ( n2395 & n2404 ) ;
  assign n2406 = ( ~n2274 & n2395 ) | ( ~n2274 & n2404 ) | ( n2395 & n2404 ) ;
  assign n2407 = ( n2274 & ~n2405 ) | ( n2274 & n2406 ) | ( ~n2405 & n2406 ) ;
  assign n2408 = n291 & n1585 ;
  assign n2409 = x88 & n295 ;
  assign n2410 = x89 | n2409 ;
  assign n2411 = ( n297 & n2409 ) | ( n297 & n2410 ) | ( n2409 & n2410 ) ;
  assign n2412 = x87 & n330 ;
  assign n2413 = n2411 | n2412 ;
  assign n2414 = ( x8 & n2408 ) | ( x8 & ~n2413 ) | ( n2408 & ~n2413 ) ;
  assign n2415 = ( ~x8 & n2413 ) | ( ~x8 & n2414 ) | ( n2413 & n2414 ) ;
  assign n2416 = ( ~n2408 & n2414 ) | ( ~n2408 & n2415 ) | ( n2414 & n2415 ) ;
  assign n2417 = ( n2277 & n2407 ) | ( n2277 & n2416 ) | ( n2407 & n2416 ) ;
  assign n2418 = ( ~n2277 & n2407 ) | ( ~n2277 & n2416 ) | ( n2407 & n2416 ) ;
  assign n2419 = ( n2277 & ~n2417 ) | ( n2277 & n2418 ) | ( ~n2417 & n2418 ) ;
  assign n2420 = n186 & n2042 ;
  assign n2421 = x91 & n190 ;
  assign n2422 = x92 | n2421 ;
  assign n2423 = ( n192 & n2421 ) | ( n192 & n2422 ) | ( n2421 & n2422 ) ;
  assign n2424 = x90 & n220 ;
  assign n2425 = n2423 | n2424 ;
  assign n2426 = ( x5 & n2420 ) | ( x5 & ~n2425 ) | ( n2420 & ~n2425 ) ;
  assign n2427 = ( ~x5 & n2425 ) | ( ~x5 & n2426 ) | ( n2425 & n2426 ) ;
  assign n2428 = ( ~n2420 & n2426 ) | ( ~n2420 & n2427 ) | ( n2426 & n2427 ) ;
  assign n2429 = ( n2289 & n2419 ) | ( n2289 & n2428 ) | ( n2419 & n2428 ) ;
  assign n2430 = ( ~n2289 & n2419 ) | ( ~n2289 & n2428 ) | ( n2419 & n2428 ) ;
  assign n2431 = ( n2289 & ~n2429 ) | ( n2289 & n2430 ) | ( ~n2429 & n2430 ) ;
  assign n2432 = ( x94 & x95 ) | ( x94 & n2292 ) | ( x95 & n2292 ) ;
  assign n2433 = ( x94 & ~x95 ) | ( x94 & n2292 ) | ( ~x95 & n2292 ) ;
  assign n2434 = ( x95 & ~n2432 ) | ( x95 & n2433 ) | ( ~n2432 & n2433 ) ;
  assign n2435 = n136 & n2434 ;
  assign n2436 = x94 & n138 ;
  assign n2437 = x95 | n2436 ;
  assign n2438 = ( n141 & n2436 ) | ( n141 & n2437 ) | ( n2436 & n2437 ) ;
  assign n2439 = x93 & n154 ;
  assign n2440 = n2438 | n2439 ;
  assign n2441 = ( x2 & n2435 ) | ( x2 & ~n2440 ) | ( n2435 & ~n2440 ) ;
  assign n2442 = ( ~x2 & n2440 ) | ( ~x2 & n2441 ) | ( n2440 & n2441 ) ;
  assign n2443 = ( ~n2435 & n2441 ) | ( ~n2435 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2444 = ( n2304 & n2431 ) | ( n2304 & n2443 ) | ( n2431 & n2443 ) ;
  assign n2445 = ( ~n2304 & n2431 ) | ( ~n2304 & n2443 ) | ( n2431 & n2443 ) ;
  assign n2446 = ( n2304 & ~n2444 ) | ( n2304 & n2445 ) | ( ~n2444 & n2445 ) ;
  assign n2447 = ( x95 & x96 ) | ( x95 & n2432 ) | ( x96 & n2432 ) ;
  assign n2448 = ( x95 & ~x96 ) | ( x95 & n2432 ) | ( ~x96 & n2432 ) ;
  assign n2449 = ( x96 & ~n2447 ) | ( x96 & n2448 ) | ( ~n2447 & n2448 ) ;
  assign n2450 = n136 & n2449 ;
  assign n2451 = x95 & n138 ;
  assign n2452 = x96 | n2451 ;
  assign n2453 = ( n141 & n2451 ) | ( n141 & n2452 ) | ( n2451 & n2452 ) ;
  assign n2454 = x94 & n154 ;
  assign n2455 = n2453 | n2454 ;
  assign n2456 = ( x2 & n2450 ) | ( x2 & ~n2455 ) | ( n2450 & ~n2455 ) ;
  assign n2457 = ( ~x2 & n2455 ) | ( ~x2 & n2456 ) | ( n2455 & n2456 ) ;
  assign n2458 = ( ~n2450 & n2456 ) | ( ~n2450 & n2457 ) | ( n2456 & n2457 ) ;
  assign n2459 = n407 & n1466 ;
  assign n2460 = x86 & n411 ;
  assign n2461 = x87 | n2460 ;
  assign n2462 = ( n413 & n2460 ) | ( n413 & n2461 ) | ( n2460 & n2461 ) ;
  assign n2463 = x85 & n491 ;
  assign n2464 = n2462 | n2463 ;
  assign n2465 = ( x11 & n2459 ) | ( x11 & ~n2464 ) | ( n2459 & ~n2464 ) ;
  assign n2466 = ( ~x11 & n2464 ) | ( ~x11 & n2465 ) | ( n2464 & n2465 ) ;
  assign n2467 = ( ~n2459 & n2465 ) | ( ~n2459 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2468 = n637 & n1016 ;
  assign n2469 = x77 & n1020 ;
  assign n2470 = x78 | n2469 ;
  assign n2471 = ( n1022 & n2469 ) | ( n1022 & n2470 ) | ( n2469 & n2470 ) ;
  assign n2472 = x76 & n1145 ;
  assign n2473 = n2471 | n2472 ;
  assign n2474 = ( x20 & n2468 ) | ( x20 & ~n2473 ) | ( n2468 & ~n2473 ) ;
  assign n2475 = ( ~x20 & n2473 ) | ( ~x20 & n2474 ) | ( n2473 & n2474 ) ;
  assign n2476 = ( ~n2468 & n2474 ) | ( ~n2468 & n2475 ) | ( n2474 & n2475 ) ;
  assign n2477 = n346 & n1617 ;
  assign n2478 = x71 & n1621 ;
  assign n2479 = x72 | n2478 ;
  assign n2480 = ( n1623 & n2478 ) | ( n1623 & n2479 ) | ( n2478 & n2479 ) ;
  assign n2481 = x70 & n1749 ;
  assign n2482 = n2480 | n2481 ;
  assign n2483 = ( x26 & n2477 ) | ( x26 & ~n2482 ) | ( n2477 & ~n2482 ) ;
  assign n2484 = ( ~x26 & n2482 ) | ( ~x26 & n2483 ) | ( n2482 & n2483 ) ;
  assign n2485 = ( ~n2477 & n2483 ) | ( ~n2477 & n2484 ) | ( n2483 & n2484 ) ;
  assign n2486 = n230 & n1949 ;
  assign n2487 = x68 & n1953 ;
  assign n2488 = x69 | n2487 ;
  assign n2489 = ( n1955 & n2487 ) | ( n1955 & n2488 ) | ( n2487 & n2488 ) ;
  assign n2490 = x67 & n2114 ;
  assign n2491 = n2489 | n2490 ;
  assign n2492 = ( ~x29 & n2486 ) | ( ~x29 & n2491 ) | ( n2486 & n2491 ) ;
  assign n2493 = ( n2486 & n2491 ) | ( n2486 & ~n2492 ) | ( n2491 & ~n2492 ) ;
  assign n2494 = ( x29 & n2492 ) | ( x29 & ~n2493 ) | ( n2492 & ~n2493 ) ;
  assign n2495 = ( x32 & n2316 ) | ( x32 & n2330 ) | ( n2316 & n2330 ) ;
  assign n2496 = ( x29 & ~x31 ) | ( x29 & n2319 ) | ( ~x31 & n2319 ) ;
  assign n2497 = ( ~n2216 & n2323 ) | ( ~n2216 & n2496 ) | ( n2323 & n2496 ) ;
  assign n2498 = x64 & n2497 ;
  assign n2499 = x65 & n2324 ;
  assign n2500 = x66 | n2499 ;
  assign n2501 = ( n2326 & n2499 ) | ( n2326 & n2500 ) | ( n2499 & n2500 ) ;
  assign n2502 = ( n151 & n152 ) | ( n151 & n2320 ) | ( n152 & n2320 ) ;
  assign n2503 = ( ~n2498 & n2501 ) | ( ~n2498 & n2502 ) | ( n2501 & n2502 ) ;
  assign n2504 = n2498 | n2503 ;
  assign n2505 = n2495 | n2504 ;
  assign n2506 = ( n2495 & n2504 ) | ( n2495 & ~n2505 ) | ( n2504 & ~n2505 ) ;
  assign n2507 = n2505 & ~n2506 ;
  assign n2508 = ( n2342 & n2494 ) | ( n2342 & n2507 ) | ( n2494 & n2507 ) ;
  assign n2509 = ( ~n2342 & n2494 ) | ( ~n2342 & n2507 ) | ( n2494 & n2507 ) ;
  assign n2510 = ( n2342 & ~n2508 ) | ( n2342 & n2509 ) | ( ~n2508 & n2509 ) ;
  assign n2511 = ( n2345 & n2485 ) | ( n2345 & n2510 ) | ( n2485 & n2510 ) ;
  assign n2512 = ( ~n2345 & n2485 ) | ( ~n2345 & n2510 ) | ( n2485 & n2510 ) ;
  assign n2513 = ( n2345 & ~n2511 ) | ( n2345 & n2512 ) | ( ~n2511 & n2512 ) ;
  assign n2514 = n461 & n1297 ;
  assign n2515 = x74 & n1301 ;
  assign n2516 = x75 | n2515 ;
  assign n2517 = ( n1303 & n2515 ) | ( n1303 & n2516 ) | ( n2515 & n2516 ) ;
  assign n2518 = x73 & n1426 ;
  assign n2519 = n2517 | n2518 ;
  assign n2520 = ( x23 & n2514 ) | ( x23 & ~n2519 ) | ( n2514 & ~n2519 ) ;
  assign n2521 = ( ~x23 & n2519 ) | ( ~x23 & n2520 ) | ( n2519 & n2520 ) ;
  assign n2522 = ( ~n2514 & n2520 ) | ( ~n2514 & n2521 ) | ( n2520 & n2521 ) ;
  assign n2523 = ( n2357 & n2513 ) | ( n2357 & n2522 ) | ( n2513 & n2522 ) ;
  assign n2524 = ( ~n2357 & n2513 ) | ( ~n2357 & n2522 ) | ( n2513 & n2522 ) ;
  assign n2525 = ( n2357 & ~n2523 ) | ( n2357 & n2524 ) | ( ~n2523 & n2524 ) ;
  assign n2526 = ( n2369 & n2476 ) | ( n2369 & n2525 ) | ( n2476 & n2525 ) ;
  assign n2527 = ( ~n2369 & n2476 ) | ( ~n2369 & n2525 ) | ( n2476 & n2525 ) ;
  assign n2528 = ( n2369 & ~n2526 ) | ( n2369 & n2527 ) | ( ~n2526 & n2527 ) ;
  assign n2529 = n810 & n910 ;
  assign n2530 = x80 & n814 ;
  assign n2531 = x81 | n2530 ;
  assign n2532 = ( n816 & n2530 ) | ( n816 & n2531 ) | ( n2530 & n2531 ) ;
  assign n2533 = x79 & n885 ;
  assign n2534 = n2532 | n2533 ;
  assign n2535 = ( x17 & n2529 ) | ( x17 & ~n2534 ) | ( n2529 & ~n2534 ) ;
  assign n2536 = ( ~x17 & n2534 ) | ( ~x17 & n2535 ) | ( n2534 & n2535 ) ;
  assign n2537 = ( ~n2529 & n2535 ) | ( ~n2529 & n2536 ) | ( n2535 & n2536 ) ;
  assign n2538 = ( n2381 & n2528 ) | ( n2381 & n2537 ) | ( n2528 & n2537 ) ;
  assign n2539 = ( ~n2381 & n2528 ) | ( ~n2381 & n2537 ) | ( n2528 & n2537 ) ;
  assign n2540 = ( n2381 & ~n2538 ) | ( n2381 & n2539 ) | ( ~n2538 & n2539 ) ;
  assign n2541 = n583 & n1097 ;
  assign n2542 = x83 & n587 ;
  assign n2543 = x84 | n2542 ;
  assign n2544 = ( n589 & n2542 ) | ( n589 & n2543 ) | ( n2542 & n2543 ) ;
  assign n2545 = x82 & n676 ;
  assign n2546 = n2544 | n2545 ;
  assign n2547 = ( x14 & n2541 ) | ( x14 & ~n2546 ) | ( n2541 & ~n2546 ) ;
  assign n2548 = ( ~x14 & n2546 ) | ( ~x14 & n2547 ) | ( n2546 & n2547 ) ;
  assign n2549 = ( ~n2541 & n2547 ) | ( ~n2541 & n2548 ) | ( n2547 & n2548 ) ;
  assign n2550 = ( n2393 & n2540 ) | ( n2393 & n2549 ) | ( n2540 & n2549 ) ;
  assign n2551 = ( ~n2393 & n2540 ) | ( ~n2393 & n2549 ) | ( n2540 & n2549 ) ;
  assign n2552 = ( n2393 & ~n2550 ) | ( n2393 & n2551 ) | ( ~n2550 & n2551 ) ;
  assign n2553 = ( n2405 & n2467 ) | ( n2405 & n2552 ) | ( n2467 & n2552 ) ;
  assign n2554 = ( ~n2405 & n2467 ) | ( ~n2405 & n2552 ) | ( n2467 & n2552 ) ;
  assign n2555 = ( n2405 & ~n2553 ) | ( n2405 & n2554 ) | ( ~n2553 & n2554 ) ;
  assign n2556 = n291 & n1701 ;
  assign n2557 = x89 & n295 ;
  assign n2558 = x90 | n2557 ;
  assign n2559 = ( n297 & n2557 ) | ( n297 & n2558 ) | ( n2557 & n2558 ) ;
  assign n2560 = x88 & n330 ;
  assign n2561 = n2559 | n2560 ;
  assign n2562 = ( x8 & n2556 ) | ( x8 & ~n2561 ) | ( n2556 & ~n2561 ) ;
  assign n2563 = ( ~x8 & n2561 ) | ( ~x8 & n2562 ) | ( n2561 & n2562 ) ;
  assign n2564 = ( ~n2556 & n2562 ) | ( ~n2556 & n2563 ) | ( n2562 & n2563 ) ;
  assign n2565 = ( n2417 & n2555 ) | ( n2417 & n2564 ) | ( n2555 & n2564 ) ;
  assign n2566 = ( ~n2417 & n2555 ) | ( ~n2417 & n2564 ) | ( n2555 & n2564 ) ;
  assign n2567 = ( n2417 & ~n2565 ) | ( n2417 & n2566 ) | ( ~n2565 & n2566 ) ;
  assign n2568 = n186 & n2057 ;
  assign n2569 = x92 & n190 ;
  assign n2570 = x93 | n2569 ;
  assign n2571 = ( n192 & n2569 ) | ( n192 & n2570 ) | ( n2569 & n2570 ) ;
  assign n2572 = x91 & n220 ;
  assign n2573 = n2571 | n2572 ;
  assign n2574 = ( x5 & n2568 ) | ( x5 & ~n2573 ) | ( n2568 & ~n2573 ) ;
  assign n2575 = ( ~x5 & n2573 ) | ( ~x5 & n2574 ) | ( n2573 & n2574 ) ;
  assign n2576 = ( ~n2568 & n2574 ) | ( ~n2568 & n2575 ) | ( n2574 & n2575 ) ;
  assign n2577 = ( n2429 & n2567 ) | ( n2429 & n2576 ) | ( n2567 & n2576 ) ;
  assign n2578 = ( ~n2429 & n2567 ) | ( ~n2429 & n2576 ) | ( n2567 & n2576 ) ;
  assign n2579 = ( n2429 & ~n2577 ) | ( n2429 & n2578 ) | ( ~n2577 & n2578 ) ;
  assign n2580 = ( n2444 & n2458 ) | ( n2444 & n2579 ) | ( n2458 & n2579 ) ;
  assign n2581 = ( ~n2444 & n2458 ) | ( ~n2444 & n2579 ) | ( n2458 & n2579 ) ;
  assign n2582 = ( n2444 & ~n2580 ) | ( n2444 & n2581 ) | ( ~n2580 & n2581 ) ;
  assign n2583 = ( x96 & x97 ) | ( x96 & n2447 ) | ( x97 & n2447 ) ;
  assign n2584 = ( x96 & ~x97 ) | ( x96 & n2447 ) | ( ~x97 & n2447 ) ;
  assign n2585 = ( x97 & ~n2583 ) | ( x97 & n2584 ) | ( ~n2583 & n2584 ) ;
  assign n2586 = n136 & n2585 ;
  assign n2587 = x96 & n138 ;
  assign n2588 = x97 | n2587 ;
  assign n2589 = ( n141 & n2587 ) | ( n141 & n2588 ) | ( n2587 & n2588 ) ;
  assign n2590 = x95 & n154 ;
  assign n2591 = n2589 | n2590 ;
  assign n2592 = ( x2 & n2586 ) | ( x2 & ~n2591 ) | ( n2586 & ~n2591 ) ;
  assign n2593 = ( ~x2 & n2591 ) | ( ~x2 & n2592 ) | ( n2591 & n2592 ) ;
  assign n2594 = ( ~n2586 & n2592 ) | ( ~n2586 & n2593 ) | ( n2592 & n2593 ) ;
  assign n2595 = n407 & n1481 ;
  assign n2596 = x87 & n411 ;
  assign n2597 = x88 | n2596 ;
  assign n2598 = ( n413 & n2596 ) | ( n413 & n2597 ) | ( n2596 & n2597 ) ;
  assign n2599 = x86 & n491 ;
  assign n2600 = n2598 | n2599 ;
  assign n2601 = ( x11 & n2595 ) | ( x11 & ~n2600 ) | ( n2595 & ~n2600 ) ;
  assign n2602 = ( ~x11 & n2600 ) | ( ~x11 & n2601 ) | ( n2600 & n2601 ) ;
  assign n2603 = ( ~n2595 & n2601 ) | ( ~n2595 & n2602 ) | ( n2601 & n2602 ) ;
  assign n2604 = n810 & n990 ;
  assign n2605 = x81 & n814 ;
  assign n2606 = x82 | n2605 ;
  assign n2607 = ( n816 & n2605 ) | ( n816 & n2606 ) | ( n2605 & n2606 ) ;
  assign n2608 = x80 & n885 ;
  assign n2609 = n2607 | n2608 ;
  assign n2610 = ( x17 & n2604 ) | ( x17 & ~n2609 ) | ( n2604 & ~n2609 ) ;
  assign n2611 = ( ~x17 & n2609 ) | ( ~x17 & n2610 ) | ( n2609 & n2610 ) ;
  assign n2612 = ( ~n2604 & n2610 ) | ( ~n2604 & n2611 ) | ( n2610 & n2611 ) ;
  assign n2613 = n390 & n1617 ;
  assign n2614 = x72 & n1621 ;
  assign n2615 = x73 | n2614 ;
  assign n2616 = ( n1623 & n2614 ) | ( n1623 & n2615 ) | ( n2614 & n2615 ) ;
  assign n2617 = x71 & n1749 ;
  assign n2618 = n2616 | n2617 ;
  assign n2619 = ( x26 & n2613 ) | ( x26 & ~n2618 ) | ( n2613 & ~n2618 ) ;
  assign n2620 = ( ~x26 & n2618 ) | ( ~x26 & n2619 ) | ( n2618 & n2619 ) ;
  assign n2621 = ( ~n2613 & n2619 ) | ( ~n2613 & n2620 ) | ( n2619 & n2620 ) ;
  assign n2622 = x66 & n2324 ;
  assign n2623 = x67 | n2622 ;
  assign n2624 = ( n2326 & n2622 ) | ( n2326 & n2623 ) | ( n2622 & n2623 ) ;
  assign n2625 = x65 & n2497 ;
  assign n2626 = n2624 | n2625 ;
  assign n2627 = n164 & n2320 ;
  assign n2628 = ( x32 & n2626 ) | ( x32 & ~n2627 ) | ( n2626 & ~n2627 ) ;
  assign n2629 = ( ~x32 & n2627 ) | ( ~x32 & n2628 ) | ( n2627 & n2628 ) ;
  assign n2630 = ( ~n2626 & n2628 ) | ( ~n2626 & n2629 ) | ( n2628 & n2629 ) ;
  assign n2631 = x32 & x33 ;
  assign n2632 = x32 | x33 ;
  assign n2633 = ~n2631 & n2632 ;
  assign n2634 = x64 & n2633 ;
  assign n2635 = x32 & ~n2505 ;
  assign n2636 = ( n2630 & n2634 ) | ( n2630 & n2635 ) | ( n2634 & n2635 ) ;
  assign n2637 = ( ~n2630 & n2634 ) | ( ~n2630 & n2635 ) | ( n2634 & n2635 ) ;
  assign n2638 = ( n2630 & ~n2636 ) | ( n2630 & n2637 ) | ( ~n2636 & n2637 ) ;
  assign n2639 = n245 & n1949 ;
  assign n2640 = x69 & n1953 ;
  assign n2641 = x70 | n2640 ;
  assign n2642 = ( n1955 & n2640 ) | ( n1955 & n2641 ) | ( n2640 & n2641 ) ;
  assign n2643 = x68 & n2114 ;
  assign n2644 = n2642 | n2643 ;
  assign n2645 = ( x29 & n2639 ) | ( x29 & ~n2644 ) | ( n2639 & ~n2644 ) ;
  assign n2646 = ( ~x29 & n2644 ) | ( ~x29 & n2645 ) | ( n2644 & n2645 ) ;
  assign n2647 = ( ~n2639 & n2645 ) | ( ~n2639 & n2646 ) | ( n2645 & n2646 ) ;
  assign n2648 = ( n2508 & n2638 ) | ( n2508 & n2647 ) | ( n2638 & n2647 ) ;
  assign n2649 = ( ~n2508 & n2638 ) | ( ~n2508 & n2647 ) | ( n2638 & n2647 ) ;
  assign n2650 = ( n2508 & ~n2648 ) | ( n2508 & n2649 ) | ( ~n2648 & n2649 ) ;
  assign n2651 = ( n2511 & n2621 ) | ( n2511 & n2650 ) | ( n2621 & n2650 ) ;
  assign n2652 = ( ~n2511 & n2621 ) | ( ~n2511 & n2650 ) | ( n2621 & n2650 ) ;
  assign n2653 = ( n2511 & ~n2651 ) | ( n2511 & n2652 ) | ( ~n2651 & n2652 ) ;
  assign n2654 = n554 & n1297 ;
  assign n2655 = x75 & n1301 ;
  assign n2656 = x76 | n2655 ;
  assign n2657 = ( n1303 & n2655 ) | ( n1303 & n2656 ) | ( n2655 & n2656 ) ;
  assign n2658 = x74 & n1426 ;
  assign n2659 = n2657 | n2658 ;
  assign n2660 = ( x23 & n2654 ) | ( x23 & ~n2659 ) | ( n2654 & ~n2659 ) ;
  assign n2661 = ( ~x23 & n2659 ) | ( ~x23 & n2660 ) | ( n2659 & n2660 ) ;
  assign n2662 = ( ~n2654 & n2660 ) | ( ~n2654 & n2661 ) | ( n2660 & n2661 ) ;
  assign n2663 = ( n2523 & n2653 ) | ( n2523 & n2662 ) | ( n2653 & n2662 ) ;
  assign n2664 = ( ~n2523 & n2653 ) | ( ~n2523 & n2662 ) | ( n2653 & n2662 ) ;
  assign n2665 = ( n2523 & ~n2663 ) | ( n2523 & n2664 ) | ( ~n2663 & n2664 ) ;
  assign n2666 = n701 & n1016 ;
  assign n2667 = x78 & n1020 ;
  assign n2668 = x79 | n2667 ;
  assign n2669 = ( n1022 & n2667 ) | ( n1022 & n2668 ) | ( n2667 & n2668 ) ;
  assign n2670 = x77 & n1145 ;
  assign n2671 = n2669 | n2670 ;
  assign n2672 = ( x20 & n2666 ) | ( x20 & ~n2671 ) | ( n2666 & ~n2671 ) ;
  assign n2673 = ( ~x20 & n2671 ) | ( ~x20 & n2672 ) | ( n2671 & n2672 ) ;
  assign n2674 = ( ~n2666 & n2672 ) | ( ~n2666 & n2673 ) | ( n2672 & n2673 ) ;
  assign n2675 = ( n2526 & n2665 ) | ( n2526 & n2674 ) | ( n2665 & n2674 ) ;
  assign n2676 = ( ~n2526 & n2665 ) | ( ~n2526 & n2674 ) | ( n2665 & n2674 ) ;
  assign n2677 = ( n2526 & ~n2675 ) | ( n2526 & n2676 ) | ( ~n2675 & n2676 ) ;
  assign n2678 = ( n2538 & n2612 ) | ( n2538 & n2677 ) | ( n2612 & n2677 ) ;
  assign n2679 = ( ~n2538 & n2612 ) | ( ~n2538 & n2677 ) | ( n2612 & n2677 ) ;
  assign n2680 = ( n2538 & ~n2678 ) | ( n2538 & n2679 ) | ( ~n2678 & n2679 ) ;
  assign n2681 = n583 & n1262 ;
  assign n2682 = x84 & n587 ;
  assign n2683 = x85 | n2682 ;
  assign n2684 = ( n589 & n2682 ) | ( n589 & n2683 ) | ( n2682 & n2683 ) ;
  assign n2685 = x83 & n676 ;
  assign n2686 = n2684 | n2685 ;
  assign n2687 = ( x14 & n2681 ) | ( x14 & ~n2686 ) | ( n2681 & ~n2686 ) ;
  assign n2688 = ( ~x14 & n2686 ) | ( ~x14 & n2687 ) | ( n2686 & n2687 ) ;
  assign n2689 = ( ~n2681 & n2687 ) | ( ~n2681 & n2688 ) | ( n2687 & n2688 ) ;
  assign n2690 = ( n2550 & n2680 ) | ( n2550 & n2689 ) | ( n2680 & n2689 ) ;
  assign n2691 = ( ~n2550 & n2680 ) | ( ~n2550 & n2689 ) | ( n2680 & n2689 ) ;
  assign n2692 = ( n2550 & ~n2690 ) | ( n2550 & n2691 ) | ( ~n2690 & n2691 ) ;
  assign n2693 = ( n2553 & n2603 ) | ( n2553 & n2692 ) | ( n2603 & n2692 ) ;
  assign n2694 = ( ~n2553 & n2603 ) | ( ~n2553 & n2692 ) | ( n2603 & n2692 ) ;
  assign n2695 = ( n2553 & ~n2693 ) | ( n2553 & n2694 ) | ( ~n2693 & n2694 ) ;
  assign n2696 = n291 & n1914 ;
  assign n2697 = x90 & n295 ;
  assign n2698 = x91 | n2697 ;
  assign n2699 = ( n297 & n2697 ) | ( n297 & n2698 ) | ( n2697 & n2698 ) ;
  assign n2700 = x89 & n330 ;
  assign n2701 = n2699 | n2700 ;
  assign n2702 = ( x8 & n2696 ) | ( x8 & ~n2701 ) | ( n2696 & ~n2701 ) ;
  assign n2703 = ( ~x8 & n2701 ) | ( ~x8 & n2702 ) | ( n2701 & n2702 ) ;
  assign n2704 = ( ~n2696 & n2702 ) | ( ~n2696 & n2703 ) | ( n2702 & n2703 ) ;
  assign n2705 = ( n2565 & n2695 ) | ( n2565 & n2704 ) | ( n2695 & n2704 ) ;
  assign n2706 = ( ~n2565 & n2695 ) | ( ~n2565 & n2704 ) | ( n2695 & n2704 ) ;
  assign n2707 = ( n2565 & ~n2705 ) | ( n2565 & n2706 ) | ( ~n2705 & n2706 ) ;
  assign n2708 = n186 & n2294 ;
  assign n2709 = x93 & n190 ;
  assign n2710 = x94 | n2709 ;
  assign n2711 = ( n192 & n2709 ) | ( n192 & n2710 ) | ( n2709 & n2710 ) ;
  assign n2712 = x92 & n220 ;
  assign n2713 = n2711 | n2712 ;
  assign n2714 = ( x5 & n2708 ) | ( x5 & ~n2713 ) | ( n2708 & ~n2713 ) ;
  assign n2715 = ( ~x5 & n2713 ) | ( ~x5 & n2714 ) | ( n2713 & n2714 ) ;
  assign n2716 = ( ~n2708 & n2714 ) | ( ~n2708 & n2715 ) | ( n2714 & n2715 ) ;
  assign n2717 = ( n2577 & n2707 ) | ( n2577 & n2716 ) | ( n2707 & n2716 ) ;
  assign n2718 = ( ~n2577 & n2707 ) | ( ~n2577 & n2716 ) | ( n2707 & n2716 ) ;
  assign n2719 = ( n2577 & ~n2717 ) | ( n2577 & n2718 ) | ( ~n2717 & n2718 ) ;
  assign n2720 = ( n2580 & n2594 ) | ( n2580 & n2719 ) | ( n2594 & n2719 ) ;
  assign n2721 = ( ~n2580 & n2594 ) | ( ~n2580 & n2719 ) | ( n2594 & n2719 ) ;
  assign n2722 = ( n2580 & ~n2720 ) | ( n2580 & n2721 ) | ( ~n2720 & n2721 ) ;
  assign n2723 = ( x97 & x98 ) | ( x97 & n2583 ) | ( x98 & n2583 ) ;
  assign n2724 = ( x97 & ~x98 ) | ( x97 & n2583 ) | ( ~x98 & n2583 ) ;
  assign n2725 = ( x98 & ~n2723 ) | ( x98 & n2724 ) | ( ~n2723 & n2724 ) ;
  assign n2726 = n136 & n2725 ;
  assign n2727 = x97 & n138 ;
  assign n2728 = x98 | n2727 ;
  assign n2729 = ( n141 & n2727 ) | ( n141 & n2728 ) | ( n2727 & n2728 ) ;
  assign n2730 = x96 & n154 ;
  assign n2731 = n2729 | n2730 ;
  assign n2732 = ( x2 & n2726 ) | ( x2 & ~n2731 ) | ( n2726 & ~n2731 ) ;
  assign n2733 = ( ~x2 & n2731 ) | ( ~x2 & n2732 ) | ( n2731 & n2732 ) ;
  assign n2734 = ( ~n2726 & n2732 ) | ( ~n2726 & n2733 ) | ( n2732 & n2733 ) ;
  assign n2735 = n291 & n2042 ;
  assign n2736 = x91 & n295 ;
  assign n2737 = x92 | n2736 ;
  assign n2738 = ( n297 & n2736 ) | ( n297 & n2737 ) | ( n2736 & n2737 ) ;
  assign n2739 = x90 & n330 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = ( x8 & n2735 ) | ( x8 & ~n2740 ) | ( n2735 & ~n2740 ) ;
  assign n2742 = ( ~x8 & n2740 ) | ( ~x8 & n2741 ) | ( n2740 & n2741 ) ;
  assign n2743 = ( ~n2735 & n2741 ) | ( ~n2735 & n2742 ) | ( n2741 & n2742 ) ;
  assign n2744 = n769 & n1016 ;
  assign n2745 = x79 & n1020 ;
  assign n2746 = x80 | n2745 ;
  assign n2747 = ( n1022 & n2745 ) | ( n1022 & n2746 ) | ( n2745 & n2746 ) ;
  assign n2748 = x78 & n1145 ;
  assign n2749 = n2747 | n2748 ;
  assign n2750 = ( x20 & n2744 ) | ( x20 & ~n2749 ) | ( n2744 & ~n2749 ) ;
  assign n2751 = ( ~x20 & n2749 ) | ( ~x20 & n2750 ) | ( n2749 & n2750 ) ;
  assign n2752 = ( ~n2744 & n2750 ) | ( ~n2744 & n2751 ) | ( n2750 & n2751 ) ;
  assign n2753 = n277 & n1949 ;
  assign n2754 = x70 & n1953 ;
  assign n2755 = x71 | n2754 ;
  assign n2756 = ( n1955 & n2754 ) | ( n1955 & n2755 ) | ( n2754 & n2755 ) ;
  assign n2757 = x69 & n2114 ;
  assign n2758 = n2756 | n2757 ;
  assign n2759 = ( x29 & n2753 ) | ( x29 & ~n2758 ) | ( n2753 & ~n2758 ) ;
  assign n2760 = ( ~x29 & n2758 ) | ( ~x29 & n2759 ) | ( n2758 & n2759 ) ;
  assign n2761 = ( ~n2753 & n2759 ) | ( ~n2753 & n2760 ) | ( n2759 & n2760 ) ;
  assign n2762 = x35 & n2634 ;
  assign n2763 = x34 | x35 ;
  assign n2764 = ( x34 & x35 ) | ( x34 & ~n2763 ) | ( x35 & ~n2763 ) ;
  assign n2765 = n2763 & ~n2764 ;
  assign n2766 = n2633 & n2765 ;
  assign n2767 = n133 & n2766 ;
  assign n2768 = ~x32 & x34 ;
  assign n2769 = x33 & x34 ;
  assign n2770 = ( n2631 & n2768 ) | ( n2631 & ~n2769 ) | ( n2768 & ~n2769 ) ;
  assign n2771 = x64 & n2770 ;
  assign n2772 = ( n2633 & ~n2763 ) | ( n2633 & n2764 ) | ( ~n2763 & n2764 ) ;
  assign n2773 = x65 | n2771 ;
  assign n2774 = ( n2771 & n2772 ) | ( n2771 & n2773 ) | ( n2772 & n2773 ) ;
  assign n2775 = ( n2762 & n2767 ) | ( n2762 & n2774 ) | ( n2767 & n2774 ) ;
  assign n2776 = n2767 | n2774 ;
  assign n2777 = ~n2762 & n2776 ;
  assign n2778 = ( n2762 & ~n2775 ) | ( n2762 & n2777 ) | ( ~n2775 & n2777 ) ;
  assign n2779 = x67 & n2324 ;
  assign n2780 = x68 | n2779 ;
  assign n2781 = ( n2326 & n2779 ) | ( n2326 & n2780 ) | ( n2779 & n2780 ) ;
  assign n2782 = x66 & n2497 ;
  assign n2783 = n2781 | n2782 ;
  assign n2784 = n201 & n2320 ;
  assign n2785 = ( x32 & n2783 ) | ( x32 & ~n2784 ) | ( n2783 & ~n2784 ) ;
  assign n2786 = ( ~x32 & n2784 ) | ( ~x32 & n2785 ) | ( n2784 & n2785 ) ;
  assign n2787 = ( ~n2783 & n2785 ) | ( ~n2783 & n2786 ) | ( n2785 & n2786 ) ;
  assign n2788 = ( n2636 & n2778 ) | ( n2636 & n2787 ) | ( n2778 & n2787 ) ;
  assign n2789 = ( ~n2636 & n2778 ) | ( ~n2636 & n2787 ) | ( n2778 & n2787 ) ;
  assign n2790 = ( n2636 & ~n2788 ) | ( n2636 & n2789 ) | ( ~n2788 & n2789 ) ;
  assign n2791 = ( n2648 & n2761 ) | ( n2648 & n2790 ) | ( n2761 & n2790 ) ;
  assign n2792 = ( ~n2648 & n2761 ) | ( ~n2648 & n2790 ) | ( n2761 & n2790 ) ;
  assign n2793 = ( n2648 & ~n2791 ) | ( n2648 & n2792 ) | ( ~n2791 & n2792 ) ;
  assign n2794 = n446 & n1617 ;
  assign n2795 = x73 & n1621 ;
  assign n2796 = x74 | n2795 ;
  assign n2797 = ( n1623 & n2795 ) | ( n1623 & n2796 ) | ( n2795 & n2796 ) ;
  assign n2798 = x72 & n1749 ;
  assign n2799 = n2797 | n2798 ;
  assign n2800 = ( x26 & n2794 ) | ( x26 & ~n2799 ) | ( n2794 & ~n2799 ) ;
  assign n2801 = ( ~x26 & n2799 ) | ( ~x26 & n2800 ) | ( n2799 & n2800 ) ;
  assign n2802 = ( ~n2794 & n2800 ) | ( ~n2794 & n2801 ) | ( n2800 & n2801 ) ;
  assign n2803 = ( n2651 & n2793 ) | ( n2651 & n2802 ) | ( n2793 & n2802 ) ;
  assign n2804 = ( ~n2651 & n2793 ) | ( ~n2651 & n2802 ) | ( n2793 & n2802 ) ;
  assign n2805 = ( n2651 & ~n2803 ) | ( n2651 & n2804 ) | ( ~n2803 & n2804 ) ;
  assign n2806 = n569 & n1297 ;
  assign n2807 = x76 & n1301 ;
  assign n2808 = x77 | n2807 ;
  assign n2809 = ( n1303 & n2807 ) | ( n1303 & n2808 ) | ( n2807 & n2808 ) ;
  assign n2810 = x75 & n1426 ;
  assign n2811 = n2809 | n2810 ;
  assign n2812 = ( x23 & n2806 ) | ( x23 & ~n2811 ) | ( n2806 & ~n2811 ) ;
  assign n2813 = ( ~x23 & n2811 ) | ( ~x23 & n2812 ) | ( n2811 & n2812 ) ;
  assign n2814 = ( ~n2806 & n2812 ) | ( ~n2806 & n2813 ) | ( n2812 & n2813 ) ;
  assign n2815 = ( n2663 & n2805 ) | ( n2663 & n2814 ) | ( n2805 & n2814 ) ;
  assign n2816 = ( ~n2663 & n2805 ) | ( ~n2663 & n2814 ) | ( n2805 & n2814 ) ;
  assign n2817 = ( n2663 & ~n2815 ) | ( n2663 & n2816 ) | ( ~n2815 & n2816 ) ;
  assign n2818 = ( n2675 & n2752 ) | ( n2675 & n2817 ) | ( n2752 & n2817 ) ;
  assign n2819 = ( ~n2675 & n2752 ) | ( ~n2675 & n2817 ) | ( n2752 & n2817 ) ;
  assign n2820 = ( n2675 & ~n2818 ) | ( n2675 & n2819 ) | ( ~n2818 & n2819 ) ;
  assign n2821 = n810 & n1082 ;
  assign n2822 = x82 & n814 ;
  assign n2823 = x83 | n2822 ;
  assign n2824 = ( n816 & n2822 ) | ( n816 & n2823 ) | ( n2822 & n2823 ) ;
  assign n2825 = x81 & n885 ;
  assign n2826 = n2824 | n2825 ;
  assign n2827 = ( x17 & n2821 ) | ( x17 & ~n2826 ) | ( n2821 & ~n2826 ) ;
  assign n2828 = ( ~x17 & n2826 ) | ( ~x17 & n2827 ) | ( n2826 & n2827 ) ;
  assign n2829 = ( ~n2821 & n2827 ) | ( ~n2821 & n2828 ) | ( n2827 & n2828 ) ;
  assign n2830 = ( n2678 & n2820 ) | ( n2678 & n2829 ) | ( n2820 & n2829 ) ;
  assign n2831 = ( ~n2678 & n2820 ) | ( ~n2678 & n2829 ) | ( n2820 & n2829 ) ;
  assign n2832 = ( n2678 & ~n2830 ) | ( n2678 & n2831 ) | ( ~n2830 & n2831 ) ;
  assign n2833 = n583 & n1366 ;
  assign n2834 = x85 & n587 ;
  assign n2835 = x86 | n2834 ;
  assign n2836 = ( n589 & n2834 ) | ( n589 & n2835 ) | ( n2834 & n2835 ) ;
  assign n2837 = x84 & n676 ;
  assign n2838 = n2836 | n2837 ;
  assign n2839 = ( x14 & n2833 ) | ( x14 & ~n2838 ) | ( n2833 & ~n2838 ) ;
  assign n2840 = ( ~x14 & n2838 ) | ( ~x14 & n2839 ) | ( n2838 & n2839 ) ;
  assign n2841 = ( ~n2833 & n2839 ) | ( ~n2833 & n2840 ) | ( n2839 & n2840 ) ;
  assign n2842 = ( n2690 & n2832 ) | ( n2690 & n2841 ) | ( n2832 & n2841 ) ;
  assign n2843 = ( ~n2690 & n2832 ) | ( ~n2690 & n2841 ) | ( n2832 & n2841 ) ;
  assign n2844 = ( n2690 & ~n2842 ) | ( n2690 & n2843 ) | ( ~n2842 & n2843 ) ;
  assign n2845 = n407 & n1585 ;
  assign n2846 = x88 & n411 ;
  assign n2847 = x89 | n2846 ;
  assign n2848 = ( n413 & n2846 ) | ( n413 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2849 = x87 & n491 ;
  assign n2850 = n2848 | n2849 ;
  assign n2851 = ( x11 & n2845 ) | ( x11 & ~n2850 ) | ( n2845 & ~n2850 ) ;
  assign n2852 = ( ~x11 & n2850 ) | ( ~x11 & n2851 ) | ( n2850 & n2851 ) ;
  assign n2853 = ( ~n2845 & n2851 ) | ( ~n2845 & n2852 ) | ( n2851 & n2852 ) ;
  assign n2854 = ( n2693 & n2844 ) | ( n2693 & n2853 ) | ( n2844 & n2853 ) ;
  assign n2855 = ( ~n2693 & n2844 ) | ( ~n2693 & n2853 ) | ( n2844 & n2853 ) ;
  assign n2856 = ( n2693 & ~n2854 ) | ( n2693 & n2855 ) | ( ~n2854 & n2855 ) ;
  assign n2857 = ( n2705 & n2743 ) | ( n2705 & n2856 ) | ( n2743 & n2856 ) ;
  assign n2858 = ( ~n2705 & n2743 ) | ( ~n2705 & n2856 ) | ( n2743 & n2856 ) ;
  assign n2859 = ( n2705 & ~n2857 ) | ( n2705 & n2858 ) | ( ~n2857 & n2858 ) ;
  assign n2860 = n186 & n2434 ;
  assign n2861 = x94 & n190 ;
  assign n2862 = x95 | n2861 ;
  assign n2863 = ( n192 & n2861 ) | ( n192 & n2862 ) | ( n2861 & n2862 ) ;
  assign n2864 = x93 & n220 ;
  assign n2865 = n2863 | n2864 ;
  assign n2866 = ( x5 & n2860 ) | ( x5 & ~n2865 ) | ( n2860 & ~n2865 ) ;
  assign n2867 = ( ~x5 & n2865 ) | ( ~x5 & n2866 ) | ( n2865 & n2866 ) ;
  assign n2868 = ( ~n2860 & n2866 ) | ( ~n2860 & n2867 ) | ( n2866 & n2867 ) ;
  assign n2869 = ( n2717 & n2859 ) | ( n2717 & n2868 ) | ( n2859 & n2868 ) ;
  assign n2870 = ( ~n2717 & n2859 ) | ( ~n2717 & n2868 ) | ( n2859 & n2868 ) ;
  assign n2871 = ( n2717 & ~n2869 ) | ( n2717 & n2870 ) | ( ~n2869 & n2870 ) ;
  assign n2872 = ( n2720 & n2734 ) | ( n2720 & n2871 ) | ( n2734 & n2871 ) ;
  assign n2873 = ( ~n2720 & n2734 ) | ( ~n2720 & n2871 ) | ( n2734 & n2871 ) ;
  assign n2874 = ( n2720 & ~n2872 ) | ( n2720 & n2873 ) | ( ~n2872 & n2873 ) ;
  assign n2875 = ( x98 & x99 ) | ( x98 & n2723 ) | ( x99 & n2723 ) ;
  assign n2876 = ( x98 & ~x99 ) | ( x98 & n2723 ) | ( ~x99 & n2723 ) ;
  assign n2877 = ( x99 & ~n2875 ) | ( x99 & n2876 ) | ( ~n2875 & n2876 ) ;
  assign n2878 = n136 & n2877 ;
  assign n2879 = x98 & n138 ;
  assign n2880 = x99 | n2879 ;
  assign n2881 = ( n141 & n2879 ) | ( n141 & n2880 ) | ( n2879 & n2880 ) ;
  assign n2882 = x97 & n154 ;
  assign n2883 = n2881 | n2882 ;
  assign n2884 = ( x2 & n2878 ) | ( x2 & ~n2883 ) | ( n2878 & ~n2883 ) ;
  assign n2885 = ( ~x2 & n2883 ) | ( ~x2 & n2884 ) | ( n2883 & n2884 ) ;
  assign n2886 = ( ~n2878 & n2884 ) | ( ~n2878 & n2885 ) | ( n2884 & n2885 ) ;
  assign n2887 = n407 & n1701 ;
  assign n2888 = x89 & n411 ;
  assign n2889 = x90 | n2888 ;
  assign n2890 = ( n413 & n2888 ) | ( n413 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2891 = x88 & n491 ;
  assign n2892 = n2890 | n2891 ;
  assign n2893 = ( x11 & n2887 ) | ( x11 & ~n2892 ) | ( n2887 & ~n2892 ) ;
  assign n2894 = ( ~x11 & n2892 ) | ( ~x11 & n2893 ) | ( n2892 & n2893 ) ;
  assign n2895 = ( ~n2887 & n2893 ) | ( ~n2887 & n2894 ) | ( n2893 & n2894 ) ;
  assign n2896 = n583 & n1466 ;
  assign n2897 = x86 & n587 ;
  assign n2898 = x87 | n2897 ;
  assign n2899 = ( n589 & n2897 ) | ( n589 & n2898 ) | ( n2897 & n2898 ) ;
  assign n2900 = x85 & n676 ;
  assign n2901 = n2899 | n2900 ;
  assign n2902 = ( x14 & n2896 ) | ( x14 & ~n2901 ) | ( n2896 & ~n2901 ) ;
  assign n2903 = ( ~x14 & n2901 ) | ( ~x14 & n2902 ) | ( n2901 & n2902 ) ;
  assign n2904 = ( ~n2896 & n2902 ) | ( ~n2896 & n2903 ) | ( n2902 & n2903 ) ;
  assign n2905 = n637 & n1297 ;
  assign n2906 = x77 & n1301 ;
  assign n2907 = x78 | n2906 ;
  assign n2908 = ( n1303 & n2906 ) | ( n1303 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2909 = x76 & n1426 ;
  assign n2910 = n2908 | n2909 ;
  assign n2911 = ( x23 & n2905 ) | ( x23 & ~n2910 ) | ( n2905 & ~n2910 ) ;
  assign n2912 = ( ~x23 & n2910 ) | ( ~x23 & n2911 ) | ( n2910 & n2911 ) ;
  assign n2913 = ( ~n2905 & n2911 ) | ( ~n2905 & n2912 ) | ( n2911 & n2912 ) ;
  assign n2914 = n461 & n1617 ;
  assign n2915 = x74 & n1621 ;
  assign n2916 = x75 | n2915 ;
  assign n2917 = ( n1623 & n2915 ) | ( n1623 & n2916 ) | ( n2915 & n2916 ) ;
  assign n2918 = x73 & n1749 ;
  assign n2919 = n2917 | n2918 ;
  assign n2920 = ( x26 & n2914 ) | ( x26 & ~n2919 ) | ( n2914 & ~n2919 ) ;
  assign n2921 = ( ~x26 & n2919 ) | ( ~x26 & n2920 ) | ( n2919 & n2920 ) ;
  assign n2922 = ( ~n2914 & n2920 ) | ( ~n2914 & n2921 ) | ( n2920 & n2921 ) ;
  assign n2923 = n346 & n1949 ;
  assign n2924 = x71 & n1953 ;
  assign n2925 = x72 | n2924 ;
  assign n2926 = ( n1955 & n2924 ) | ( n1955 & n2925 ) | ( n2924 & n2925 ) ;
  assign n2927 = x70 & n2114 ;
  assign n2928 = n2926 | n2927 ;
  assign n2929 = ( x29 & n2923 ) | ( x29 & ~n2928 ) | ( n2923 & ~n2928 ) ;
  assign n2930 = ( ~x29 & n2928 ) | ( ~x29 & n2929 ) | ( n2928 & n2929 ) ;
  assign n2931 = ( ~n2923 & n2929 ) | ( ~n2923 & n2930 ) | ( n2929 & n2930 ) ;
  assign n2932 = n230 & n2320 ;
  assign n2933 = x68 & n2324 ;
  assign n2934 = x69 | n2933 ;
  assign n2935 = ( n2326 & n2933 ) | ( n2326 & n2934 ) | ( n2933 & n2934 ) ;
  assign n2936 = x67 & n2497 ;
  assign n2937 = n2935 | n2936 ;
  assign n2938 = ( ~x32 & n2932 ) | ( ~x32 & n2937 ) | ( n2932 & n2937 ) ;
  assign n2939 = ( n2932 & n2937 ) | ( n2932 & ~n2938 ) | ( n2937 & ~n2938 ) ;
  assign n2940 = ( x32 & n2938 ) | ( x32 & ~n2939 ) | ( n2938 & ~n2939 ) ;
  assign n2941 = ( x35 & n2762 ) | ( x35 & n2776 ) | ( n2762 & n2776 ) ;
  assign n2942 = ( x32 & ~x34 ) | ( x32 & n2765 ) | ( ~x34 & n2765 ) ;
  assign n2943 = ( ~n2632 & n2769 ) | ( ~n2632 & n2942 ) | ( n2769 & n2942 ) ;
  assign n2944 = x64 & n2943 ;
  assign n2945 = x65 & n2770 ;
  assign n2946 = x66 | n2945 ;
  assign n2947 = ( n2772 & n2945 ) | ( n2772 & n2946 ) | ( n2945 & n2946 ) ;
  assign n2948 = ( n151 & n152 ) | ( n151 & n2766 ) | ( n152 & n2766 ) ;
  assign n2949 = ( ~n2944 & n2947 ) | ( ~n2944 & n2948 ) | ( n2947 & n2948 ) ;
  assign n2950 = n2944 | n2949 ;
  assign n2951 = n2941 | n2950 ;
  assign n2952 = ( n2941 & n2950 ) | ( n2941 & ~n2951 ) | ( n2950 & ~n2951 ) ;
  assign n2953 = n2951 & ~n2952 ;
  assign n2954 = ( n2788 & n2940 ) | ( n2788 & n2953 ) | ( n2940 & n2953 ) ;
  assign n2955 = ( ~n2788 & n2940 ) | ( ~n2788 & n2953 ) | ( n2940 & n2953 ) ;
  assign n2956 = ( n2788 & ~n2954 ) | ( n2788 & n2955 ) | ( ~n2954 & n2955 ) ;
  assign n2957 = ( n2791 & n2931 ) | ( n2791 & n2956 ) | ( n2931 & n2956 ) ;
  assign n2958 = ( ~n2791 & n2931 ) | ( ~n2791 & n2956 ) | ( n2931 & n2956 ) ;
  assign n2959 = ( n2791 & ~n2957 ) | ( n2791 & n2958 ) | ( ~n2957 & n2958 ) ;
  assign n2960 = ( n2803 & n2922 ) | ( n2803 & n2959 ) | ( n2922 & n2959 ) ;
  assign n2961 = ( ~n2803 & n2922 ) | ( ~n2803 & n2959 ) | ( n2922 & n2959 ) ;
  assign n2962 = ( n2803 & ~n2960 ) | ( n2803 & n2961 ) | ( ~n2960 & n2961 ) ;
  assign n2963 = ( n2815 & n2913 ) | ( n2815 & n2962 ) | ( n2913 & n2962 ) ;
  assign n2964 = ( ~n2815 & n2913 ) | ( ~n2815 & n2962 ) | ( n2913 & n2962 ) ;
  assign n2965 = ( n2815 & ~n2963 ) | ( n2815 & n2964 ) | ( ~n2963 & n2964 ) ;
  assign n2966 = n910 & n1016 ;
  assign n2967 = x80 & n1020 ;
  assign n2968 = x81 | n2967 ;
  assign n2969 = ( n1022 & n2967 ) | ( n1022 & n2968 ) | ( n2967 & n2968 ) ;
  assign n2970 = x79 & n1145 ;
  assign n2971 = n2969 | n2970 ;
  assign n2972 = ( x20 & n2966 ) | ( x20 & ~n2971 ) | ( n2966 & ~n2971 ) ;
  assign n2973 = ( ~x20 & n2971 ) | ( ~x20 & n2972 ) | ( n2971 & n2972 ) ;
  assign n2974 = ( ~n2966 & n2972 ) | ( ~n2966 & n2973 ) | ( n2972 & n2973 ) ;
  assign n2975 = ( n2818 & n2965 ) | ( n2818 & n2974 ) | ( n2965 & n2974 ) ;
  assign n2976 = ( ~n2818 & n2965 ) | ( ~n2818 & n2974 ) | ( n2965 & n2974 ) ;
  assign n2977 = ( n2818 & ~n2975 ) | ( n2818 & n2976 ) | ( ~n2975 & n2976 ) ;
  assign n2978 = n810 & n1097 ;
  assign n2979 = x83 & n814 ;
  assign n2980 = x84 | n2979 ;
  assign n2981 = ( n816 & n2979 ) | ( n816 & n2980 ) | ( n2979 & n2980 ) ;
  assign n2982 = x82 & n885 ;
  assign n2983 = n2981 | n2982 ;
  assign n2984 = ( x17 & n2978 ) | ( x17 & ~n2983 ) | ( n2978 & ~n2983 ) ;
  assign n2985 = ( ~x17 & n2983 ) | ( ~x17 & n2984 ) | ( n2983 & n2984 ) ;
  assign n2986 = ( ~n2978 & n2984 ) | ( ~n2978 & n2985 ) | ( n2984 & n2985 ) ;
  assign n2987 = ( n2830 & n2977 ) | ( n2830 & n2986 ) | ( n2977 & n2986 ) ;
  assign n2988 = ( ~n2830 & n2977 ) | ( ~n2830 & n2986 ) | ( n2977 & n2986 ) ;
  assign n2989 = ( n2830 & ~n2987 ) | ( n2830 & n2988 ) | ( ~n2987 & n2988 ) ;
  assign n2990 = ( n2842 & n2904 ) | ( n2842 & n2989 ) | ( n2904 & n2989 ) ;
  assign n2991 = ( ~n2842 & n2904 ) | ( ~n2842 & n2989 ) | ( n2904 & n2989 ) ;
  assign n2992 = ( n2842 & ~n2990 ) | ( n2842 & n2991 ) | ( ~n2990 & n2991 ) ;
  assign n2993 = ( n2854 & n2895 ) | ( n2854 & n2992 ) | ( n2895 & n2992 ) ;
  assign n2994 = ( ~n2854 & n2895 ) | ( ~n2854 & n2992 ) | ( n2895 & n2992 ) ;
  assign n2995 = ( n2854 & ~n2993 ) | ( n2854 & n2994 ) | ( ~n2993 & n2994 ) ;
  assign n2996 = n291 & n2057 ;
  assign n2997 = x92 & n295 ;
  assign n2998 = x93 | n2997 ;
  assign n2999 = ( n297 & n2997 ) | ( n297 & n2998 ) | ( n2997 & n2998 ) ;
  assign n3000 = x91 & n330 ;
  assign n3001 = n2999 | n3000 ;
  assign n3002 = ( x8 & n2996 ) | ( x8 & ~n3001 ) | ( n2996 & ~n3001 ) ;
  assign n3003 = ( ~x8 & n3001 ) | ( ~x8 & n3002 ) | ( n3001 & n3002 ) ;
  assign n3004 = ( ~n2996 & n3002 ) | ( ~n2996 & n3003 ) | ( n3002 & n3003 ) ;
  assign n3005 = ( n2857 & n2995 ) | ( n2857 & n3004 ) | ( n2995 & n3004 ) ;
  assign n3006 = ( ~n2857 & n2995 ) | ( ~n2857 & n3004 ) | ( n2995 & n3004 ) ;
  assign n3007 = ( n2857 & ~n3005 ) | ( n2857 & n3006 ) | ( ~n3005 & n3006 ) ;
  assign n3008 = n186 & n2449 ;
  assign n3009 = x95 & n190 ;
  assign n3010 = x96 | n3009 ;
  assign n3011 = ( n192 & n3009 ) | ( n192 & n3010 ) | ( n3009 & n3010 ) ;
  assign n3012 = x94 & n220 ;
  assign n3013 = n3011 | n3012 ;
  assign n3014 = ( x5 & n3008 ) | ( x5 & ~n3013 ) | ( n3008 & ~n3013 ) ;
  assign n3015 = ( ~x5 & n3013 ) | ( ~x5 & n3014 ) | ( n3013 & n3014 ) ;
  assign n3016 = ( ~n3008 & n3014 ) | ( ~n3008 & n3015 ) | ( n3014 & n3015 ) ;
  assign n3017 = ( n2869 & n3007 ) | ( n2869 & n3016 ) | ( n3007 & n3016 ) ;
  assign n3018 = ( ~n2869 & n3007 ) | ( ~n2869 & n3016 ) | ( n3007 & n3016 ) ;
  assign n3019 = ( n2869 & ~n3017 ) | ( n2869 & n3018 ) | ( ~n3017 & n3018 ) ;
  assign n3020 = ( n2872 & n2886 ) | ( n2872 & n3019 ) | ( n2886 & n3019 ) ;
  assign n3021 = ( ~n2872 & n2886 ) | ( ~n2872 & n3019 ) | ( n2886 & n3019 ) ;
  assign n3022 = ( n2872 & ~n3020 ) | ( n2872 & n3021 ) | ( ~n3020 & n3021 ) ;
  assign n3023 = n186 & n2585 ;
  assign n3024 = x96 & n190 ;
  assign n3025 = x97 | n3024 ;
  assign n3026 = ( n192 & n3024 ) | ( n192 & n3025 ) | ( n3024 & n3025 ) ;
  assign n3027 = x95 & n220 ;
  assign n3028 = n3026 | n3027 ;
  assign n3029 = ( x5 & n3023 ) | ( x5 & ~n3028 ) | ( n3023 & ~n3028 ) ;
  assign n3030 = ( ~x5 & n3028 ) | ( ~x5 & n3029 ) | ( n3028 & n3029 ) ;
  assign n3031 = ( ~n3023 & n3029 ) | ( ~n3023 & n3030 ) | ( n3029 & n3030 ) ;
  assign n3032 = n291 & n2294 ;
  assign n3033 = x93 & n295 ;
  assign n3034 = x94 | n3033 ;
  assign n3035 = ( n297 & n3033 ) | ( n297 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3036 = x92 & n330 ;
  assign n3037 = n3035 | n3036 ;
  assign n3038 = ( x8 & n3032 ) | ( x8 & ~n3037 ) | ( n3032 & ~n3037 ) ;
  assign n3039 = ( ~x8 & n3037 ) | ( ~x8 & n3038 ) | ( n3037 & n3038 ) ;
  assign n3040 = ( ~n3032 & n3038 ) | ( ~n3032 & n3039 ) | ( n3038 & n3039 ) ;
  assign n3041 = n583 & n1481 ;
  assign n3042 = x87 & n587 ;
  assign n3043 = x88 | n3042 ;
  assign n3044 = ( n589 & n3042 ) | ( n589 & n3043 ) | ( n3042 & n3043 ) ;
  assign n3045 = x86 & n676 ;
  assign n3046 = n3044 | n3045 ;
  assign n3047 = ( x14 & n3041 ) | ( x14 & ~n3046 ) | ( n3041 & ~n3046 ) ;
  assign n3048 = ( ~x14 & n3046 ) | ( ~x14 & n3047 ) | ( n3046 & n3047 ) ;
  assign n3049 = ( ~n3041 & n3047 ) | ( ~n3041 & n3048 ) | ( n3047 & n3048 ) ;
  assign n3050 = n990 & n1016 ;
  assign n3051 = x81 & n1020 ;
  assign n3052 = x82 | n3051 ;
  assign n3053 = ( n1022 & n3051 ) | ( n1022 & n3052 ) | ( n3051 & n3052 ) ;
  assign n3054 = x80 & n1145 ;
  assign n3055 = n3053 | n3054 ;
  assign n3056 = ( x20 & n3050 ) | ( x20 & ~n3055 ) | ( n3050 & ~n3055 ) ;
  assign n3057 = ( ~x20 & n3055 ) | ( ~x20 & n3056 ) | ( n3055 & n3056 ) ;
  assign n3058 = ( ~n3050 & n3056 ) | ( ~n3050 & n3057 ) | ( n3056 & n3057 ) ;
  assign n3059 = n390 & n1949 ;
  assign n3060 = x72 & n1953 ;
  assign n3061 = x73 | n3060 ;
  assign n3062 = ( n1955 & n3060 ) | ( n1955 & n3061 ) | ( n3060 & n3061 ) ;
  assign n3063 = x71 & n2114 ;
  assign n3064 = n3062 | n3063 ;
  assign n3065 = ( x29 & n3059 ) | ( x29 & ~n3064 ) | ( n3059 & ~n3064 ) ;
  assign n3066 = ( ~x29 & n3064 ) | ( ~x29 & n3065 ) | ( n3064 & n3065 ) ;
  assign n3067 = ( ~n3059 & n3065 ) | ( ~n3059 & n3066 ) | ( n3065 & n3066 ) ;
  assign n3068 = x66 & n2770 ;
  assign n3069 = x67 | n3068 ;
  assign n3070 = ( n2772 & n3068 ) | ( n2772 & n3069 ) | ( n3068 & n3069 ) ;
  assign n3071 = x65 & n2943 ;
  assign n3072 = n3070 | n3071 ;
  assign n3073 = n164 & n2766 ;
  assign n3074 = ( x35 & n3072 ) | ( x35 & ~n3073 ) | ( n3072 & ~n3073 ) ;
  assign n3075 = ( ~x35 & n3073 ) | ( ~x35 & n3074 ) | ( n3073 & n3074 ) ;
  assign n3076 = ( ~n3072 & n3074 ) | ( ~n3072 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3077 = x35 & x36 ;
  assign n3078 = x35 | x36 ;
  assign n3079 = ~n3077 & n3078 ;
  assign n3080 = x64 & n3079 ;
  assign n3081 = x35 & ~n2951 ;
  assign n3082 = ( n3076 & n3080 ) | ( n3076 & n3081 ) | ( n3080 & n3081 ) ;
  assign n3083 = ( ~n3076 & n3080 ) | ( ~n3076 & n3081 ) | ( n3080 & n3081 ) ;
  assign n3084 = ( n3076 & ~n3082 ) | ( n3076 & n3083 ) | ( ~n3082 & n3083 ) ;
  assign n3085 = n245 & n2320 ;
  assign n3086 = x69 & n2324 ;
  assign n3087 = x70 | n3086 ;
  assign n3088 = ( n2326 & n3086 ) | ( n2326 & n3087 ) | ( n3086 & n3087 ) ;
  assign n3089 = x68 & n2497 ;
  assign n3090 = n3088 | n3089 ;
  assign n3091 = ( x32 & n3085 ) | ( x32 & ~n3090 ) | ( n3085 & ~n3090 ) ;
  assign n3092 = ( ~x32 & n3090 ) | ( ~x32 & n3091 ) | ( n3090 & n3091 ) ;
  assign n3093 = ( ~n3085 & n3091 ) | ( ~n3085 & n3092 ) | ( n3091 & n3092 ) ;
  assign n3094 = ( n2954 & n3084 ) | ( n2954 & n3093 ) | ( n3084 & n3093 ) ;
  assign n3095 = ( ~n2954 & n3084 ) | ( ~n2954 & n3093 ) | ( n3084 & n3093 ) ;
  assign n3096 = ( n2954 & ~n3094 ) | ( n2954 & n3095 ) | ( ~n3094 & n3095 ) ;
  assign n3097 = ( n2957 & n3067 ) | ( n2957 & n3096 ) | ( n3067 & n3096 ) ;
  assign n3098 = ( ~n2957 & n3067 ) | ( ~n2957 & n3096 ) | ( n3067 & n3096 ) ;
  assign n3099 = ( n2957 & ~n3097 ) | ( n2957 & n3098 ) | ( ~n3097 & n3098 ) ;
  assign n3100 = n554 & n1617 ;
  assign n3101 = x75 & n1621 ;
  assign n3102 = x76 | n3101 ;
  assign n3103 = ( n1623 & n3101 ) | ( n1623 & n3102 ) | ( n3101 & n3102 ) ;
  assign n3104 = x74 & n1749 ;
  assign n3105 = n3103 | n3104 ;
  assign n3106 = ( x26 & n3100 ) | ( x26 & ~n3105 ) | ( n3100 & ~n3105 ) ;
  assign n3107 = ( ~x26 & n3105 ) | ( ~x26 & n3106 ) | ( n3105 & n3106 ) ;
  assign n3108 = ( ~n3100 & n3106 ) | ( ~n3100 & n3107 ) | ( n3106 & n3107 ) ;
  assign n3109 = ( n2960 & n3099 ) | ( n2960 & n3108 ) | ( n3099 & n3108 ) ;
  assign n3110 = ( n2960 & ~n3099 ) | ( n2960 & n3108 ) | ( ~n3099 & n3108 ) ;
  assign n3111 = ( n3099 & ~n3109 ) | ( n3099 & n3110 ) | ( ~n3109 & n3110 ) ;
  assign n3112 = n701 & n1297 ;
  assign n3113 = x78 & n1301 ;
  assign n3114 = x79 | n3113 ;
  assign n3115 = ( n1303 & n3113 ) | ( n1303 & n3114 ) | ( n3113 & n3114 ) ;
  assign n3116 = x77 & n1426 ;
  assign n3117 = n3115 | n3116 ;
  assign n3118 = ( x23 & n3112 ) | ( x23 & ~n3117 ) | ( n3112 & ~n3117 ) ;
  assign n3119 = ( ~x23 & n3117 ) | ( ~x23 & n3118 ) | ( n3117 & n3118 ) ;
  assign n3120 = ( ~n3112 & n3118 ) | ( ~n3112 & n3119 ) | ( n3118 & n3119 ) ;
  assign n3121 = ( n2963 & n3111 ) | ( n2963 & n3120 ) | ( n3111 & n3120 ) ;
  assign n3122 = ( ~n2963 & n3111 ) | ( ~n2963 & n3120 ) | ( n3111 & n3120 ) ;
  assign n3123 = ( n2963 & ~n3121 ) | ( n2963 & n3122 ) | ( ~n3121 & n3122 ) ;
  assign n3124 = ( n2975 & n3058 ) | ( n2975 & n3123 ) | ( n3058 & n3123 ) ;
  assign n3125 = ( ~n2975 & n3058 ) | ( ~n2975 & n3123 ) | ( n3058 & n3123 ) ;
  assign n3126 = ( n2975 & ~n3124 ) | ( n2975 & n3125 ) | ( ~n3124 & n3125 ) ;
  assign n3127 = n810 & n1262 ;
  assign n3128 = x84 & n814 ;
  assign n3129 = x85 | n3128 ;
  assign n3130 = ( n816 & n3128 ) | ( n816 & n3129 ) | ( n3128 & n3129 ) ;
  assign n3131 = x83 & n885 ;
  assign n3132 = n3130 | n3131 ;
  assign n3133 = ( x17 & n3127 ) | ( x17 & ~n3132 ) | ( n3127 & ~n3132 ) ;
  assign n3134 = ( ~x17 & n3132 ) | ( ~x17 & n3133 ) | ( n3132 & n3133 ) ;
  assign n3135 = ( ~n3127 & n3133 ) | ( ~n3127 & n3134 ) | ( n3133 & n3134 ) ;
  assign n3136 = ( n2987 & n3126 ) | ( n2987 & n3135 ) | ( n3126 & n3135 ) ;
  assign n3137 = ( ~n2987 & n3126 ) | ( ~n2987 & n3135 ) | ( n3126 & n3135 ) ;
  assign n3138 = ( n2987 & ~n3136 ) | ( n2987 & n3137 ) | ( ~n3136 & n3137 ) ;
  assign n3139 = ( n2990 & n3049 ) | ( n2990 & n3138 ) | ( n3049 & n3138 ) ;
  assign n3140 = ( ~n2990 & n3049 ) | ( ~n2990 & n3138 ) | ( n3049 & n3138 ) ;
  assign n3141 = ( n2990 & ~n3139 ) | ( n2990 & n3140 ) | ( ~n3139 & n3140 ) ;
  assign n3142 = n407 & n1914 ;
  assign n3143 = x90 & n411 ;
  assign n3144 = x91 | n3143 ;
  assign n3145 = ( n413 & n3143 ) | ( n413 & n3144 ) | ( n3143 & n3144 ) ;
  assign n3146 = x89 & n491 ;
  assign n3147 = n3145 | n3146 ;
  assign n3148 = ( x11 & n3142 ) | ( x11 & ~n3147 ) | ( n3142 & ~n3147 ) ;
  assign n3149 = ( ~x11 & n3147 ) | ( ~x11 & n3148 ) | ( n3147 & n3148 ) ;
  assign n3150 = ( ~n3142 & n3148 ) | ( ~n3142 & n3149 ) | ( n3148 & n3149 ) ;
  assign n3151 = ( n2993 & n3141 ) | ( n2993 & n3150 ) | ( n3141 & n3150 ) ;
  assign n3152 = ( ~n2993 & n3141 ) | ( ~n2993 & n3150 ) | ( n3141 & n3150 ) ;
  assign n3153 = ( n2993 & ~n3151 ) | ( n2993 & n3152 ) | ( ~n3151 & n3152 ) ;
  assign n3154 = ( n3005 & n3040 ) | ( n3005 & n3153 ) | ( n3040 & n3153 ) ;
  assign n3155 = ( ~n3005 & n3040 ) | ( ~n3005 & n3153 ) | ( n3040 & n3153 ) ;
  assign n3156 = ( n3005 & ~n3154 ) | ( n3005 & n3155 ) | ( ~n3154 & n3155 ) ;
  assign n3157 = ( n3017 & n3031 ) | ( n3017 & n3156 ) | ( n3031 & n3156 ) ;
  assign n3158 = ( ~n3017 & n3031 ) | ( ~n3017 & n3156 ) | ( n3031 & n3156 ) ;
  assign n3159 = ( n3017 & ~n3157 ) | ( n3017 & n3158 ) | ( ~n3157 & n3158 ) ;
  assign n3160 = ( x99 & x100 ) | ( x99 & n2875 ) | ( x100 & n2875 ) ;
  assign n3161 = ( x99 & ~x100 ) | ( x99 & n2875 ) | ( ~x100 & n2875 ) ;
  assign n3162 = ( x100 & ~n3160 ) | ( x100 & n3161 ) | ( ~n3160 & n3161 ) ;
  assign n3163 = n136 & n3162 ;
  assign n3164 = x99 & n138 ;
  assign n3165 = x100 | n3164 ;
  assign n3166 = ( n141 & n3164 ) | ( n141 & n3165 ) | ( n3164 & n3165 ) ;
  assign n3167 = x98 & n154 ;
  assign n3168 = n3166 | n3167 ;
  assign n3169 = ( x2 & n3163 ) | ( x2 & ~n3168 ) | ( n3163 & ~n3168 ) ;
  assign n3170 = ( ~x2 & n3168 ) | ( ~x2 & n3169 ) | ( n3168 & n3169 ) ;
  assign n3171 = ( ~n3163 & n3169 ) | ( ~n3163 & n3170 ) | ( n3169 & n3170 ) ;
  assign n3172 = ( n3020 & n3159 ) | ( n3020 & n3171 ) | ( n3159 & n3171 ) ;
  assign n3173 = ( ~n3020 & n3159 ) | ( ~n3020 & n3171 ) | ( n3159 & n3171 ) ;
  assign n3174 = ( n3020 & ~n3172 ) | ( n3020 & n3173 ) | ( ~n3172 & n3173 ) ;
  assign n3175 = n291 & n2434 ;
  assign n3176 = x94 & n295 ;
  assign n3177 = x95 | n3176 ;
  assign n3178 = ( n297 & n3176 ) | ( n297 & n3177 ) | ( n3176 & n3177 ) ;
  assign n3179 = x93 & n330 ;
  assign n3180 = n3178 | n3179 ;
  assign n3181 = ( x8 & n3175 ) | ( x8 & ~n3180 ) | ( n3175 & ~n3180 ) ;
  assign n3182 = ( ~x8 & n3180 ) | ( ~x8 & n3181 ) | ( n3180 & n3181 ) ;
  assign n3183 = ( ~n3175 & n3181 ) | ( ~n3175 & n3182 ) | ( n3181 & n3182 ) ;
  assign n3184 = n407 & n2042 ;
  assign n3185 = x91 & n411 ;
  assign n3186 = x92 | n3185 ;
  assign n3187 = ( n413 & n3185 ) | ( n413 & n3186 ) | ( n3185 & n3186 ) ;
  assign n3188 = x90 & n491 ;
  assign n3189 = n3187 | n3188 ;
  assign n3190 = ( x11 & n3184 ) | ( x11 & ~n3189 ) | ( n3184 & ~n3189 ) ;
  assign n3191 = ( ~x11 & n3189 ) | ( ~x11 & n3190 ) | ( n3189 & n3190 ) ;
  assign n3192 = ( ~n3184 & n3190 ) | ( ~n3184 & n3191 ) | ( n3190 & n3191 ) ;
  assign n3193 = n569 & n1617 ;
  assign n3194 = x76 & n1621 ;
  assign n3195 = x77 | n3194 ;
  assign n3196 = ( n1623 & n3194 ) | ( n1623 & n3195 ) | ( n3194 & n3195 ) ;
  assign n3197 = x75 & n1749 ;
  assign n3198 = n3196 | n3197 ;
  assign n3199 = ( x26 & n3193 ) | ( x26 & ~n3198 ) | ( n3193 & ~n3198 ) ;
  assign n3200 = ( ~x26 & n3198 ) | ( ~x26 & n3199 ) | ( n3198 & n3199 ) ;
  assign n3201 = ( ~n3193 & n3199 ) | ( ~n3193 & n3200 ) | ( n3199 & n3200 ) ;
  assign n3202 = n446 & n1949 ;
  assign n3203 = x73 & n1953 ;
  assign n3204 = x74 | n3203 ;
  assign n3205 = ( n1955 & n3203 ) | ( n1955 & n3204 ) | ( n3203 & n3204 ) ;
  assign n3206 = x72 & n2114 ;
  assign n3207 = n3205 | n3206 ;
  assign n3208 = ( x29 & n3202 ) | ( x29 & ~n3207 ) | ( n3202 & ~n3207 ) ;
  assign n3209 = ( ~x29 & n3207 ) | ( ~x29 & n3208 ) | ( n3207 & n3208 ) ;
  assign n3210 = ( ~n3202 & n3208 ) | ( ~n3202 & n3209 ) | ( n3208 & n3209 ) ;
  assign n3211 = n277 & n2320 ;
  assign n3212 = x70 & n2324 ;
  assign n3213 = x71 | n3212 ;
  assign n3214 = ( n2326 & n3212 ) | ( n2326 & n3213 ) | ( n3212 & n3213 ) ;
  assign n3215 = x69 & n2497 ;
  assign n3216 = n3214 | n3215 ;
  assign n3217 = ( x32 & n3211 ) | ( x32 & ~n3216 ) | ( n3211 & ~n3216 ) ;
  assign n3218 = ( ~x32 & n3216 ) | ( ~x32 & n3217 ) | ( n3216 & n3217 ) ;
  assign n3219 = ( ~n3211 & n3217 ) | ( ~n3211 & n3218 ) | ( n3217 & n3218 ) ;
  assign n3220 = x38 & n3080 ;
  assign n3221 = x37 | x38 ;
  assign n3222 = ( x37 & x38 ) | ( x37 & ~n3221 ) | ( x38 & ~n3221 ) ;
  assign n3223 = n3221 & ~n3222 ;
  assign n3224 = n3079 & n3223 ;
  assign n3225 = n133 & n3224 ;
  assign n3226 = ~x35 & x37 ;
  assign n3227 = x36 & x37 ;
  assign n3228 = ( n3077 & n3226 ) | ( n3077 & ~n3227 ) | ( n3226 & ~n3227 ) ;
  assign n3229 = x64 & n3228 ;
  assign n3230 = ( n3079 & ~n3221 ) | ( n3079 & n3222 ) | ( ~n3221 & n3222 ) ;
  assign n3231 = x65 | n3229 ;
  assign n3232 = ( n3229 & n3230 ) | ( n3229 & n3231 ) | ( n3230 & n3231 ) ;
  assign n3233 = ( n3220 & n3225 ) | ( n3220 & n3232 ) | ( n3225 & n3232 ) ;
  assign n3234 = n3225 | n3232 ;
  assign n3235 = ~n3220 & n3234 ;
  assign n3236 = ( n3220 & ~n3233 ) | ( n3220 & n3235 ) | ( ~n3233 & n3235 ) ;
  assign n3237 = x67 & n2770 ;
  assign n3238 = x68 | n3237 ;
  assign n3239 = ( n2772 & n3237 ) | ( n2772 & n3238 ) | ( n3237 & n3238 ) ;
  assign n3240 = x66 & n2943 ;
  assign n3241 = n3239 | n3240 ;
  assign n3242 = n201 & n2766 ;
  assign n3243 = ( x35 & n3241 ) | ( x35 & ~n3242 ) | ( n3241 & ~n3242 ) ;
  assign n3244 = ( ~x35 & n3242 ) | ( ~x35 & n3243 ) | ( n3242 & n3243 ) ;
  assign n3245 = ( ~n3241 & n3243 ) | ( ~n3241 & n3244 ) | ( n3243 & n3244 ) ;
  assign n3246 = ( n3082 & n3236 ) | ( n3082 & n3245 ) | ( n3236 & n3245 ) ;
  assign n3247 = ( ~n3082 & n3236 ) | ( ~n3082 & n3245 ) | ( n3236 & n3245 ) ;
  assign n3248 = ( n3082 & ~n3246 ) | ( n3082 & n3247 ) | ( ~n3246 & n3247 ) ;
  assign n3249 = ( n3094 & n3219 ) | ( n3094 & n3248 ) | ( n3219 & n3248 ) ;
  assign n3250 = ( ~n3094 & n3219 ) | ( ~n3094 & n3248 ) | ( n3219 & n3248 ) ;
  assign n3251 = ( n3094 & ~n3249 ) | ( n3094 & n3250 ) | ( ~n3249 & n3250 ) ;
  assign n3252 = ( n3097 & n3210 ) | ( n3097 & n3251 ) | ( n3210 & n3251 ) ;
  assign n3253 = ( ~n3097 & n3210 ) | ( ~n3097 & n3251 ) | ( n3210 & n3251 ) ;
  assign n3254 = ( n3097 & ~n3252 ) | ( n3097 & n3253 ) | ( ~n3252 & n3253 ) ;
  assign n3255 = ( n3109 & n3201 ) | ( n3109 & n3254 ) | ( n3201 & n3254 ) ;
  assign n3256 = ( ~n3109 & n3201 ) | ( ~n3109 & n3254 ) | ( n3201 & n3254 ) ;
  assign n3257 = ( n3109 & ~n3255 ) | ( n3109 & n3256 ) | ( ~n3255 & n3256 ) ;
  assign n3258 = n769 & n1297 ;
  assign n3259 = x79 & n1301 ;
  assign n3260 = x80 | n3259 ;
  assign n3261 = ( n1303 & n3259 ) | ( n1303 & n3260 ) | ( n3259 & n3260 ) ;
  assign n3262 = x78 & n1426 ;
  assign n3263 = n3261 | n3262 ;
  assign n3264 = ( x23 & n3258 ) | ( x23 & ~n3263 ) | ( n3258 & ~n3263 ) ;
  assign n3265 = ( ~x23 & n3263 ) | ( ~x23 & n3264 ) | ( n3263 & n3264 ) ;
  assign n3266 = ( ~n3258 & n3264 ) | ( ~n3258 & n3265 ) | ( n3264 & n3265 ) ;
  assign n3267 = ( n3121 & n3257 ) | ( n3121 & n3266 ) | ( n3257 & n3266 ) ;
  assign n3268 = ( ~n3121 & n3257 ) | ( ~n3121 & n3266 ) | ( n3257 & n3266 ) ;
  assign n3269 = ( n3121 & ~n3267 ) | ( n3121 & n3268 ) | ( ~n3267 & n3268 ) ;
  assign n3270 = n1016 & n1082 ;
  assign n3271 = x82 & n1020 ;
  assign n3272 = x83 | n3271 ;
  assign n3273 = ( n1022 & n3271 ) | ( n1022 & n3272 ) | ( n3271 & n3272 ) ;
  assign n3274 = x81 & n1145 ;
  assign n3275 = n3273 | n3274 ;
  assign n3276 = ( x20 & n3270 ) | ( x20 & ~n3275 ) | ( n3270 & ~n3275 ) ;
  assign n3277 = ( ~x20 & n3275 ) | ( ~x20 & n3276 ) | ( n3275 & n3276 ) ;
  assign n3278 = ( ~n3270 & n3276 ) | ( ~n3270 & n3277 ) | ( n3276 & n3277 ) ;
  assign n3279 = ( n3124 & n3269 ) | ( n3124 & n3278 ) | ( n3269 & n3278 ) ;
  assign n3280 = ( ~n3124 & n3269 ) | ( ~n3124 & n3278 ) | ( n3269 & n3278 ) ;
  assign n3281 = ( n3124 & ~n3279 ) | ( n3124 & n3280 ) | ( ~n3279 & n3280 ) ;
  assign n3282 = n810 & n1366 ;
  assign n3283 = x85 & n814 ;
  assign n3284 = x86 | n3283 ;
  assign n3285 = ( n816 & n3283 ) | ( n816 & n3284 ) | ( n3283 & n3284 ) ;
  assign n3286 = x84 & n885 ;
  assign n3287 = n3285 | n3286 ;
  assign n3288 = ( x17 & n3282 ) | ( x17 & ~n3287 ) | ( n3282 & ~n3287 ) ;
  assign n3289 = ( ~x17 & n3287 ) | ( ~x17 & n3288 ) | ( n3287 & n3288 ) ;
  assign n3290 = ( ~n3282 & n3288 ) | ( ~n3282 & n3289 ) | ( n3288 & n3289 ) ;
  assign n3291 = ( n3136 & n3281 ) | ( n3136 & n3290 ) | ( n3281 & n3290 ) ;
  assign n3292 = ( ~n3136 & n3281 ) | ( ~n3136 & n3290 ) | ( n3281 & n3290 ) ;
  assign n3293 = ( n3136 & ~n3291 ) | ( n3136 & n3292 ) | ( ~n3291 & n3292 ) ;
  assign n3294 = n583 & n1585 ;
  assign n3295 = x88 & n587 ;
  assign n3296 = x89 | n3295 ;
  assign n3297 = ( n589 & n3295 ) | ( n589 & n3296 ) | ( n3295 & n3296 ) ;
  assign n3298 = x87 & n676 ;
  assign n3299 = n3297 | n3298 ;
  assign n3300 = ( x14 & n3294 ) | ( x14 & ~n3299 ) | ( n3294 & ~n3299 ) ;
  assign n3301 = ( ~x14 & n3299 ) | ( ~x14 & n3300 ) | ( n3299 & n3300 ) ;
  assign n3302 = ( ~n3294 & n3300 ) | ( ~n3294 & n3301 ) | ( n3300 & n3301 ) ;
  assign n3303 = ( n3139 & n3293 ) | ( n3139 & n3302 ) | ( n3293 & n3302 ) ;
  assign n3304 = ( ~n3139 & n3293 ) | ( ~n3139 & n3302 ) | ( n3293 & n3302 ) ;
  assign n3305 = ( n3139 & ~n3303 ) | ( n3139 & n3304 ) | ( ~n3303 & n3304 ) ;
  assign n3306 = ( n3151 & n3192 ) | ( n3151 & n3305 ) | ( n3192 & n3305 ) ;
  assign n3307 = ( ~n3151 & n3192 ) | ( ~n3151 & n3305 ) | ( n3192 & n3305 ) ;
  assign n3308 = ( n3151 & ~n3306 ) | ( n3151 & n3307 ) | ( ~n3306 & n3307 ) ;
  assign n3309 = ( n3154 & n3183 ) | ( n3154 & n3308 ) | ( n3183 & n3308 ) ;
  assign n3310 = ( ~n3154 & n3183 ) | ( ~n3154 & n3308 ) | ( n3183 & n3308 ) ;
  assign n3311 = ( n3154 & ~n3309 ) | ( n3154 & n3310 ) | ( ~n3309 & n3310 ) ;
  assign n3312 = n186 & n2725 ;
  assign n3313 = x97 & n190 ;
  assign n3314 = x98 | n3313 ;
  assign n3315 = ( n192 & n3313 ) | ( n192 & n3314 ) | ( n3313 & n3314 ) ;
  assign n3316 = x96 & n220 ;
  assign n3317 = n3315 | n3316 ;
  assign n3318 = ( x5 & n3312 ) | ( x5 & ~n3317 ) | ( n3312 & ~n3317 ) ;
  assign n3319 = ( ~x5 & n3317 ) | ( ~x5 & n3318 ) | ( n3317 & n3318 ) ;
  assign n3320 = ( ~n3312 & n3318 ) | ( ~n3312 & n3319 ) | ( n3318 & n3319 ) ;
  assign n3321 = ( n3157 & n3311 ) | ( n3157 & n3320 ) | ( n3311 & n3320 ) ;
  assign n3322 = ( ~n3157 & n3311 ) | ( ~n3157 & n3320 ) | ( n3311 & n3320 ) ;
  assign n3323 = ( n3157 & ~n3321 ) | ( n3157 & n3322 ) | ( ~n3321 & n3322 ) ;
  assign n3324 = ( x100 & x101 ) | ( x100 & n3160 ) | ( x101 & n3160 ) ;
  assign n3325 = ( x100 & ~x101 ) | ( x100 & n3160 ) | ( ~x101 & n3160 ) ;
  assign n3326 = ( x101 & ~n3324 ) | ( x101 & n3325 ) | ( ~n3324 & n3325 ) ;
  assign n3327 = n136 & n3326 ;
  assign n3328 = x100 & n138 ;
  assign n3329 = x101 | n3328 ;
  assign n3330 = ( n141 & n3328 ) | ( n141 & n3329 ) | ( n3328 & n3329 ) ;
  assign n3331 = x99 & n154 ;
  assign n3332 = n3330 | n3331 ;
  assign n3333 = ( x2 & n3327 ) | ( x2 & ~n3332 ) | ( n3327 & ~n3332 ) ;
  assign n3334 = ( ~x2 & n3332 ) | ( ~x2 & n3333 ) | ( n3332 & n3333 ) ;
  assign n3335 = ( ~n3327 & n3333 ) | ( ~n3327 & n3334 ) | ( n3333 & n3334 ) ;
  assign n3336 = ( n3172 & n3323 ) | ( n3172 & n3335 ) | ( n3323 & n3335 ) ;
  assign n3337 = ( ~n3172 & n3323 ) | ( ~n3172 & n3335 ) | ( n3323 & n3335 ) ;
  assign n3338 = ( n3172 & ~n3336 ) | ( n3172 & n3337 ) | ( ~n3336 & n3337 ) ;
  assign n3339 = n186 & n2877 ;
  assign n3340 = x98 & n190 ;
  assign n3341 = x99 | n3340 ;
  assign n3342 = ( n192 & n3340 ) | ( n192 & n3341 ) | ( n3340 & n3341 ) ;
  assign n3343 = x97 & n220 ;
  assign n3344 = n3342 | n3343 ;
  assign n3345 = ( x5 & n3339 ) | ( x5 & ~n3344 ) | ( n3339 & ~n3344 ) ;
  assign n3346 = ( ~x5 & n3344 ) | ( ~x5 & n3345 ) | ( n3344 & n3345 ) ;
  assign n3347 = ( ~n3339 & n3345 ) | ( ~n3339 & n3346 ) | ( n3345 & n3346 ) ;
  assign n3348 = n291 & n2449 ;
  assign n3349 = x95 & n295 ;
  assign n3350 = x96 | n3349 ;
  assign n3351 = ( n297 & n3349 ) | ( n297 & n3350 ) | ( n3349 & n3350 ) ;
  assign n3352 = x94 & n330 ;
  assign n3353 = n3351 | n3352 ;
  assign n3354 = ( x8 & n3348 ) | ( x8 & ~n3353 ) | ( n3348 & ~n3353 ) ;
  assign n3355 = ( ~x8 & n3353 ) | ( ~x8 & n3354 ) | ( n3353 & n3354 ) ;
  assign n3356 = ( ~n3348 & n3354 ) | ( ~n3348 & n3355 ) | ( n3354 & n3355 ) ;
  assign n3357 = n407 & n2057 ;
  assign n3358 = x92 & n411 ;
  assign n3359 = x93 | n3358 ;
  assign n3360 = ( n413 & n3358 ) | ( n413 & n3359 ) | ( n3358 & n3359 ) ;
  assign n3361 = x91 & n491 ;
  assign n3362 = n3360 | n3361 ;
  assign n3363 = ( x11 & n3357 ) | ( x11 & ~n3362 ) | ( n3357 & ~n3362 ) ;
  assign n3364 = ( ~x11 & n3362 ) | ( ~x11 & n3363 ) | ( n3362 & n3363 ) ;
  assign n3365 = ( ~n3357 & n3363 ) | ( ~n3357 & n3364 ) | ( n3363 & n3364 ) ;
  assign n3366 = n583 & n1701 ;
  assign n3367 = x89 & n587 ;
  assign n3368 = x90 | n3367 ;
  assign n3369 = ( n589 & n3367 ) | ( n589 & n3368 ) | ( n3367 & n3368 ) ;
  assign n3370 = x88 & n676 ;
  assign n3371 = n3369 | n3370 ;
  assign n3372 = ( x14 & n3366 ) | ( x14 & ~n3371 ) | ( n3366 & ~n3371 ) ;
  assign n3373 = ( ~x14 & n3371 ) | ( ~x14 & n3372 ) | ( n3371 & n3372 ) ;
  assign n3374 = ( ~n3366 & n3372 ) | ( ~n3366 & n3373 ) | ( n3372 & n3373 ) ;
  assign n3375 = n637 & n1617 ;
  assign n3376 = x77 & n1621 ;
  assign n3377 = x78 | n3376 ;
  assign n3378 = ( n1623 & n3376 ) | ( n1623 & n3377 ) | ( n3376 & n3377 ) ;
  assign n3379 = x76 & n1749 ;
  assign n3380 = n3378 | n3379 ;
  assign n3381 = ( x26 & n3375 ) | ( x26 & ~n3380 ) | ( n3375 & ~n3380 ) ;
  assign n3382 = ( ~x26 & n3380 ) | ( ~x26 & n3381 ) | ( n3380 & n3381 ) ;
  assign n3383 = ( ~n3375 & n3381 ) | ( ~n3375 & n3382 ) | ( n3381 & n3382 ) ;
  assign n3384 = n461 & n1949 ;
  assign n3385 = x74 & n1953 ;
  assign n3386 = x75 | n3385 ;
  assign n3387 = ( n1955 & n3385 ) | ( n1955 & n3386 ) | ( n3385 & n3386 ) ;
  assign n3388 = x73 & n2114 ;
  assign n3389 = n3387 | n3388 ;
  assign n3390 = ( x29 & n3384 ) | ( x29 & ~n3389 ) | ( n3384 & ~n3389 ) ;
  assign n3391 = ( ~x29 & n3389 ) | ( ~x29 & n3390 ) | ( n3389 & n3390 ) ;
  assign n3392 = ( ~n3384 & n3390 ) | ( ~n3384 & n3391 ) | ( n3390 & n3391 ) ;
  assign n3393 = n346 & n2320 ;
  assign n3394 = x71 & n2324 ;
  assign n3395 = x72 | n3394 ;
  assign n3396 = ( n2326 & n3394 ) | ( n2326 & n3395 ) | ( n3394 & n3395 ) ;
  assign n3397 = x70 & n2497 ;
  assign n3398 = n3396 | n3397 ;
  assign n3399 = ( x32 & n3393 ) | ( x32 & ~n3398 ) | ( n3393 & ~n3398 ) ;
  assign n3400 = ( ~x32 & n3398 ) | ( ~x32 & n3399 ) | ( n3398 & n3399 ) ;
  assign n3401 = ( ~n3393 & n3399 ) | ( ~n3393 & n3400 ) | ( n3399 & n3400 ) ;
  assign n3402 = n230 & n2766 ;
  assign n3403 = x68 & n2770 ;
  assign n3404 = x69 | n3403 ;
  assign n3405 = ( n2772 & n3403 ) | ( n2772 & n3404 ) | ( n3403 & n3404 ) ;
  assign n3406 = x67 & n2943 ;
  assign n3407 = n3405 | n3406 ;
  assign n3408 = ( ~x35 & n3402 ) | ( ~x35 & n3407 ) | ( n3402 & n3407 ) ;
  assign n3409 = ( n3402 & n3407 ) | ( n3402 & ~n3408 ) | ( n3407 & ~n3408 ) ;
  assign n3410 = ( x35 & n3408 ) | ( x35 & ~n3409 ) | ( n3408 & ~n3409 ) ;
  assign n3411 = ( x38 & n3220 ) | ( x38 & n3234 ) | ( n3220 & n3234 ) ;
  assign n3412 = ( x35 & ~x37 ) | ( x35 & n3223 ) | ( ~x37 & n3223 ) ;
  assign n3413 = ( ~n3078 & n3227 ) | ( ~n3078 & n3412 ) | ( n3227 & n3412 ) ;
  assign n3414 = x64 & n3413 ;
  assign n3415 = x65 & n3228 ;
  assign n3416 = x66 | n3415 ;
  assign n3417 = ( n3230 & n3415 ) | ( n3230 & n3416 ) | ( n3415 & n3416 ) ;
  assign n3418 = ( n151 & n152 ) | ( n151 & n3224 ) | ( n152 & n3224 ) ;
  assign n3419 = ( ~n3414 & n3417 ) | ( ~n3414 & n3418 ) | ( n3417 & n3418 ) ;
  assign n3420 = n3414 | n3419 ;
  assign n3421 = n3411 | n3420 ;
  assign n3422 = ( n3411 & n3420 ) | ( n3411 & ~n3421 ) | ( n3420 & ~n3421 ) ;
  assign n3423 = n3421 & ~n3422 ;
  assign n3424 = ( n3246 & n3410 ) | ( n3246 & n3423 ) | ( n3410 & n3423 ) ;
  assign n3425 = ( ~n3246 & n3410 ) | ( ~n3246 & n3423 ) | ( n3410 & n3423 ) ;
  assign n3426 = ( n3246 & ~n3424 ) | ( n3246 & n3425 ) | ( ~n3424 & n3425 ) ;
  assign n3427 = ( n3249 & n3401 ) | ( n3249 & n3426 ) | ( n3401 & n3426 ) ;
  assign n3428 = ( ~n3249 & n3401 ) | ( ~n3249 & n3426 ) | ( n3401 & n3426 ) ;
  assign n3429 = ( n3249 & ~n3427 ) | ( n3249 & n3428 ) | ( ~n3427 & n3428 ) ;
  assign n3430 = ( n3252 & n3392 ) | ( n3252 & n3429 ) | ( n3392 & n3429 ) ;
  assign n3431 = ( ~n3252 & n3392 ) | ( ~n3252 & n3429 ) | ( n3392 & n3429 ) ;
  assign n3432 = ( n3252 & ~n3430 ) | ( n3252 & n3431 ) | ( ~n3430 & n3431 ) ;
  assign n3433 = ( n3255 & n3383 ) | ( n3255 & n3432 ) | ( n3383 & n3432 ) ;
  assign n3434 = ( ~n3255 & n3383 ) | ( ~n3255 & n3432 ) | ( n3383 & n3432 ) ;
  assign n3435 = ( n3255 & ~n3433 ) | ( n3255 & n3434 ) | ( ~n3433 & n3434 ) ;
  assign n3436 = n910 & n1297 ;
  assign n3437 = x80 & n1301 ;
  assign n3438 = x81 | n3437 ;
  assign n3439 = ( n1303 & n3437 ) | ( n1303 & n3438 ) | ( n3437 & n3438 ) ;
  assign n3440 = x79 & n1426 ;
  assign n3441 = n3439 | n3440 ;
  assign n3442 = ( x23 & n3436 ) | ( x23 & ~n3441 ) | ( n3436 & ~n3441 ) ;
  assign n3443 = ( ~x23 & n3441 ) | ( ~x23 & n3442 ) | ( n3441 & n3442 ) ;
  assign n3444 = ( ~n3436 & n3442 ) | ( ~n3436 & n3443 ) | ( n3442 & n3443 ) ;
  assign n3445 = ( n3267 & n3435 ) | ( n3267 & n3444 ) | ( n3435 & n3444 ) ;
  assign n3446 = ( ~n3267 & n3435 ) | ( ~n3267 & n3444 ) | ( n3435 & n3444 ) ;
  assign n3447 = ( n3267 & ~n3445 ) | ( n3267 & n3446 ) | ( ~n3445 & n3446 ) ;
  assign n3448 = n1016 & n1097 ;
  assign n3449 = x83 & n1020 ;
  assign n3450 = x84 | n3449 ;
  assign n3451 = ( n1022 & n3449 ) | ( n1022 & n3450 ) | ( n3449 & n3450 ) ;
  assign n3452 = x82 & n1145 ;
  assign n3453 = n3451 | n3452 ;
  assign n3454 = ( x20 & n3448 ) | ( x20 & ~n3453 ) | ( n3448 & ~n3453 ) ;
  assign n3455 = ( ~x20 & n3453 ) | ( ~x20 & n3454 ) | ( n3453 & n3454 ) ;
  assign n3456 = ( ~n3448 & n3454 ) | ( ~n3448 & n3455 ) | ( n3454 & n3455 ) ;
  assign n3457 = ( n3279 & n3447 ) | ( n3279 & n3456 ) | ( n3447 & n3456 ) ;
  assign n3458 = ( ~n3279 & n3447 ) | ( ~n3279 & n3456 ) | ( n3447 & n3456 ) ;
  assign n3459 = ( n3279 & ~n3457 ) | ( n3279 & n3458 ) | ( ~n3457 & n3458 ) ;
  assign n3460 = n810 & n1466 ;
  assign n3461 = x86 & n814 ;
  assign n3462 = x87 | n3461 ;
  assign n3463 = ( n816 & n3461 ) | ( n816 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3464 = x85 & n885 ;
  assign n3465 = n3463 | n3464 ;
  assign n3466 = ( x17 & n3460 ) | ( x17 & ~n3465 ) | ( n3460 & ~n3465 ) ;
  assign n3467 = ( ~x17 & n3465 ) | ( ~x17 & n3466 ) | ( n3465 & n3466 ) ;
  assign n3468 = ( ~n3460 & n3466 ) | ( ~n3460 & n3467 ) | ( n3466 & n3467 ) ;
  assign n3469 = ( n3291 & n3459 ) | ( n3291 & n3468 ) | ( n3459 & n3468 ) ;
  assign n3470 = ( ~n3291 & n3459 ) | ( ~n3291 & n3468 ) | ( n3459 & n3468 ) ;
  assign n3471 = ( n3291 & ~n3469 ) | ( n3291 & n3470 ) | ( ~n3469 & n3470 ) ;
  assign n3472 = ( n3303 & n3374 ) | ( n3303 & n3471 ) | ( n3374 & n3471 ) ;
  assign n3473 = ( ~n3303 & n3374 ) | ( ~n3303 & n3471 ) | ( n3374 & n3471 ) ;
  assign n3474 = ( n3303 & ~n3472 ) | ( n3303 & n3473 ) | ( ~n3472 & n3473 ) ;
  assign n3475 = ( n3306 & n3365 ) | ( n3306 & n3474 ) | ( n3365 & n3474 ) ;
  assign n3476 = ( ~n3306 & n3365 ) | ( ~n3306 & n3474 ) | ( n3365 & n3474 ) ;
  assign n3477 = ( n3306 & ~n3475 ) | ( n3306 & n3476 ) | ( ~n3475 & n3476 ) ;
  assign n3478 = ( n3309 & n3356 ) | ( n3309 & n3477 ) | ( n3356 & n3477 ) ;
  assign n3479 = ( ~n3309 & n3356 ) | ( ~n3309 & n3477 ) | ( n3356 & n3477 ) ;
  assign n3480 = ( n3309 & ~n3478 ) | ( n3309 & n3479 ) | ( ~n3478 & n3479 ) ;
  assign n3481 = ( n3321 & n3347 ) | ( n3321 & n3480 ) | ( n3347 & n3480 ) ;
  assign n3482 = ( ~n3321 & n3347 ) | ( ~n3321 & n3480 ) | ( n3347 & n3480 ) ;
  assign n3483 = ( n3321 & ~n3481 ) | ( n3321 & n3482 ) | ( ~n3481 & n3482 ) ;
  assign n3484 = ( x101 & x102 ) | ( x101 & n3324 ) | ( x102 & n3324 ) ;
  assign n3485 = ( x101 & ~x102 ) | ( x101 & n3324 ) | ( ~x102 & n3324 ) ;
  assign n3486 = ( x102 & ~n3484 ) | ( x102 & n3485 ) | ( ~n3484 & n3485 ) ;
  assign n3487 = n136 & n3486 ;
  assign n3488 = x101 & n138 ;
  assign n3489 = x102 | n3488 ;
  assign n3490 = ( n141 & n3488 ) | ( n141 & n3489 ) | ( n3488 & n3489 ) ;
  assign n3491 = x100 & n154 ;
  assign n3492 = n3490 | n3491 ;
  assign n3493 = ( x2 & n3487 ) | ( x2 & ~n3492 ) | ( n3487 & ~n3492 ) ;
  assign n3494 = ( ~x2 & n3492 ) | ( ~x2 & n3493 ) | ( n3492 & n3493 ) ;
  assign n3495 = ( ~n3487 & n3493 ) | ( ~n3487 & n3494 ) | ( n3493 & n3494 ) ;
  assign n3496 = ( n3336 & n3483 ) | ( n3336 & n3495 ) | ( n3483 & n3495 ) ;
  assign n3497 = ( ~n3336 & n3483 ) | ( ~n3336 & n3495 ) | ( n3483 & n3495 ) ;
  assign n3498 = ( n3336 & ~n3496 ) | ( n3336 & n3497 ) | ( ~n3496 & n3497 ) ;
  assign n3499 = n186 & n3162 ;
  assign n3500 = x99 & n190 ;
  assign n3501 = x100 | n3500 ;
  assign n3502 = ( n192 & n3500 ) | ( n192 & n3501 ) | ( n3500 & n3501 ) ;
  assign n3503 = x98 & n220 ;
  assign n3504 = n3502 | n3503 ;
  assign n3505 = ( x5 & n3499 ) | ( x5 & ~n3504 ) | ( n3499 & ~n3504 ) ;
  assign n3506 = ( ~x5 & n3504 ) | ( ~x5 & n3505 ) | ( n3504 & n3505 ) ;
  assign n3507 = ( ~n3499 & n3505 ) | ( ~n3499 & n3506 ) | ( n3505 & n3506 ) ;
  assign n3508 = n407 & n2294 ;
  assign n3509 = x93 & n411 ;
  assign n3510 = x94 | n3509 ;
  assign n3511 = ( n413 & n3509 ) | ( n413 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3512 = x92 & n491 ;
  assign n3513 = n3511 | n3512 ;
  assign n3514 = ( x11 & n3508 ) | ( x11 & ~n3513 ) | ( n3508 & ~n3513 ) ;
  assign n3515 = ( ~x11 & n3513 ) | ( ~x11 & n3514 ) | ( n3513 & n3514 ) ;
  assign n3516 = ( ~n3508 & n3514 ) | ( ~n3508 & n3515 ) | ( n3514 & n3515 ) ;
  assign n3517 = n990 & n1297 ;
  assign n3518 = x81 & n1301 ;
  assign n3519 = x82 | n3518 ;
  assign n3520 = ( n1303 & n3518 ) | ( n1303 & n3519 ) | ( n3518 & n3519 ) ;
  assign n3521 = x80 & n1426 ;
  assign n3522 = n3520 | n3521 ;
  assign n3523 = ( x23 & n3517 ) | ( x23 & ~n3522 ) | ( n3517 & ~n3522 ) ;
  assign n3524 = ( ~x23 & n3522 ) | ( ~x23 & n3523 ) | ( n3522 & n3523 ) ;
  assign n3525 = ( ~n3517 & n3523 ) | ( ~n3517 & n3524 ) | ( n3523 & n3524 ) ;
  assign n3526 = x66 & n3228 ;
  assign n3527 = x67 | n3526 ;
  assign n3528 = ( n3230 & n3526 ) | ( n3230 & n3527 ) | ( n3526 & n3527 ) ;
  assign n3529 = x65 & n3413 ;
  assign n3530 = n3528 | n3529 ;
  assign n3531 = n164 & n3224 ;
  assign n3532 = ( x38 & n3530 ) | ( x38 & ~n3531 ) | ( n3530 & ~n3531 ) ;
  assign n3533 = ( ~x38 & n3531 ) | ( ~x38 & n3532 ) | ( n3531 & n3532 ) ;
  assign n3534 = ( ~n3530 & n3532 ) | ( ~n3530 & n3533 ) | ( n3532 & n3533 ) ;
  assign n3535 = x38 & x39 ;
  assign n3536 = x38 | x39 ;
  assign n3537 = ~n3535 & n3536 ;
  assign n3538 = x64 & n3537 ;
  assign n3539 = x38 & ~n3421 ;
  assign n3540 = ( n3534 & n3538 ) | ( n3534 & n3539 ) | ( n3538 & n3539 ) ;
  assign n3541 = ( ~n3534 & n3538 ) | ( ~n3534 & n3539 ) | ( n3538 & n3539 ) ;
  assign n3542 = ( n3534 & ~n3540 ) | ( n3534 & n3541 ) | ( ~n3540 & n3541 ) ;
  assign n3543 = n245 & n2766 ;
  assign n3544 = x69 & n2770 ;
  assign n3545 = x70 | n3544 ;
  assign n3546 = ( n2772 & n3544 ) | ( n2772 & n3545 ) | ( n3544 & n3545 ) ;
  assign n3547 = x68 & n2943 ;
  assign n3548 = n3546 | n3547 ;
  assign n3549 = ( x35 & n3543 ) | ( x35 & ~n3548 ) | ( n3543 & ~n3548 ) ;
  assign n3550 = ( ~x35 & n3548 ) | ( ~x35 & n3549 ) | ( n3548 & n3549 ) ;
  assign n3551 = ( ~n3543 & n3549 ) | ( ~n3543 & n3550 ) | ( n3549 & n3550 ) ;
  assign n3552 = ( n3424 & n3542 ) | ( n3424 & n3551 ) | ( n3542 & n3551 ) ;
  assign n3553 = ( ~n3424 & n3542 ) | ( ~n3424 & n3551 ) | ( n3542 & n3551 ) ;
  assign n3554 = ( n3424 & ~n3552 ) | ( n3424 & n3553 ) | ( ~n3552 & n3553 ) ;
  assign n3555 = n390 & n2320 ;
  assign n3556 = x72 & n2324 ;
  assign n3557 = x73 | n3556 ;
  assign n3558 = ( n2326 & n3556 ) | ( n2326 & n3557 ) | ( n3556 & n3557 ) ;
  assign n3559 = x71 & n2497 ;
  assign n3560 = n3558 | n3559 ;
  assign n3561 = ( x32 & n3555 ) | ( x32 & ~n3560 ) | ( n3555 & ~n3560 ) ;
  assign n3562 = ( ~x32 & n3560 ) | ( ~x32 & n3561 ) | ( n3560 & n3561 ) ;
  assign n3563 = ( ~n3555 & n3561 ) | ( ~n3555 & n3562 ) | ( n3561 & n3562 ) ;
  assign n3564 = ( n3427 & n3554 ) | ( n3427 & n3563 ) | ( n3554 & n3563 ) ;
  assign n3565 = ( ~n3427 & n3554 ) | ( ~n3427 & n3563 ) | ( n3554 & n3563 ) ;
  assign n3566 = ( n3427 & ~n3564 ) | ( n3427 & n3565 ) | ( ~n3564 & n3565 ) ;
  assign n3567 = n554 & n1949 ;
  assign n3568 = x75 & n1953 ;
  assign n3569 = x76 | n3568 ;
  assign n3570 = ( n1955 & n3568 ) | ( n1955 & n3569 ) | ( n3568 & n3569 ) ;
  assign n3571 = x74 & n2114 ;
  assign n3572 = n3570 | n3571 ;
  assign n3573 = ( x29 & n3567 ) | ( x29 & ~n3572 ) | ( n3567 & ~n3572 ) ;
  assign n3574 = ( ~x29 & n3572 ) | ( ~x29 & n3573 ) | ( n3572 & n3573 ) ;
  assign n3575 = ( ~n3567 & n3573 ) | ( ~n3567 & n3574 ) | ( n3573 & n3574 ) ;
  assign n3576 = ( n3430 & n3566 ) | ( n3430 & n3575 ) | ( n3566 & n3575 ) ;
  assign n3577 = ( n3430 & ~n3566 ) | ( n3430 & n3575 ) | ( ~n3566 & n3575 ) ;
  assign n3578 = ( n3566 & ~n3576 ) | ( n3566 & n3577 ) | ( ~n3576 & n3577 ) ;
  assign n3579 = n701 & n1617 ;
  assign n3580 = x78 & n1621 ;
  assign n3581 = x79 | n3580 ;
  assign n3582 = ( n1623 & n3580 ) | ( n1623 & n3581 ) | ( n3580 & n3581 ) ;
  assign n3583 = x77 & n1749 ;
  assign n3584 = n3582 | n3583 ;
  assign n3585 = ( x26 & n3579 ) | ( x26 & ~n3584 ) | ( n3579 & ~n3584 ) ;
  assign n3586 = ( ~x26 & n3584 ) | ( ~x26 & n3585 ) | ( n3584 & n3585 ) ;
  assign n3587 = ( ~n3579 & n3585 ) | ( ~n3579 & n3586 ) | ( n3585 & n3586 ) ;
  assign n3588 = ( n3433 & n3578 ) | ( n3433 & n3587 ) | ( n3578 & n3587 ) ;
  assign n3589 = ( ~n3433 & n3578 ) | ( ~n3433 & n3587 ) | ( n3578 & n3587 ) ;
  assign n3590 = ( n3433 & ~n3588 ) | ( n3433 & n3589 ) | ( ~n3588 & n3589 ) ;
  assign n3591 = ( n3445 & n3525 ) | ( n3445 & n3590 ) | ( n3525 & n3590 ) ;
  assign n3592 = ( ~n3445 & n3525 ) | ( ~n3445 & n3590 ) | ( n3525 & n3590 ) ;
  assign n3593 = ( n3445 & ~n3591 ) | ( n3445 & n3592 ) | ( ~n3591 & n3592 ) ;
  assign n3594 = n1016 & n1262 ;
  assign n3595 = x84 & n1020 ;
  assign n3596 = x85 | n3595 ;
  assign n3597 = ( n1022 & n3595 ) | ( n1022 & n3596 ) | ( n3595 & n3596 ) ;
  assign n3598 = x83 & n1145 ;
  assign n3599 = n3597 | n3598 ;
  assign n3600 = ( x20 & n3594 ) | ( x20 & ~n3599 ) | ( n3594 & ~n3599 ) ;
  assign n3601 = ( ~x20 & n3599 ) | ( ~x20 & n3600 ) | ( n3599 & n3600 ) ;
  assign n3602 = ( ~n3594 & n3600 ) | ( ~n3594 & n3601 ) | ( n3600 & n3601 ) ;
  assign n3603 = ( n3457 & n3593 ) | ( n3457 & n3602 ) | ( n3593 & n3602 ) ;
  assign n3604 = ( ~n3457 & n3593 ) | ( ~n3457 & n3602 ) | ( n3593 & n3602 ) ;
  assign n3605 = ( n3457 & ~n3603 ) | ( n3457 & n3604 ) | ( ~n3603 & n3604 ) ;
  assign n3606 = n810 & n1481 ;
  assign n3607 = x87 & n814 ;
  assign n3608 = x88 | n3607 ;
  assign n3609 = ( n816 & n3607 ) | ( n816 & n3608 ) | ( n3607 & n3608 ) ;
  assign n3610 = x86 & n885 ;
  assign n3611 = n3609 | n3610 ;
  assign n3612 = ( x17 & n3606 ) | ( x17 & ~n3611 ) | ( n3606 & ~n3611 ) ;
  assign n3613 = ( ~x17 & n3611 ) | ( ~x17 & n3612 ) | ( n3611 & n3612 ) ;
  assign n3614 = ( ~n3606 & n3612 ) | ( ~n3606 & n3613 ) | ( n3612 & n3613 ) ;
  assign n3615 = ( n3469 & n3605 ) | ( n3469 & n3614 ) | ( n3605 & n3614 ) ;
  assign n3616 = ( ~n3469 & n3605 ) | ( ~n3469 & n3614 ) | ( n3605 & n3614 ) ;
  assign n3617 = ( n3469 & ~n3615 ) | ( n3469 & n3616 ) | ( ~n3615 & n3616 ) ;
  assign n3618 = n583 & n1914 ;
  assign n3619 = x90 & n587 ;
  assign n3620 = x91 | n3619 ;
  assign n3621 = ( n589 & n3619 ) | ( n589 & n3620 ) | ( n3619 & n3620 ) ;
  assign n3622 = x89 & n676 ;
  assign n3623 = n3621 | n3622 ;
  assign n3624 = ( x14 & n3618 ) | ( x14 & ~n3623 ) | ( n3618 & ~n3623 ) ;
  assign n3625 = ( ~x14 & n3623 ) | ( ~x14 & n3624 ) | ( n3623 & n3624 ) ;
  assign n3626 = ( ~n3618 & n3624 ) | ( ~n3618 & n3625 ) | ( n3624 & n3625 ) ;
  assign n3627 = ( n3472 & n3617 ) | ( n3472 & n3626 ) | ( n3617 & n3626 ) ;
  assign n3628 = ( ~n3472 & n3617 ) | ( ~n3472 & n3626 ) | ( n3617 & n3626 ) ;
  assign n3629 = ( n3472 & ~n3627 ) | ( n3472 & n3628 ) | ( ~n3627 & n3628 ) ;
  assign n3630 = ( n3475 & n3516 ) | ( n3475 & n3629 ) | ( n3516 & n3629 ) ;
  assign n3631 = ( ~n3475 & n3516 ) | ( ~n3475 & n3629 ) | ( n3516 & n3629 ) ;
  assign n3632 = ( n3475 & ~n3630 ) | ( n3475 & n3631 ) | ( ~n3630 & n3631 ) ;
  assign n3633 = n291 & n2585 ;
  assign n3634 = x96 & n295 ;
  assign n3635 = x97 | n3634 ;
  assign n3636 = ( n297 & n3634 ) | ( n297 & n3635 ) | ( n3634 & n3635 ) ;
  assign n3637 = x95 & n330 ;
  assign n3638 = n3636 | n3637 ;
  assign n3639 = ( x8 & n3633 ) | ( x8 & ~n3638 ) | ( n3633 & ~n3638 ) ;
  assign n3640 = ( ~x8 & n3638 ) | ( ~x8 & n3639 ) | ( n3638 & n3639 ) ;
  assign n3641 = ( ~n3633 & n3639 ) | ( ~n3633 & n3640 ) | ( n3639 & n3640 ) ;
  assign n3642 = ( n3478 & n3632 ) | ( n3478 & n3641 ) | ( n3632 & n3641 ) ;
  assign n3643 = ( ~n3478 & n3632 ) | ( ~n3478 & n3641 ) | ( n3632 & n3641 ) ;
  assign n3644 = ( n3478 & ~n3642 ) | ( n3478 & n3643 ) | ( ~n3642 & n3643 ) ;
  assign n3645 = ( n3481 & n3507 ) | ( n3481 & n3644 ) | ( n3507 & n3644 ) ;
  assign n3646 = ( ~n3481 & n3507 ) | ( ~n3481 & n3644 ) | ( n3507 & n3644 ) ;
  assign n3647 = ( n3481 & ~n3645 ) | ( n3481 & n3646 ) | ( ~n3645 & n3646 ) ;
  assign n3648 = ( x102 & x103 ) | ( x102 & n3484 ) | ( x103 & n3484 ) ;
  assign n3649 = ( x102 & ~x103 ) | ( x102 & n3484 ) | ( ~x103 & n3484 ) ;
  assign n3650 = ( x103 & ~n3648 ) | ( x103 & n3649 ) | ( ~n3648 & n3649 ) ;
  assign n3651 = n136 & n3650 ;
  assign n3652 = x102 & n138 ;
  assign n3653 = x103 | n3652 ;
  assign n3654 = ( n141 & n3652 ) | ( n141 & n3653 ) | ( n3652 & n3653 ) ;
  assign n3655 = x101 & n154 ;
  assign n3656 = n3654 | n3655 ;
  assign n3657 = ( x2 & n3651 ) | ( x2 & ~n3656 ) | ( n3651 & ~n3656 ) ;
  assign n3658 = ( ~x2 & n3656 ) | ( ~x2 & n3657 ) | ( n3656 & n3657 ) ;
  assign n3659 = ( ~n3651 & n3657 ) | ( ~n3651 & n3658 ) | ( n3657 & n3658 ) ;
  assign n3660 = ( n3496 & n3647 ) | ( n3496 & n3659 ) | ( n3647 & n3659 ) ;
  assign n3661 = ( ~n3496 & n3647 ) | ( ~n3496 & n3659 ) | ( n3647 & n3659 ) ;
  assign n3662 = ( n3496 & ~n3660 ) | ( n3496 & n3661 ) | ( ~n3660 & n3661 ) ;
  assign n3663 = ( x103 & x104 ) | ( x103 & n3648 ) | ( x104 & n3648 ) ;
  assign n3664 = ( x103 & ~x104 ) | ( x103 & n3648 ) | ( ~x104 & n3648 ) ;
  assign n3665 = ( x104 & ~n3663 ) | ( x104 & n3664 ) | ( ~n3663 & n3664 ) ;
  assign n3666 = n136 & n3665 ;
  assign n3667 = x103 & n138 ;
  assign n3668 = x104 | n3667 ;
  assign n3669 = ( n141 & n3667 ) | ( n141 & n3668 ) | ( n3667 & n3668 ) ;
  assign n3670 = x102 & n154 ;
  assign n3671 = n3669 | n3670 ;
  assign n3672 = ( x2 & n3666 ) | ( x2 & ~n3671 ) | ( n3666 & ~n3671 ) ;
  assign n3673 = ( ~x2 & n3671 ) | ( ~x2 & n3672 ) | ( n3671 & n3672 ) ;
  assign n3674 = ( ~n3666 & n3672 ) | ( ~n3666 & n3673 ) | ( n3672 & n3673 ) ;
  assign n3675 = n291 & n2725 ;
  assign n3676 = x97 & n295 ;
  assign n3677 = x98 | n3676 ;
  assign n3678 = ( n297 & n3676 ) | ( n297 & n3677 ) | ( n3676 & n3677 ) ;
  assign n3679 = x96 & n330 ;
  assign n3680 = n3678 | n3679 ;
  assign n3681 = ( x8 & n3675 ) | ( x8 & ~n3680 ) | ( n3675 & ~n3680 ) ;
  assign n3682 = ( ~x8 & n3680 ) | ( ~x8 & n3681 ) | ( n3680 & n3681 ) ;
  assign n3683 = ( ~n3675 & n3681 ) | ( ~n3675 & n3682 ) | ( n3681 & n3682 ) ;
  assign n3684 = n407 & n2434 ;
  assign n3685 = x94 & n411 ;
  assign n3686 = x95 | n3685 ;
  assign n3687 = ( n413 & n3685 ) | ( n413 & n3686 ) | ( n3685 & n3686 ) ;
  assign n3688 = x93 & n491 ;
  assign n3689 = n3687 | n3688 ;
  assign n3690 = ( x11 & n3684 ) | ( x11 & ~n3689 ) | ( n3684 & ~n3689 ) ;
  assign n3691 = ( ~x11 & n3689 ) | ( ~x11 & n3690 ) | ( n3689 & n3690 ) ;
  assign n3692 = ( ~n3684 & n3690 ) | ( ~n3684 & n3691 ) | ( n3690 & n3691 ) ;
  assign n3693 = n583 & n2042 ;
  assign n3694 = x91 & n587 ;
  assign n3695 = x92 | n3694 ;
  assign n3696 = ( n589 & n3694 ) | ( n589 & n3695 ) | ( n3694 & n3695 ) ;
  assign n3697 = x90 & n676 ;
  assign n3698 = n3696 | n3697 ;
  assign n3699 = ( x14 & n3693 ) | ( x14 & ~n3698 ) | ( n3693 & ~n3698 ) ;
  assign n3700 = ( ~x14 & n3698 ) | ( ~x14 & n3699 ) | ( n3698 & n3699 ) ;
  assign n3701 = ( ~n3693 & n3699 ) | ( ~n3693 & n3700 ) | ( n3699 & n3700 ) ;
  assign n3702 = n569 & n1949 ;
  assign n3703 = x76 & n1953 ;
  assign n3704 = x77 | n3703 ;
  assign n3705 = ( n1955 & n3703 ) | ( n1955 & n3704 ) | ( n3703 & n3704 ) ;
  assign n3706 = x75 & n2114 ;
  assign n3707 = n3705 | n3706 ;
  assign n3708 = ( x29 & n3702 ) | ( x29 & ~n3707 ) | ( n3702 & ~n3707 ) ;
  assign n3709 = ( ~x29 & n3707 ) | ( ~x29 & n3708 ) | ( n3707 & n3708 ) ;
  assign n3710 = ( ~n3702 & n3708 ) | ( ~n3702 & n3709 ) | ( n3708 & n3709 ) ;
  assign n3711 = x41 & n3538 ;
  assign n3712 = x40 | x41 ;
  assign n3713 = ( x40 & x41 ) | ( x40 & ~n3712 ) | ( x41 & ~n3712 ) ;
  assign n3714 = n3712 & ~n3713 ;
  assign n3715 = n3537 & n3714 ;
  assign n3716 = n133 & n3715 ;
  assign n3717 = ~x38 & x40 ;
  assign n3718 = x39 & x40 ;
  assign n3719 = ( n3535 & n3717 ) | ( n3535 & ~n3718 ) | ( n3717 & ~n3718 ) ;
  assign n3720 = x64 & n3719 ;
  assign n3721 = ( n3537 & ~n3712 ) | ( n3537 & n3713 ) | ( ~n3712 & n3713 ) ;
  assign n3722 = x65 | n3720 ;
  assign n3723 = ( n3720 & n3721 ) | ( n3720 & n3722 ) | ( n3721 & n3722 ) ;
  assign n3724 = ( n3711 & n3716 ) | ( n3711 & n3723 ) | ( n3716 & n3723 ) ;
  assign n3725 = n3716 | n3723 ;
  assign n3726 = ~n3711 & n3725 ;
  assign n3727 = ( n3711 & ~n3724 ) | ( n3711 & n3726 ) | ( ~n3724 & n3726 ) ;
  assign n3728 = x67 & n3228 ;
  assign n3729 = x68 | n3728 ;
  assign n3730 = ( n3230 & n3728 ) | ( n3230 & n3729 ) | ( n3728 & n3729 ) ;
  assign n3731 = x66 & n3413 ;
  assign n3732 = n3730 | n3731 ;
  assign n3733 = n201 & n3224 ;
  assign n3734 = ( x38 & n3732 ) | ( x38 & ~n3733 ) | ( n3732 & ~n3733 ) ;
  assign n3735 = ( ~x38 & n3733 ) | ( ~x38 & n3734 ) | ( n3733 & n3734 ) ;
  assign n3736 = ( ~n3732 & n3734 ) | ( ~n3732 & n3735 ) | ( n3734 & n3735 ) ;
  assign n3737 = ( n3540 & n3727 ) | ( n3540 & n3736 ) | ( n3727 & n3736 ) ;
  assign n3738 = ( ~n3540 & n3727 ) | ( ~n3540 & n3736 ) | ( n3727 & n3736 ) ;
  assign n3739 = ( n3540 & ~n3737 ) | ( n3540 & n3738 ) | ( ~n3737 & n3738 ) ;
  assign n3740 = n277 & n2766 ;
  assign n3741 = x70 & n2770 ;
  assign n3742 = x71 | n3741 ;
  assign n3743 = ( n2772 & n3741 ) | ( n2772 & n3742 ) | ( n3741 & n3742 ) ;
  assign n3744 = x69 & n2943 ;
  assign n3745 = n3743 | n3744 ;
  assign n3746 = ( x35 & n3740 ) | ( x35 & ~n3745 ) | ( n3740 & ~n3745 ) ;
  assign n3747 = ( ~x35 & n3745 ) | ( ~x35 & n3746 ) | ( n3745 & n3746 ) ;
  assign n3748 = ( ~n3740 & n3746 ) | ( ~n3740 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3749 = ( n3552 & n3739 ) | ( n3552 & n3748 ) | ( n3739 & n3748 ) ;
  assign n3750 = ( ~n3552 & n3739 ) | ( ~n3552 & n3748 ) | ( n3739 & n3748 ) ;
  assign n3751 = ( n3552 & ~n3749 ) | ( n3552 & n3750 ) | ( ~n3749 & n3750 ) ;
  assign n3752 = n446 & n2320 ;
  assign n3753 = x73 & n2324 ;
  assign n3754 = x74 | n3753 ;
  assign n3755 = ( n2326 & n3753 ) | ( n2326 & n3754 ) | ( n3753 & n3754 ) ;
  assign n3756 = x72 & n2497 ;
  assign n3757 = n3755 | n3756 ;
  assign n3758 = ( x32 & n3752 ) | ( x32 & ~n3757 ) | ( n3752 & ~n3757 ) ;
  assign n3759 = ( ~x32 & n3757 ) | ( ~x32 & n3758 ) | ( n3757 & n3758 ) ;
  assign n3760 = ( ~n3752 & n3758 ) | ( ~n3752 & n3759 ) | ( n3758 & n3759 ) ;
  assign n3761 = ( n3564 & n3751 ) | ( n3564 & n3760 ) | ( n3751 & n3760 ) ;
  assign n3762 = ( ~n3564 & n3751 ) | ( ~n3564 & n3760 ) | ( n3751 & n3760 ) ;
  assign n3763 = ( n3564 & ~n3761 ) | ( n3564 & n3762 ) | ( ~n3761 & n3762 ) ;
  assign n3764 = ( n3576 & n3710 ) | ( n3576 & n3763 ) | ( n3710 & n3763 ) ;
  assign n3765 = ( ~n3576 & n3710 ) | ( ~n3576 & n3763 ) | ( n3710 & n3763 ) ;
  assign n3766 = ( n3576 & ~n3764 ) | ( n3576 & n3765 ) | ( ~n3764 & n3765 ) ;
  assign n3767 = n769 & n1617 ;
  assign n3768 = x79 & n1621 ;
  assign n3769 = x80 | n3768 ;
  assign n3770 = ( n1623 & n3768 ) | ( n1623 & n3769 ) | ( n3768 & n3769 ) ;
  assign n3771 = x78 & n1749 ;
  assign n3772 = n3770 | n3771 ;
  assign n3773 = ( x26 & n3767 ) | ( x26 & ~n3772 ) | ( n3767 & ~n3772 ) ;
  assign n3774 = ( ~x26 & n3772 ) | ( ~x26 & n3773 ) | ( n3772 & n3773 ) ;
  assign n3775 = ( ~n3767 & n3773 ) | ( ~n3767 & n3774 ) | ( n3773 & n3774 ) ;
  assign n3776 = ( n3588 & n3766 ) | ( n3588 & n3775 ) | ( n3766 & n3775 ) ;
  assign n3777 = ( ~n3588 & n3766 ) | ( ~n3588 & n3775 ) | ( n3766 & n3775 ) ;
  assign n3778 = ( n3588 & ~n3776 ) | ( n3588 & n3777 ) | ( ~n3776 & n3777 ) ;
  assign n3779 = n1082 & n1297 ;
  assign n3780 = x82 & n1301 ;
  assign n3781 = x83 | n3780 ;
  assign n3782 = ( n1303 & n3780 ) | ( n1303 & n3781 ) | ( n3780 & n3781 ) ;
  assign n3783 = x81 & n1426 ;
  assign n3784 = n3782 | n3783 ;
  assign n3785 = ( x23 & n3779 ) | ( x23 & ~n3784 ) | ( n3779 & ~n3784 ) ;
  assign n3786 = ( ~x23 & n3784 ) | ( ~x23 & n3785 ) | ( n3784 & n3785 ) ;
  assign n3787 = ( ~n3779 & n3785 ) | ( ~n3779 & n3786 ) | ( n3785 & n3786 ) ;
  assign n3788 = ( n3591 & n3778 ) | ( n3591 & n3787 ) | ( n3778 & n3787 ) ;
  assign n3789 = ( ~n3591 & n3778 ) | ( ~n3591 & n3787 ) | ( n3778 & n3787 ) ;
  assign n3790 = ( n3591 & ~n3788 ) | ( n3591 & n3789 ) | ( ~n3788 & n3789 ) ;
  assign n3791 = n1016 & n1366 ;
  assign n3792 = x85 & n1020 ;
  assign n3793 = x86 | n3792 ;
  assign n3794 = ( n1022 & n3792 ) | ( n1022 & n3793 ) | ( n3792 & n3793 ) ;
  assign n3795 = x84 & n1145 ;
  assign n3796 = n3794 | n3795 ;
  assign n3797 = ( x20 & n3791 ) | ( x20 & ~n3796 ) | ( n3791 & ~n3796 ) ;
  assign n3798 = ( ~x20 & n3796 ) | ( ~x20 & n3797 ) | ( n3796 & n3797 ) ;
  assign n3799 = ( ~n3791 & n3797 ) | ( ~n3791 & n3798 ) | ( n3797 & n3798 ) ;
  assign n3800 = ( n3603 & n3790 ) | ( n3603 & n3799 ) | ( n3790 & n3799 ) ;
  assign n3801 = ( ~n3603 & n3790 ) | ( ~n3603 & n3799 ) | ( n3790 & n3799 ) ;
  assign n3802 = ( n3603 & ~n3800 ) | ( n3603 & n3801 ) | ( ~n3800 & n3801 ) ;
  assign n3803 = n810 & n1585 ;
  assign n3804 = x88 & n814 ;
  assign n3805 = x89 | n3804 ;
  assign n3806 = ( n816 & n3804 ) | ( n816 & n3805 ) | ( n3804 & n3805 ) ;
  assign n3807 = x87 & n885 ;
  assign n3808 = n3806 | n3807 ;
  assign n3809 = ( x17 & n3803 ) | ( x17 & ~n3808 ) | ( n3803 & ~n3808 ) ;
  assign n3810 = ( ~x17 & n3808 ) | ( ~x17 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3811 = ( ~n3803 & n3809 ) | ( ~n3803 & n3810 ) | ( n3809 & n3810 ) ;
  assign n3812 = ( n3615 & n3802 ) | ( n3615 & n3811 ) | ( n3802 & n3811 ) ;
  assign n3813 = ( ~n3615 & n3802 ) | ( ~n3615 & n3811 ) | ( n3802 & n3811 ) ;
  assign n3814 = ( n3615 & ~n3812 ) | ( n3615 & n3813 ) | ( ~n3812 & n3813 ) ;
  assign n3815 = ( n3627 & n3701 ) | ( n3627 & n3814 ) | ( n3701 & n3814 ) ;
  assign n3816 = ( ~n3627 & n3701 ) | ( ~n3627 & n3814 ) | ( n3701 & n3814 ) ;
  assign n3817 = ( n3627 & ~n3815 ) | ( n3627 & n3816 ) | ( ~n3815 & n3816 ) ;
  assign n3818 = ( n3630 & n3692 ) | ( n3630 & n3817 ) | ( n3692 & n3817 ) ;
  assign n3819 = ( ~n3630 & n3692 ) | ( ~n3630 & n3817 ) | ( n3692 & n3817 ) ;
  assign n3820 = ( n3630 & ~n3818 ) | ( n3630 & n3819 ) | ( ~n3818 & n3819 ) ;
  assign n3821 = ( n3642 & n3683 ) | ( n3642 & n3820 ) | ( n3683 & n3820 ) ;
  assign n3822 = ( ~n3642 & n3683 ) | ( ~n3642 & n3820 ) | ( n3683 & n3820 ) ;
  assign n3823 = ( n3642 & ~n3821 ) | ( n3642 & n3822 ) | ( ~n3821 & n3822 ) ;
  assign n3824 = n186 & n3326 ;
  assign n3825 = x100 & n190 ;
  assign n3826 = x101 | n3825 ;
  assign n3827 = ( n192 & n3825 ) | ( n192 & n3826 ) | ( n3825 & n3826 ) ;
  assign n3828 = x99 & n220 ;
  assign n3829 = n3827 | n3828 ;
  assign n3830 = ( x5 & n3824 ) | ( x5 & ~n3829 ) | ( n3824 & ~n3829 ) ;
  assign n3831 = ( ~x5 & n3829 ) | ( ~x5 & n3830 ) | ( n3829 & n3830 ) ;
  assign n3832 = ( ~n3824 & n3830 ) | ( ~n3824 & n3831 ) | ( n3830 & n3831 ) ;
  assign n3833 = ( n3645 & n3823 ) | ( n3645 & n3832 ) | ( n3823 & n3832 ) ;
  assign n3834 = ( ~n3645 & n3823 ) | ( ~n3645 & n3832 ) | ( n3823 & n3832 ) ;
  assign n3835 = ( n3645 & ~n3833 ) | ( n3645 & n3834 ) | ( ~n3833 & n3834 ) ;
  assign n3836 = ( n3660 & n3674 ) | ( n3660 & n3835 ) | ( n3674 & n3835 ) ;
  assign n3837 = ( ~n3660 & n3674 ) | ( ~n3660 & n3835 ) | ( n3674 & n3835 ) ;
  assign n3838 = ( n3660 & ~n3836 ) | ( n3660 & n3837 ) | ( ~n3836 & n3837 ) ;
  assign n3839 = n186 & n3486 ;
  assign n3840 = x101 & n190 ;
  assign n3841 = x102 | n3840 ;
  assign n3842 = ( n192 & n3840 ) | ( n192 & n3841 ) | ( n3840 & n3841 ) ;
  assign n3843 = x100 & n220 ;
  assign n3844 = n3842 | n3843 ;
  assign n3845 = ( x5 & n3839 ) | ( x5 & ~n3844 ) | ( n3839 & ~n3844 ) ;
  assign n3846 = ( ~x5 & n3844 ) | ( ~x5 & n3845 ) | ( n3844 & n3845 ) ;
  assign n3847 = ( ~n3839 & n3845 ) | ( ~n3839 & n3846 ) | ( n3845 & n3846 ) ;
  assign n3848 = n407 & n2449 ;
  assign n3849 = x95 & n411 ;
  assign n3850 = x96 | n3849 ;
  assign n3851 = ( n413 & n3849 ) | ( n413 & n3850 ) | ( n3849 & n3850 ) ;
  assign n3852 = x94 & n491 ;
  assign n3853 = n3851 | n3852 ;
  assign n3854 = ( x11 & n3848 ) | ( x11 & ~n3853 ) | ( n3848 & ~n3853 ) ;
  assign n3855 = ( ~x11 & n3853 ) | ( ~x11 & n3854 ) | ( n3853 & n3854 ) ;
  assign n3856 = ( ~n3848 & n3854 ) | ( ~n3848 & n3855 ) | ( n3854 & n3855 ) ;
  assign n3857 = n583 & n2057 ;
  assign n3858 = x92 & n587 ;
  assign n3859 = x93 | n3858 ;
  assign n3860 = ( n589 & n3858 ) | ( n589 & n3859 ) | ( n3858 & n3859 ) ;
  assign n3861 = x91 & n676 ;
  assign n3862 = n3860 | n3861 ;
  assign n3863 = ( x14 & n3857 ) | ( x14 & ~n3862 ) | ( n3857 & ~n3862 ) ;
  assign n3864 = ( ~x14 & n3862 ) | ( ~x14 & n3863 ) | ( n3862 & n3863 ) ;
  assign n3865 = ( ~n3857 & n3863 ) | ( ~n3857 & n3864 ) | ( n3863 & n3864 ) ;
  assign n3866 = n810 & n1701 ;
  assign n3867 = x89 & n814 ;
  assign n3868 = x90 | n3867 ;
  assign n3869 = ( n816 & n3867 ) | ( n816 & n3868 ) | ( n3867 & n3868 ) ;
  assign n3870 = x88 & n885 ;
  assign n3871 = n3869 | n3870 ;
  assign n3872 = ( x17 & n3866 ) | ( x17 & ~n3871 ) | ( n3866 & ~n3871 ) ;
  assign n3873 = ( ~x17 & n3871 ) | ( ~x17 & n3872 ) | ( n3871 & n3872 ) ;
  assign n3874 = ( ~n3866 & n3872 ) | ( ~n3866 & n3873 ) | ( n3872 & n3873 ) ;
  assign n3875 = n910 & n1617 ;
  assign n3876 = x80 & n1621 ;
  assign n3877 = x81 | n3876 ;
  assign n3878 = ( n1623 & n3876 ) | ( n1623 & n3877 ) | ( n3876 & n3877 ) ;
  assign n3879 = x79 & n1749 ;
  assign n3880 = n3878 | n3879 ;
  assign n3881 = ( x26 & n3875 ) | ( x26 & ~n3880 ) | ( n3875 & ~n3880 ) ;
  assign n3882 = ( ~x26 & n3880 ) | ( ~x26 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3883 = ( ~n3875 & n3881 ) | ( ~n3875 & n3882 ) | ( n3881 & n3882 ) ;
  assign n3884 = n637 & n1949 ;
  assign n3885 = x77 & n1953 ;
  assign n3886 = x78 | n3885 ;
  assign n3887 = ( n1955 & n3885 ) | ( n1955 & n3886 ) | ( n3885 & n3886 ) ;
  assign n3888 = x76 & n2114 ;
  assign n3889 = n3887 | n3888 ;
  assign n3890 = ( x29 & n3884 ) | ( x29 & ~n3889 ) | ( n3884 & ~n3889 ) ;
  assign n3891 = ( ~x29 & n3889 ) | ( ~x29 & n3890 ) | ( n3889 & n3890 ) ;
  assign n3892 = ( ~n3884 & n3890 ) | ( ~n3884 & n3891 ) | ( n3890 & n3891 ) ;
  assign n3893 = n461 & n2320 ;
  assign n3894 = x74 & n2324 ;
  assign n3895 = x75 | n3894 ;
  assign n3896 = ( n2326 & n3894 ) | ( n2326 & n3895 ) | ( n3894 & n3895 ) ;
  assign n3897 = x73 & n2497 ;
  assign n3898 = n3896 | n3897 ;
  assign n3899 = ( x32 & n3893 ) | ( x32 & ~n3898 ) | ( n3893 & ~n3898 ) ;
  assign n3900 = ( ~x32 & n3898 ) | ( ~x32 & n3899 ) | ( n3898 & n3899 ) ;
  assign n3901 = ( ~n3893 & n3899 ) | ( ~n3893 & n3900 ) | ( n3899 & n3900 ) ;
  assign n3902 = n346 & n2766 ;
  assign n3903 = x71 & n2770 ;
  assign n3904 = x72 | n3903 ;
  assign n3905 = ( n2772 & n3903 ) | ( n2772 & n3904 ) | ( n3903 & n3904 ) ;
  assign n3906 = x70 & n2943 ;
  assign n3907 = n3905 | n3906 ;
  assign n3908 = ( x35 & n3902 ) | ( x35 & ~n3907 ) | ( n3902 & ~n3907 ) ;
  assign n3909 = ( ~x35 & n3907 ) | ( ~x35 & n3908 ) | ( n3907 & n3908 ) ;
  assign n3910 = ( ~n3902 & n3908 ) | ( ~n3902 & n3909 ) | ( n3908 & n3909 ) ;
  assign n3911 = n230 & n3224 ;
  assign n3912 = x68 & n3228 ;
  assign n3913 = x69 | n3912 ;
  assign n3914 = ( n3230 & n3912 ) | ( n3230 & n3913 ) | ( n3912 & n3913 ) ;
  assign n3915 = x67 & n3413 ;
  assign n3916 = n3914 | n3915 ;
  assign n3917 = ( ~x38 & n3911 ) | ( ~x38 & n3916 ) | ( n3911 & n3916 ) ;
  assign n3918 = ( n3911 & n3916 ) | ( n3911 & ~n3917 ) | ( n3916 & ~n3917 ) ;
  assign n3919 = ( x38 & n3917 ) | ( x38 & ~n3918 ) | ( n3917 & ~n3918 ) ;
  assign n3920 = ( x41 & n3711 ) | ( x41 & n3725 ) | ( n3711 & n3725 ) ;
  assign n3921 = ( x38 & ~x40 ) | ( x38 & n3714 ) | ( ~x40 & n3714 ) ;
  assign n3922 = ( ~n3536 & n3718 ) | ( ~n3536 & n3921 ) | ( n3718 & n3921 ) ;
  assign n3923 = x64 & n3922 ;
  assign n3924 = x65 & n3719 ;
  assign n3925 = x66 | n3924 ;
  assign n3926 = ( n3721 & n3924 ) | ( n3721 & n3925 ) | ( n3924 & n3925 ) ;
  assign n3927 = ( n151 & n152 ) | ( n151 & n3715 ) | ( n152 & n3715 ) ;
  assign n3928 = ( ~n3923 & n3926 ) | ( ~n3923 & n3927 ) | ( n3926 & n3927 ) ;
  assign n3929 = n3923 | n3928 ;
  assign n3930 = n3920 | n3929 ;
  assign n3931 = ( n3920 & n3929 ) | ( n3920 & ~n3930 ) | ( n3929 & ~n3930 ) ;
  assign n3932 = n3930 & ~n3931 ;
  assign n3933 = ( n3737 & n3919 ) | ( n3737 & n3932 ) | ( n3919 & n3932 ) ;
  assign n3934 = ( ~n3737 & n3919 ) | ( ~n3737 & n3932 ) | ( n3919 & n3932 ) ;
  assign n3935 = ( n3737 & ~n3933 ) | ( n3737 & n3934 ) | ( ~n3933 & n3934 ) ;
  assign n3936 = ( n3749 & n3910 ) | ( n3749 & n3935 ) | ( n3910 & n3935 ) ;
  assign n3937 = ( ~n3749 & n3910 ) | ( ~n3749 & n3935 ) | ( n3910 & n3935 ) ;
  assign n3938 = ( n3749 & ~n3936 ) | ( n3749 & n3937 ) | ( ~n3936 & n3937 ) ;
  assign n3939 = ( n3761 & n3901 ) | ( n3761 & n3938 ) | ( n3901 & n3938 ) ;
  assign n3940 = ( ~n3761 & n3901 ) | ( ~n3761 & n3938 ) | ( n3901 & n3938 ) ;
  assign n3941 = ( n3761 & ~n3939 ) | ( n3761 & n3940 ) | ( ~n3939 & n3940 ) ;
  assign n3942 = ( n3764 & n3892 ) | ( n3764 & n3941 ) | ( n3892 & n3941 ) ;
  assign n3943 = ( ~n3764 & n3892 ) | ( ~n3764 & n3941 ) | ( n3892 & n3941 ) ;
  assign n3944 = ( n3764 & ~n3942 ) | ( n3764 & n3943 ) | ( ~n3942 & n3943 ) ;
  assign n3945 = ( n3776 & n3883 ) | ( n3776 & n3944 ) | ( n3883 & n3944 ) ;
  assign n3946 = ( ~n3776 & n3883 ) | ( ~n3776 & n3944 ) | ( n3883 & n3944 ) ;
  assign n3947 = ( n3776 & ~n3945 ) | ( n3776 & n3946 ) | ( ~n3945 & n3946 ) ;
  assign n3948 = n1097 & n1297 ;
  assign n3949 = x83 & n1301 ;
  assign n3950 = x84 | n3949 ;
  assign n3951 = ( n1303 & n3949 ) | ( n1303 & n3950 ) | ( n3949 & n3950 ) ;
  assign n3952 = x82 & n1426 ;
  assign n3953 = n3951 | n3952 ;
  assign n3954 = ( x23 & n3948 ) | ( x23 & ~n3953 ) | ( n3948 & ~n3953 ) ;
  assign n3955 = ( ~x23 & n3953 ) | ( ~x23 & n3954 ) | ( n3953 & n3954 ) ;
  assign n3956 = ( ~n3948 & n3954 ) | ( ~n3948 & n3955 ) | ( n3954 & n3955 ) ;
  assign n3957 = ( n3788 & n3947 ) | ( n3788 & n3956 ) | ( n3947 & n3956 ) ;
  assign n3958 = ( ~n3788 & n3947 ) | ( ~n3788 & n3956 ) | ( n3947 & n3956 ) ;
  assign n3959 = ( n3788 & ~n3957 ) | ( n3788 & n3958 ) | ( ~n3957 & n3958 ) ;
  assign n3960 = n1016 & n1466 ;
  assign n3961 = x86 & n1020 ;
  assign n3962 = x87 | n3961 ;
  assign n3963 = ( n1022 & n3961 ) | ( n1022 & n3962 ) | ( n3961 & n3962 ) ;
  assign n3964 = x85 & n1145 ;
  assign n3965 = n3963 | n3964 ;
  assign n3966 = ( x20 & n3960 ) | ( x20 & ~n3965 ) | ( n3960 & ~n3965 ) ;
  assign n3967 = ( ~x20 & n3965 ) | ( ~x20 & n3966 ) | ( n3965 & n3966 ) ;
  assign n3968 = ( ~n3960 & n3966 ) | ( ~n3960 & n3967 ) | ( n3966 & n3967 ) ;
  assign n3969 = ( n3800 & n3959 ) | ( n3800 & n3968 ) | ( n3959 & n3968 ) ;
  assign n3970 = ( ~n3800 & n3959 ) | ( ~n3800 & n3968 ) | ( n3959 & n3968 ) ;
  assign n3971 = ( n3800 & ~n3969 ) | ( n3800 & n3970 ) | ( ~n3969 & n3970 ) ;
  assign n3972 = ( n3812 & n3874 ) | ( n3812 & n3971 ) | ( n3874 & n3971 ) ;
  assign n3973 = ( ~n3812 & n3874 ) | ( ~n3812 & n3971 ) | ( n3874 & n3971 ) ;
  assign n3974 = ( n3812 & ~n3972 ) | ( n3812 & n3973 ) | ( ~n3972 & n3973 ) ;
  assign n3975 = ( n3815 & n3865 ) | ( n3815 & n3974 ) | ( n3865 & n3974 ) ;
  assign n3976 = ( ~n3815 & n3865 ) | ( ~n3815 & n3974 ) | ( n3865 & n3974 ) ;
  assign n3977 = ( n3815 & ~n3975 ) | ( n3815 & n3976 ) | ( ~n3975 & n3976 ) ;
  assign n3978 = ( n3818 & n3856 ) | ( n3818 & n3977 ) | ( n3856 & n3977 ) ;
  assign n3979 = ( ~n3818 & n3856 ) | ( ~n3818 & n3977 ) | ( n3856 & n3977 ) ;
  assign n3980 = ( n3818 & ~n3978 ) | ( n3818 & n3979 ) | ( ~n3978 & n3979 ) ;
  assign n3981 = n291 & n2877 ;
  assign n3982 = x98 & n295 ;
  assign n3983 = x99 | n3982 ;
  assign n3984 = ( n297 & n3982 ) | ( n297 & n3983 ) | ( n3982 & n3983 ) ;
  assign n3985 = x97 & n330 ;
  assign n3986 = n3984 | n3985 ;
  assign n3987 = ( x8 & n3981 ) | ( x8 & ~n3986 ) | ( n3981 & ~n3986 ) ;
  assign n3988 = ( ~x8 & n3986 ) | ( ~x8 & n3987 ) | ( n3986 & n3987 ) ;
  assign n3989 = ( ~n3981 & n3987 ) | ( ~n3981 & n3988 ) | ( n3987 & n3988 ) ;
  assign n3990 = ( n3821 & n3980 ) | ( n3821 & n3989 ) | ( n3980 & n3989 ) ;
  assign n3991 = ( ~n3821 & n3980 ) | ( ~n3821 & n3989 ) | ( n3980 & n3989 ) ;
  assign n3992 = ( n3821 & ~n3990 ) | ( n3821 & n3991 ) | ( ~n3990 & n3991 ) ;
  assign n3993 = ( n3833 & n3847 ) | ( n3833 & n3992 ) | ( n3847 & n3992 ) ;
  assign n3994 = ( ~n3833 & n3847 ) | ( ~n3833 & n3992 ) | ( n3847 & n3992 ) ;
  assign n3995 = ( n3833 & ~n3993 ) | ( n3833 & n3994 ) | ( ~n3993 & n3994 ) ;
  assign n3996 = ( x104 & x105 ) | ( x104 & n3663 ) | ( x105 & n3663 ) ;
  assign n3997 = ( x104 & ~x105 ) | ( x104 & n3663 ) | ( ~x105 & n3663 ) ;
  assign n3998 = ( x105 & ~n3996 ) | ( x105 & n3997 ) | ( ~n3996 & n3997 ) ;
  assign n3999 = n136 & n3998 ;
  assign n4000 = x104 & n138 ;
  assign n4001 = x105 | n4000 ;
  assign n4002 = ( n141 & n4000 ) | ( n141 & n4001 ) | ( n4000 & n4001 ) ;
  assign n4003 = x103 & n154 ;
  assign n4004 = n4002 | n4003 ;
  assign n4005 = ( x2 & n3999 ) | ( x2 & ~n4004 ) | ( n3999 & ~n4004 ) ;
  assign n4006 = ( ~x2 & n4004 ) | ( ~x2 & n4005 ) | ( n4004 & n4005 ) ;
  assign n4007 = ( ~n3999 & n4005 ) | ( ~n3999 & n4006 ) | ( n4005 & n4006 ) ;
  assign n4008 = ( n3836 & n3995 ) | ( n3836 & n4007 ) | ( n3995 & n4007 ) ;
  assign n4009 = ( ~n3836 & n3995 ) | ( ~n3836 & n4007 ) | ( n3995 & n4007 ) ;
  assign n4010 = ( n3836 & ~n4008 ) | ( n3836 & n4009 ) | ( ~n4008 & n4009 ) ;
  assign n4011 = ( x105 & x106 ) | ( x105 & n3996 ) | ( x106 & n3996 ) ;
  assign n4012 = ( x105 & ~x106 ) | ( x105 & n3996 ) | ( ~x106 & n3996 ) ;
  assign n4013 = ( x106 & ~n4011 ) | ( x106 & n4012 ) | ( ~n4011 & n4012 ) ;
  assign n4014 = n136 & n4013 ;
  assign n4015 = x105 & n138 ;
  assign n4016 = x106 | n4015 ;
  assign n4017 = ( n141 & n4015 ) | ( n141 & n4016 ) | ( n4015 & n4016 ) ;
  assign n4018 = x104 & n154 ;
  assign n4019 = n4017 | n4018 ;
  assign n4020 = ( x2 & n4014 ) | ( x2 & ~n4019 ) | ( n4014 & ~n4019 ) ;
  assign n4021 = ( ~x2 & n4019 ) | ( ~x2 & n4020 ) | ( n4019 & n4020 ) ;
  assign n4022 = ( ~n4014 & n4020 ) | ( ~n4014 & n4021 ) | ( n4020 & n4021 ) ;
  assign n4023 = n186 & n3650 ;
  assign n4024 = x102 & n190 ;
  assign n4025 = x103 | n4024 ;
  assign n4026 = ( n192 & n4024 ) | ( n192 & n4025 ) | ( n4024 & n4025 ) ;
  assign n4027 = x101 & n220 ;
  assign n4028 = n4026 | n4027 ;
  assign n4029 = ( x5 & n4023 ) | ( x5 & ~n4028 ) | ( n4023 & ~n4028 ) ;
  assign n4030 = ( ~x5 & n4028 ) | ( ~x5 & n4029 ) | ( n4028 & n4029 ) ;
  assign n4031 = ( ~n4023 & n4029 ) | ( ~n4023 & n4030 ) | ( n4029 & n4030 ) ;
  assign n4032 = n291 & n3162 ;
  assign n4033 = x99 & n295 ;
  assign n4034 = x100 | n4033 ;
  assign n4035 = ( n297 & n4033 ) | ( n297 & n4034 ) | ( n4033 & n4034 ) ;
  assign n4036 = x98 & n330 ;
  assign n4037 = n4035 | n4036 ;
  assign n4038 = ( x8 & n4032 ) | ( x8 & ~n4037 ) | ( n4032 & ~n4037 ) ;
  assign n4039 = ( ~x8 & n4037 ) | ( ~x8 & n4038 ) | ( n4037 & n4038 ) ;
  assign n4040 = ( ~n4032 & n4038 ) | ( ~n4032 & n4039 ) | ( n4038 & n4039 ) ;
  assign n4041 = n583 & n2294 ;
  assign n4042 = x93 & n587 ;
  assign n4043 = x94 | n4042 ;
  assign n4044 = ( n589 & n4042 ) | ( n589 & n4043 ) | ( n4042 & n4043 ) ;
  assign n4045 = x92 & n676 ;
  assign n4046 = n4044 | n4045 ;
  assign n4047 = ( x14 & n4041 ) | ( x14 & ~n4046 ) | ( n4041 & ~n4046 ) ;
  assign n4048 = ( ~x14 & n4046 ) | ( ~x14 & n4047 ) | ( n4046 & n4047 ) ;
  assign n4049 = ( ~n4041 & n4047 ) | ( ~n4041 & n4048 ) | ( n4047 & n4048 ) ;
  assign n4050 = n990 & n1617 ;
  assign n4051 = x81 & n1621 ;
  assign n4052 = x82 | n4051 ;
  assign n4053 = ( n1623 & n4051 ) | ( n1623 & n4052 ) | ( n4051 & n4052 ) ;
  assign n4054 = x80 & n1749 ;
  assign n4055 = n4053 | n4054 ;
  assign n4056 = ( x26 & n4050 ) | ( x26 & ~n4055 ) | ( n4050 & ~n4055 ) ;
  assign n4057 = ( ~x26 & n4055 ) | ( ~x26 & n4056 ) | ( n4055 & n4056 ) ;
  assign n4058 = ( ~n4050 & n4056 ) | ( ~n4050 & n4057 ) | ( n4056 & n4057 ) ;
  assign n4059 = n701 & n1949 ;
  assign n4060 = x78 & n1953 ;
  assign n4061 = x79 | n4060 ;
  assign n4062 = ( n1955 & n4060 ) | ( n1955 & n4061 ) | ( n4060 & n4061 ) ;
  assign n4063 = x77 & n2114 ;
  assign n4064 = n4062 | n4063 ;
  assign n4065 = ( x29 & n4059 ) | ( x29 & ~n4064 ) | ( n4059 & ~n4064 ) ;
  assign n4066 = ( ~x29 & n4064 ) | ( ~x29 & n4065 ) | ( n4064 & n4065 ) ;
  assign n4067 = ( ~n4059 & n4065 ) | ( ~n4059 & n4066 ) | ( n4065 & n4066 ) ;
  assign n4068 = n554 & n2320 ;
  assign n4069 = x75 & n2324 ;
  assign n4070 = x76 | n4069 ;
  assign n4071 = ( n2326 & n4069 ) | ( n2326 & n4070 ) | ( n4069 & n4070 ) ;
  assign n4072 = x74 & n2497 ;
  assign n4073 = n4071 | n4072 ;
  assign n4074 = ( x32 & n4068 ) | ( x32 & ~n4073 ) | ( n4068 & ~n4073 ) ;
  assign n4075 = ( ~x32 & n4073 ) | ( ~x32 & n4074 ) | ( n4073 & n4074 ) ;
  assign n4076 = ( ~n4068 & n4074 ) | ( ~n4068 & n4075 ) | ( n4074 & n4075 ) ;
  assign n4077 = x66 & n3719 ;
  assign n4078 = x67 | n4077 ;
  assign n4079 = ( n3721 & n4077 ) | ( n3721 & n4078 ) | ( n4077 & n4078 ) ;
  assign n4080 = x65 & n3922 ;
  assign n4081 = n4079 | n4080 ;
  assign n4082 = n164 & n3715 ;
  assign n4083 = ( x41 & n4081 ) | ( x41 & ~n4082 ) | ( n4081 & ~n4082 ) ;
  assign n4084 = ( ~x41 & n4082 ) | ( ~x41 & n4083 ) | ( n4082 & n4083 ) ;
  assign n4085 = ( ~n4081 & n4083 ) | ( ~n4081 & n4084 ) | ( n4083 & n4084 ) ;
  assign n4086 = x41 & x42 ;
  assign n4087 = x41 | x42 ;
  assign n4088 = ~n4086 & n4087 ;
  assign n4089 = x64 & n4088 ;
  assign n4090 = x41 & ~n3930 ;
  assign n4091 = ( n4085 & n4089 ) | ( n4085 & n4090 ) | ( n4089 & n4090 ) ;
  assign n4092 = ( ~n4085 & n4089 ) | ( ~n4085 & n4090 ) | ( n4089 & n4090 ) ;
  assign n4093 = ( n4085 & ~n4091 ) | ( n4085 & n4092 ) | ( ~n4091 & n4092 ) ;
  assign n4094 = n245 & n3224 ;
  assign n4095 = x69 & n3228 ;
  assign n4096 = x70 | n4095 ;
  assign n4097 = ( n3230 & n4095 ) | ( n3230 & n4096 ) | ( n4095 & n4096 ) ;
  assign n4098 = x68 & n3413 ;
  assign n4099 = n4097 | n4098 ;
  assign n4100 = ( x38 & n4094 ) | ( x38 & ~n4099 ) | ( n4094 & ~n4099 ) ;
  assign n4101 = ( ~x38 & n4099 ) | ( ~x38 & n4100 ) | ( n4099 & n4100 ) ;
  assign n4102 = ( ~n4094 & n4100 ) | ( ~n4094 & n4101 ) | ( n4100 & n4101 ) ;
  assign n4103 = ( n3933 & n4093 ) | ( n3933 & n4102 ) | ( n4093 & n4102 ) ;
  assign n4104 = ( ~n3933 & n4093 ) | ( ~n3933 & n4102 ) | ( n4093 & n4102 ) ;
  assign n4105 = ( n3933 & ~n4103 ) | ( n3933 & n4104 ) | ( ~n4103 & n4104 ) ;
  assign n4106 = n390 & n2766 ;
  assign n4107 = x72 & n2770 ;
  assign n4108 = x73 | n4107 ;
  assign n4109 = ( n2772 & n4107 ) | ( n2772 & n4108 ) | ( n4107 & n4108 ) ;
  assign n4110 = x71 & n2943 ;
  assign n4111 = n4109 | n4110 ;
  assign n4112 = ( x35 & n4106 ) | ( x35 & ~n4111 ) | ( n4106 & ~n4111 ) ;
  assign n4113 = ( ~x35 & n4111 ) | ( ~x35 & n4112 ) | ( n4111 & n4112 ) ;
  assign n4114 = ( ~n4106 & n4112 ) | ( ~n4106 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4115 = ( n3936 & n4105 ) | ( n3936 & n4114 ) | ( n4105 & n4114 ) ;
  assign n4116 = ( ~n3936 & n4105 ) | ( ~n3936 & n4114 ) | ( n4105 & n4114 ) ;
  assign n4117 = ( n3936 & ~n4115 ) | ( n3936 & n4116 ) | ( ~n4115 & n4116 ) ;
  assign n4118 = ( n3939 & n4076 ) | ( n3939 & n4117 ) | ( n4076 & n4117 ) ;
  assign n4119 = ( ~n3939 & n4076 ) | ( ~n3939 & n4117 ) | ( n4076 & n4117 ) ;
  assign n4120 = ( n3939 & ~n4118 ) | ( n3939 & n4119 ) | ( ~n4118 & n4119 ) ;
  assign n4121 = ( n3942 & n4067 ) | ( n3942 & n4120 ) | ( n4067 & n4120 ) ;
  assign n4122 = ( ~n3942 & n4067 ) | ( ~n3942 & n4120 ) | ( n4067 & n4120 ) ;
  assign n4123 = ( n3942 & ~n4121 ) | ( n3942 & n4122 ) | ( ~n4121 & n4122 ) ;
  assign n4124 = ( n3945 & n4058 ) | ( n3945 & n4123 ) | ( n4058 & n4123 ) ;
  assign n4125 = ( ~n3945 & n4058 ) | ( ~n3945 & n4123 ) | ( n4058 & n4123 ) ;
  assign n4126 = ( n3945 & ~n4124 ) | ( n3945 & n4125 ) | ( ~n4124 & n4125 ) ;
  assign n4127 = n1262 & n1297 ;
  assign n4128 = x84 & n1301 ;
  assign n4129 = x85 | n4128 ;
  assign n4130 = ( n1303 & n4128 ) | ( n1303 & n4129 ) | ( n4128 & n4129 ) ;
  assign n4131 = x83 & n1426 ;
  assign n4132 = n4130 | n4131 ;
  assign n4133 = ( x23 & n4127 ) | ( x23 & ~n4132 ) | ( n4127 & ~n4132 ) ;
  assign n4134 = ( ~x23 & n4132 ) | ( ~x23 & n4133 ) | ( n4132 & n4133 ) ;
  assign n4135 = ( ~n4127 & n4133 ) | ( ~n4127 & n4134 ) | ( n4133 & n4134 ) ;
  assign n4136 = ( n3957 & n4126 ) | ( n3957 & n4135 ) | ( n4126 & n4135 ) ;
  assign n4137 = ( ~n3957 & n4126 ) | ( ~n3957 & n4135 ) | ( n4126 & n4135 ) ;
  assign n4138 = ( n3957 & ~n4136 ) | ( n3957 & n4137 ) | ( ~n4136 & n4137 ) ;
  assign n4139 = n1016 & n1481 ;
  assign n4140 = x87 & n1020 ;
  assign n4141 = x88 | n4140 ;
  assign n4142 = ( n1022 & n4140 ) | ( n1022 & n4141 ) | ( n4140 & n4141 ) ;
  assign n4143 = x86 & n1145 ;
  assign n4144 = n4142 | n4143 ;
  assign n4145 = ( x20 & n4139 ) | ( x20 & ~n4144 ) | ( n4139 & ~n4144 ) ;
  assign n4146 = ( ~x20 & n4144 ) | ( ~x20 & n4145 ) | ( n4144 & n4145 ) ;
  assign n4147 = ( ~n4139 & n4145 ) | ( ~n4139 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4148 = ( n3969 & n4138 ) | ( n3969 & n4147 ) | ( n4138 & n4147 ) ;
  assign n4149 = ( ~n3969 & n4138 ) | ( ~n3969 & n4147 ) | ( n4138 & n4147 ) ;
  assign n4150 = ( n3969 & ~n4148 ) | ( n3969 & n4149 ) | ( ~n4148 & n4149 ) ;
  assign n4151 = n810 & n1914 ;
  assign n4152 = x90 & n814 ;
  assign n4153 = x91 | n4152 ;
  assign n4154 = ( n816 & n4152 ) | ( n816 & n4153 ) | ( n4152 & n4153 ) ;
  assign n4155 = x89 & n885 ;
  assign n4156 = n4154 | n4155 ;
  assign n4157 = ( x17 & n4151 ) | ( x17 & ~n4156 ) | ( n4151 & ~n4156 ) ;
  assign n4158 = ( ~x17 & n4156 ) | ( ~x17 & n4157 ) | ( n4156 & n4157 ) ;
  assign n4159 = ( ~n4151 & n4157 ) | ( ~n4151 & n4158 ) | ( n4157 & n4158 ) ;
  assign n4160 = ( n3972 & n4150 ) | ( n3972 & n4159 ) | ( n4150 & n4159 ) ;
  assign n4161 = ( ~n3972 & n4150 ) | ( ~n3972 & n4159 ) | ( n4150 & n4159 ) ;
  assign n4162 = ( n3972 & ~n4160 ) | ( n3972 & n4161 ) | ( ~n4160 & n4161 ) ;
  assign n4163 = ( n3975 & n4049 ) | ( n3975 & n4162 ) | ( n4049 & n4162 ) ;
  assign n4164 = ( ~n3975 & n4049 ) | ( ~n3975 & n4162 ) | ( n4049 & n4162 ) ;
  assign n4165 = ( n3975 & ~n4163 ) | ( n3975 & n4164 ) | ( ~n4163 & n4164 ) ;
  assign n4166 = n407 & n2585 ;
  assign n4167 = x96 & n411 ;
  assign n4168 = x97 | n4167 ;
  assign n4169 = ( n413 & n4167 ) | ( n413 & n4168 ) | ( n4167 & n4168 ) ;
  assign n4170 = x95 & n491 ;
  assign n4171 = n4169 | n4170 ;
  assign n4172 = ( x11 & n4166 ) | ( x11 & ~n4171 ) | ( n4166 & ~n4171 ) ;
  assign n4173 = ( ~x11 & n4171 ) | ( ~x11 & n4172 ) | ( n4171 & n4172 ) ;
  assign n4174 = ( ~n4166 & n4172 ) | ( ~n4166 & n4173 ) | ( n4172 & n4173 ) ;
  assign n4175 = ( n3978 & n4165 ) | ( n3978 & n4174 ) | ( n4165 & n4174 ) ;
  assign n4176 = ( ~n3978 & n4165 ) | ( ~n3978 & n4174 ) | ( n4165 & n4174 ) ;
  assign n4177 = ( n3978 & ~n4175 ) | ( n3978 & n4176 ) | ( ~n4175 & n4176 ) ;
  assign n4178 = ( n3990 & n4040 ) | ( n3990 & n4177 ) | ( n4040 & n4177 ) ;
  assign n4179 = ( ~n3990 & n4040 ) | ( ~n3990 & n4177 ) | ( n4040 & n4177 ) ;
  assign n4180 = ( n3990 & ~n4178 ) | ( n3990 & n4179 ) | ( ~n4178 & n4179 ) ;
  assign n4181 = ( n3993 & n4031 ) | ( n3993 & n4180 ) | ( n4031 & n4180 ) ;
  assign n4182 = ( ~n3993 & n4031 ) | ( ~n3993 & n4180 ) | ( n4031 & n4180 ) ;
  assign n4183 = ( n3993 & ~n4181 ) | ( n3993 & n4182 ) | ( ~n4181 & n4182 ) ;
  assign n4184 = ( n4008 & n4022 ) | ( n4008 & n4183 ) | ( n4022 & n4183 ) ;
  assign n4185 = ( ~n4008 & n4022 ) | ( ~n4008 & n4183 ) | ( n4022 & n4183 ) ;
  assign n4186 = ( n4008 & ~n4184 ) | ( n4008 & n4185 ) | ( ~n4184 & n4185 ) ;
  assign n4187 = n186 & n3665 ;
  assign n4188 = x103 & n190 ;
  assign n4189 = x104 | n4188 ;
  assign n4190 = ( n192 & n4188 ) | ( n192 & n4189 ) | ( n4188 & n4189 ) ;
  assign n4191 = x102 & n220 ;
  assign n4192 = n4190 | n4191 ;
  assign n4193 = ( x5 & n4187 ) | ( x5 & ~n4192 ) | ( n4187 & ~n4192 ) ;
  assign n4194 = ( ~x5 & n4192 ) | ( ~x5 & n4193 ) | ( n4192 & n4193 ) ;
  assign n4195 = ( ~n4187 & n4193 ) | ( ~n4187 & n4194 ) | ( n4193 & n4194 ) ;
  assign n4196 = n583 & n2434 ;
  assign n4197 = x94 & n587 ;
  assign n4198 = x95 | n4197 ;
  assign n4199 = ( n589 & n4197 ) | ( n589 & n4198 ) | ( n4197 & n4198 ) ;
  assign n4200 = x93 & n676 ;
  assign n4201 = n4199 | n4200 ;
  assign n4202 = ( x14 & n4196 ) | ( x14 & ~n4201 ) | ( n4196 & ~n4201 ) ;
  assign n4203 = ( ~x14 & n4201 ) | ( ~x14 & n4202 ) | ( n4201 & n4202 ) ;
  assign n4204 = ( ~n4196 & n4202 ) | ( ~n4196 & n4203 ) | ( n4202 & n4203 ) ;
  assign n4205 = n810 & n2042 ;
  assign n4206 = x91 & n814 ;
  assign n4207 = x92 | n4206 ;
  assign n4208 = ( n816 & n4206 ) | ( n816 & n4207 ) | ( n4206 & n4207 ) ;
  assign n4209 = x90 & n885 ;
  assign n4210 = n4208 | n4209 ;
  assign n4211 = ( x17 & n4205 ) | ( x17 & ~n4210 ) | ( n4205 & ~n4210 ) ;
  assign n4212 = ( ~x17 & n4210 ) | ( ~x17 & n4211 ) | ( n4210 & n4211 ) ;
  assign n4213 = ( ~n4205 & n4211 ) | ( ~n4205 & n4212 ) | ( n4211 & n4212 ) ;
  assign n4214 = n569 & n2320 ;
  assign n4215 = x76 & n2324 ;
  assign n4216 = x77 | n4215 ;
  assign n4217 = ( n2326 & n4215 ) | ( n2326 & n4216 ) | ( n4215 & n4216 ) ;
  assign n4218 = x75 & n2497 ;
  assign n4219 = n4217 | n4218 ;
  assign n4220 = ( x32 & n4214 ) | ( x32 & ~n4219 ) | ( n4214 & ~n4219 ) ;
  assign n4221 = ( ~x32 & n4219 ) | ( ~x32 & n4220 ) | ( n4219 & n4220 ) ;
  assign n4222 = ( ~n4214 & n4220 ) | ( ~n4214 & n4221 ) | ( n4220 & n4221 ) ;
  assign n4223 = x44 & n4089 ;
  assign n4224 = x43 | x44 ;
  assign n4225 = ( x43 & x44 ) | ( x43 & ~n4224 ) | ( x44 & ~n4224 ) ;
  assign n4226 = n4224 & ~n4225 ;
  assign n4227 = n4088 & n4226 ;
  assign n4228 = n133 & n4227 ;
  assign n4229 = ~x41 & x43 ;
  assign n4230 = x42 & x43 ;
  assign n4231 = ( n4086 & n4229 ) | ( n4086 & ~n4230 ) | ( n4229 & ~n4230 ) ;
  assign n4232 = x64 & n4231 ;
  assign n4233 = ( n4088 & ~n4224 ) | ( n4088 & n4225 ) | ( ~n4224 & n4225 ) ;
  assign n4234 = x65 | n4232 ;
  assign n4235 = ( n4232 & n4233 ) | ( n4232 & n4234 ) | ( n4233 & n4234 ) ;
  assign n4236 = ( n4223 & n4228 ) | ( n4223 & n4235 ) | ( n4228 & n4235 ) ;
  assign n4237 = n4228 | n4235 ;
  assign n4238 = ~n4223 & n4237 ;
  assign n4239 = ( n4223 & ~n4236 ) | ( n4223 & n4238 ) | ( ~n4236 & n4238 ) ;
  assign n4240 = x67 & n3719 ;
  assign n4241 = x68 | n4240 ;
  assign n4242 = ( n3721 & n4240 ) | ( n3721 & n4241 ) | ( n4240 & n4241 ) ;
  assign n4243 = x66 & n3922 ;
  assign n4244 = n4242 | n4243 ;
  assign n4245 = n201 & n3715 ;
  assign n4246 = ( x41 & n4244 ) | ( x41 & ~n4245 ) | ( n4244 & ~n4245 ) ;
  assign n4247 = ( ~x41 & n4245 ) | ( ~x41 & n4246 ) | ( n4245 & n4246 ) ;
  assign n4248 = ( ~n4244 & n4246 ) | ( ~n4244 & n4247 ) | ( n4246 & n4247 ) ;
  assign n4249 = ( n4091 & n4239 ) | ( n4091 & n4248 ) | ( n4239 & n4248 ) ;
  assign n4250 = ( ~n4091 & n4239 ) | ( ~n4091 & n4248 ) | ( n4239 & n4248 ) ;
  assign n4251 = ( n4091 & ~n4249 ) | ( n4091 & n4250 ) | ( ~n4249 & n4250 ) ;
  assign n4252 = n277 & n3224 ;
  assign n4253 = x70 & n3228 ;
  assign n4254 = x71 | n4253 ;
  assign n4255 = ( n3230 & n4253 ) | ( n3230 & n4254 ) | ( n4253 & n4254 ) ;
  assign n4256 = x69 & n3413 ;
  assign n4257 = n4255 | n4256 ;
  assign n4258 = ( x38 & n4252 ) | ( x38 & ~n4257 ) | ( n4252 & ~n4257 ) ;
  assign n4259 = ( ~x38 & n4257 ) | ( ~x38 & n4258 ) | ( n4257 & n4258 ) ;
  assign n4260 = ( ~n4252 & n4258 ) | ( ~n4252 & n4259 ) | ( n4258 & n4259 ) ;
  assign n4261 = ( n4103 & n4251 ) | ( n4103 & n4260 ) | ( n4251 & n4260 ) ;
  assign n4262 = ( ~n4103 & n4251 ) | ( ~n4103 & n4260 ) | ( n4251 & n4260 ) ;
  assign n4263 = ( n4103 & ~n4261 ) | ( n4103 & n4262 ) | ( ~n4261 & n4262 ) ;
  assign n4264 = n446 & n2766 ;
  assign n4265 = x73 & n2770 ;
  assign n4266 = x74 | n4265 ;
  assign n4267 = ( n2772 & n4265 ) | ( n2772 & n4266 ) | ( n4265 & n4266 ) ;
  assign n4268 = x72 & n2943 ;
  assign n4269 = n4267 | n4268 ;
  assign n4270 = ( x35 & n4264 ) | ( x35 & ~n4269 ) | ( n4264 & ~n4269 ) ;
  assign n4271 = ( ~x35 & n4269 ) | ( ~x35 & n4270 ) | ( n4269 & n4270 ) ;
  assign n4272 = ( ~n4264 & n4270 ) | ( ~n4264 & n4271 ) | ( n4270 & n4271 ) ;
  assign n4273 = ( n4115 & n4263 ) | ( n4115 & n4272 ) | ( n4263 & n4272 ) ;
  assign n4274 = ( ~n4115 & n4263 ) | ( ~n4115 & n4272 ) | ( n4263 & n4272 ) ;
  assign n4275 = ( n4115 & ~n4273 ) | ( n4115 & n4274 ) | ( ~n4273 & n4274 ) ;
  assign n4276 = ( n4118 & n4222 ) | ( n4118 & n4275 ) | ( n4222 & n4275 ) ;
  assign n4277 = ( ~n4118 & n4222 ) | ( ~n4118 & n4275 ) | ( n4222 & n4275 ) ;
  assign n4278 = ( n4118 & ~n4276 ) | ( n4118 & n4277 ) | ( ~n4276 & n4277 ) ;
  assign n4279 = n769 & n1949 ;
  assign n4280 = x79 & n1953 ;
  assign n4281 = x80 | n4280 ;
  assign n4282 = ( n1955 & n4280 ) | ( n1955 & n4281 ) | ( n4280 & n4281 ) ;
  assign n4283 = x78 & n2114 ;
  assign n4284 = n4282 | n4283 ;
  assign n4285 = ( x29 & n4279 ) | ( x29 & ~n4284 ) | ( n4279 & ~n4284 ) ;
  assign n4286 = ( ~x29 & n4284 ) | ( ~x29 & n4285 ) | ( n4284 & n4285 ) ;
  assign n4287 = ( ~n4279 & n4285 ) | ( ~n4279 & n4286 ) | ( n4285 & n4286 ) ;
  assign n4288 = ( n4121 & n4278 ) | ( n4121 & n4287 ) | ( n4278 & n4287 ) ;
  assign n4289 = ( ~n4121 & n4278 ) | ( ~n4121 & n4287 ) | ( n4278 & n4287 ) ;
  assign n4290 = ( n4121 & ~n4288 ) | ( n4121 & n4289 ) | ( ~n4288 & n4289 ) ;
  assign n4291 = n1082 & n1617 ;
  assign n4292 = x82 & n1621 ;
  assign n4293 = x83 | n4292 ;
  assign n4294 = ( n1623 & n4292 ) | ( n1623 & n4293 ) | ( n4292 & n4293 ) ;
  assign n4295 = x81 & n1749 ;
  assign n4296 = n4294 | n4295 ;
  assign n4297 = ( x26 & n4291 ) | ( x26 & ~n4296 ) | ( n4291 & ~n4296 ) ;
  assign n4298 = ( ~x26 & n4296 ) | ( ~x26 & n4297 ) | ( n4296 & n4297 ) ;
  assign n4299 = ( ~n4291 & n4297 ) | ( ~n4291 & n4298 ) | ( n4297 & n4298 ) ;
  assign n4300 = ( n4124 & n4290 ) | ( n4124 & n4299 ) | ( n4290 & n4299 ) ;
  assign n4301 = ( ~n4124 & n4290 ) | ( ~n4124 & n4299 ) | ( n4290 & n4299 ) ;
  assign n4302 = ( n4124 & ~n4300 ) | ( n4124 & n4301 ) | ( ~n4300 & n4301 ) ;
  assign n4303 = n1297 & n1366 ;
  assign n4304 = x85 & n1301 ;
  assign n4305 = x86 | n4304 ;
  assign n4306 = ( n1303 & n4304 ) | ( n1303 & n4305 ) | ( n4304 & n4305 ) ;
  assign n4307 = x84 & n1426 ;
  assign n4308 = n4306 | n4307 ;
  assign n4309 = ( x23 & n4303 ) | ( x23 & ~n4308 ) | ( n4303 & ~n4308 ) ;
  assign n4310 = ( ~x23 & n4308 ) | ( ~x23 & n4309 ) | ( n4308 & n4309 ) ;
  assign n4311 = ( ~n4303 & n4309 ) | ( ~n4303 & n4310 ) | ( n4309 & n4310 ) ;
  assign n4312 = ( n4136 & n4302 ) | ( n4136 & n4311 ) | ( n4302 & n4311 ) ;
  assign n4313 = ( ~n4136 & n4302 ) | ( ~n4136 & n4311 ) | ( n4302 & n4311 ) ;
  assign n4314 = ( n4136 & ~n4312 ) | ( n4136 & n4313 ) | ( ~n4312 & n4313 ) ;
  assign n4315 = n1016 & n1585 ;
  assign n4316 = x88 & n1020 ;
  assign n4317 = x89 | n4316 ;
  assign n4318 = ( n1022 & n4316 ) | ( n1022 & n4317 ) | ( n4316 & n4317 ) ;
  assign n4319 = x87 & n1145 ;
  assign n4320 = n4318 | n4319 ;
  assign n4321 = ( x20 & n4315 ) | ( x20 & ~n4320 ) | ( n4315 & ~n4320 ) ;
  assign n4322 = ( ~x20 & n4320 ) | ( ~x20 & n4321 ) | ( n4320 & n4321 ) ;
  assign n4323 = ( ~n4315 & n4321 ) | ( ~n4315 & n4322 ) | ( n4321 & n4322 ) ;
  assign n4324 = ( n4148 & n4314 ) | ( n4148 & n4323 ) | ( n4314 & n4323 ) ;
  assign n4325 = ( ~n4148 & n4314 ) | ( ~n4148 & n4323 ) | ( n4314 & n4323 ) ;
  assign n4326 = ( n4148 & ~n4324 ) | ( n4148 & n4325 ) | ( ~n4324 & n4325 ) ;
  assign n4327 = ( n4160 & n4213 ) | ( n4160 & n4326 ) | ( n4213 & n4326 ) ;
  assign n4328 = ( ~n4160 & n4213 ) | ( ~n4160 & n4326 ) | ( n4213 & n4326 ) ;
  assign n4329 = ( n4160 & ~n4327 ) | ( n4160 & n4328 ) | ( ~n4327 & n4328 ) ;
  assign n4330 = ( n4163 & n4204 ) | ( n4163 & n4329 ) | ( n4204 & n4329 ) ;
  assign n4331 = ( ~n4163 & n4204 ) | ( ~n4163 & n4329 ) | ( n4204 & n4329 ) ;
  assign n4332 = ( n4163 & ~n4330 ) | ( n4163 & n4331 ) | ( ~n4330 & n4331 ) ;
  assign n4333 = n407 & n2725 ;
  assign n4334 = x97 & n411 ;
  assign n4335 = x98 | n4334 ;
  assign n4336 = ( n413 & n4334 ) | ( n413 & n4335 ) | ( n4334 & n4335 ) ;
  assign n4337 = x96 & n491 ;
  assign n4338 = n4336 | n4337 ;
  assign n4339 = ( x11 & n4333 ) | ( x11 & ~n4338 ) | ( n4333 & ~n4338 ) ;
  assign n4340 = ( ~x11 & n4338 ) | ( ~x11 & n4339 ) | ( n4338 & n4339 ) ;
  assign n4341 = ( ~n4333 & n4339 ) | ( ~n4333 & n4340 ) | ( n4339 & n4340 ) ;
  assign n4342 = ( n4175 & n4332 ) | ( n4175 & n4341 ) | ( n4332 & n4341 ) ;
  assign n4343 = ( ~n4175 & n4332 ) | ( ~n4175 & n4341 ) | ( n4332 & n4341 ) ;
  assign n4344 = ( n4175 & ~n4342 ) | ( n4175 & n4343 ) | ( ~n4342 & n4343 ) ;
  assign n4345 = n291 & n3326 ;
  assign n4346 = x100 & n295 ;
  assign n4347 = x101 | n4346 ;
  assign n4348 = ( n297 & n4346 ) | ( n297 & n4347 ) | ( n4346 & n4347 ) ;
  assign n4349 = x99 & n330 ;
  assign n4350 = n4348 | n4349 ;
  assign n4351 = ( x8 & n4345 ) | ( x8 & ~n4350 ) | ( n4345 & ~n4350 ) ;
  assign n4352 = ( ~x8 & n4350 ) | ( ~x8 & n4351 ) | ( n4350 & n4351 ) ;
  assign n4353 = ( ~n4345 & n4351 ) | ( ~n4345 & n4352 ) | ( n4351 & n4352 ) ;
  assign n4354 = ( n4178 & n4344 ) | ( n4178 & n4353 ) | ( n4344 & n4353 ) ;
  assign n4355 = ( ~n4178 & n4344 ) | ( ~n4178 & n4353 ) | ( n4344 & n4353 ) ;
  assign n4356 = ( n4178 & ~n4354 ) | ( n4178 & n4355 ) | ( ~n4354 & n4355 ) ;
  assign n4357 = ( n4181 & n4195 ) | ( n4181 & n4356 ) | ( n4195 & n4356 ) ;
  assign n4358 = ( ~n4181 & n4195 ) | ( ~n4181 & n4356 ) | ( n4195 & n4356 ) ;
  assign n4359 = ( n4181 & ~n4357 ) | ( n4181 & n4358 ) | ( ~n4357 & n4358 ) ;
  assign n4360 = ( x106 & x107 ) | ( x106 & n4011 ) | ( x107 & n4011 ) ;
  assign n4361 = ( x106 & ~x107 ) | ( x106 & n4011 ) | ( ~x107 & n4011 ) ;
  assign n4362 = ( x107 & ~n4360 ) | ( x107 & n4361 ) | ( ~n4360 & n4361 ) ;
  assign n4363 = n136 & n4362 ;
  assign n4364 = x106 & n138 ;
  assign n4365 = x107 | n4364 ;
  assign n4366 = ( n141 & n4364 ) | ( n141 & n4365 ) | ( n4364 & n4365 ) ;
  assign n4367 = x105 & n154 ;
  assign n4368 = n4366 | n4367 ;
  assign n4369 = ( x2 & n4363 ) | ( x2 & ~n4368 ) | ( n4363 & ~n4368 ) ;
  assign n4370 = ( ~x2 & n4368 ) | ( ~x2 & n4369 ) | ( n4368 & n4369 ) ;
  assign n4371 = ( ~n4363 & n4369 ) | ( ~n4363 & n4370 ) | ( n4369 & n4370 ) ;
  assign n4372 = ( n4184 & n4359 ) | ( n4184 & n4371 ) | ( n4359 & n4371 ) ;
  assign n4373 = ( ~n4184 & n4359 ) | ( ~n4184 & n4371 ) | ( n4359 & n4371 ) ;
  assign n4374 = ( n4184 & ~n4372 ) | ( n4184 & n4373 ) | ( ~n4372 & n4373 ) ;
  assign n4375 = ( x107 & x108 ) | ( x107 & n4360 ) | ( x108 & n4360 ) ;
  assign n4376 = ( x107 & ~x108 ) | ( x107 & n4360 ) | ( ~x108 & n4360 ) ;
  assign n4377 = ( x108 & ~n4375 ) | ( x108 & n4376 ) | ( ~n4375 & n4376 ) ;
  assign n4378 = n136 & n4377 ;
  assign n4379 = x107 & n138 ;
  assign n4380 = x108 | n4379 ;
  assign n4381 = ( n141 & n4379 ) | ( n141 & n4380 ) | ( n4379 & n4380 ) ;
  assign n4382 = x106 & n154 ;
  assign n4383 = n4381 | n4382 ;
  assign n4384 = ( x2 & n4378 ) | ( x2 & ~n4383 ) | ( n4378 & ~n4383 ) ;
  assign n4385 = ( ~x2 & n4383 ) | ( ~x2 & n4384 ) | ( n4383 & n4384 ) ;
  assign n4386 = ( ~n4378 & n4384 ) | ( ~n4378 & n4385 ) | ( n4384 & n4385 ) ;
  assign n4387 = n186 & n3998 ;
  assign n4388 = x104 & n190 ;
  assign n4389 = x105 | n4388 ;
  assign n4390 = ( n192 & n4388 ) | ( n192 & n4389 ) | ( n4388 & n4389 ) ;
  assign n4391 = x103 & n220 ;
  assign n4392 = n4390 | n4391 ;
  assign n4393 = ( x5 & n4387 ) | ( x5 & ~n4392 ) | ( n4387 & ~n4392 ) ;
  assign n4394 = ( ~x5 & n4392 ) | ( ~x5 & n4393 ) | ( n4392 & n4393 ) ;
  assign n4395 = ( ~n4387 & n4393 ) | ( ~n4387 & n4394 ) | ( n4393 & n4394 ) ;
  assign n4396 = n583 & n2449 ;
  assign n4397 = x95 & n587 ;
  assign n4398 = x96 | n4397 ;
  assign n4399 = ( n589 & n4397 ) | ( n589 & n4398 ) | ( n4397 & n4398 ) ;
  assign n4400 = x94 & n676 ;
  assign n4401 = n4399 | n4400 ;
  assign n4402 = ( x14 & n4396 ) | ( x14 & ~n4401 ) | ( n4396 & ~n4401 ) ;
  assign n4403 = ( ~x14 & n4401 ) | ( ~x14 & n4402 ) | ( n4401 & n4402 ) ;
  assign n4404 = ( ~n4396 & n4402 ) | ( ~n4396 & n4403 ) | ( n4402 & n4403 ) ;
  assign n4405 = n810 & n2057 ;
  assign n4406 = x92 & n814 ;
  assign n4407 = x93 | n4406 ;
  assign n4408 = ( n816 & n4406 ) | ( n816 & n4407 ) | ( n4406 & n4407 ) ;
  assign n4409 = x91 & n885 ;
  assign n4410 = n4408 | n4409 ;
  assign n4411 = ( x17 & n4405 ) | ( x17 & ~n4410 ) | ( n4405 & ~n4410 ) ;
  assign n4412 = ( ~x17 & n4410 ) | ( ~x17 & n4411 ) | ( n4410 & n4411 ) ;
  assign n4413 = ( ~n4405 & n4411 ) | ( ~n4405 & n4412 ) | ( n4411 & n4412 ) ;
  assign n4414 = n1016 & n1701 ;
  assign n4415 = x89 & n1020 ;
  assign n4416 = x90 | n4415 ;
  assign n4417 = ( n1022 & n4415 ) | ( n1022 & n4416 ) | ( n4415 & n4416 ) ;
  assign n4418 = x88 & n1145 ;
  assign n4419 = n4417 | n4418 ;
  assign n4420 = ( x20 & n4414 ) | ( x20 & ~n4419 ) | ( n4414 & ~n4419 ) ;
  assign n4421 = ( ~x20 & n4419 ) | ( ~x20 & n4420 ) | ( n4419 & n4420 ) ;
  assign n4422 = ( ~n4414 & n4420 ) | ( ~n4414 & n4421 ) | ( n4420 & n4421 ) ;
  assign n4423 = n910 & n1949 ;
  assign n4424 = x80 & n1953 ;
  assign n4425 = x81 | n4424 ;
  assign n4426 = ( n1955 & n4424 ) | ( n1955 & n4425 ) | ( n4424 & n4425 ) ;
  assign n4427 = x79 & n2114 ;
  assign n4428 = n4426 | n4427 ;
  assign n4429 = ( x29 & n4423 ) | ( x29 & ~n4428 ) | ( n4423 & ~n4428 ) ;
  assign n4430 = ( ~x29 & n4428 ) | ( ~x29 & n4429 ) | ( n4428 & n4429 ) ;
  assign n4431 = ( ~n4423 & n4429 ) | ( ~n4423 & n4430 ) | ( n4429 & n4430 ) ;
  assign n4432 = n637 & n2320 ;
  assign n4433 = x77 & n2324 ;
  assign n4434 = x78 | n4433 ;
  assign n4435 = ( n2326 & n4433 ) | ( n2326 & n4434 ) | ( n4433 & n4434 ) ;
  assign n4436 = x76 & n2497 ;
  assign n4437 = n4435 | n4436 ;
  assign n4438 = ( x32 & n4432 ) | ( x32 & ~n4437 ) | ( n4432 & ~n4437 ) ;
  assign n4439 = ( ~x32 & n4437 ) | ( ~x32 & n4438 ) | ( n4437 & n4438 ) ;
  assign n4440 = ( ~n4432 & n4438 ) | ( ~n4432 & n4439 ) | ( n4438 & n4439 ) ;
  assign n4441 = n461 & n2766 ;
  assign n4442 = x74 & n2770 ;
  assign n4443 = x75 | n4442 ;
  assign n4444 = ( n2772 & n4442 ) | ( n2772 & n4443 ) | ( n4442 & n4443 ) ;
  assign n4445 = x73 & n2943 ;
  assign n4446 = n4444 | n4445 ;
  assign n4447 = ( x35 & n4441 ) | ( x35 & ~n4446 ) | ( n4441 & ~n4446 ) ;
  assign n4448 = ( ~x35 & n4446 ) | ( ~x35 & n4447 ) | ( n4446 & n4447 ) ;
  assign n4449 = ( ~n4441 & n4447 ) | ( ~n4441 & n4448 ) | ( n4447 & n4448 ) ;
  assign n4450 = n346 & n3224 ;
  assign n4451 = x71 & n3228 ;
  assign n4452 = x72 | n4451 ;
  assign n4453 = ( n3230 & n4451 ) | ( n3230 & n4452 ) | ( n4451 & n4452 ) ;
  assign n4454 = x70 & n3413 ;
  assign n4455 = n4453 | n4454 ;
  assign n4456 = ( x38 & n4450 ) | ( x38 & ~n4455 ) | ( n4450 & ~n4455 ) ;
  assign n4457 = ( ~x38 & n4455 ) | ( ~x38 & n4456 ) | ( n4455 & n4456 ) ;
  assign n4458 = ( ~n4450 & n4456 ) | ( ~n4450 & n4457 ) | ( n4456 & n4457 ) ;
  assign n4459 = n230 & n3715 ;
  assign n4460 = x68 & n3719 ;
  assign n4461 = x69 | n4460 ;
  assign n4462 = ( n3721 & n4460 ) | ( n3721 & n4461 ) | ( n4460 & n4461 ) ;
  assign n4463 = x67 & n3922 ;
  assign n4464 = n4462 | n4463 ;
  assign n4465 = ( ~x41 & n4459 ) | ( ~x41 & n4464 ) | ( n4459 & n4464 ) ;
  assign n4466 = ( n4459 & n4464 ) | ( n4459 & ~n4465 ) | ( n4464 & ~n4465 ) ;
  assign n4467 = ( x41 & n4465 ) | ( x41 & ~n4466 ) | ( n4465 & ~n4466 ) ;
  assign n4468 = ( x44 & n4223 ) | ( x44 & n4237 ) | ( n4223 & n4237 ) ;
  assign n4469 = ( x41 & ~x43 ) | ( x41 & n4226 ) | ( ~x43 & n4226 ) ;
  assign n4470 = ( ~n4087 & n4230 ) | ( ~n4087 & n4469 ) | ( n4230 & n4469 ) ;
  assign n4471 = x64 & n4470 ;
  assign n4472 = x65 & n4231 ;
  assign n4473 = x66 | n4472 ;
  assign n4474 = ( n4233 & n4472 ) | ( n4233 & n4473 ) | ( n4472 & n4473 ) ;
  assign n4475 = ( n151 & n152 ) | ( n151 & n4227 ) | ( n152 & n4227 ) ;
  assign n4476 = ( ~n4471 & n4474 ) | ( ~n4471 & n4475 ) | ( n4474 & n4475 ) ;
  assign n4477 = n4471 | n4476 ;
  assign n4478 = n4468 | n4477 ;
  assign n4479 = ( n4468 & n4477 ) | ( n4468 & ~n4478 ) | ( n4477 & ~n4478 ) ;
  assign n4480 = n4478 & ~n4479 ;
  assign n4481 = ( n4249 & n4467 ) | ( n4249 & n4480 ) | ( n4467 & n4480 ) ;
  assign n4482 = ( ~n4249 & n4467 ) | ( ~n4249 & n4480 ) | ( n4467 & n4480 ) ;
  assign n4483 = ( n4249 & ~n4481 ) | ( n4249 & n4482 ) | ( ~n4481 & n4482 ) ;
  assign n4484 = ( n4261 & n4458 ) | ( n4261 & n4483 ) | ( n4458 & n4483 ) ;
  assign n4485 = ( ~n4261 & n4458 ) | ( ~n4261 & n4483 ) | ( n4458 & n4483 ) ;
  assign n4486 = ( n4261 & ~n4484 ) | ( n4261 & n4485 ) | ( ~n4484 & n4485 ) ;
  assign n4487 = ( n4273 & n4449 ) | ( n4273 & n4486 ) | ( n4449 & n4486 ) ;
  assign n4488 = ( ~n4273 & n4449 ) | ( ~n4273 & n4486 ) | ( n4449 & n4486 ) ;
  assign n4489 = ( n4273 & ~n4487 ) | ( n4273 & n4488 ) | ( ~n4487 & n4488 ) ;
  assign n4490 = ( n4276 & n4440 ) | ( n4276 & n4489 ) | ( n4440 & n4489 ) ;
  assign n4491 = ( ~n4276 & n4440 ) | ( ~n4276 & n4489 ) | ( n4440 & n4489 ) ;
  assign n4492 = ( n4276 & ~n4490 ) | ( n4276 & n4491 ) | ( ~n4490 & n4491 ) ;
  assign n4493 = ( n4288 & n4431 ) | ( n4288 & n4492 ) | ( n4431 & n4492 ) ;
  assign n4494 = ( ~n4288 & n4431 ) | ( ~n4288 & n4492 ) | ( n4431 & n4492 ) ;
  assign n4495 = ( n4288 & ~n4493 ) | ( n4288 & n4494 ) | ( ~n4493 & n4494 ) ;
  assign n4496 = n1097 & n1617 ;
  assign n4497 = x83 & n1621 ;
  assign n4498 = x84 | n4497 ;
  assign n4499 = ( n1623 & n4497 ) | ( n1623 & n4498 ) | ( n4497 & n4498 ) ;
  assign n4500 = x82 & n1749 ;
  assign n4501 = n4499 | n4500 ;
  assign n4502 = ( x26 & n4496 ) | ( x26 & ~n4501 ) | ( n4496 & ~n4501 ) ;
  assign n4503 = ( ~x26 & n4501 ) | ( ~x26 & n4502 ) | ( n4501 & n4502 ) ;
  assign n4504 = ( ~n4496 & n4502 ) | ( ~n4496 & n4503 ) | ( n4502 & n4503 ) ;
  assign n4505 = ( n4300 & n4495 ) | ( n4300 & n4504 ) | ( n4495 & n4504 ) ;
  assign n4506 = ( ~n4300 & n4495 ) | ( ~n4300 & n4504 ) | ( n4495 & n4504 ) ;
  assign n4507 = ( n4300 & ~n4505 ) | ( n4300 & n4506 ) | ( ~n4505 & n4506 ) ;
  assign n4508 = n1297 & n1466 ;
  assign n4509 = x86 & n1301 ;
  assign n4510 = x87 | n4509 ;
  assign n4511 = ( n1303 & n4509 ) | ( n1303 & n4510 ) | ( n4509 & n4510 ) ;
  assign n4512 = x85 & n1426 ;
  assign n4513 = n4511 | n4512 ;
  assign n4514 = ( x23 & n4508 ) | ( x23 & ~n4513 ) | ( n4508 & ~n4513 ) ;
  assign n4515 = ( ~x23 & n4513 ) | ( ~x23 & n4514 ) | ( n4513 & n4514 ) ;
  assign n4516 = ( ~n4508 & n4514 ) | ( ~n4508 & n4515 ) | ( n4514 & n4515 ) ;
  assign n4517 = ( n4312 & n4507 ) | ( n4312 & n4516 ) | ( n4507 & n4516 ) ;
  assign n4518 = ( ~n4312 & n4507 ) | ( ~n4312 & n4516 ) | ( n4507 & n4516 ) ;
  assign n4519 = ( n4312 & ~n4517 ) | ( n4312 & n4518 ) | ( ~n4517 & n4518 ) ;
  assign n4520 = ( n4324 & n4422 ) | ( n4324 & n4519 ) | ( n4422 & n4519 ) ;
  assign n4521 = ( ~n4324 & n4422 ) | ( ~n4324 & n4519 ) | ( n4422 & n4519 ) ;
  assign n4522 = ( n4324 & ~n4520 ) | ( n4324 & n4521 ) | ( ~n4520 & n4521 ) ;
  assign n4523 = ( n4327 & n4413 ) | ( n4327 & n4522 ) | ( n4413 & n4522 ) ;
  assign n4524 = ( ~n4327 & n4413 ) | ( ~n4327 & n4522 ) | ( n4413 & n4522 ) ;
  assign n4525 = ( n4327 & ~n4523 ) | ( n4327 & n4524 ) | ( ~n4523 & n4524 ) ;
  assign n4526 = ( n4330 & n4404 ) | ( n4330 & n4525 ) | ( n4404 & n4525 ) ;
  assign n4527 = ( ~n4330 & n4404 ) | ( ~n4330 & n4525 ) | ( n4404 & n4525 ) ;
  assign n4528 = ( n4330 & ~n4526 ) | ( n4330 & n4527 ) | ( ~n4526 & n4527 ) ;
  assign n4529 = n407 & n2877 ;
  assign n4530 = x98 & n411 ;
  assign n4531 = x99 | n4530 ;
  assign n4532 = ( n413 & n4530 ) | ( n413 & n4531 ) | ( n4530 & n4531 ) ;
  assign n4533 = x97 & n491 ;
  assign n4534 = n4532 | n4533 ;
  assign n4535 = ( x11 & n4529 ) | ( x11 & ~n4534 ) | ( n4529 & ~n4534 ) ;
  assign n4536 = ( ~x11 & n4534 ) | ( ~x11 & n4535 ) | ( n4534 & n4535 ) ;
  assign n4537 = ( ~n4529 & n4535 ) | ( ~n4529 & n4536 ) | ( n4535 & n4536 ) ;
  assign n4538 = ( n4342 & n4528 ) | ( n4342 & n4537 ) | ( n4528 & n4537 ) ;
  assign n4539 = ( ~n4342 & n4528 ) | ( ~n4342 & n4537 ) | ( n4528 & n4537 ) ;
  assign n4540 = ( n4342 & ~n4538 ) | ( n4342 & n4539 ) | ( ~n4538 & n4539 ) ;
  assign n4541 = n291 & n3486 ;
  assign n4542 = x101 & n295 ;
  assign n4543 = x102 | n4542 ;
  assign n4544 = ( n297 & n4542 ) | ( n297 & n4543 ) | ( n4542 & n4543 ) ;
  assign n4545 = x100 & n330 ;
  assign n4546 = n4544 | n4545 ;
  assign n4547 = ( x8 & n4541 ) | ( x8 & ~n4546 ) | ( n4541 & ~n4546 ) ;
  assign n4548 = ( ~x8 & n4546 ) | ( ~x8 & n4547 ) | ( n4546 & n4547 ) ;
  assign n4549 = ( ~n4541 & n4547 ) | ( ~n4541 & n4548 ) | ( n4547 & n4548 ) ;
  assign n4550 = ( n4354 & n4540 ) | ( n4354 & n4549 ) | ( n4540 & n4549 ) ;
  assign n4551 = ( ~n4354 & n4540 ) | ( ~n4354 & n4549 ) | ( n4540 & n4549 ) ;
  assign n4552 = ( n4354 & ~n4550 ) | ( n4354 & n4551 ) | ( ~n4550 & n4551 ) ;
  assign n4553 = ( n4357 & n4395 ) | ( n4357 & n4552 ) | ( n4395 & n4552 ) ;
  assign n4554 = ( ~n4357 & n4395 ) | ( ~n4357 & n4552 ) | ( n4395 & n4552 ) ;
  assign n4555 = ( n4357 & ~n4553 ) | ( n4357 & n4554 ) | ( ~n4553 & n4554 ) ;
  assign n4556 = ( n4372 & n4386 ) | ( n4372 & n4555 ) | ( n4386 & n4555 ) ;
  assign n4557 = ( ~n4372 & n4386 ) | ( ~n4372 & n4555 ) | ( n4386 & n4555 ) ;
  assign n4558 = ( n4372 & ~n4556 ) | ( n4372 & n4557 ) | ( ~n4556 & n4557 ) ;
  assign n4559 = n407 & n3162 ;
  assign n4560 = x99 & n411 ;
  assign n4561 = x100 | n4560 ;
  assign n4562 = ( n413 & n4560 ) | ( n413 & n4561 ) | ( n4560 & n4561 ) ;
  assign n4563 = x98 & n491 ;
  assign n4564 = n4562 | n4563 ;
  assign n4565 = ( x11 & n4559 ) | ( x11 & ~n4564 ) | ( n4559 & ~n4564 ) ;
  assign n4566 = ( ~x11 & n4564 ) | ( ~x11 & n4565 ) | ( n4564 & n4565 ) ;
  assign n4567 = ( ~n4559 & n4565 ) | ( ~n4559 & n4566 ) | ( n4565 & n4566 ) ;
  assign n4568 = n810 & n2294 ;
  assign n4569 = x93 & n814 ;
  assign n4570 = x94 | n4569 ;
  assign n4571 = ( n816 & n4569 ) | ( n816 & n4570 ) | ( n4569 & n4570 ) ;
  assign n4572 = x92 & n885 ;
  assign n4573 = n4571 | n4572 ;
  assign n4574 = ( x17 & n4568 ) | ( x17 & ~n4573 ) | ( n4568 & ~n4573 ) ;
  assign n4575 = ( ~x17 & n4573 ) | ( ~x17 & n4574 ) | ( n4573 & n4574 ) ;
  assign n4576 = ( ~n4568 & n4574 ) | ( ~n4568 & n4575 ) | ( n4574 & n4575 ) ;
  assign n4577 = n990 & n1949 ;
  assign n4578 = x81 & n1953 ;
  assign n4579 = x82 | n4578 ;
  assign n4580 = ( n1955 & n4578 ) | ( n1955 & n4579 ) | ( n4578 & n4579 ) ;
  assign n4581 = x80 & n2114 ;
  assign n4582 = n4580 | n4581 ;
  assign n4583 = ( x29 & n4577 ) | ( x29 & ~n4582 ) | ( n4577 & ~n4582 ) ;
  assign n4584 = ( ~x29 & n4582 ) | ( ~x29 & n4583 ) | ( n4582 & n4583 ) ;
  assign n4585 = ( ~n4577 & n4583 ) | ( ~n4577 & n4584 ) | ( n4583 & n4584 ) ;
  assign n4586 = n701 & n2320 ;
  assign n4587 = x78 & n2324 ;
  assign n4588 = x79 | n4587 ;
  assign n4589 = ( n2326 & n4587 ) | ( n2326 & n4588 ) | ( n4587 & n4588 ) ;
  assign n4590 = x77 & n2497 ;
  assign n4591 = n4589 | n4590 ;
  assign n4592 = ( x32 & n4586 ) | ( x32 & ~n4591 ) | ( n4586 & ~n4591 ) ;
  assign n4593 = ( ~x32 & n4591 ) | ( ~x32 & n4592 ) | ( n4591 & n4592 ) ;
  assign n4594 = ( ~n4586 & n4592 ) | ( ~n4586 & n4593 ) | ( n4592 & n4593 ) ;
  assign n4595 = n554 & n2766 ;
  assign n4596 = x75 & n2770 ;
  assign n4597 = x76 | n4596 ;
  assign n4598 = ( n2772 & n4596 ) | ( n2772 & n4597 ) | ( n4596 & n4597 ) ;
  assign n4599 = x74 & n2943 ;
  assign n4600 = n4598 | n4599 ;
  assign n4601 = ( x35 & n4595 ) | ( x35 & ~n4600 ) | ( n4595 & ~n4600 ) ;
  assign n4602 = ( ~x35 & n4600 ) | ( ~x35 & n4601 ) | ( n4600 & n4601 ) ;
  assign n4603 = ( ~n4595 & n4601 ) | ( ~n4595 & n4602 ) | ( n4601 & n4602 ) ;
  assign n4604 = x66 & n4231 ;
  assign n4605 = x67 | n4604 ;
  assign n4606 = ( n4233 & n4604 ) | ( n4233 & n4605 ) | ( n4604 & n4605 ) ;
  assign n4607 = x65 & n4470 ;
  assign n4608 = n4606 | n4607 ;
  assign n4609 = n164 & n4227 ;
  assign n4610 = ( x44 & n4608 ) | ( x44 & ~n4609 ) | ( n4608 & ~n4609 ) ;
  assign n4611 = ( ~x44 & n4609 ) | ( ~x44 & n4610 ) | ( n4609 & n4610 ) ;
  assign n4612 = ( ~n4608 & n4610 ) | ( ~n4608 & n4611 ) | ( n4610 & n4611 ) ;
  assign n4613 = x44 & x45 ;
  assign n4614 = x44 | x45 ;
  assign n4615 = ~n4613 & n4614 ;
  assign n4616 = x64 & n4615 ;
  assign n4617 = x44 & ~n4478 ;
  assign n4618 = ( n4612 & n4616 ) | ( n4612 & n4617 ) | ( n4616 & n4617 ) ;
  assign n4619 = ( ~n4612 & n4616 ) | ( ~n4612 & n4617 ) | ( n4616 & n4617 ) ;
  assign n4620 = ( n4612 & ~n4618 ) | ( n4612 & n4619 ) | ( ~n4618 & n4619 ) ;
  assign n4621 = n245 & n3715 ;
  assign n4622 = x69 & n3719 ;
  assign n4623 = x70 | n4622 ;
  assign n4624 = ( n3721 & n4622 ) | ( n3721 & n4623 ) | ( n4622 & n4623 ) ;
  assign n4625 = x68 & n3922 ;
  assign n4626 = n4624 | n4625 ;
  assign n4627 = ( x41 & n4621 ) | ( x41 & ~n4626 ) | ( n4621 & ~n4626 ) ;
  assign n4628 = ( ~x41 & n4626 ) | ( ~x41 & n4627 ) | ( n4626 & n4627 ) ;
  assign n4629 = ( ~n4621 & n4627 ) | ( ~n4621 & n4628 ) | ( n4627 & n4628 ) ;
  assign n4630 = ( n4481 & n4620 ) | ( n4481 & n4629 ) | ( n4620 & n4629 ) ;
  assign n4631 = ( ~n4481 & n4620 ) | ( ~n4481 & n4629 ) | ( n4620 & n4629 ) ;
  assign n4632 = ( n4481 & ~n4630 ) | ( n4481 & n4631 ) | ( ~n4630 & n4631 ) ;
  assign n4633 = n390 & n3224 ;
  assign n4634 = x72 & n3228 ;
  assign n4635 = x73 | n4634 ;
  assign n4636 = ( n3230 & n4634 ) | ( n3230 & n4635 ) | ( n4634 & n4635 ) ;
  assign n4637 = x71 & n3413 ;
  assign n4638 = n4636 | n4637 ;
  assign n4639 = ( x38 & n4633 ) | ( x38 & ~n4638 ) | ( n4633 & ~n4638 ) ;
  assign n4640 = ( ~x38 & n4638 ) | ( ~x38 & n4639 ) | ( n4638 & n4639 ) ;
  assign n4641 = ( ~n4633 & n4639 ) | ( ~n4633 & n4640 ) | ( n4639 & n4640 ) ;
  assign n4642 = ( n4484 & n4632 ) | ( n4484 & n4641 ) | ( n4632 & n4641 ) ;
  assign n4643 = ( ~n4484 & n4632 ) | ( ~n4484 & n4641 ) | ( n4632 & n4641 ) ;
  assign n4644 = ( n4484 & ~n4642 ) | ( n4484 & n4643 ) | ( ~n4642 & n4643 ) ;
  assign n4645 = ( n4487 & n4603 ) | ( n4487 & n4644 ) | ( n4603 & n4644 ) ;
  assign n4646 = ( ~n4487 & n4603 ) | ( ~n4487 & n4644 ) | ( n4603 & n4644 ) ;
  assign n4647 = ( n4487 & ~n4645 ) | ( n4487 & n4646 ) | ( ~n4645 & n4646 ) ;
  assign n4648 = ( n4490 & n4594 ) | ( n4490 & n4647 ) | ( n4594 & n4647 ) ;
  assign n4649 = ( ~n4490 & n4594 ) | ( ~n4490 & n4647 ) | ( n4594 & n4647 ) ;
  assign n4650 = ( n4490 & ~n4648 ) | ( n4490 & n4649 ) | ( ~n4648 & n4649 ) ;
  assign n4651 = ( n4493 & n4585 ) | ( n4493 & n4650 ) | ( n4585 & n4650 ) ;
  assign n4652 = ( ~n4493 & n4585 ) | ( ~n4493 & n4650 ) | ( n4585 & n4650 ) ;
  assign n4653 = ( n4493 & ~n4651 ) | ( n4493 & n4652 ) | ( ~n4651 & n4652 ) ;
  assign n4654 = n1262 & n1617 ;
  assign n4655 = x84 & n1621 ;
  assign n4656 = x85 | n4655 ;
  assign n4657 = ( n1623 & n4655 ) | ( n1623 & n4656 ) | ( n4655 & n4656 ) ;
  assign n4658 = x83 & n1749 ;
  assign n4659 = n4657 | n4658 ;
  assign n4660 = ( x26 & n4654 ) | ( x26 & ~n4659 ) | ( n4654 & ~n4659 ) ;
  assign n4661 = ( ~x26 & n4659 ) | ( ~x26 & n4660 ) | ( n4659 & n4660 ) ;
  assign n4662 = ( ~n4654 & n4660 ) | ( ~n4654 & n4661 ) | ( n4660 & n4661 ) ;
  assign n4663 = ( n4505 & n4653 ) | ( n4505 & n4662 ) | ( n4653 & n4662 ) ;
  assign n4664 = ( ~n4505 & n4653 ) | ( ~n4505 & n4662 ) | ( n4653 & n4662 ) ;
  assign n4665 = ( n4505 & ~n4663 ) | ( n4505 & n4664 ) | ( ~n4663 & n4664 ) ;
  assign n4666 = n1297 & n1481 ;
  assign n4667 = x87 & n1301 ;
  assign n4668 = x88 | n4667 ;
  assign n4669 = ( n1303 & n4667 ) | ( n1303 & n4668 ) | ( n4667 & n4668 ) ;
  assign n4670 = x86 & n1426 ;
  assign n4671 = n4669 | n4670 ;
  assign n4672 = ( x23 & n4666 ) | ( x23 & ~n4671 ) | ( n4666 & ~n4671 ) ;
  assign n4673 = ( ~x23 & n4671 ) | ( ~x23 & n4672 ) | ( n4671 & n4672 ) ;
  assign n4674 = ( ~n4666 & n4672 ) | ( ~n4666 & n4673 ) | ( n4672 & n4673 ) ;
  assign n4675 = ( n4517 & n4665 ) | ( n4517 & n4674 ) | ( n4665 & n4674 ) ;
  assign n4676 = ( ~n4517 & n4665 ) | ( ~n4517 & n4674 ) | ( n4665 & n4674 ) ;
  assign n4677 = ( n4517 & ~n4675 ) | ( n4517 & n4676 ) | ( ~n4675 & n4676 ) ;
  assign n4678 = n1016 & n1914 ;
  assign n4679 = x90 & n1020 ;
  assign n4680 = x91 | n4679 ;
  assign n4681 = ( n1022 & n4679 ) | ( n1022 & n4680 ) | ( n4679 & n4680 ) ;
  assign n4682 = x89 & n1145 ;
  assign n4683 = n4681 | n4682 ;
  assign n4684 = ( x20 & n4678 ) | ( x20 & ~n4683 ) | ( n4678 & ~n4683 ) ;
  assign n4685 = ( ~x20 & n4683 ) | ( ~x20 & n4684 ) | ( n4683 & n4684 ) ;
  assign n4686 = ( ~n4678 & n4684 ) | ( ~n4678 & n4685 ) | ( n4684 & n4685 ) ;
  assign n4687 = ( n4520 & n4677 ) | ( n4520 & n4686 ) | ( n4677 & n4686 ) ;
  assign n4688 = ( ~n4520 & n4677 ) | ( ~n4520 & n4686 ) | ( n4677 & n4686 ) ;
  assign n4689 = ( n4520 & ~n4687 ) | ( n4520 & n4688 ) | ( ~n4687 & n4688 ) ;
  assign n4690 = ( n4523 & n4576 ) | ( n4523 & n4689 ) | ( n4576 & n4689 ) ;
  assign n4691 = ( ~n4523 & n4576 ) | ( ~n4523 & n4689 ) | ( n4576 & n4689 ) ;
  assign n4692 = ( n4523 & ~n4690 ) | ( n4523 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n4693 = n583 & n2585 ;
  assign n4694 = x96 & n587 ;
  assign n4695 = x97 | n4694 ;
  assign n4696 = ( n589 & n4694 ) | ( n589 & n4695 ) | ( n4694 & n4695 ) ;
  assign n4697 = x95 & n676 ;
  assign n4698 = n4696 | n4697 ;
  assign n4699 = ( x14 & n4693 ) | ( x14 & ~n4698 ) | ( n4693 & ~n4698 ) ;
  assign n4700 = ( ~x14 & n4698 ) | ( ~x14 & n4699 ) | ( n4698 & n4699 ) ;
  assign n4701 = ( ~n4693 & n4699 ) | ( ~n4693 & n4700 ) | ( n4699 & n4700 ) ;
  assign n4702 = ( n4526 & n4692 ) | ( n4526 & n4701 ) | ( n4692 & n4701 ) ;
  assign n4703 = ( ~n4526 & n4692 ) | ( ~n4526 & n4701 ) | ( n4692 & n4701 ) ;
  assign n4704 = ( n4526 & ~n4702 ) | ( n4526 & n4703 ) | ( ~n4702 & n4703 ) ;
  assign n4705 = ( n4538 & n4567 ) | ( n4538 & n4704 ) | ( n4567 & n4704 ) ;
  assign n4706 = ( ~n4538 & n4567 ) | ( ~n4538 & n4704 ) | ( n4567 & n4704 ) ;
  assign n4707 = ( n4538 & ~n4705 ) | ( n4538 & n4706 ) | ( ~n4705 & n4706 ) ;
  assign n4708 = n291 & n3650 ;
  assign n4709 = x102 & n295 ;
  assign n4710 = x103 | n4709 ;
  assign n4711 = ( n297 & n4709 ) | ( n297 & n4710 ) | ( n4709 & n4710 ) ;
  assign n4712 = x101 & n330 ;
  assign n4713 = n4711 | n4712 ;
  assign n4714 = ( x8 & n4708 ) | ( x8 & ~n4713 ) | ( n4708 & ~n4713 ) ;
  assign n4715 = ( ~x8 & n4713 ) | ( ~x8 & n4714 ) | ( n4713 & n4714 ) ;
  assign n4716 = ( ~n4708 & n4714 ) | ( ~n4708 & n4715 ) | ( n4714 & n4715 ) ;
  assign n4717 = ( n4550 & n4707 ) | ( n4550 & n4716 ) | ( n4707 & n4716 ) ;
  assign n4718 = ( ~n4550 & n4707 ) | ( ~n4550 & n4716 ) | ( n4707 & n4716 ) ;
  assign n4719 = ( n4550 & ~n4717 ) | ( n4550 & n4718 ) | ( ~n4717 & n4718 ) ;
  assign n4720 = n186 & n4013 ;
  assign n4721 = x105 & n190 ;
  assign n4722 = x106 | n4721 ;
  assign n4723 = ( n192 & n4721 ) | ( n192 & n4722 ) | ( n4721 & n4722 ) ;
  assign n4724 = x104 & n220 ;
  assign n4725 = n4723 | n4724 ;
  assign n4726 = ( x5 & n4720 ) | ( x5 & ~n4725 ) | ( n4720 & ~n4725 ) ;
  assign n4727 = ( ~x5 & n4725 ) | ( ~x5 & n4726 ) | ( n4725 & n4726 ) ;
  assign n4728 = ( ~n4720 & n4726 ) | ( ~n4720 & n4727 ) | ( n4726 & n4727 ) ;
  assign n4729 = ( n4553 & n4719 ) | ( n4553 & n4728 ) | ( n4719 & n4728 ) ;
  assign n4730 = ( ~n4553 & n4719 ) | ( ~n4553 & n4728 ) | ( n4719 & n4728 ) ;
  assign n4731 = ( n4553 & ~n4729 ) | ( n4553 & n4730 ) | ( ~n4729 & n4730 ) ;
  assign n4732 = ( x108 & x109 ) | ( x108 & n4375 ) | ( x109 & n4375 ) ;
  assign n4733 = ( x108 & ~x109 ) | ( x108 & n4375 ) | ( ~x109 & n4375 ) ;
  assign n4734 = ( x109 & ~n4732 ) | ( x109 & n4733 ) | ( ~n4732 & n4733 ) ;
  assign n4735 = n136 & n4734 ;
  assign n4736 = x108 & n138 ;
  assign n4737 = x109 | n4736 ;
  assign n4738 = ( n141 & n4736 ) | ( n141 & n4737 ) | ( n4736 & n4737 ) ;
  assign n4739 = x107 & n154 ;
  assign n4740 = n4738 | n4739 ;
  assign n4741 = ( x2 & n4735 ) | ( x2 & ~n4740 ) | ( n4735 & ~n4740 ) ;
  assign n4742 = ( ~x2 & n4740 ) | ( ~x2 & n4741 ) | ( n4740 & n4741 ) ;
  assign n4743 = ( ~n4735 & n4741 ) | ( ~n4735 & n4742 ) | ( n4741 & n4742 ) ;
  assign n4744 = ( n4556 & n4731 ) | ( n4556 & n4743 ) | ( n4731 & n4743 ) ;
  assign n4745 = ( ~n4556 & n4731 ) | ( ~n4556 & n4743 ) | ( n4731 & n4743 ) ;
  assign n4746 = ( n4556 & ~n4744 ) | ( n4556 & n4745 ) | ( ~n4744 & n4745 ) ;
  assign n4747 = n186 & n4362 ;
  assign n4748 = x106 & n190 ;
  assign n4749 = x107 | n4748 ;
  assign n4750 = ( n192 & n4748 ) | ( n192 & n4749 ) | ( n4748 & n4749 ) ;
  assign n4751 = x105 & n220 ;
  assign n4752 = n4750 | n4751 ;
  assign n4753 = ( x5 & n4747 ) | ( x5 & ~n4752 ) | ( n4747 & ~n4752 ) ;
  assign n4754 = ( ~x5 & n4752 ) | ( ~x5 & n4753 ) | ( n4752 & n4753 ) ;
  assign n4755 = ( ~n4747 & n4753 ) | ( ~n4747 & n4754 ) | ( n4753 & n4754 ) ;
  assign n4756 = n810 & n2434 ;
  assign n4757 = x94 & n814 ;
  assign n4758 = x95 | n4757 ;
  assign n4759 = ( n816 & n4757 ) | ( n816 & n4758 ) | ( n4757 & n4758 ) ;
  assign n4760 = x93 & n885 ;
  assign n4761 = n4759 | n4760 ;
  assign n4762 = ( x17 & n4756 ) | ( x17 & ~n4761 ) | ( n4756 & ~n4761 ) ;
  assign n4763 = ( ~x17 & n4761 ) | ( ~x17 & n4762 ) | ( n4761 & n4762 ) ;
  assign n4764 = ( ~n4756 & n4762 ) | ( ~n4756 & n4763 ) | ( n4762 & n4763 ) ;
  assign n4765 = n1016 & n2042 ;
  assign n4766 = x91 & n1020 ;
  assign n4767 = x92 | n4766 ;
  assign n4768 = ( n1022 & n4766 ) | ( n1022 & n4767 ) | ( n4766 & n4767 ) ;
  assign n4769 = x90 & n1145 ;
  assign n4770 = n4768 | n4769 ;
  assign n4771 = ( x20 & n4765 ) | ( x20 & ~n4770 ) | ( n4765 & ~n4770 ) ;
  assign n4772 = ( ~x20 & n4770 ) | ( ~x20 & n4771 ) | ( n4770 & n4771 ) ;
  assign n4773 = ( ~n4765 & n4771 ) | ( ~n4765 & n4772 ) | ( n4771 & n4772 ) ;
  assign n4774 = n569 & n2766 ;
  assign n4775 = x76 & n2770 ;
  assign n4776 = x77 | n4775 ;
  assign n4777 = ( n2772 & n4775 ) | ( n2772 & n4776 ) | ( n4775 & n4776 ) ;
  assign n4778 = x75 & n2943 ;
  assign n4779 = n4777 | n4778 ;
  assign n4780 = ( x35 & n4774 ) | ( x35 & ~n4779 ) | ( n4774 & ~n4779 ) ;
  assign n4781 = ( ~x35 & n4779 ) | ( ~x35 & n4780 ) | ( n4779 & n4780 ) ;
  assign n4782 = ( ~n4774 & n4780 ) | ( ~n4774 & n4781 ) | ( n4780 & n4781 ) ;
  assign n4783 = x47 & n4616 ;
  assign n4784 = x46 | x47 ;
  assign n4785 = ( x46 & x47 ) | ( x46 & ~n4784 ) | ( x47 & ~n4784 ) ;
  assign n4786 = n4784 & ~n4785 ;
  assign n4787 = n4615 & n4786 ;
  assign n4788 = n133 & n4787 ;
  assign n4789 = ~x44 & x46 ;
  assign n4790 = x45 & x46 ;
  assign n4791 = ( n4613 & n4789 ) | ( n4613 & ~n4790 ) | ( n4789 & ~n4790 ) ;
  assign n4792 = x64 & n4791 ;
  assign n4793 = ( n4615 & ~n4784 ) | ( n4615 & n4785 ) | ( ~n4784 & n4785 ) ;
  assign n4794 = x65 | n4792 ;
  assign n4795 = ( n4792 & n4793 ) | ( n4792 & n4794 ) | ( n4793 & n4794 ) ;
  assign n4796 = ( n4783 & n4788 ) | ( n4783 & n4795 ) | ( n4788 & n4795 ) ;
  assign n4797 = n4788 | n4795 ;
  assign n4798 = ~n4783 & n4797 ;
  assign n4799 = ( n4783 & ~n4796 ) | ( n4783 & n4798 ) | ( ~n4796 & n4798 ) ;
  assign n4800 = x67 & n4231 ;
  assign n4801 = x68 | n4800 ;
  assign n4802 = ( n4233 & n4800 ) | ( n4233 & n4801 ) | ( n4800 & n4801 ) ;
  assign n4803 = x66 & n4470 ;
  assign n4804 = n4802 | n4803 ;
  assign n4805 = n201 & n4227 ;
  assign n4806 = ( x44 & n4804 ) | ( x44 & ~n4805 ) | ( n4804 & ~n4805 ) ;
  assign n4807 = ( ~x44 & n4805 ) | ( ~x44 & n4806 ) | ( n4805 & n4806 ) ;
  assign n4808 = ( ~n4804 & n4806 ) | ( ~n4804 & n4807 ) | ( n4806 & n4807 ) ;
  assign n4809 = ( n4618 & n4799 ) | ( n4618 & n4808 ) | ( n4799 & n4808 ) ;
  assign n4810 = ( ~n4618 & n4799 ) | ( ~n4618 & n4808 ) | ( n4799 & n4808 ) ;
  assign n4811 = ( n4618 & ~n4809 ) | ( n4618 & n4810 ) | ( ~n4809 & n4810 ) ;
  assign n4812 = n277 & n3715 ;
  assign n4813 = x70 & n3719 ;
  assign n4814 = x71 | n4813 ;
  assign n4815 = ( n3721 & n4813 ) | ( n3721 & n4814 ) | ( n4813 & n4814 ) ;
  assign n4816 = x69 & n3922 ;
  assign n4817 = n4815 | n4816 ;
  assign n4818 = ( x41 & n4812 ) | ( x41 & ~n4817 ) | ( n4812 & ~n4817 ) ;
  assign n4819 = ( ~x41 & n4817 ) | ( ~x41 & n4818 ) | ( n4817 & n4818 ) ;
  assign n4820 = ( ~n4812 & n4818 ) | ( ~n4812 & n4819 ) | ( n4818 & n4819 ) ;
  assign n4821 = ( n4630 & n4811 ) | ( n4630 & n4820 ) | ( n4811 & n4820 ) ;
  assign n4822 = ( ~n4630 & n4811 ) | ( ~n4630 & n4820 ) | ( n4811 & n4820 ) ;
  assign n4823 = ( n4630 & ~n4821 ) | ( n4630 & n4822 ) | ( ~n4821 & n4822 ) ;
  assign n4824 = n446 & n3224 ;
  assign n4825 = x73 & n3228 ;
  assign n4826 = x74 | n4825 ;
  assign n4827 = ( n3230 & n4825 ) | ( n3230 & n4826 ) | ( n4825 & n4826 ) ;
  assign n4828 = x72 & n3413 ;
  assign n4829 = n4827 | n4828 ;
  assign n4830 = ( x38 & n4824 ) | ( x38 & ~n4829 ) | ( n4824 & ~n4829 ) ;
  assign n4831 = ( ~x38 & n4829 ) | ( ~x38 & n4830 ) | ( n4829 & n4830 ) ;
  assign n4832 = ( ~n4824 & n4830 ) | ( ~n4824 & n4831 ) | ( n4830 & n4831 ) ;
  assign n4833 = ( n4642 & n4823 ) | ( n4642 & n4832 ) | ( n4823 & n4832 ) ;
  assign n4834 = ( ~n4642 & n4823 ) | ( ~n4642 & n4832 ) | ( n4823 & n4832 ) ;
  assign n4835 = ( n4642 & ~n4833 ) | ( n4642 & n4834 ) | ( ~n4833 & n4834 ) ;
  assign n4836 = ( n4645 & n4782 ) | ( n4645 & n4835 ) | ( n4782 & n4835 ) ;
  assign n4837 = ( ~n4645 & n4782 ) | ( ~n4645 & n4835 ) | ( n4782 & n4835 ) ;
  assign n4838 = ( n4645 & ~n4836 ) | ( n4645 & n4837 ) | ( ~n4836 & n4837 ) ;
  assign n4839 = n769 & n2320 ;
  assign n4840 = x79 & n2324 ;
  assign n4841 = x80 | n4840 ;
  assign n4842 = ( n2326 & n4840 ) | ( n2326 & n4841 ) | ( n4840 & n4841 ) ;
  assign n4843 = x78 & n2497 ;
  assign n4844 = n4842 | n4843 ;
  assign n4845 = ( x32 & n4839 ) | ( x32 & ~n4844 ) | ( n4839 & ~n4844 ) ;
  assign n4846 = ( ~x32 & n4844 ) | ( ~x32 & n4845 ) | ( n4844 & n4845 ) ;
  assign n4847 = ( ~n4839 & n4845 ) | ( ~n4839 & n4846 ) | ( n4845 & n4846 ) ;
  assign n4848 = ( n4648 & n4838 ) | ( n4648 & n4847 ) | ( n4838 & n4847 ) ;
  assign n4849 = ( ~n4648 & n4838 ) | ( ~n4648 & n4847 ) | ( n4838 & n4847 ) ;
  assign n4850 = ( n4648 & ~n4848 ) | ( n4648 & n4849 ) | ( ~n4848 & n4849 ) ;
  assign n4851 = n1082 & n1949 ;
  assign n4852 = x82 & n1953 ;
  assign n4853 = x83 | n4852 ;
  assign n4854 = ( n1955 & n4852 ) | ( n1955 & n4853 ) | ( n4852 & n4853 ) ;
  assign n4855 = x81 & n2114 ;
  assign n4856 = n4854 | n4855 ;
  assign n4857 = ( x29 & n4851 ) | ( x29 & ~n4856 ) | ( n4851 & ~n4856 ) ;
  assign n4858 = ( ~x29 & n4856 ) | ( ~x29 & n4857 ) | ( n4856 & n4857 ) ;
  assign n4859 = ( ~n4851 & n4857 ) | ( ~n4851 & n4858 ) | ( n4857 & n4858 ) ;
  assign n4860 = ( n4651 & n4850 ) | ( n4651 & n4859 ) | ( n4850 & n4859 ) ;
  assign n4861 = ( ~n4651 & n4850 ) | ( ~n4651 & n4859 ) | ( n4850 & n4859 ) ;
  assign n4862 = ( n4651 & ~n4860 ) | ( n4651 & n4861 ) | ( ~n4860 & n4861 ) ;
  assign n4863 = n1366 & n1617 ;
  assign n4864 = x85 & n1621 ;
  assign n4865 = x86 | n4864 ;
  assign n4866 = ( n1623 & n4864 ) | ( n1623 & n4865 ) | ( n4864 & n4865 ) ;
  assign n4867 = x84 & n1749 ;
  assign n4868 = n4866 | n4867 ;
  assign n4869 = ( x26 & n4863 ) | ( x26 & ~n4868 ) | ( n4863 & ~n4868 ) ;
  assign n4870 = ( ~x26 & n4868 ) | ( ~x26 & n4869 ) | ( n4868 & n4869 ) ;
  assign n4871 = ( ~n4863 & n4869 ) | ( ~n4863 & n4870 ) | ( n4869 & n4870 ) ;
  assign n4872 = ( n4663 & n4862 ) | ( n4663 & n4871 ) | ( n4862 & n4871 ) ;
  assign n4873 = ( ~n4663 & n4862 ) | ( ~n4663 & n4871 ) | ( n4862 & n4871 ) ;
  assign n4874 = ( n4663 & ~n4872 ) | ( n4663 & n4873 ) | ( ~n4872 & n4873 ) ;
  assign n4875 = n1297 & n1585 ;
  assign n4876 = x88 & n1301 ;
  assign n4877 = x89 | n4876 ;
  assign n4878 = ( n1303 & n4876 ) | ( n1303 & n4877 ) | ( n4876 & n4877 ) ;
  assign n4879 = x87 & n1426 ;
  assign n4880 = n4878 | n4879 ;
  assign n4881 = ( x23 & n4875 ) | ( x23 & ~n4880 ) | ( n4875 & ~n4880 ) ;
  assign n4882 = ( ~x23 & n4880 ) | ( ~x23 & n4881 ) | ( n4880 & n4881 ) ;
  assign n4883 = ( ~n4875 & n4881 ) | ( ~n4875 & n4882 ) | ( n4881 & n4882 ) ;
  assign n4884 = ( n4675 & n4874 ) | ( n4675 & n4883 ) | ( n4874 & n4883 ) ;
  assign n4885 = ( ~n4675 & n4874 ) | ( ~n4675 & n4883 ) | ( n4874 & n4883 ) ;
  assign n4886 = ( n4675 & ~n4884 ) | ( n4675 & n4885 ) | ( ~n4884 & n4885 ) ;
  assign n4887 = ( n4687 & n4773 ) | ( n4687 & n4886 ) | ( n4773 & n4886 ) ;
  assign n4888 = ( ~n4687 & n4773 ) | ( ~n4687 & n4886 ) | ( n4773 & n4886 ) ;
  assign n4889 = ( n4687 & ~n4887 ) | ( n4687 & n4888 ) | ( ~n4887 & n4888 ) ;
  assign n4890 = ( n4690 & n4764 ) | ( n4690 & n4889 ) | ( n4764 & n4889 ) ;
  assign n4891 = ( ~n4690 & n4764 ) | ( ~n4690 & n4889 ) | ( n4764 & n4889 ) ;
  assign n4892 = ( n4690 & ~n4890 ) | ( n4690 & n4891 ) | ( ~n4890 & n4891 ) ;
  assign n4893 = n583 & n2725 ;
  assign n4894 = x97 & n587 ;
  assign n4895 = x98 | n4894 ;
  assign n4896 = ( n589 & n4894 ) | ( n589 & n4895 ) | ( n4894 & n4895 ) ;
  assign n4897 = x96 & n676 ;
  assign n4898 = n4896 | n4897 ;
  assign n4899 = ( x14 & n4893 ) | ( x14 & ~n4898 ) | ( n4893 & ~n4898 ) ;
  assign n4900 = ( ~x14 & n4898 ) | ( ~x14 & n4899 ) | ( n4898 & n4899 ) ;
  assign n4901 = ( ~n4893 & n4899 ) | ( ~n4893 & n4900 ) | ( n4899 & n4900 ) ;
  assign n4902 = ( n4702 & n4892 ) | ( n4702 & n4901 ) | ( n4892 & n4901 ) ;
  assign n4903 = ( ~n4702 & n4892 ) | ( ~n4702 & n4901 ) | ( n4892 & n4901 ) ;
  assign n4904 = ( n4702 & ~n4902 ) | ( n4702 & n4903 ) | ( ~n4902 & n4903 ) ;
  assign n4905 = n407 & n3326 ;
  assign n4906 = x100 & n411 ;
  assign n4907 = x101 | n4906 ;
  assign n4908 = ( n413 & n4906 ) | ( n413 & n4907 ) | ( n4906 & n4907 ) ;
  assign n4909 = x99 & n491 ;
  assign n4910 = n4908 | n4909 ;
  assign n4911 = ( x11 & n4905 ) | ( x11 & ~n4910 ) | ( n4905 & ~n4910 ) ;
  assign n4912 = ( ~x11 & n4910 ) | ( ~x11 & n4911 ) | ( n4910 & n4911 ) ;
  assign n4913 = ( ~n4905 & n4911 ) | ( ~n4905 & n4912 ) | ( n4911 & n4912 ) ;
  assign n4914 = ( n4705 & n4904 ) | ( n4705 & n4913 ) | ( n4904 & n4913 ) ;
  assign n4915 = ( ~n4705 & n4904 ) | ( ~n4705 & n4913 ) | ( n4904 & n4913 ) ;
  assign n4916 = ( n4705 & ~n4914 ) | ( n4705 & n4915 ) | ( ~n4914 & n4915 ) ;
  assign n4917 = n291 & n3665 ;
  assign n4918 = x103 & n295 ;
  assign n4919 = x104 | n4918 ;
  assign n4920 = ( n297 & n4918 ) | ( n297 & n4919 ) | ( n4918 & n4919 ) ;
  assign n4921 = x102 & n330 ;
  assign n4922 = n4920 | n4921 ;
  assign n4923 = ( x8 & n4917 ) | ( x8 & ~n4922 ) | ( n4917 & ~n4922 ) ;
  assign n4924 = ( ~x8 & n4922 ) | ( ~x8 & n4923 ) | ( n4922 & n4923 ) ;
  assign n4925 = ( ~n4917 & n4923 ) | ( ~n4917 & n4924 ) | ( n4923 & n4924 ) ;
  assign n4926 = ( n4717 & n4916 ) | ( n4717 & n4925 ) | ( n4916 & n4925 ) ;
  assign n4927 = ( ~n4717 & n4916 ) | ( ~n4717 & n4925 ) | ( n4916 & n4925 ) ;
  assign n4928 = ( n4717 & ~n4926 ) | ( n4717 & n4927 ) | ( ~n4926 & n4927 ) ;
  assign n4929 = ( n4729 & n4755 ) | ( n4729 & n4928 ) | ( n4755 & n4928 ) ;
  assign n4930 = ( ~n4729 & n4755 ) | ( ~n4729 & n4928 ) | ( n4755 & n4928 ) ;
  assign n4931 = ( n4729 & ~n4929 ) | ( n4729 & n4930 ) | ( ~n4929 & n4930 ) ;
  assign n4932 = ( x109 & x110 ) | ( x109 & n4732 ) | ( x110 & n4732 ) ;
  assign n4933 = ( x109 & ~x110 ) | ( x109 & n4732 ) | ( ~x110 & n4732 ) ;
  assign n4934 = ( x110 & ~n4932 ) | ( x110 & n4933 ) | ( ~n4932 & n4933 ) ;
  assign n4935 = n136 & n4934 ;
  assign n4936 = x109 & n138 ;
  assign n4937 = x110 | n4936 ;
  assign n4938 = ( n141 & n4936 ) | ( n141 & n4937 ) | ( n4936 & n4937 ) ;
  assign n4939 = x108 & n154 ;
  assign n4940 = n4938 | n4939 ;
  assign n4941 = ( x2 & n4935 ) | ( x2 & ~n4940 ) | ( n4935 & ~n4940 ) ;
  assign n4942 = ( ~x2 & n4940 ) | ( ~x2 & n4941 ) | ( n4940 & n4941 ) ;
  assign n4943 = ( ~n4935 & n4941 ) | ( ~n4935 & n4942 ) | ( n4941 & n4942 ) ;
  assign n4944 = ( n4744 & n4931 ) | ( n4744 & n4943 ) | ( n4931 & n4943 ) ;
  assign n4945 = ( ~n4744 & n4931 ) | ( ~n4744 & n4943 ) | ( n4931 & n4943 ) ;
  assign n4946 = ( n4744 & ~n4944 ) | ( n4744 & n4945 ) | ( ~n4944 & n4945 ) ;
  assign n4947 = n186 & n4377 ;
  assign n4948 = x107 & n190 ;
  assign n4949 = x108 | n4948 ;
  assign n4950 = ( n192 & n4948 ) | ( n192 & n4949 ) | ( n4948 & n4949 ) ;
  assign n4951 = x106 & n220 ;
  assign n4952 = n4950 | n4951 ;
  assign n4953 = ( x5 & n4947 ) | ( x5 & ~n4952 ) | ( n4947 & ~n4952 ) ;
  assign n4954 = ( ~x5 & n4952 ) | ( ~x5 & n4953 ) | ( n4952 & n4953 ) ;
  assign n4955 = ( ~n4947 & n4953 ) | ( ~n4947 & n4954 ) | ( n4953 & n4954 ) ;
  assign n4956 = n810 & n2449 ;
  assign n4957 = x95 & n814 ;
  assign n4958 = x96 | n4957 ;
  assign n4959 = ( n816 & n4957 ) | ( n816 & n4958 ) | ( n4957 & n4958 ) ;
  assign n4960 = x94 & n885 ;
  assign n4961 = n4959 | n4960 ;
  assign n4962 = ( x17 & n4956 ) | ( x17 & ~n4961 ) | ( n4956 & ~n4961 ) ;
  assign n4963 = ( ~x17 & n4961 ) | ( ~x17 & n4962 ) | ( n4961 & n4962 ) ;
  assign n4964 = ( ~n4956 & n4962 ) | ( ~n4956 & n4963 ) | ( n4962 & n4963 ) ;
  assign n4965 = n1016 & n2057 ;
  assign n4966 = x92 & n1020 ;
  assign n4967 = x93 | n4966 ;
  assign n4968 = ( n1022 & n4966 ) | ( n1022 & n4967 ) | ( n4966 & n4967 ) ;
  assign n4969 = x91 & n1145 ;
  assign n4970 = n4968 | n4969 ;
  assign n4971 = ( x20 & n4965 ) | ( x20 & ~n4970 ) | ( n4965 & ~n4970 ) ;
  assign n4972 = ( ~x20 & n4970 ) | ( ~x20 & n4971 ) | ( n4970 & n4971 ) ;
  assign n4973 = ( ~n4965 & n4971 ) | ( ~n4965 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4974 = n1297 & n1701 ;
  assign n4975 = x89 & n1301 ;
  assign n4976 = x90 | n4975 ;
  assign n4977 = ( n1303 & n4975 ) | ( n1303 & n4976 ) | ( n4975 & n4976 ) ;
  assign n4978 = x88 & n1426 ;
  assign n4979 = n4977 | n4978 ;
  assign n4980 = ( x23 & n4974 ) | ( x23 & ~n4979 ) | ( n4974 & ~n4979 ) ;
  assign n4981 = ( ~x23 & n4979 ) | ( ~x23 & n4980 ) | ( n4979 & n4980 ) ;
  assign n4982 = ( ~n4974 & n4980 ) | ( ~n4974 & n4981 ) | ( n4980 & n4981 ) ;
  assign n4983 = n1097 & n1949 ;
  assign n4984 = x83 & n1953 ;
  assign n4985 = x84 | n4984 ;
  assign n4986 = ( n1955 & n4984 ) | ( n1955 & n4985 ) | ( n4984 & n4985 ) ;
  assign n4987 = x82 & n2114 ;
  assign n4988 = n4986 | n4987 ;
  assign n4989 = ( x29 & n4983 ) | ( x29 & ~n4988 ) | ( n4983 & ~n4988 ) ;
  assign n4990 = ( ~x29 & n4988 ) | ( ~x29 & n4989 ) | ( n4988 & n4989 ) ;
  assign n4991 = ( ~n4983 & n4989 ) | ( ~n4983 & n4990 ) | ( n4989 & n4990 ) ;
  assign n4992 = n910 & n2320 ;
  assign n4993 = x80 & n2324 ;
  assign n4994 = x81 | n4993 ;
  assign n4995 = ( n2326 & n4993 ) | ( n2326 & n4994 ) | ( n4993 & n4994 ) ;
  assign n4996 = x79 & n2497 ;
  assign n4997 = n4995 | n4996 ;
  assign n4998 = ( x32 & n4992 ) | ( x32 & ~n4997 ) | ( n4992 & ~n4997 ) ;
  assign n4999 = ( ~x32 & n4997 ) | ( ~x32 & n4998 ) | ( n4997 & n4998 ) ;
  assign n5000 = ( ~n4992 & n4998 ) | ( ~n4992 & n4999 ) | ( n4998 & n4999 ) ;
  assign n5001 = n461 & n3224 ;
  assign n5002 = x74 & n3228 ;
  assign n5003 = x75 | n5002 ;
  assign n5004 = ( n3230 & n5002 ) | ( n3230 & n5003 ) | ( n5002 & n5003 ) ;
  assign n5005 = x73 & n3413 ;
  assign n5006 = n5004 | n5005 ;
  assign n5007 = ( x38 & n5001 ) | ( x38 & ~n5006 ) | ( n5001 & ~n5006 ) ;
  assign n5008 = ( ~x38 & n5006 ) | ( ~x38 & n5007 ) | ( n5006 & n5007 ) ;
  assign n5009 = ( ~n5001 & n5007 ) | ( ~n5001 & n5008 ) | ( n5007 & n5008 ) ;
  assign n5010 = n346 & n3715 ;
  assign n5011 = x71 & n3719 ;
  assign n5012 = x72 | n5011 ;
  assign n5013 = ( n3721 & n5011 ) | ( n3721 & n5012 ) | ( n5011 & n5012 ) ;
  assign n5014 = x70 & n3922 ;
  assign n5015 = n5013 | n5014 ;
  assign n5016 = ( x41 & n5010 ) | ( x41 & ~n5015 ) | ( n5010 & ~n5015 ) ;
  assign n5017 = ( ~x41 & n5015 ) | ( ~x41 & n5016 ) | ( n5015 & n5016 ) ;
  assign n5018 = ( ~n5010 & n5016 ) | ( ~n5010 & n5017 ) | ( n5016 & n5017 ) ;
  assign n5019 = n230 & n4227 ;
  assign n5020 = x68 & n4231 ;
  assign n5021 = x69 | n5020 ;
  assign n5022 = ( n4233 & n5020 ) | ( n4233 & n5021 ) | ( n5020 & n5021 ) ;
  assign n5023 = x67 & n4470 ;
  assign n5024 = n5022 | n5023 ;
  assign n5025 = ( ~x44 & n5019 ) | ( ~x44 & n5024 ) | ( n5019 & n5024 ) ;
  assign n5026 = ( n5019 & n5024 ) | ( n5019 & ~n5025 ) | ( n5024 & ~n5025 ) ;
  assign n5027 = ( x44 & n5025 ) | ( x44 & ~n5026 ) | ( n5025 & ~n5026 ) ;
  assign n5028 = ( x47 & n4783 ) | ( x47 & n4797 ) | ( n4783 & n4797 ) ;
  assign n5029 = ( x44 & ~x46 ) | ( x44 & n4786 ) | ( ~x46 & n4786 ) ;
  assign n5030 = ( ~n4614 & n4790 ) | ( ~n4614 & n5029 ) | ( n4790 & n5029 ) ;
  assign n5031 = x64 & n5030 ;
  assign n5032 = x65 & n4791 ;
  assign n5033 = x66 | n5032 ;
  assign n5034 = ( n4793 & n5032 ) | ( n4793 & n5033 ) | ( n5032 & n5033 ) ;
  assign n5035 = ( n151 & n152 ) | ( n151 & n4787 ) | ( n152 & n4787 ) ;
  assign n5036 = ( ~n5031 & n5034 ) | ( ~n5031 & n5035 ) | ( n5034 & n5035 ) ;
  assign n5037 = n5031 | n5036 ;
  assign n5038 = n5028 | n5037 ;
  assign n5039 = ( n5028 & n5037 ) | ( n5028 & ~n5038 ) | ( n5037 & ~n5038 ) ;
  assign n5040 = n5038 & ~n5039 ;
  assign n5041 = ( n4809 & n5027 ) | ( n4809 & n5040 ) | ( n5027 & n5040 ) ;
  assign n5042 = ( ~n4809 & n5027 ) | ( ~n4809 & n5040 ) | ( n5027 & n5040 ) ;
  assign n5043 = ( n4809 & ~n5041 ) | ( n4809 & n5042 ) | ( ~n5041 & n5042 ) ;
  assign n5044 = ( n4821 & n5018 ) | ( n4821 & n5043 ) | ( n5018 & n5043 ) ;
  assign n5045 = ( ~n4821 & n5018 ) | ( ~n4821 & n5043 ) | ( n5018 & n5043 ) ;
  assign n5046 = ( n4821 & ~n5044 ) | ( n4821 & n5045 ) | ( ~n5044 & n5045 ) ;
  assign n5047 = ( n4833 & n5009 ) | ( n4833 & n5046 ) | ( n5009 & n5046 ) ;
  assign n5048 = ( ~n4833 & n5009 ) | ( ~n4833 & n5046 ) | ( n5009 & n5046 ) ;
  assign n5049 = ( n4833 & ~n5047 ) | ( n4833 & n5048 ) | ( ~n5047 & n5048 ) ;
  assign n5050 = n637 & n2766 ;
  assign n5051 = x77 & n2770 ;
  assign n5052 = x78 | n5051 ;
  assign n5053 = ( n2772 & n5051 ) | ( n2772 & n5052 ) | ( n5051 & n5052 ) ;
  assign n5054 = x76 & n2943 ;
  assign n5055 = n5053 | n5054 ;
  assign n5056 = ( x35 & n5050 ) | ( x35 & ~n5055 ) | ( n5050 & ~n5055 ) ;
  assign n5057 = ( ~x35 & n5055 ) | ( ~x35 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5058 = ( ~n5050 & n5056 ) | ( ~n5050 & n5057 ) | ( n5056 & n5057 ) ;
  assign n5059 = ( n4836 & n5049 ) | ( n4836 & n5058 ) | ( n5049 & n5058 ) ;
  assign n5060 = ( ~n4836 & n5049 ) | ( ~n4836 & n5058 ) | ( n5049 & n5058 ) ;
  assign n5061 = ( n4836 & ~n5059 ) | ( n4836 & n5060 ) | ( ~n5059 & n5060 ) ;
  assign n5062 = ( n4848 & n5000 ) | ( n4848 & n5061 ) | ( n5000 & n5061 ) ;
  assign n5063 = ( ~n4848 & n5000 ) | ( ~n4848 & n5061 ) | ( n5000 & n5061 ) ;
  assign n5064 = ( n4848 & ~n5062 ) | ( n4848 & n5063 ) | ( ~n5062 & n5063 ) ;
  assign n5065 = ( n4860 & n4991 ) | ( n4860 & n5064 ) | ( n4991 & n5064 ) ;
  assign n5066 = ( ~n4860 & n4991 ) | ( ~n4860 & n5064 ) | ( n4991 & n5064 ) ;
  assign n5067 = ( n4860 & ~n5065 ) | ( n4860 & n5066 ) | ( ~n5065 & n5066 ) ;
  assign n5068 = n1466 & n1617 ;
  assign n5069 = x86 & n1621 ;
  assign n5070 = x87 | n5069 ;
  assign n5071 = ( n1623 & n5069 ) | ( n1623 & n5070 ) | ( n5069 & n5070 ) ;
  assign n5072 = x85 & n1749 ;
  assign n5073 = n5071 | n5072 ;
  assign n5074 = ( x26 & n5068 ) | ( x26 & ~n5073 ) | ( n5068 & ~n5073 ) ;
  assign n5075 = ( ~x26 & n5073 ) | ( ~x26 & n5074 ) | ( n5073 & n5074 ) ;
  assign n5076 = ( ~n5068 & n5074 ) | ( ~n5068 & n5075 ) | ( n5074 & n5075 ) ;
  assign n5077 = ( n4872 & n5067 ) | ( n4872 & n5076 ) | ( n5067 & n5076 ) ;
  assign n5078 = ( ~n4872 & n5067 ) | ( ~n4872 & n5076 ) | ( n5067 & n5076 ) ;
  assign n5079 = ( n4872 & ~n5077 ) | ( n4872 & n5078 ) | ( ~n5077 & n5078 ) ;
  assign n5080 = ( n4884 & n4982 ) | ( n4884 & n5079 ) | ( n4982 & n5079 ) ;
  assign n5081 = ( ~n4884 & n4982 ) | ( ~n4884 & n5079 ) | ( n4982 & n5079 ) ;
  assign n5082 = ( n4884 & ~n5080 ) | ( n4884 & n5081 ) | ( ~n5080 & n5081 ) ;
  assign n5083 = ( n4887 & n4973 ) | ( n4887 & n5082 ) | ( n4973 & n5082 ) ;
  assign n5084 = ( ~n4887 & n4973 ) | ( ~n4887 & n5082 ) | ( n4973 & n5082 ) ;
  assign n5085 = ( n4887 & ~n5083 ) | ( n4887 & n5084 ) | ( ~n5083 & n5084 ) ;
  assign n5086 = ( n4890 & n4964 ) | ( n4890 & n5085 ) | ( n4964 & n5085 ) ;
  assign n5087 = ( ~n4890 & n4964 ) | ( ~n4890 & n5085 ) | ( n4964 & n5085 ) ;
  assign n5088 = ( n4890 & ~n5086 ) | ( n4890 & n5087 ) | ( ~n5086 & n5087 ) ;
  assign n5089 = n583 & n2877 ;
  assign n5090 = x98 & n587 ;
  assign n5091 = x99 | n5090 ;
  assign n5092 = ( n589 & n5090 ) | ( n589 & n5091 ) | ( n5090 & n5091 ) ;
  assign n5093 = x97 & n676 ;
  assign n5094 = n5092 | n5093 ;
  assign n5095 = ( x14 & n5089 ) | ( x14 & ~n5094 ) | ( n5089 & ~n5094 ) ;
  assign n5096 = ( ~x14 & n5094 ) | ( ~x14 & n5095 ) | ( n5094 & n5095 ) ;
  assign n5097 = ( ~n5089 & n5095 ) | ( ~n5089 & n5096 ) | ( n5095 & n5096 ) ;
  assign n5098 = ( n4902 & n5088 ) | ( n4902 & n5097 ) | ( n5088 & n5097 ) ;
  assign n5099 = ( ~n4902 & n5088 ) | ( ~n4902 & n5097 ) | ( n5088 & n5097 ) ;
  assign n5100 = ( n4902 & ~n5098 ) | ( n4902 & n5099 ) | ( ~n5098 & n5099 ) ;
  assign n5101 = n407 & n3486 ;
  assign n5102 = x101 & n411 ;
  assign n5103 = x102 | n5102 ;
  assign n5104 = ( n413 & n5102 ) | ( n413 & n5103 ) | ( n5102 & n5103 ) ;
  assign n5105 = x100 & n491 ;
  assign n5106 = n5104 | n5105 ;
  assign n5107 = ( x11 & n5101 ) | ( x11 & ~n5106 ) | ( n5101 & ~n5106 ) ;
  assign n5108 = ( ~x11 & n5106 ) | ( ~x11 & n5107 ) | ( n5106 & n5107 ) ;
  assign n5109 = ( ~n5101 & n5107 ) | ( ~n5101 & n5108 ) | ( n5107 & n5108 ) ;
  assign n5110 = ( n4914 & n5100 ) | ( n4914 & n5109 ) | ( n5100 & n5109 ) ;
  assign n5111 = ( ~n4914 & n5100 ) | ( ~n4914 & n5109 ) | ( n5100 & n5109 ) ;
  assign n5112 = ( n4914 & ~n5110 ) | ( n4914 & n5111 ) | ( ~n5110 & n5111 ) ;
  assign n5113 = n291 & n3998 ;
  assign n5114 = x104 & n295 ;
  assign n5115 = x105 | n5114 ;
  assign n5116 = ( n297 & n5114 ) | ( n297 & n5115 ) | ( n5114 & n5115 ) ;
  assign n5117 = x103 & n330 ;
  assign n5118 = n5116 | n5117 ;
  assign n5119 = ( x8 & n5113 ) | ( x8 & ~n5118 ) | ( n5113 & ~n5118 ) ;
  assign n5120 = ( ~x8 & n5118 ) | ( ~x8 & n5119 ) | ( n5118 & n5119 ) ;
  assign n5121 = ( ~n5113 & n5119 ) | ( ~n5113 & n5120 ) | ( n5119 & n5120 ) ;
  assign n5122 = ( n4926 & n5112 ) | ( n4926 & n5121 ) | ( n5112 & n5121 ) ;
  assign n5123 = ( ~n4926 & n5112 ) | ( ~n4926 & n5121 ) | ( n5112 & n5121 ) ;
  assign n5124 = ( n4926 & ~n5122 ) | ( n4926 & n5123 ) | ( ~n5122 & n5123 ) ;
  assign n5125 = ( n4929 & n4955 ) | ( n4929 & n5124 ) | ( n4955 & n5124 ) ;
  assign n5126 = ( ~n4929 & n4955 ) | ( ~n4929 & n5124 ) | ( n4955 & n5124 ) ;
  assign n5127 = ( n4929 & ~n5125 ) | ( n4929 & n5126 ) | ( ~n5125 & n5126 ) ;
  assign n5128 = ( x110 & x111 ) | ( x110 & n4932 ) | ( x111 & n4932 ) ;
  assign n5129 = ( x110 & ~x111 ) | ( x110 & n4932 ) | ( ~x111 & n4932 ) ;
  assign n5130 = ( x111 & ~n5128 ) | ( x111 & n5129 ) | ( ~n5128 & n5129 ) ;
  assign n5131 = n136 & n5130 ;
  assign n5132 = x110 & n138 ;
  assign n5133 = x111 | n5132 ;
  assign n5134 = ( n141 & n5132 ) | ( n141 & n5133 ) | ( n5132 & n5133 ) ;
  assign n5135 = x109 & n154 ;
  assign n5136 = n5134 | n5135 ;
  assign n5137 = ( x2 & n5131 ) | ( x2 & ~n5136 ) | ( n5131 & ~n5136 ) ;
  assign n5138 = ( ~x2 & n5136 ) | ( ~x2 & n5137 ) | ( n5136 & n5137 ) ;
  assign n5139 = ( ~n5131 & n5137 ) | ( ~n5131 & n5138 ) | ( n5137 & n5138 ) ;
  assign n5140 = ( n4944 & n5127 ) | ( n4944 & n5139 ) | ( n5127 & n5139 ) ;
  assign n5141 = ( ~n4944 & n5127 ) | ( ~n4944 & n5139 ) | ( n5127 & n5139 ) ;
  assign n5142 = ( n4944 & ~n5140 ) | ( n4944 & n5141 ) | ( ~n5140 & n5141 ) ;
  assign n5143 = ( x111 & x112 ) | ( x111 & n5128 ) | ( x112 & n5128 ) ;
  assign n5144 = ( x111 & ~x112 ) | ( x111 & n5128 ) | ( ~x112 & n5128 ) ;
  assign n5145 = ( x112 & ~n5143 ) | ( x112 & n5144 ) | ( ~n5143 & n5144 ) ;
  assign n5146 = n136 & n5145 ;
  assign n5147 = x111 & n138 ;
  assign n5148 = x112 | n5147 ;
  assign n5149 = ( n141 & n5147 ) | ( n141 & n5148 ) | ( n5147 & n5148 ) ;
  assign n5150 = x110 & n154 ;
  assign n5151 = n5149 | n5150 ;
  assign n5152 = ( x2 & n5146 ) | ( x2 & ~n5151 ) | ( n5146 & ~n5151 ) ;
  assign n5153 = ( ~x2 & n5151 ) | ( ~x2 & n5152 ) | ( n5151 & n5152 ) ;
  assign n5154 = ( ~n5146 & n5152 ) | ( ~n5146 & n5153 ) | ( n5152 & n5153 ) ;
  assign n5155 = n186 & n4734 ;
  assign n5156 = x108 & n190 ;
  assign n5157 = x109 | n5156 ;
  assign n5158 = ( n192 & n5156 ) | ( n192 & n5157 ) | ( n5156 & n5157 ) ;
  assign n5159 = x107 & n220 ;
  assign n5160 = n5158 | n5159 ;
  assign n5161 = ( x5 & n5155 ) | ( x5 & ~n5160 ) | ( n5155 & ~n5160 ) ;
  assign n5162 = ( ~x5 & n5160 ) | ( ~x5 & n5161 ) | ( n5160 & n5161 ) ;
  assign n5163 = ( ~n5155 & n5161 ) | ( ~n5155 & n5162 ) | ( n5161 & n5162 ) ;
  assign n5164 = n583 & n3162 ;
  assign n5165 = x99 & n587 ;
  assign n5166 = x100 | n5165 ;
  assign n5167 = ( n589 & n5165 ) | ( n589 & n5166 ) | ( n5165 & n5166 ) ;
  assign n5168 = x98 & n676 ;
  assign n5169 = n5167 | n5168 ;
  assign n5170 = ( x14 & n5164 ) | ( x14 & ~n5169 ) | ( n5164 & ~n5169 ) ;
  assign n5171 = ( ~x14 & n5169 ) | ( ~x14 & n5170 ) | ( n5169 & n5170 ) ;
  assign n5172 = ( ~n5164 & n5170 ) | ( ~n5164 & n5171 ) | ( n5170 & n5171 ) ;
  assign n5173 = n1016 & n2294 ;
  assign n5174 = x93 & n1020 ;
  assign n5175 = x94 | n5174 ;
  assign n5176 = ( n1022 & n5174 ) | ( n1022 & n5175 ) | ( n5174 & n5175 ) ;
  assign n5177 = x92 & n1145 ;
  assign n5178 = n5176 | n5177 ;
  assign n5179 = ( x20 & n5173 ) | ( x20 & ~n5178 ) | ( n5173 & ~n5178 ) ;
  assign n5180 = ( ~x20 & n5178 ) | ( ~x20 & n5179 ) | ( n5178 & n5179 ) ;
  assign n5181 = ( ~n5173 & n5179 ) | ( ~n5173 & n5180 ) | ( n5179 & n5180 ) ;
  assign n5182 = n701 & n2766 ;
  assign n5183 = x78 & n2770 ;
  assign n5184 = x79 | n5183 ;
  assign n5185 = ( n2772 & n5183 ) | ( n2772 & n5184 ) | ( n5183 & n5184 ) ;
  assign n5186 = x77 & n2943 ;
  assign n5187 = n5185 | n5186 ;
  assign n5188 = ( x35 & n5182 ) | ( x35 & ~n5187 ) | ( n5182 & ~n5187 ) ;
  assign n5189 = ( ~x35 & n5187 ) | ( ~x35 & n5188 ) | ( n5187 & n5188 ) ;
  assign n5190 = ( ~n5182 & n5188 ) | ( ~n5182 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5191 = n554 & n3224 ;
  assign n5192 = x75 & n3228 ;
  assign n5193 = x76 | n5192 ;
  assign n5194 = ( n3230 & n5192 ) | ( n3230 & n5193 ) | ( n5192 & n5193 ) ;
  assign n5195 = x74 & n3413 ;
  assign n5196 = n5194 | n5195 ;
  assign n5197 = ( x38 & n5191 ) | ( x38 & ~n5196 ) | ( n5191 & ~n5196 ) ;
  assign n5198 = ( ~x38 & n5196 ) | ( ~x38 & n5197 ) | ( n5196 & n5197 ) ;
  assign n5199 = ( ~n5191 & n5197 ) | ( ~n5191 & n5198 ) | ( n5197 & n5198 ) ;
  assign n5200 = x66 & n4791 ;
  assign n5201 = x67 | n5200 ;
  assign n5202 = ( n4793 & n5200 ) | ( n4793 & n5201 ) | ( n5200 & n5201 ) ;
  assign n5203 = x65 & n5030 ;
  assign n5204 = n5202 | n5203 ;
  assign n5205 = n164 & n4787 ;
  assign n5206 = ( x47 & n5204 ) | ( x47 & ~n5205 ) | ( n5204 & ~n5205 ) ;
  assign n5207 = ( ~x47 & n5205 ) | ( ~x47 & n5206 ) | ( n5205 & n5206 ) ;
  assign n5208 = ( ~n5204 & n5206 ) | ( ~n5204 & n5207 ) | ( n5206 & n5207 ) ;
  assign n5209 = x47 & x48 ;
  assign n5210 = x47 | x48 ;
  assign n5211 = ~n5209 & n5210 ;
  assign n5212 = x64 & n5211 ;
  assign n5213 = x47 & ~n5038 ;
  assign n5214 = ( n5208 & n5212 ) | ( n5208 & n5213 ) | ( n5212 & n5213 ) ;
  assign n5215 = ( ~n5208 & n5212 ) | ( ~n5208 & n5213 ) | ( n5212 & n5213 ) ;
  assign n5216 = ( n5208 & ~n5214 ) | ( n5208 & n5215 ) | ( ~n5214 & n5215 ) ;
  assign n5217 = n245 & n4227 ;
  assign n5218 = x69 & n4231 ;
  assign n5219 = x70 | n5218 ;
  assign n5220 = ( n4233 & n5218 ) | ( n4233 & n5219 ) | ( n5218 & n5219 ) ;
  assign n5221 = x68 & n4470 ;
  assign n5222 = n5220 | n5221 ;
  assign n5223 = ( x44 & n5217 ) | ( x44 & ~n5222 ) | ( n5217 & ~n5222 ) ;
  assign n5224 = ( ~x44 & n5222 ) | ( ~x44 & n5223 ) | ( n5222 & n5223 ) ;
  assign n5225 = ( ~n5217 & n5223 ) | ( ~n5217 & n5224 ) | ( n5223 & n5224 ) ;
  assign n5226 = ( n5041 & n5216 ) | ( n5041 & n5225 ) | ( n5216 & n5225 ) ;
  assign n5227 = ( ~n5041 & n5216 ) | ( ~n5041 & n5225 ) | ( n5216 & n5225 ) ;
  assign n5228 = ( n5041 & ~n5226 ) | ( n5041 & n5227 ) | ( ~n5226 & n5227 ) ;
  assign n5229 = n390 & n3715 ;
  assign n5230 = x72 & n3719 ;
  assign n5231 = x73 | n5230 ;
  assign n5232 = ( n3721 & n5230 ) | ( n3721 & n5231 ) | ( n5230 & n5231 ) ;
  assign n5233 = x71 & n3922 ;
  assign n5234 = n5232 | n5233 ;
  assign n5235 = ( x41 & n5229 ) | ( x41 & ~n5234 ) | ( n5229 & ~n5234 ) ;
  assign n5236 = ( ~x41 & n5234 ) | ( ~x41 & n5235 ) | ( n5234 & n5235 ) ;
  assign n5237 = ( ~n5229 & n5235 ) | ( ~n5229 & n5236 ) | ( n5235 & n5236 ) ;
  assign n5238 = ( n5044 & n5228 ) | ( n5044 & n5237 ) | ( n5228 & n5237 ) ;
  assign n5239 = ( ~n5044 & n5228 ) | ( ~n5044 & n5237 ) | ( n5228 & n5237 ) ;
  assign n5240 = ( n5044 & ~n5238 ) | ( n5044 & n5239 ) | ( ~n5238 & n5239 ) ;
  assign n5241 = ( n5047 & n5199 ) | ( n5047 & n5240 ) | ( n5199 & n5240 ) ;
  assign n5242 = ( ~n5047 & n5199 ) | ( ~n5047 & n5240 ) | ( n5199 & n5240 ) ;
  assign n5243 = ( n5047 & ~n5241 ) | ( n5047 & n5242 ) | ( ~n5241 & n5242 ) ;
  assign n5244 = ( n5059 & n5190 ) | ( n5059 & n5243 ) | ( n5190 & n5243 ) ;
  assign n5245 = ( ~n5059 & n5190 ) | ( ~n5059 & n5243 ) | ( n5190 & n5243 ) ;
  assign n5246 = ( n5059 & ~n5244 ) | ( n5059 & n5245 ) | ( ~n5244 & n5245 ) ;
  assign n5247 = n990 & n2320 ;
  assign n5248 = x81 & n2324 ;
  assign n5249 = x82 | n5248 ;
  assign n5250 = ( n2326 & n5248 ) | ( n2326 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5251 = x80 & n2497 ;
  assign n5252 = n5250 | n5251 ;
  assign n5253 = ( x32 & n5247 ) | ( x32 & ~n5252 ) | ( n5247 & ~n5252 ) ;
  assign n5254 = ( ~x32 & n5252 ) | ( ~x32 & n5253 ) | ( n5252 & n5253 ) ;
  assign n5255 = ( ~n5247 & n5253 ) | ( ~n5247 & n5254 ) | ( n5253 & n5254 ) ;
  assign n5256 = ( n5062 & n5246 ) | ( n5062 & n5255 ) | ( n5246 & n5255 ) ;
  assign n5257 = ( ~n5062 & n5246 ) | ( ~n5062 & n5255 ) | ( n5246 & n5255 ) ;
  assign n5258 = ( n5062 & ~n5256 ) | ( n5062 & n5257 ) | ( ~n5256 & n5257 ) ;
  assign n5259 = n1262 & n1949 ;
  assign n5260 = x84 & n1953 ;
  assign n5261 = x85 | n5260 ;
  assign n5262 = ( n1955 & n5260 ) | ( n1955 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5263 = x83 & n2114 ;
  assign n5264 = n5262 | n5263 ;
  assign n5265 = ( x29 & n5259 ) | ( x29 & ~n5264 ) | ( n5259 & ~n5264 ) ;
  assign n5266 = ( ~x29 & n5264 ) | ( ~x29 & n5265 ) | ( n5264 & n5265 ) ;
  assign n5267 = ( ~n5259 & n5265 ) | ( ~n5259 & n5266 ) | ( n5265 & n5266 ) ;
  assign n5268 = ( n5065 & n5258 ) | ( n5065 & n5267 ) | ( n5258 & n5267 ) ;
  assign n5269 = ( ~n5065 & n5258 ) | ( ~n5065 & n5267 ) | ( n5258 & n5267 ) ;
  assign n5270 = ( n5065 & ~n5268 ) | ( n5065 & n5269 ) | ( ~n5268 & n5269 ) ;
  assign n5271 = n1481 & n1617 ;
  assign n5272 = x87 & n1621 ;
  assign n5273 = x88 | n5272 ;
  assign n5274 = ( n1623 & n5272 ) | ( n1623 & n5273 ) | ( n5272 & n5273 ) ;
  assign n5275 = x86 & n1749 ;
  assign n5276 = n5274 | n5275 ;
  assign n5277 = ( x26 & n5271 ) | ( x26 & ~n5276 ) | ( n5271 & ~n5276 ) ;
  assign n5278 = ( ~x26 & n5276 ) | ( ~x26 & n5277 ) | ( n5276 & n5277 ) ;
  assign n5279 = ( ~n5271 & n5277 ) | ( ~n5271 & n5278 ) | ( n5277 & n5278 ) ;
  assign n5280 = ( n5077 & n5270 ) | ( n5077 & n5279 ) | ( n5270 & n5279 ) ;
  assign n5281 = ( ~n5077 & n5270 ) | ( ~n5077 & n5279 ) | ( n5270 & n5279 ) ;
  assign n5282 = ( n5077 & ~n5280 ) | ( n5077 & n5281 ) | ( ~n5280 & n5281 ) ;
  assign n5283 = n1297 & n1914 ;
  assign n5284 = x90 & n1301 ;
  assign n5285 = x91 | n5284 ;
  assign n5286 = ( n1303 & n5284 ) | ( n1303 & n5285 ) | ( n5284 & n5285 ) ;
  assign n5287 = x89 & n1426 ;
  assign n5288 = n5286 | n5287 ;
  assign n5289 = ( x23 & n5283 ) | ( x23 & ~n5288 ) | ( n5283 & ~n5288 ) ;
  assign n5290 = ( ~x23 & n5288 ) | ( ~x23 & n5289 ) | ( n5288 & n5289 ) ;
  assign n5291 = ( ~n5283 & n5289 ) | ( ~n5283 & n5290 ) | ( n5289 & n5290 ) ;
  assign n5292 = ( n5080 & n5282 ) | ( n5080 & n5291 ) | ( n5282 & n5291 ) ;
  assign n5293 = ( ~n5080 & n5282 ) | ( ~n5080 & n5291 ) | ( n5282 & n5291 ) ;
  assign n5294 = ( n5080 & ~n5292 ) | ( n5080 & n5293 ) | ( ~n5292 & n5293 ) ;
  assign n5295 = ( n5083 & n5181 ) | ( n5083 & n5294 ) | ( n5181 & n5294 ) ;
  assign n5296 = ( ~n5083 & n5181 ) | ( ~n5083 & n5294 ) | ( n5181 & n5294 ) ;
  assign n5297 = ( n5083 & ~n5295 ) | ( n5083 & n5296 ) | ( ~n5295 & n5296 ) ;
  assign n5298 = n810 & n2585 ;
  assign n5299 = x96 & n814 ;
  assign n5300 = x97 | n5299 ;
  assign n5301 = ( n816 & n5299 ) | ( n816 & n5300 ) | ( n5299 & n5300 ) ;
  assign n5302 = x95 & n885 ;
  assign n5303 = n5301 | n5302 ;
  assign n5304 = ( x17 & n5298 ) | ( x17 & ~n5303 ) | ( n5298 & ~n5303 ) ;
  assign n5305 = ( ~x17 & n5303 ) | ( ~x17 & n5304 ) | ( n5303 & n5304 ) ;
  assign n5306 = ( ~n5298 & n5304 ) | ( ~n5298 & n5305 ) | ( n5304 & n5305 ) ;
  assign n5307 = ( n5086 & n5297 ) | ( n5086 & n5306 ) | ( n5297 & n5306 ) ;
  assign n5308 = ( ~n5086 & n5297 ) | ( ~n5086 & n5306 ) | ( n5297 & n5306 ) ;
  assign n5309 = ( n5086 & ~n5307 ) | ( n5086 & n5308 ) | ( ~n5307 & n5308 ) ;
  assign n5310 = ( n5098 & n5172 ) | ( n5098 & n5309 ) | ( n5172 & n5309 ) ;
  assign n5311 = ( ~n5098 & n5172 ) | ( ~n5098 & n5309 ) | ( n5172 & n5309 ) ;
  assign n5312 = ( n5098 & ~n5310 ) | ( n5098 & n5311 ) | ( ~n5310 & n5311 ) ;
  assign n5313 = n407 & n3650 ;
  assign n5314 = x102 & n411 ;
  assign n5315 = x103 | n5314 ;
  assign n5316 = ( n413 & n5314 ) | ( n413 & n5315 ) | ( n5314 & n5315 ) ;
  assign n5317 = x101 & n491 ;
  assign n5318 = n5316 | n5317 ;
  assign n5319 = ( x11 & n5313 ) | ( x11 & ~n5318 ) | ( n5313 & ~n5318 ) ;
  assign n5320 = ( ~x11 & n5318 ) | ( ~x11 & n5319 ) | ( n5318 & n5319 ) ;
  assign n5321 = ( ~n5313 & n5319 ) | ( ~n5313 & n5320 ) | ( n5319 & n5320 ) ;
  assign n5322 = ( n5110 & n5312 ) | ( n5110 & n5321 ) | ( n5312 & n5321 ) ;
  assign n5323 = ( ~n5110 & n5312 ) | ( ~n5110 & n5321 ) | ( n5312 & n5321 ) ;
  assign n5324 = ( n5110 & ~n5322 ) | ( n5110 & n5323 ) | ( ~n5322 & n5323 ) ;
  assign n5325 = n291 & n4013 ;
  assign n5326 = x105 & n295 ;
  assign n5327 = x106 | n5326 ;
  assign n5328 = ( n297 & n5326 ) | ( n297 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5329 = x104 & n330 ;
  assign n5330 = n5328 | n5329 ;
  assign n5331 = ( x8 & n5325 ) | ( x8 & ~n5330 ) | ( n5325 & ~n5330 ) ;
  assign n5332 = ( ~x8 & n5330 ) | ( ~x8 & n5331 ) | ( n5330 & n5331 ) ;
  assign n5333 = ( ~n5325 & n5331 ) | ( ~n5325 & n5332 ) | ( n5331 & n5332 ) ;
  assign n5334 = ( n5122 & n5324 ) | ( n5122 & n5333 ) | ( n5324 & n5333 ) ;
  assign n5335 = ( ~n5122 & n5324 ) | ( ~n5122 & n5333 ) | ( n5324 & n5333 ) ;
  assign n5336 = ( n5122 & ~n5334 ) | ( n5122 & n5335 ) | ( ~n5334 & n5335 ) ;
  assign n5337 = ( n5125 & n5163 ) | ( n5125 & n5336 ) | ( n5163 & n5336 ) ;
  assign n5338 = ( ~n5125 & n5163 ) | ( ~n5125 & n5336 ) | ( n5163 & n5336 ) ;
  assign n5339 = ( n5125 & ~n5337 ) | ( n5125 & n5338 ) | ( ~n5337 & n5338 ) ;
  assign n5340 = ( n5140 & n5154 ) | ( n5140 & n5339 ) | ( n5154 & n5339 ) ;
  assign n5341 = ( ~n5140 & n5154 ) | ( ~n5140 & n5339 ) | ( n5154 & n5339 ) ;
  assign n5342 = ( n5140 & ~n5340 ) | ( n5140 & n5341 ) | ( ~n5340 & n5341 ) ;
  assign n5343 = n1016 & n2434 ;
  assign n5344 = x94 & n1020 ;
  assign n5345 = x95 | n5344 ;
  assign n5346 = ( n1022 & n5344 ) | ( n1022 & n5345 ) | ( n5344 & n5345 ) ;
  assign n5347 = x93 & n1145 ;
  assign n5348 = n5346 | n5347 ;
  assign n5349 = ( x20 & n5343 ) | ( x20 & ~n5348 ) | ( n5343 & ~n5348 ) ;
  assign n5350 = ( ~x20 & n5348 ) | ( ~x20 & n5349 ) | ( n5348 & n5349 ) ;
  assign n5351 = ( ~n5343 & n5349 ) | ( ~n5343 & n5350 ) | ( n5349 & n5350 ) ;
  assign n5352 = n1297 & n2042 ;
  assign n5353 = x91 & n1301 ;
  assign n5354 = x92 | n5353 ;
  assign n5355 = ( n1303 & n5353 ) | ( n1303 & n5354 ) | ( n5353 & n5354 ) ;
  assign n5356 = x90 & n1426 ;
  assign n5357 = n5355 | n5356 ;
  assign n5358 = ( x23 & n5352 ) | ( x23 & ~n5357 ) | ( n5352 & ~n5357 ) ;
  assign n5359 = ( ~x23 & n5357 ) | ( ~x23 & n5358 ) | ( n5357 & n5358 ) ;
  assign n5360 = ( ~n5352 & n5358 ) | ( ~n5352 & n5359 ) | ( n5358 & n5359 ) ;
  assign n5361 = n569 & n3224 ;
  assign n5362 = x76 & n3228 ;
  assign n5363 = x77 | n5362 ;
  assign n5364 = ( n3230 & n5362 ) | ( n3230 & n5363 ) | ( n5362 & n5363 ) ;
  assign n5365 = x75 & n3413 ;
  assign n5366 = n5364 | n5365 ;
  assign n5367 = ( x38 & n5361 ) | ( x38 & ~n5366 ) | ( n5361 & ~n5366 ) ;
  assign n5368 = ( ~x38 & n5366 ) | ( ~x38 & n5367 ) | ( n5366 & n5367 ) ;
  assign n5369 = ( ~n5361 & n5367 ) | ( ~n5361 & n5368 ) | ( n5367 & n5368 ) ;
  assign n5370 = x50 & n5212 ;
  assign n5371 = x49 | x50 ;
  assign n5372 = ( x49 & x50 ) | ( x49 & ~n5371 ) | ( x50 & ~n5371 ) ;
  assign n5373 = n5371 & ~n5372 ;
  assign n5374 = n5211 & n5373 ;
  assign n5375 = n133 & n5374 ;
  assign n5376 = ~x47 & x49 ;
  assign n5377 = x48 & x49 ;
  assign n5378 = ( n5209 & n5376 ) | ( n5209 & ~n5377 ) | ( n5376 & ~n5377 ) ;
  assign n5379 = x64 & n5378 ;
  assign n5380 = ( n5211 & ~n5371 ) | ( n5211 & n5372 ) | ( ~n5371 & n5372 ) ;
  assign n5381 = x65 | n5379 ;
  assign n5382 = ( n5379 & n5380 ) | ( n5379 & n5381 ) | ( n5380 & n5381 ) ;
  assign n5383 = ( n5370 & n5375 ) | ( n5370 & n5382 ) | ( n5375 & n5382 ) ;
  assign n5384 = n5375 | n5382 ;
  assign n5385 = ~n5370 & n5384 ;
  assign n5386 = ( n5370 & ~n5383 ) | ( n5370 & n5385 ) | ( ~n5383 & n5385 ) ;
  assign n5387 = x67 & n4791 ;
  assign n5388 = x68 | n5387 ;
  assign n5389 = ( n4793 & n5387 ) | ( n4793 & n5388 ) | ( n5387 & n5388 ) ;
  assign n5390 = x66 & n5030 ;
  assign n5391 = n5389 | n5390 ;
  assign n5392 = n201 & n4787 ;
  assign n5393 = ( x47 & n5391 ) | ( x47 & ~n5392 ) | ( n5391 & ~n5392 ) ;
  assign n5394 = ( ~x47 & n5392 ) | ( ~x47 & n5393 ) | ( n5392 & n5393 ) ;
  assign n5395 = ( ~n5391 & n5393 ) | ( ~n5391 & n5394 ) | ( n5393 & n5394 ) ;
  assign n5396 = ( n5214 & n5386 ) | ( n5214 & n5395 ) | ( n5386 & n5395 ) ;
  assign n5397 = ( ~n5214 & n5386 ) | ( ~n5214 & n5395 ) | ( n5386 & n5395 ) ;
  assign n5398 = ( n5214 & ~n5396 ) | ( n5214 & n5397 ) | ( ~n5396 & n5397 ) ;
  assign n5399 = n277 & n4227 ;
  assign n5400 = x70 & n4231 ;
  assign n5401 = x71 | n5400 ;
  assign n5402 = ( n4233 & n5400 ) | ( n4233 & n5401 ) | ( n5400 & n5401 ) ;
  assign n5403 = x69 & n4470 ;
  assign n5404 = n5402 | n5403 ;
  assign n5405 = ( x44 & n5399 ) | ( x44 & ~n5404 ) | ( n5399 & ~n5404 ) ;
  assign n5406 = ( ~x44 & n5404 ) | ( ~x44 & n5405 ) | ( n5404 & n5405 ) ;
  assign n5407 = ( ~n5399 & n5405 ) | ( ~n5399 & n5406 ) | ( n5405 & n5406 ) ;
  assign n5408 = ( n5226 & n5398 ) | ( n5226 & n5407 ) | ( n5398 & n5407 ) ;
  assign n5409 = ( ~n5226 & n5398 ) | ( ~n5226 & n5407 ) | ( n5398 & n5407 ) ;
  assign n5410 = ( n5226 & ~n5408 ) | ( n5226 & n5409 ) | ( ~n5408 & n5409 ) ;
  assign n5411 = n446 & n3715 ;
  assign n5412 = x73 & n3719 ;
  assign n5413 = x74 | n5412 ;
  assign n5414 = ( n3721 & n5412 ) | ( n3721 & n5413 ) | ( n5412 & n5413 ) ;
  assign n5415 = x72 & n3922 ;
  assign n5416 = n5414 | n5415 ;
  assign n5417 = ( x41 & n5411 ) | ( x41 & ~n5416 ) | ( n5411 & ~n5416 ) ;
  assign n5418 = ( ~x41 & n5416 ) | ( ~x41 & n5417 ) | ( n5416 & n5417 ) ;
  assign n5419 = ( ~n5411 & n5417 ) | ( ~n5411 & n5418 ) | ( n5417 & n5418 ) ;
  assign n5420 = ( n5238 & n5410 ) | ( n5238 & n5419 ) | ( n5410 & n5419 ) ;
  assign n5421 = ( ~n5238 & n5410 ) | ( ~n5238 & n5419 ) | ( n5410 & n5419 ) ;
  assign n5422 = ( n5238 & ~n5420 ) | ( n5238 & n5421 ) | ( ~n5420 & n5421 ) ;
  assign n5423 = ( n5241 & n5369 ) | ( n5241 & n5422 ) | ( n5369 & n5422 ) ;
  assign n5424 = ( ~n5241 & n5369 ) | ( ~n5241 & n5422 ) | ( n5369 & n5422 ) ;
  assign n5425 = ( n5241 & ~n5423 ) | ( n5241 & n5424 ) | ( ~n5423 & n5424 ) ;
  assign n5426 = n769 & n2766 ;
  assign n5427 = x79 & n2770 ;
  assign n5428 = x80 | n5427 ;
  assign n5429 = ( n2772 & n5427 ) | ( n2772 & n5428 ) | ( n5427 & n5428 ) ;
  assign n5430 = x78 & n2943 ;
  assign n5431 = n5429 | n5430 ;
  assign n5432 = ( x35 & n5426 ) | ( x35 & ~n5431 ) | ( n5426 & ~n5431 ) ;
  assign n5433 = ( ~x35 & n5431 ) | ( ~x35 & n5432 ) | ( n5431 & n5432 ) ;
  assign n5434 = ( ~n5426 & n5432 ) | ( ~n5426 & n5433 ) | ( n5432 & n5433 ) ;
  assign n5435 = ( n5244 & n5425 ) | ( n5244 & n5434 ) | ( n5425 & n5434 ) ;
  assign n5436 = ( ~n5244 & n5425 ) | ( ~n5244 & n5434 ) | ( n5425 & n5434 ) ;
  assign n5437 = ( n5244 & ~n5435 ) | ( n5244 & n5436 ) | ( ~n5435 & n5436 ) ;
  assign n5438 = n1082 & n2320 ;
  assign n5439 = x82 & n2324 ;
  assign n5440 = x83 | n5439 ;
  assign n5441 = ( n2326 & n5439 ) | ( n2326 & n5440 ) | ( n5439 & n5440 ) ;
  assign n5442 = x81 & n2497 ;
  assign n5443 = n5441 | n5442 ;
  assign n5444 = ( x32 & n5438 ) | ( x32 & ~n5443 ) | ( n5438 & ~n5443 ) ;
  assign n5445 = ( ~x32 & n5443 ) | ( ~x32 & n5444 ) | ( n5443 & n5444 ) ;
  assign n5446 = ( ~n5438 & n5444 ) | ( ~n5438 & n5445 ) | ( n5444 & n5445 ) ;
  assign n5447 = ( n5256 & n5437 ) | ( n5256 & n5446 ) | ( n5437 & n5446 ) ;
  assign n5448 = ( ~n5256 & n5437 ) | ( ~n5256 & n5446 ) | ( n5437 & n5446 ) ;
  assign n5449 = ( n5256 & ~n5447 ) | ( n5256 & n5448 ) | ( ~n5447 & n5448 ) ;
  assign n5450 = n1366 & n1949 ;
  assign n5451 = x85 & n1953 ;
  assign n5452 = x86 | n5451 ;
  assign n5453 = ( n1955 & n5451 ) | ( n1955 & n5452 ) | ( n5451 & n5452 ) ;
  assign n5454 = x84 & n2114 ;
  assign n5455 = n5453 | n5454 ;
  assign n5456 = ( x29 & n5450 ) | ( x29 & ~n5455 ) | ( n5450 & ~n5455 ) ;
  assign n5457 = ( ~x29 & n5455 ) | ( ~x29 & n5456 ) | ( n5455 & n5456 ) ;
  assign n5458 = ( ~n5450 & n5456 ) | ( ~n5450 & n5457 ) | ( n5456 & n5457 ) ;
  assign n5459 = ( n5268 & n5449 ) | ( n5268 & n5458 ) | ( n5449 & n5458 ) ;
  assign n5460 = ( ~n5268 & n5449 ) | ( ~n5268 & n5458 ) | ( n5449 & n5458 ) ;
  assign n5461 = ( n5268 & ~n5459 ) | ( n5268 & n5460 ) | ( ~n5459 & n5460 ) ;
  assign n5462 = n1585 & n1617 ;
  assign n5463 = x88 & n1621 ;
  assign n5464 = x89 | n5463 ;
  assign n5465 = ( n1623 & n5463 ) | ( n1623 & n5464 ) | ( n5463 & n5464 ) ;
  assign n5466 = x87 & n1749 ;
  assign n5467 = n5465 | n5466 ;
  assign n5468 = ( x26 & n5462 ) | ( x26 & ~n5467 ) | ( n5462 & ~n5467 ) ;
  assign n5469 = ( ~x26 & n5467 ) | ( ~x26 & n5468 ) | ( n5467 & n5468 ) ;
  assign n5470 = ( ~n5462 & n5468 ) | ( ~n5462 & n5469 ) | ( n5468 & n5469 ) ;
  assign n5471 = ( n5280 & n5461 ) | ( n5280 & n5470 ) | ( n5461 & n5470 ) ;
  assign n5472 = ( ~n5280 & n5461 ) | ( ~n5280 & n5470 ) | ( n5461 & n5470 ) ;
  assign n5473 = ( n5280 & ~n5471 ) | ( n5280 & n5472 ) | ( ~n5471 & n5472 ) ;
  assign n5474 = ( n5292 & n5360 ) | ( n5292 & n5473 ) | ( n5360 & n5473 ) ;
  assign n5475 = ( ~n5292 & n5360 ) | ( ~n5292 & n5473 ) | ( n5360 & n5473 ) ;
  assign n5476 = ( n5292 & ~n5474 ) | ( n5292 & n5475 ) | ( ~n5474 & n5475 ) ;
  assign n5477 = ( n5295 & n5351 ) | ( n5295 & n5476 ) | ( n5351 & n5476 ) ;
  assign n5478 = ( ~n5295 & n5351 ) | ( ~n5295 & n5476 ) | ( n5351 & n5476 ) ;
  assign n5479 = ( n5295 & ~n5477 ) | ( n5295 & n5478 ) | ( ~n5477 & n5478 ) ;
  assign n5480 = n810 & n2725 ;
  assign n5481 = x97 & n814 ;
  assign n5482 = x98 | n5481 ;
  assign n5483 = ( n816 & n5481 ) | ( n816 & n5482 ) | ( n5481 & n5482 ) ;
  assign n5484 = x96 & n885 ;
  assign n5485 = n5483 | n5484 ;
  assign n5486 = ( x17 & n5480 ) | ( x17 & ~n5485 ) | ( n5480 & ~n5485 ) ;
  assign n5487 = ( ~x17 & n5485 ) | ( ~x17 & n5486 ) | ( n5485 & n5486 ) ;
  assign n5488 = ( ~n5480 & n5486 ) | ( ~n5480 & n5487 ) | ( n5486 & n5487 ) ;
  assign n5489 = ( n5307 & n5479 ) | ( n5307 & n5488 ) | ( n5479 & n5488 ) ;
  assign n5490 = ( ~n5307 & n5479 ) | ( ~n5307 & n5488 ) | ( n5479 & n5488 ) ;
  assign n5491 = ( n5307 & ~n5489 ) | ( n5307 & n5490 ) | ( ~n5489 & n5490 ) ;
  assign n5492 = n583 & n3326 ;
  assign n5493 = x100 & n587 ;
  assign n5494 = x101 | n5493 ;
  assign n5495 = ( n589 & n5493 ) | ( n589 & n5494 ) | ( n5493 & n5494 ) ;
  assign n5496 = x99 & n676 ;
  assign n5497 = n5495 | n5496 ;
  assign n5498 = ( x14 & n5492 ) | ( x14 & ~n5497 ) | ( n5492 & ~n5497 ) ;
  assign n5499 = ( ~x14 & n5497 ) | ( ~x14 & n5498 ) | ( n5497 & n5498 ) ;
  assign n5500 = ( ~n5492 & n5498 ) | ( ~n5492 & n5499 ) | ( n5498 & n5499 ) ;
  assign n5501 = ( n5310 & n5491 ) | ( n5310 & n5500 ) | ( n5491 & n5500 ) ;
  assign n5502 = ( ~n5310 & n5491 ) | ( ~n5310 & n5500 ) | ( n5491 & n5500 ) ;
  assign n5503 = ( n5310 & ~n5501 ) | ( n5310 & n5502 ) | ( ~n5501 & n5502 ) ;
  assign n5504 = n407 & n3665 ;
  assign n5505 = x103 & n411 ;
  assign n5506 = x104 | n5505 ;
  assign n5507 = ( n413 & n5505 ) | ( n413 & n5506 ) | ( n5505 & n5506 ) ;
  assign n5508 = x102 & n491 ;
  assign n5509 = n5507 | n5508 ;
  assign n5510 = ( x11 & n5504 ) | ( x11 & ~n5509 ) | ( n5504 & ~n5509 ) ;
  assign n5511 = ( ~x11 & n5509 ) | ( ~x11 & n5510 ) | ( n5509 & n5510 ) ;
  assign n5512 = ( ~n5504 & n5510 ) | ( ~n5504 & n5511 ) | ( n5510 & n5511 ) ;
  assign n5513 = ( n5322 & n5503 ) | ( n5322 & n5512 ) | ( n5503 & n5512 ) ;
  assign n5514 = ( ~n5322 & n5503 ) | ( ~n5322 & n5512 ) | ( n5503 & n5512 ) ;
  assign n5515 = ( n5322 & ~n5513 ) | ( n5322 & n5514 ) | ( ~n5513 & n5514 ) ;
  assign n5516 = n291 & n4362 ;
  assign n5517 = x106 & n295 ;
  assign n5518 = x107 | n5517 ;
  assign n5519 = ( n297 & n5517 ) | ( n297 & n5518 ) | ( n5517 & n5518 ) ;
  assign n5520 = x105 & n330 ;
  assign n5521 = n5519 | n5520 ;
  assign n5522 = ( x8 & n5516 ) | ( x8 & ~n5521 ) | ( n5516 & ~n5521 ) ;
  assign n5523 = ( ~x8 & n5521 ) | ( ~x8 & n5522 ) | ( n5521 & n5522 ) ;
  assign n5524 = ( ~n5516 & n5522 ) | ( ~n5516 & n5523 ) | ( n5522 & n5523 ) ;
  assign n5525 = ( n5334 & n5515 ) | ( n5334 & n5524 ) | ( n5515 & n5524 ) ;
  assign n5526 = ( ~n5334 & n5515 ) | ( ~n5334 & n5524 ) | ( n5515 & n5524 ) ;
  assign n5527 = ( n5334 & ~n5525 ) | ( n5334 & n5526 ) | ( ~n5525 & n5526 ) ;
  assign n5528 = n186 & n4934 ;
  assign n5529 = x109 & n190 ;
  assign n5530 = x110 | n5529 ;
  assign n5531 = ( n192 & n5529 ) | ( n192 & n5530 ) | ( n5529 & n5530 ) ;
  assign n5532 = x108 & n220 ;
  assign n5533 = n5531 | n5532 ;
  assign n5534 = ( x5 & n5528 ) | ( x5 & ~n5533 ) | ( n5528 & ~n5533 ) ;
  assign n5535 = ( ~x5 & n5533 ) | ( ~x5 & n5534 ) | ( n5533 & n5534 ) ;
  assign n5536 = ( ~n5528 & n5534 ) | ( ~n5528 & n5535 ) | ( n5534 & n5535 ) ;
  assign n5537 = ( n5337 & n5527 ) | ( n5337 & n5536 ) | ( n5527 & n5536 ) ;
  assign n5538 = ( ~n5337 & n5527 ) | ( ~n5337 & n5536 ) | ( n5527 & n5536 ) ;
  assign n5539 = ( n5337 & ~n5537 ) | ( n5337 & n5538 ) | ( ~n5537 & n5538 ) ;
  assign n5540 = ( x112 & x113 ) | ( x112 & n5143 ) | ( x113 & n5143 ) ;
  assign n5541 = ( x112 & ~x113 ) | ( x112 & n5143 ) | ( ~x113 & n5143 ) ;
  assign n5542 = ( x113 & ~n5540 ) | ( x113 & n5541 ) | ( ~n5540 & n5541 ) ;
  assign n5543 = n136 & n5542 ;
  assign n5544 = x112 & n138 ;
  assign n5545 = x113 | n5544 ;
  assign n5546 = ( n141 & n5544 ) | ( n141 & n5545 ) | ( n5544 & n5545 ) ;
  assign n5547 = x111 & n154 ;
  assign n5548 = n5546 | n5547 ;
  assign n5549 = ( x2 & n5543 ) | ( x2 & ~n5548 ) | ( n5543 & ~n5548 ) ;
  assign n5550 = ( ~x2 & n5548 ) | ( ~x2 & n5549 ) | ( n5548 & n5549 ) ;
  assign n5551 = ( ~n5543 & n5549 ) | ( ~n5543 & n5550 ) | ( n5549 & n5550 ) ;
  assign n5552 = ( n5340 & n5539 ) | ( n5340 & n5551 ) | ( n5539 & n5551 ) ;
  assign n5553 = ( ~n5340 & n5539 ) | ( ~n5340 & n5551 ) | ( n5539 & n5551 ) ;
  assign n5554 = ( n5340 & ~n5552 ) | ( n5340 & n5553 ) | ( ~n5552 & n5553 ) ;
  assign n5555 = n186 & n5130 ;
  assign n5556 = x110 & n190 ;
  assign n5557 = x111 | n5556 ;
  assign n5558 = ( n192 & n5556 ) | ( n192 & n5557 ) | ( n5556 & n5557 ) ;
  assign n5559 = x109 & n220 ;
  assign n5560 = n5558 | n5559 ;
  assign n5561 = ( x5 & n5555 ) | ( x5 & ~n5560 ) | ( n5555 & ~n5560 ) ;
  assign n5562 = ( ~x5 & n5560 ) | ( ~x5 & n5561 ) | ( n5560 & n5561 ) ;
  assign n5563 = ( ~n5555 & n5561 ) | ( ~n5555 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5564 = n1016 & n2449 ;
  assign n5565 = x95 & n1020 ;
  assign n5566 = x96 | n5565 ;
  assign n5567 = ( n1022 & n5565 ) | ( n1022 & n5566 ) | ( n5565 & n5566 ) ;
  assign n5568 = x94 & n1145 ;
  assign n5569 = n5567 | n5568 ;
  assign n5570 = ( x20 & n5564 ) | ( x20 & ~n5569 ) | ( n5564 & ~n5569 ) ;
  assign n5571 = ( ~x20 & n5569 ) | ( ~x20 & n5570 ) | ( n5569 & n5570 ) ;
  assign n5572 = ( ~n5564 & n5570 ) | ( ~n5564 & n5571 ) | ( n5570 & n5571 ) ;
  assign n5573 = n1297 & n2057 ;
  assign n5574 = x92 & n1301 ;
  assign n5575 = x93 | n5574 ;
  assign n5576 = ( n1303 & n5574 ) | ( n1303 & n5575 ) | ( n5574 & n5575 ) ;
  assign n5577 = x91 & n1426 ;
  assign n5578 = n5576 | n5577 ;
  assign n5579 = ( x23 & n5573 ) | ( x23 & ~n5578 ) | ( n5573 & ~n5578 ) ;
  assign n5580 = ( ~x23 & n5578 ) | ( ~x23 & n5579 ) | ( n5578 & n5579 ) ;
  assign n5581 = ( ~n5573 & n5579 ) | ( ~n5573 & n5580 ) | ( n5579 & n5580 ) ;
  assign n5582 = n1617 & n1701 ;
  assign n5583 = x89 & n1621 ;
  assign n5584 = x90 | n5583 ;
  assign n5585 = ( n1623 & n5583 ) | ( n1623 & n5584 ) | ( n5583 & n5584 ) ;
  assign n5586 = x88 & n1749 ;
  assign n5587 = n5585 | n5586 ;
  assign n5588 = ( x26 & n5582 ) | ( x26 & ~n5587 ) | ( n5582 & ~n5587 ) ;
  assign n5589 = ( ~x26 & n5587 ) | ( ~x26 & n5588 ) | ( n5587 & n5588 ) ;
  assign n5590 = ( ~n5582 & n5588 ) | ( ~n5582 & n5589 ) | ( n5588 & n5589 ) ;
  assign n5591 = n1097 & n2320 ;
  assign n5592 = x83 & n2324 ;
  assign n5593 = x84 | n5592 ;
  assign n5594 = ( n2326 & n5592 ) | ( n2326 & n5593 ) | ( n5592 & n5593 ) ;
  assign n5595 = x82 & n2497 ;
  assign n5596 = n5594 | n5595 ;
  assign n5597 = ( x32 & n5591 ) | ( x32 & ~n5596 ) | ( n5591 & ~n5596 ) ;
  assign n5598 = ( ~x32 & n5596 ) | ( ~x32 & n5597 ) | ( n5596 & n5597 ) ;
  assign n5599 = ( ~n5591 & n5597 ) | ( ~n5591 & n5598 ) | ( n5597 & n5598 ) ;
  assign n5600 = n910 & n2766 ;
  assign n5601 = x80 & n2770 ;
  assign n5602 = x81 | n5601 ;
  assign n5603 = ( n2772 & n5601 ) | ( n2772 & n5602 ) | ( n5601 & n5602 ) ;
  assign n5604 = x79 & n2943 ;
  assign n5605 = n5603 | n5604 ;
  assign n5606 = ( x35 & n5600 ) | ( x35 & ~n5605 ) | ( n5600 & ~n5605 ) ;
  assign n5607 = ( ~x35 & n5605 ) | ( ~x35 & n5606 ) | ( n5605 & n5606 ) ;
  assign n5608 = ( ~n5600 & n5606 ) | ( ~n5600 & n5607 ) | ( n5606 & n5607 ) ;
  assign n5609 = n461 & n3715 ;
  assign n5610 = x74 & n3719 ;
  assign n5611 = x75 | n5610 ;
  assign n5612 = ( n3721 & n5610 ) | ( n3721 & n5611 ) | ( n5610 & n5611 ) ;
  assign n5613 = x73 & n3922 ;
  assign n5614 = n5612 | n5613 ;
  assign n5615 = ( x41 & n5609 ) | ( x41 & ~n5614 ) | ( n5609 & ~n5614 ) ;
  assign n5616 = ( ~x41 & n5614 ) | ( ~x41 & n5615 ) | ( n5614 & n5615 ) ;
  assign n5617 = ( ~n5609 & n5615 ) | ( ~n5609 & n5616 ) | ( n5615 & n5616 ) ;
  assign n5618 = n346 & n4227 ;
  assign n5619 = x71 & n4231 ;
  assign n5620 = x72 | n5619 ;
  assign n5621 = ( n4233 & n5619 ) | ( n4233 & n5620 ) | ( n5619 & n5620 ) ;
  assign n5622 = x70 & n4470 ;
  assign n5623 = n5621 | n5622 ;
  assign n5624 = ( x44 & n5618 ) | ( x44 & ~n5623 ) | ( n5618 & ~n5623 ) ;
  assign n5625 = ( ~x44 & n5623 ) | ( ~x44 & n5624 ) | ( n5623 & n5624 ) ;
  assign n5626 = ( ~n5618 & n5624 ) | ( ~n5618 & n5625 ) | ( n5624 & n5625 ) ;
  assign n5627 = n230 & n4787 ;
  assign n5628 = x68 & n4791 ;
  assign n5629 = x69 | n5628 ;
  assign n5630 = ( n4793 & n5628 ) | ( n4793 & n5629 ) | ( n5628 & n5629 ) ;
  assign n5631 = x67 & n5030 ;
  assign n5632 = n5630 | n5631 ;
  assign n5633 = ( ~x47 & n5627 ) | ( ~x47 & n5632 ) | ( n5627 & n5632 ) ;
  assign n5634 = ( n5627 & n5632 ) | ( n5627 & ~n5633 ) | ( n5632 & ~n5633 ) ;
  assign n5635 = ( x47 & n5633 ) | ( x47 & ~n5634 ) | ( n5633 & ~n5634 ) ;
  assign n5636 = ( x50 & n5370 ) | ( x50 & n5384 ) | ( n5370 & n5384 ) ;
  assign n5637 = ( x47 & ~x49 ) | ( x47 & n5373 ) | ( ~x49 & n5373 ) ;
  assign n5638 = ( ~n5210 & n5377 ) | ( ~n5210 & n5637 ) | ( n5377 & n5637 ) ;
  assign n5639 = x64 & n5638 ;
  assign n5640 = x65 & n5378 ;
  assign n5641 = x66 | n5640 ;
  assign n5642 = ( n5380 & n5640 ) | ( n5380 & n5641 ) | ( n5640 & n5641 ) ;
  assign n5643 = ( n151 & n152 ) | ( n151 & n5374 ) | ( n152 & n5374 ) ;
  assign n5644 = ( ~n5639 & n5642 ) | ( ~n5639 & n5643 ) | ( n5642 & n5643 ) ;
  assign n5645 = n5639 | n5644 ;
  assign n5646 = n5636 | n5645 ;
  assign n5647 = ( n5636 & n5645 ) | ( n5636 & ~n5646 ) | ( n5645 & ~n5646 ) ;
  assign n5648 = n5646 & ~n5647 ;
  assign n5649 = ( n5396 & n5635 ) | ( n5396 & n5648 ) | ( n5635 & n5648 ) ;
  assign n5650 = ( ~n5396 & n5635 ) | ( ~n5396 & n5648 ) | ( n5635 & n5648 ) ;
  assign n5651 = ( n5396 & ~n5649 ) | ( n5396 & n5650 ) | ( ~n5649 & n5650 ) ;
  assign n5652 = ( n5408 & n5626 ) | ( n5408 & n5651 ) | ( n5626 & n5651 ) ;
  assign n5653 = ( ~n5408 & n5626 ) | ( ~n5408 & n5651 ) | ( n5626 & n5651 ) ;
  assign n5654 = ( n5408 & ~n5652 ) | ( n5408 & n5653 ) | ( ~n5652 & n5653 ) ;
  assign n5655 = ( n5420 & n5617 ) | ( n5420 & n5654 ) | ( n5617 & n5654 ) ;
  assign n5656 = ( ~n5420 & n5617 ) | ( ~n5420 & n5654 ) | ( n5617 & n5654 ) ;
  assign n5657 = ( n5420 & ~n5655 ) | ( n5420 & n5656 ) | ( ~n5655 & n5656 ) ;
  assign n5658 = n637 & n3224 ;
  assign n5659 = x77 & n3228 ;
  assign n5660 = x78 | n5659 ;
  assign n5661 = ( n3230 & n5659 ) | ( n3230 & n5660 ) | ( n5659 & n5660 ) ;
  assign n5662 = x76 & n3413 ;
  assign n5663 = n5661 | n5662 ;
  assign n5664 = ( x38 & n5658 ) | ( x38 & ~n5663 ) | ( n5658 & ~n5663 ) ;
  assign n5665 = ( ~x38 & n5663 ) | ( ~x38 & n5664 ) | ( n5663 & n5664 ) ;
  assign n5666 = ( ~n5658 & n5664 ) | ( ~n5658 & n5665 ) | ( n5664 & n5665 ) ;
  assign n5667 = ( n5423 & n5657 ) | ( n5423 & n5666 ) | ( n5657 & n5666 ) ;
  assign n5668 = ( ~n5423 & n5657 ) | ( ~n5423 & n5666 ) | ( n5657 & n5666 ) ;
  assign n5669 = ( n5423 & ~n5667 ) | ( n5423 & n5668 ) | ( ~n5667 & n5668 ) ;
  assign n5670 = ( n5435 & n5608 ) | ( n5435 & n5669 ) | ( n5608 & n5669 ) ;
  assign n5671 = ( ~n5435 & n5608 ) | ( ~n5435 & n5669 ) | ( n5608 & n5669 ) ;
  assign n5672 = ( n5435 & ~n5670 ) | ( n5435 & n5671 ) | ( ~n5670 & n5671 ) ;
  assign n5673 = ( n5447 & n5599 ) | ( n5447 & n5672 ) | ( n5599 & n5672 ) ;
  assign n5674 = ( ~n5447 & n5599 ) | ( ~n5447 & n5672 ) | ( n5599 & n5672 ) ;
  assign n5675 = ( n5447 & ~n5673 ) | ( n5447 & n5674 ) | ( ~n5673 & n5674 ) ;
  assign n5676 = n1466 & n1949 ;
  assign n5677 = x86 & n1953 ;
  assign n5678 = x87 | n5677 ;
  assign n5679 = ( n1955 & n5677 ) | ( n1955 & n5678 ) | ( n5677 & n5678 ) ;
  assign n5680 = x85 & n2114 ;
  assign n5681 = n5679 | n5680 ;
  assign n5682 = ( x29 & n5676 ) | ( x29 & ~n5681 ) | ( n5676 & ~n5681 ) ;
  assign n5683 = ( ~x29 & n5681 ) | ( ~x29 & n5682 ) | ( n5681 & n5682 ) ;
  assign n5684 = ( ~n5676 & n5682 ) | ( ~n5676 & n5683 ) | ( n5682 & n5683 ) ;
  assign n5685 = ( n5459 & n5675 ) | ( n5459 & n5684 ) | ( n5675 & n5684 ) ;
  assign n5686 = ( ~n5459 & n5675 ) | ( ~n5459 & n5684 ) | ( n5675 & n5684 ) ;
  assign n5687 = ( n5459 & ~n5685 ) | ( n5459 & n5686 ) | ( ~n5685 & n5686 ) ;
  assign n5688 = ( n5471 & n5590 ) | ( n5471 & n5687 ) | ( n5590 & n5687 ) ;
  assign n5689 = ( ~n5471 & n5590 ) | ( ~n5471 & n5687 ) | ( n5590 & n5687 ) ;
  assign n5690 = ( n5471 & ~n5688 ) | ( n5471 & n5689 ) | ( ~n5688 & n5689 ) ;
  assign n5691 = ( n5474 & n5581 ) | ( n5474 & n5690 ) | ( n5581 & n5690 ) ;
  assign n5692 = ( ~n5474 & n5581 ) | ( ~n5474 & n5690 ) | ( n5581 & n5690 ) ;
  assign n5693 = ( n5474 & ~n5691 ) | ( n5474 & n5692 ) | ( ~n5691 & n5692 ) ;
  assign n5694 = ( n5477 & n5572 ) | ( n5477 & n5693 ) | ( n5572 & n5693 ) ;
  assign n5695 = ( ~n5477 & n5572 ) | ( ~n5477 & n5693 ) | ( n5572 & n5693 ) ;
  assign n5696 = ( n5477 & ~n5694 ) | ( n5477 & n5695 ) | ( ~n5694 & n5695 ) ;
  assign n5697 = n810 & n2877 ;
  assign n5698 = x98 & n814 ;
  assign n5699 = x99 | n5698 ;
  assign n5700 = ( n816 & n5698 ) | ( n816 & n5699 ) | ( n5698 & n5699 ) ;
  assign n5701 = x97 & n885 ;
  assign n5702 = n5700 | n5701 ;
  assign n5703 = ( x17 & n5697 ) | ( x17 & ~n5702 ) | ( n5697 & ~n5702 ) ;
  assign n5704 = ( ~x17 & n5702 ) | ( ~x17 & n5703 ) | ( n5702 & n5703 ) ;
  assign n5705 = ( ~n5697 & n5703 ) | ( ~n5697 & n5704 ) | ( n5703 & n5704 ) ;
  assign n5706 = ( n5489 & n5696 ) | ( n5489 & n5705 ) | ( n5696 & n5705 ) ;
  assign n5707 = ( ~n5489 & n5696 ) | ( ~n5489 & n5705 ) | ( n5696 & n5705 ) ;
  assign n5708 = ( n5489 & ~n5706 ) | ( n5489 & n5707 ) | ( ~n5706 & n5707 ) ;
  assign n5709 = n583 & n3486 ;
  assign n5710 = x101 & n587 ;
  assign n5711 = x102 | n5710 ;
  assign n5712 = ( n589 & n5710 ) | ( n589 & n5711 ) | ( n5710 & n5711 ) ;
  assign n5713 = x100 & n676 ;
  assign n5714 = n5712 | n5713 ;
  assign n5715 = ( x14 & n5709 ) | ( x14 & ~n5714 ) | ( n5709 & ~n5714 ) ;
  assign n5716 = ( ~x14 & n5714 ) | ( ~x14 & n5715 ) | ( n5714 & n5715 ) ;
  assign n5717 = ( ~n5709 & n5715 ) | ( ~n5709 & n5716 ) | ( n5715 & n5716 ) ;
  assign n5718 = ( n5501 & n5708 ) | ( n5501 & n5717 ) | ( n5708 & n5717 ) ;
  assign n5719 = ( ~n5501 & n5708 ) | ( ~n5501 & n5717 ) | ( n5708 & n5717 ) ;
  assign n5720 = ( n5501 & ~n5718 ) | ( n5501 & n5719 ) | ( ~n5718 & n5719 ) ;
  assign n5721 = n407 & n3998 ;
  assign n5722 = x104 & n411 ;
  assign n5723 = x105 | n5722 ;
  assign n5724 = ( n413 & n5722 ) | ( n413 & n5723 ) | ( n5722 & n5723 ) ;
  assign n5725 = x103 & n491 ;
  assign n5726 = n5724 | n5725 ;
  assign n5727 = ( x11 & n5721 ) | ( x11 & ~n5726 ) | ( n5721 & ~n5726 ) ;
  assign n5728 = ( ~x11 & n5726 ) | ( ~x11 & n5727 ) | ( n5726 & n5727 ) ;
  assign n5729 = ( ~n5721 & n5727 ) | ( ~n5721 & n5728 ) | ( n5727 & n5728 ) ;
  assign n5730 = ( n5513 & n5720 ) | ( n5513 & n5729 ) | ( n5720 & n5729 ) ;
  assign n5731 = ( ~n5513 & n5720 ) | ( ~n5513 & n5729 ) | ( n5720 & n5729 ) ;
  assign n5732 = ( n5513 & ~n5730 ) | ( n5513 & n5731 ) | ( ~n5730 & n5731 ) ;
  assign n5733 = n291 & n4377 ;
  assign n5734 = x107 & n295 ;
  assign n5735 = x108 | n5734 ;
  assign n5736 = ( n297 & n5734 ) | ( n297 & n5735 ) | ( n5734 & n5735 ) ;
  assign n5737 = x106 & n330 ;
  assign n5738 = n5736 | n5737 ;
  assign n5739 = ( x8 & n5733 ) | ( x8 & ~n5738 ) | ( n5733 & ~n5738 ) ;
  assign n5740 = ( ~x8 & n5738 ) | ( ~x8 & n5739 ) | ( n5738 & n5739 ) ;
  assign n5741 = ( ~n5733 & n5739 ) | ( ~n5733 & n5740 ) | ( n5739 & n5740 ) ;
  assign n5742 = ( n5525 & n5732 ) | ( n5525 & n5741 ) | ( n5732 & n5741 ) ;
  assign n5743 = ( ~n5525 & n5732 ) | ( ~n5525 & n5741 ) | ( n5732 & n5741 ) ;
  assign n5744 = ( n5525 & ~n5742 ) | ( n5525 & n5743 ) | ( ~n5742 & n5743 ) ;
  assign n5745 = ( n5537 & n5563 ) | ( n5537 & n5744 ) | ( n5563 & n5744 ) ;
  assign n5746 = ( ~n5537 & n5563 ) | ( ~n5537 & n5744 ) | ( n5563 & n5744 ) ;
  assign n5747 = ( n5537 & ~n5745 ) | ( n5537 & n5746 ) | ( ~n5745 & n5746 ) ;
  assign n5748 = ( x113 & x114 ) | ( x113 & n5540 ) | ( x114 & n5540 ) ;
  assign n5749 = ( x113 & ~x114 ) | ( x113 & n5540 ) | ( ~x114 & n5540 ) ;
  assign n5750 = ( x114 & ~n5748 ) | ( x114 & n5749 ) | ( ~n5748 & n5749 ) ;
  assign n5751 = n136 & n5750 ;
  assign n5752 = x113 & n138 ;
  assign n5753 = x114 | n5752 ;
  assign n5754 = ( n141 & n5752 ) | ( n141 & n5753 ) | ( n5752 & n5753 ) ;
  assign n5755 = x112 & n154 ;
  assign n5756 = n5754 | n5755 ;
  assign n5757 = ( x2 & n5751 ) | ( x2 & ~n5756 ) | ( n5751 & ~n5756 ) ;
  assign n5758 = ( ~x2 & n5756 ) | ( ~x2 & n5757 ) | ( n5756 & n5757 ) ;
  assign n5759 = ( ~n5751 & n5757 ) | ( ~n5751 & n5758 ) | ( n5757 & n5758 ) ;
  assign n5760 = ( n5552 & n5747 ) | ( n5552 & n5759 ) | ( n5747 & n5759 ) ;
  assign n5761 = ( ~n5552 & n5747 ) | ( ~n5552 & n5759 ) | ( n5747 & n5759 ) ;
  assign n5762 = ( n5552 & ~n5760 ) | ( n5552 & n5761 ) | ( ~n5760 & n5761 ) ;
  assign n5763 = ( x114 & x115 ) | ( x114 & n5748 ) | ( x115 & n5748 ) ;
  assign n5764 = ( x114 & ~x115 ) | ( x114 & n5748 ) | ( ~x115 & n5748 ) ;
  assign n5765 = ( x115 & ~n5763 ) | ( x115 & n5764 ) | ( ~n5763 & n5764 ) ;
  assign n5766 = n136 & n5765 ;
  assign n5767 = x114 & n138 ;
  assign n5768 = x115 | n5767 ;
  assign n5769 = ( n141 & n5767 ) | ( n141 & n5768 ) | ( n5767 & n5768 ) ;
  assign n5770 = x113 & n154 ;
  assign n5771 = n5769 | n5770 ;
  assign n5772 = ( x2 & n5766 ) | ( x2 & ~n5771 ) | ( n5766 & ~n5771 ) ;
  assign n5773 = ( ~x2 & n5771 ) | ( ~x2 & n5772 ) | ( n5771 & n5772 ) ;
  assign n5774 = ( ~n5766 & n5772 ) | ( ~n5766 & n5773 ) | ( n5772 & n5773 ) ;
  assign n5775 = n186 & n5145 ;
  assign n5776 = x111 & n190 ;
  assign n5777 = x112 | n5776 ;
  assign n5778 = ( n192 & n5776 ) | ( n192 & n5777 ) | ( n5776 & n5777 ) ;
  assign n5779 = x110 & n220 ;
  assign n5780 = n5778 | n5779 ;
  assign n5781 = ( x5 & n5775 ) | ( x5 & ~n5780 ) | ( n5775 & ~n5780 ) ;
  assign n5782 = ( ~x5 & n5780 ) | ( ~x5 & n5781 ) | ( n5780 & n5781 ) ;
  assign n5783 = ( ~n5775 & n5781 ) | ( ~n5775 & n5782 ) | ( n5781 & n5782 ) ;
  assign n5784 = n810 & n3162 ;
  assign n5785 = x99 & n814 ;
  assign n5786 = x100 | n5785 ;
  assign n5787 = ( n816 & n5785 ) | ( n816 & n5786 ) | ( n5785 & n5786 ) ;
  assign n5788 = x98 & n885 ;
  assign n5789 = n5787 | n5788 ;
  assign n5790 = ( x17 & n5784 ) | ( x17 & ~n5789 ) | ( n5784 & ~n5789 ) ;
  assign n5791 = ( ~x17 & n5789 ) | ( ~x17 & n5790 ) | ( n5789 & n5790 ) ;
  assign n5792 = ( ~n5784 & n5790 ) | ( ~n5784 & n5791 ) | ( n5790 & n5791 ) ;
  assign n5793 = n1297 & n2294 ;
  assign n5794 = x93 & n1301 ;
  assign n5795 = x94 | n5794 ;
  assign n5796 = ( n1303 & n5794 ) | ( n1303 & n5795 ) | ( n5794 & n5795 ) ;
  assign n5797 = x92 & n1426 ;
  assign n5798 = n5796 | n5797 ;
  assign n5799 = ( x23 & n5793 ) | ( x23 & ~n5798 ) | ( n5793 & ~n5798 ) ;
  assign n5800 = ( ~x23 & n5798 ) | ( ~x23 & n5799 ) | ( n5798 & n5799 ) ;
  assign n5801 = ( ~n5793 & n5799 ) | ( ~n5793 & n5800 ) | ( n5799 & n5800 ) ;
  assign n5802 = n990 & n2766 ;
  assign n5803 = x81 & n2770 ;
  assign n5804 = x82 | n5803 ;
  assign n5805 = ( n2772 & n5803 ) | ( n2772 & n5804 ) | ( n5803 & n5804 ) ;
  assign n5806 = x80 & n2943 ;
  assign n5807 = n5805 | n5806 ;
  assign n5808 = ( x35 & n5802 ) | ( x35 & ~n5807 ) | ( n5802 & ~n5807 ) ;
  assign n5809 = ( ~x35 & n5807 ) | ( ~x35 & n5808 ) | ( n5807 & n5808 ) ;
  assign n5810 = ( ~n5802 & n5808 ) | ( ~n5802 & n5809 ) | ( n5808 & n5809 ) ;
  assign n5811 = n701 & n3224 ;
  assign n5812 = x78 & n3228 ;
  assign n5813 = x79 | n5812 ;
  assign n5814 = ( n3230 & n5812 ) | ( n3230 & n5813 ) | ( n5812 & n5813 ) ;
  assign n5815 = x77 & n3413 ;
  assign n5816 = n5814 | n5815 ;
  assign n5817 = ( x38 & n5811 ) | ( x38 & ~n5816 ) | ( n5811 & ~n5816 ) ;
  assign n5818 = ( ~x38 & n5816 ) | ( ~x38 & n5817 ) | ( n5816 & n5817 ) ;
  assign n5819 = ( ~n5811 & n5817 ) | ( ~n5811 & n5818 ) | ( n5817 & n5818 ) ;
  assign n5820 = n554 & n3715 ;
  assign n5821 = x75 & n3719 ;
  assign n5822 = x76 | n5821 ;
  assign n5823 = ( n3721 & n5821 ) | ( n3721 & n5822 ) | ( n5821 & n5822 ) ;
  assign n5824 = x74 & n3922 ;
  assign n5825 = n5823 | n5824 ;
  assign n5826 = ( x41 & n5820 ) | ( x41 & ~n5825 ) | ( n5820 & ~n5825 ) ;
  assign n5827 = ( ~x41 & n5825 ) | ( ~x41 & n5826 ) | ( n5825 & n5826 ) ;
  assign n5828 = ( ~n5820 & n5826 ) | ( ~n5820 & n5827 ) | ( n5826 & n5827 ) ;
  assign n5829 = x66 & n5378 ;
  assign n5830 = x67 | n5829 ;
  assign n5831 = ( n5380 & n5829 ) | ( n5380 & n5830 ) | ( n5829 & n5830 ) ;
  assign n5832 = x65 & n5638 ;
  assign n5833 = n5831 | n5832 ;
  assign n5834 = n164 & n5374 ;
  assign n5835 = ( x50 & n5833 ) | ( x50 & ~n5834 ) | ( n5833 & ~n5834 ) ;
  assign n5836 = ( ~x50 & n5834 ) | ( ~x50 & n5835 ) | ( n5834 & n5835 ) ;
  assign n5837 = ( ~n5833 & n5835 ) | ( ~n5833 & n5836 ) | ( n5835 & n5836 ) ;
  assign n5838 = x50 & x51 ;
  assign n5839 = x50 | x51 ;
  assign n5840 = ~n5838 & n5839 ;
  assign n5841 = x64 & n5840 ;
  assign n5842 = x50 & ~n5646 ;
  assign n5843 = ( n5837 & n5841 ) | ( n5837 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5844 = ( ~n5837 & n5841 ) | ( ~n5837 & n5842 ) | ( n5841 & n5842 ) ;
  assign n5845 = ( n5837 & ~n5843 ) | ( n5837 & n5844 ) | ( ~n5843 & n5844 ) ;
  assign n5846 = n245 & n4787 ;
  assign n5847 = x69 & n4791 ;
  assign n5848 = x70 | n5847 ;
  assign n5849 = ( n4793 & n5847 ) | ( n4793 & n5848 ) | ( n5847 & n5848 ) ;
  assign n5850 = x68 & n5030 ;
  assign n5851 = n5849 | n5850 ;
  assign n5852 = ( x47 & n5846 ) | ( x47 & ~n5851 ) | ( n5846 & ~n5851 ) ;
  assign n5853 = ( ~x47 & n5851 ) | ( ~x47 & n5852 ) | ( n5851 & n5852 ) ;
  assign n5854 = ( ~n5846 & n5852 ) | ( ~n5846 & n5853 ) | ( n5852 & n5853 ) ;
  assign n5855 = ( n5649 & n5845 ) | ( n5649 & n5854 ) | ( n5845 & n5854 ) ;
  assign n5856 = ( ~n5649 & n5845 ) | ( ~n5649 & n5854 ) | ( n5845 & n5854 ) ;
  assign n5857 = ( n5649 & ~n5855 ) | ( n5649 & n5856 ) | ( ~n5855 & n5856 ) ;
  assign n5858 = n390 & n4227 ;
  assign n5859 = x72 & n4231 ;
  assign n5860 = x73 | n5859 ;
  assign n5861 = ( n4233 & n5859 ) | ( n4233 & n5860 ) | ( n5859 & n5860 ) ;
  assign n5862 = x71 & n4470 ;
  assign n5863 = n5861 | n5862 ;
  assign n5864 = ( x44 & n5858 ) | ( x44 & ~n5863 ) | ( n5858 & ~n5863 ) ;
  assign n5865 = ( ~x44 & n5863 ) | ( ~x44 & n5864 ) | ( n5863 & n5864 ) ;
  assign n5866 = ( ~n5858 & n5864 ) | ( ~n5858 & n5865 ) | ( n5864 & n5865 ) ;
  assign n5867 = ( n5652 & n5857 ) | ( n5652 & n5866 ) | ( n5857 & n5866 ) ;
  assign n5868 = ( ~n5652 & n5857 ) | ( ~n5652 & n5866 ) | ( n5857 & n5866 ) ;
  assign n5869 = ( n5652 & ~n5867 ) | ( n5652 & n5868 ) | ( ~n5867 & n5868 ) ;
  assign n5870 = ( n5655 & n5828 ) | ( n5655 & n5869 ) | ( n5828 & n5869 ) ;
  assign n5871 = ( ~n5655 & n5828 ) | ( ~n5655 & n5869 ) | ( n5828 & n5869 ) ;
  assign n5872 = ( n5655 & ~n5870 ) | ( n5655 & n5871 ) | ( ~n5870 & n5871 ) ;
  assign n5873 = ( n5667 & n5819 ) | ( n5667 & n5872 ) | ( n5819 & n5872 ) ;
  assign n5874 = ( ~n5667 & n5819 ) | ( ~n5667 & n5872 ) | ( n5819 & n5872 ) ;
  assign n5875 = ( n5667 & ~n5873 ) | ( n5667 & n5874 ) | ( ~n5873 & n5874 ) ;
  assign n5876 = ( n5670 & n5810 ) | ( n5670 & n5875 ) | ( n5810 & n5875 ) ;
  assign n5877 = ( ~n5670 & n5810 ) | ( ~n5670 & n5875 ) | ( n5810 & n5875 ) ;
  assign n5878 = ( n5670 & ~n5876 ) | ( n5670 & n5877 ) | ( ~n5876 & n5877 ) ;
  assign n5879 = n1262 & n2320 ;
  assign n5880 = x84 & n2324 ;
  assign n5881 = x85 | n5880 ;
  assign n5882 = ( n2326 & n5880 ) | ( n2326 & n5881 ) | ( n5880 & n5881 ) ;
  assign n5883 = x83 & n2497 ;
  assign n5884 = n5882 | n5883 ;
  assign n5885 = ( x32 & n5879 ) | ( x32 & ~n5884 ) | ( n5879 & ~n5884 ) ;
  assign n5886 = ( ~x32 & n5884 ) | ( ~x32 & n5885 ) | ( n5884 & n5885 ) ;
  assign n5887 = ( ~n5879 & n5885 ) | ( ~n5879 & n5886 ) | ( n5885 & n5886 ) ;
  assign n5888 = ( n5673 & n5878 ) | ( n5673 & n5887 ) | ( n5878 & n5887 ) ;
  assign n5889 = ( ~n5673 & n5878 ) | ( ~n5673 & n5887 ) | ( n5878 & n5887 ) ;
  assign n5890 = ( n5673 & ~n5888 ) | ( n5673 & n5889 ) | ( ~n5888 & n5889 ) ;
  assign n5891 = n1481 & n1949 ;
  assign n5892 = x87 & n1953 ;
  assign n5893 = x88 | n5892 ;
  assign n5894 = ( n1955 & n5892 ) | ( n1955 & n5893 ) | ( n5892 & n5893 ) ;
  assign n5895 = x86 & n2114 ;
  assign n5896 = n5894 | n5895 ;
  assign n5897 = ( x29 & n5891 ) | ( x29 & ~n5896 ) | ( n5891 & ~n5896 ) ;
  assign n5898 = ( ~x29 & n5896 ) | ( ~x29 & n5897 ) | ( n5896 & n5897 ) ;
  assign n5899 = ( ~n5891 & n5897 ) | ( ~n5891 & n5898 ) | ( n5897 & n5898 ) ;
  assign n5900 = ( n5685 & n5890 ) | ( n5685 & n5899 ) | ( n5890 & n5899 ) ;
  assign n5901 = ( ~n5685 & n5890 ) | ( ~n5685 & n5899 ) | ( n5890 & n5899 ) ;
  assign n5902 = ( n5685 & ~n5900 ) | ( n5685 & n5901 ) | ( ~n5900 & n5901 ) ;
  assign n5903 = n1617 & n1914 ;
  assign n5904 = x90 & n1621 ;
  assign n5905 = x91 | n5904 ;
  assign n5906 = ( n1623 & n5904 ) | ( n1623 & n5905 ) | ( n5904 & n5905 ) ;
  assign n5907 = x89 & n1749 ;
  assign n5908 = n5906 | n5907 ;
  assign n5909 = ( x26 & n5903 ) | ( x26 & ~n5908 ) | ( n5903 & ~n5908 ) ;
  assign n5910 = ( ~x26 & n5908 ) | ( ~x26 & n5909 ) | ( n5908 & n5909 ) ;
  assign n5911 = ( ~n5903 & n5909 ) | ( ~n5903 & n5910 ) | ( n5909 & n5910 ) ;
  assign n5912 = ( n5688 & n5902 ) | ( n5688 & n5911 ) | ( n5902 & n5911 ) ;
  assign n5913 = ( ~n5688 & n5902 ) | ( ~n5688 & n5911 ) | ( n5902 & n5911 ) ;
  assign n5914 = ( n5688 & ~n5912 ) | ( n5688 & n5913 ) | ( ~n5912 & n5913 ) ;
  assign n5915 = ( n5691 & n5801 ) | ( n5691 & n5914 ) | ( n5801 & n5914 ) ;
  assign n5916 = ( ~n5691 & n5801 ) | ( ~n5691 & n5914 ) | ( n5801 & n5914 ) ;
  assign n5917 = ( n5691 & ~n5915 ) | ( n5691 & n5916 ) | ( ~n5915 & n5916 ) ;
  assign n5918 = n1016 & n2585 ;
  assign n5919 = x96 & n1020 ;
  assign n5920 = x97 | n5919 ;
  assign n5921 = ( n1022 & n5919 ) | ( n1022 & n5920 ) | ( n5919 & n5920 ) ;
  assign n5922 = x95 & n1145 ;
  assign n5923 = n5921 | n5922 ;
  assign n5924 = ( x20 & n5918 ) | ( x20 & ~n5923 ) | ( n5918 & ~n5923 ) ;
  assign n5925 = ( ~x20 & n5923 ) | ( ~x20 & n5924 ) | ( n5923 & n5924 ) ;
  assign n5926 = ( ~n5918 & n5924 ) | ( ~n5918 & n5925 ) | ( n5924 & n5925 ) ;
  assign n5927 = ( n5694 & n5917 ) | ( n5694 & n5926 ) | ( n5917 & n5926 ) ;
  assign n5928 = ( ~n5694 & n5917 ) | ( ~n5694 & n5926 ) | ( n5917 & n5926 ) ;
  assign n5929 = ( n5694 & ~n5927 ) | ( n5694 & n5928 ) | ( ~n5927 & n5928 ) ;
  assign n5930 = ( n5706 & n5792 ) | ( n5706 & n5929 ) | ( n5792 & n5929 ) ;
  assign n5931 = ( ~n5706 & n5792 ) | ( ~n5706 & n5929 ) | ( n5792 & n5929 ) ;
  assign n5932 = ( n5706 & ~n5930 ) | ( n5706 & n5931 ) | ( ~n5930 & n5931 ) ;
  assign n5933 = n583 & n3650 ;
  assign n5934 = x102 & n587 ;
  assign n5935 = x103 | n5934 ;
  assign n5936 = ( n589 & n5934 ) | ( n589 & n5935 ) | ( n5934 & n5935 ) ;
  assign n5937 = x101 & n676 ;
  assign n5938 = n5936 | n5937 ;
  assign n5939 = ( x14 & n5933 ) | ( x14 & ~n5938 ) | ( n5933 & ~n5938 ) ;
  assign n5940 = ( ~x14 & n5938 ) | ( ~x14 & n5939 ) | ( n5938 & n5939 ) ;
  assign n5941 = ( ~n5933 & n5939 ) | ( ~n5933 & n5940 ) | ( n5939 & n5940 ) ;
  assign n5942 = ( n5718 & n5932 ) | ( n5718 & n5941 ) | ( n5932 & n5941 ) ;
  assign n5943 = ( ~n5718 & n5932 ) | ( ~n5718 & n5941 ) | ( n5932 & n5941 ) ;
  assign n5944 = ( n5718 & ~n5942 ) | ( n5718 & n5943 ) | ( ~n5942 & n5943 ) ;
  assign n5945 = n407 & n4013 ;
  assign n5946 = x105 & n411 ;
  assign n5947 = x106 | n5946 ;
  assign n5948 = ( n413 & n5946 ) | ( n413 & n5947 ) | ( n5946 & n5947 ) ;
  assign n5949 = x104 & n491 ;
  assign n5950 = n5948 | n5949 ;
  assign n5951 = ( x11 & n5945 ) | ( x11 & ~n5950 ) | ( n5945 & ~n5950 ) ;
  assign n5952 = ( ~x11 & n5950 ) | ( ~x11 & n5951 ) | ( n5950 & n5951 ) ;
  assign n5953 = ( ~n5945 & n5951 ) | ( ~n5945 & n5952 ) | ( n5951 & n5952 ) ;
  assign n5954 = ( n5730 & n5944 ) | ( n5730 & n5953 ) | ( n5944 & n5953 ) ;
  assign n5955 = ( n5730 & ~n5944 ) | ( n5730 & n5953 ) | ( ~n5944 & n5953 ) ;
  assign n5956 = ( n5944 & ~n5954 ) | ( n5944 & n5955 ) | ( ~n5954 & n5955 ) ;
  assign n5957 = n291 & n4734 ;
  assign n5958 = x108 & n295 ;
  assign n5959 = x109 | n5958 ;
  assign n5960 = ( n297 & n5958 ) | ( n297 & n5959 ) | ( n5958 & n5959 ) ;
  assign n5961 = x107 & n330 ;
  assign n5962 = n5960 | n5961 ;
  assign n5963 = ( x8 & n5957 ) | ( x8 & ~n5962 ) | ( n5957 & ~n5962 ) ;
  assign n5964 = ( ~x8 & n5962 ) | ( ~x8 & n5963 ) | ( n5962 & n5963 ) ;
  assign n5965 = ( ~n5957 & n5963 ) | ( ~n5957 & n5964 ) | ( n5963 & n5964 ) ;
  assign n5966 = ( n5742 & n5956 ) | ( n5742 & n5965 ) | ( n5956 & n5965 ) ;
  assign n5967 = ( ~n5742 & n5956 ) | ( ~n5742 & n5965 ) | ( n5956 & n5965 ) ;
  assign n5968 = ( n5742 & ~n5966 ) | ( n5742 & n5967 ) | ( ~n5966 & n5967 ) ;
  assign n5969 = ( n5745 & n5783 ) | ( n5745 & n5968 ) | ( n5783 & n5968 ) ;
  assign n5970 = ( ~n5745 & n5783 ) | ( ~n5745 & n5968 ) | ( n5783 & n5968 ) ;
  assign n5971 = ( n5745 & ~n5969 ) | ( n5745 & n5970 ) | ( ~n5969 & n5970 ) ;
  assign n5972 = ( n5760 & n5774 ) | ( n5760 & n5971 ) | ( n5774 & n5971 ) ;
  assign n5973 = ( ~n5760 & n5774 ) | ( ~n5760 & n5971 ) | ( n5774 & n5971 ) ;
  assign n5974 = ( n5760 & ~n5972 ) | ( n5760 & n5973 ) | ( ~n5972 & n5973 ) ;
  assign n5975 = ( x115 & x116 ) | ( x115 & n5763 ) | ( x116 & n5763 ) ;
  assign n5976 = ( x115 & ~x116 ) | ( x115 & n5763 ) | ( ~x116 & n5763 ) ;
  assign n5977 = ( x116 & ~n5975 ) | ( x116 & n5976 ) | ( ~n5975 & n5976 ) ;
  assign n5978 = n136 & n5977 ;
  assign n5979 = x115 & n138 ;
  assign n5980 = x116 | n5979 ;
  assign n5981 = ( n141 & n5979 ) | ( n141 & n5980 ) | ( n5979 & n5980 ) ;
  assign n5982 = x114 & n154 ;
  assign n5983 = n5981 | n5982 ;
  assign n5984 = ( x2 & n5978 ) | ( x2 & ~n5983 ) | ( n5978 & ~n5983 ) ;
  assign n5985 = ( ~x2 & n5983 ) | ( ~x2 & n5984 ) | ( n5983 & n5984 ) ;
  assign n5986 = ( ~n5978 & n5984 ) | ( ~n5978 & n5985 ) | ( n5984 & n5985 ) ;
  assign n5987 = n291 & n4934 ;
  assign n5988 = x109 & n295 ;
  assign n5989 = x110 | n5988 ;
  assign n5990 = ( n297 & n5988 ) | ( n297 & n5989 ) | ( n5988 & n5989 ) ;
  assign n5991 = x108 & n330 ;
  assign n5992 = n5990 | n5991 ;
  assign n5993 = ( x8 & n5987 ) | ( x8 & ~n5992 ) | ( n5987 & ~n5992 ) ;
  assign n5994 = ( ~x8 & n5992 ) | ( ~x8 & n5993 ) | ( n5992 & n5993 ) ;
  assign n5995 = ( ~n5987 & n5993 ) | ( ~n5987 & n5994 ) | ( n5993 & n5994 ) ;
  assign n5996 = n1617 & n2042 ;
  assign n5997 = x91 & n1621 ;
  assign n5998 = x92 | n5997 ;
  assign n5999 = ( n1623 & n5997 ) | ( n1623 & n5998 ) | ( n5997 & n5998 ) ;
  assign n6000 = x90 & n1749 ;
  assign n6001 = n5999 | n6000 ;
  assign n6002 = ( x26 & n5996 ) | ( x26 & ~n6001 ) | ( n5996 & ~n6001 ) ;
  assign n6003 = ( ~x26 & n6001 ) | ( ~x26 & n6002 ) | ( n6001 & n6002 ) ;
  assign n6004 = ( ~n5996 & n6002 ) | ( ~n5996 & n6003 ) | ( n6002 & n6003 ) ;
  assign n6005 = n1366 & n2320 ;
  assign n6006 = x85 & n2324 ;
  assign n6007 = x86 | n6006 ;
  assign n6008 = ( n2326 & n6006 ) | ( n2326 & n6007 ) | ( n6006 & n6007 ) ;
  assign n6009 = x84 & n2497 ;
  assign n6010 = n6008 | n6009 ;
  assign n6011 = ( x32 & n6005 ) | ( x32 & ~n6010 ) | ( n6005 & ~n6010 ) ;
  assign n6012 = ( ~x32 & n6010 ) | ( ~x32 & n6011 ) | ( n6010 & n6011 ) ;
  assign n6013 = ( ~n6005 & n6011 ) | ( ~n6005 & n6012 ) | ( n6011 & n6012 ) ;
  assign n6014 = n569 & n3715 ;
  assign n6015 = x76 & n3719 ;
  assign n6016 = x77 | n6015 ;
  assign n6017 = ( n3721 & n6015 ) | ( n3721 & n6016 ) | ( n6015 & n6016 ) ;
  assign n6018 = x75 & n3922 ;
  assign n6019 = n6017 | n6018 ;
  assign n6020 = ( x41 & n6014 ) | ( x41 & ~n6019 ) | ( n6014 & ~n6019 ) ;
  assign n6021 = ( ~x41 & n6019 ) | ( ~x41 & n6020 ) | ( n6019 & n6020 ) ;
  assign n6022 = ( ~n6014 & n6020 ) | ( ~n6014 & n6021 ) | ( n6020 & n6021 ) ;
  assign n6023 = x53 & n5841 ;
  assign n6024 = x52 | x53 ;
  assign n6025 = ( x52 & x53 ) | ( x52 & ~n6024 ) | ( x53 & ~n6024 ) ;
  assign n6026 = n6024 & ~n6025 ;
  assign n6027 = n5840 & n6026 ;
  assign n6028 = n133 & n6027 ;
  assign n6029 = ~x50 & x52 ;
  assign n6030 = x51 & x52 ;
  assign n6031 = ( n5838 & n6029 ) | ( n5838 & ~n6030 ) | ( n6029 & ~n6030 ) ;
  assign n6032 = x64 & n6031 ;
  assign n6033 = ( n5840 & ~n6024 ) | ( n5840 & n6025 ) | ( ~n6024 & n6025 ) ;
  assign n6034 = x65 | n6032 ;
  assign n6035 = ( n6032 & n6033 ) | ( n6032 & n6034 ) | ( n6033 & n6034 ) ;
  assign n6036 = ( n6023 & n6028 ) | ( n6023 & n6035 ) | ( n6028 & n6035 ) ;
  assign n6037 = n6028 | n6035 ;
  assign n6038 = ~n6023 & n6037 ;
  assign n6039 = ( n6023 & ~n6036 ) | ( n6023 & n6038 ) | ( ~n6036 & n6038 ) ;
  assign n6040 = x67 & n5378 ;
  assign n6041 = x68 | n6040 ;
  assign n6042 = ( n5380 & n6040 ) | ( n5380 & n6041 ) | ( n6040 & n6041 ) ;
  assign n6043 = x66 & n5638 ;
  assign n6044 = n6042 | n6043 ;
  assign n6045 = n201 & n5374 ;
  assign n6046 = ( x50 & n6044 ) | ( x50 & ~n6045 ) | ( n6044 & ~n6045 ) ;
  assign n6047 = ( ~x50 & n6045 ) | ( ~x50 & n6046 ) | ( n6045 & n6046 ) ;
  assign n6048 = ( ~n6044 & n6046 ) | ( ~n6044 & n6047 ) | ( n6046 & n6047 ) ;
  assign n6049 = ( n5843 & n6039 ) | ( n5843 & n6048 ) | ( n6039 & n6048 ) ;
  assign n6050 = ( ~n5843 & n6039 ) | ( ~n5843 & n6048 ) | ( n6039 & n6048 ) ;
  assign n6051 = ( n5843 & ~n6049 ) | ( n5843 & n6050 ) | ( ~n6049 & n6050 ) ;
  assign n6052 = n277 & n4787 ;
  assign n6053 = x70 & n4791 ;
  assign n6054 = x71 | n6053 ;
  assign n6055 = ( n4793 & n6053 ) | ( n4793 & n6054 ) | ( n6053 & n6054 ) ;
  assign n6056 = x69 & n5030 ;
  assign n6057 = n6055 | n6056 ;
  assign n6058 = ( x47 & n6052 ) | ( x47 & ~n6057 ) | ( n6052 & ~n6057 ) ;
  assign n6059 = ( ~x47 & n6057 ) | ( ~x47 & n6058 ) | ( n6057 & n6058 ) ;
  assign n6060 = ( ~n6052 & n6058 ) | ( ~n6052 & n6059 ) | ( n6058 & n6059 ) ;
  assign n6061 = ( n5855 & n6051 ) | ( n5855 & n6060 ) | ( n6051 & n6060 ) ;
  assign n6062 = ( ~n5855 & n6051 ) | ( ~n5855 & n6060 ) | ( n6051 & n6060 ) ;
  assign n6063 = ( n5855 & ~n6061 ) | ( n5855 & n6062 ) | ( ~n6061 & n6062 ) ;
  assign n6064 = n446 & n4227 ;
  assign n6065 = x73 & n4231 ;
  assign n6066 = x74 | n6065 ;
  assign n6067 = ( n4233 & n6065 ) | ( n4233 & n6066 ) | ( n6065 & n6066 ) ;
  assign n6068 = x72 & n4470 ;
  assign n6069 = n6067 | n6068 ;
  assign n6070 = ( x44 & n6064 ) | ( x44 & ~n6069 ) | ( n6064 & ~n6069 ) ;
  assign n6071 = ( ~x44 & n6069 ) | ( ~x44 & n6070 ) | ( n6069 & n6070 ) ;
  assign n6072 = ( ~n6064 & n6070 ) | ( ~n6064 & n6071 ) | ( n6070 & n6071 ) ;
  assign n6073 = ( n5867 & n6063 ) | ( n5867 & n6072 ) | ( n6063 & n6072 ) ;
  assign n6074 = ( ~n5867 & n6063 ) | ( ~n5867 & n6072 ) | ( n6063 & n6072 ) ;
  assign n6075 = ( n5867 & ~n6073 ) | ( n5867 & n6074 ) | ( ~n6073 & n6074 ) ;
  assign n6076 = ( n5870 & n6022 ) | ( n5870 & n6075 ) | ( n6022 & n6075 ) ;
  assign n6077 = ( ~n5870 & n6022 ) | ( ~n5870 & n6075 ) | ( n6022 & n6075 ) ;
  assign n6078 = ( n5870 & ~n6076 ) | ( n5870 & n6077 ) | ( ~n6076 & n6077 ) ;
  assign n6079 = n769 & n3224 ;
  assign n6080 = x79 & n3228 ;
  assign n6081 = x80 | n6080 ;
  assign n6082 = ( n3230 & n6080 ) | ( n3230 & n6081 ) | ( n6080 & n6081 ) ;
  assign n6083 = x78 & n3413 ;
  assign n6084 = n6082 | n6083 ;
  assign n6085 = ( x38 & n6079 ) | ( x38 & ~n6084 ) | ( n6079 & ~n6084 ) ;
  assign n6086 = ( ~x38 & n6084 ) | ( ~x38 & n6085 ) | ( n6084 & n6085 ) ;
  assign n6087 = ( ~n6079 & n6085 ) | ( ~n6079 & n6086 ) | ( n6085 & n6086 ) ;
  assign n6088 = ( n5873 & n6078 ) | ( n5873 & n6087 ) | ( n6078 & n6087 ) ;
  assign n6089 = ( ~n5873 & n6078 ) | ( ~n5873 & n6087 ) | ( n6078 & n6087 ) ;
  assign n6090 = ( n5873 & ~n6088 ) | ( n5873 & n6089 ) | ( ~n6088 & n6089 ) ;
  assign n6091 = n1082 & n2766 ;
  assign n6092 = x82 & n2770 ;
  assign n6093 = x83 | n6092 ;
  assign n6094 = ( n2772 & n6092 ) | ( n2772 & n6093 ) | ( n6092 & n6093 ) ;
  assign n6095 = x81 & n2943 ;
  assign n6096 = n6094 | n6095 ;
  assign n6097 = ( x35 & n6091 ) | ( x35 & ~n6096 ) | ( n6091 & ~n6096 ) ;
  assign n6098 = ( ~x35 & n6096 ) | ( ~x35 & n6097 ) | ( n6096 & n6097 ) ;
  assign n6099 = ( ~n6091 & n6097 ) | ( ~n6091 & n6098 ) | ( n6097 & n6098 ) ;
  assign n6100 = ( n5876 & n6090 ) | ( n5876 & n6099 ) | ( n6090 & n6099 ) ;
  assign n6101 = ( ~n5876 & n6090 ) | ( ~n5876 & n6099 ) | ( n6090 & n6099 ) ;
  assign n6102 = ( n5876 & ~n6100 ) | ( n5876 & n6101 ) | ( ~n6100 & n6101 ) ;
  assign n6103 = ( n5888 & n6013 ) | ( n5888 & n6102 ) | ( n6013 & n6102 ) ;
  assign n6104 = ( ~n5888 & n6013 ) | ( ~n5888 & n6102 ) | ( n6013 & n6102 ) ;
  assign n6105 = ( n5888 & ~n6103 ) | ( n5888 & n6104 ) | ( ~n6103 & n6104 ) ;
  assign n6106 = n1585 & n1949 ;
  assign n6107 = x88 & n1953 ;
  assign n6108 = x89 | n6107 ;
  assign n6109 = ( n1955 & n6107 ) | ( n1955 & n6108 ) | ( n6107 & n6108 ) ;
  assign n6110 = x87 & n2114 ;
  assign n6111 = n6109 | n6110 ;
  assign n6112 = ( x29 & n6106 ) | ( x29 & ~n6111 ) | ( n6106 & ~n6111 ) ;
  assign n6113 = ( ~x29 & n6111 ) | ( ~x29 & n6112 ) | ( n6111 & n6112 ) ;
  assign n6114 = ( ~n6106 & n6112 ) | ( ~n6106 & n6113 ) | ( n6112 & n6113 ) ;
  assign n6115 = ( n5900 & n6105 ) | ( n5900 & n6114 ) | ( n6105 & n6114 ) ;
  assign n6116 = ( ~n5900 & n6105 ) | ( ~n5900 & n6114 ) | ( n6105 & n6114 ) ;
  assign n6117 = ( n5900 & ~n6115 ) | ( n5900 & n6116 ) | ( ~n6115 & n6116 ) ;
  assign n6118 = ( n5912 & n6004 ) | ( n5912 & n6117 ) | ( n6004 & n6117 ) ;
  assign n6119 = ( ~n5912 & n6004 ) | ( ~n5912 & n6117 ) | ( n6004 & n6117 ) ;
  assign n6120 = ( n5912 & ~n6118 ) | ( n5912 & n6119 ) | ( ~n6118 & n6119 ) ;
  assign n6121 = n1297 & n2434 ;
  assign n6122 = x94 & n1301 ;
  assign n6123 = x95 | n6122 ;
  assign n6124 = ( n1303 & n6122 ) | ( n1303 & n6123 ) | ( n6122 & n6123 ) ;
  assign n6125 = x93 & n1426 ;
  assign n6126 = n6124 | n6125 ;
  assign n6127 = ( x23 & n6121 ) | ( x23 & ~n6126 ) | ( n6121 & ~n6126 ) ;
  assign n6128 = ( ~x23 & n6126 ) | ( ~x23 & n6127 ) | ( n6126 & n6127 ) ;
  assign n6129 = ( ~n6121 & n6127 ) | ( ~n6121 & n6128 ) | ( n6127 & n6128 ) ;
  assign n6130 = ( n5915 & n6120 ) | ( n5915 & n6129 ) | ( n6120 & n6129 ) ;
  assign n6131 = ( ~n5915 & n6120 ) | ( ~n5915 & n6129 ) | ( n6120 & n6129 ) ;
  assign n6132 = ( n5915 & ~n6130 ) | ( n5915 & n6131 ) | ( ~n6130 & n6131 ) ;
  assign n6133 = n1016 & n2725 ;
  assign n6134 = x97 & n1020 ;
  assign n6135 = x98 | n6134 ;
  assign n6136 = ( n1022 & n6134 ) | ( n1022 & n6135 ) | ( n6134 & n6135 ) ;
  assign n6137 = x96 & n1145 ;
  assign n6138 = n6136 | n6137 ;
  assign n6139 = ( x20 & n6133 ) | ( x20 & ~n6138 ) | ( n6133 & ~n6138 ) ;
  assign n6140 = ( ~x20 & n6138 ) | ( ~x20 & n6139 ) | ( n6138 & n6139 ) ;
  assign n6141 = ( ~n6133 & n6139 ) | ( ~n6133 & n6140 ) | ( n6139 & n6140 ) ;
  assign n6142 = ( n5927 & n6132 ) | ( n5927 & n6141 ) | ( n6132 & n6141 ) ;
  assign n6143 = ( ~n5927 & n6132 ) | ( ~n5927 & n6141 ) | ( n6132 & n6141 ) ;
  assign n6144 = ( n5927 & ~n6142 ) | ( n5927 & n6143 ) | ( ~n6142 & n6143 ) ;
  assign n6145 = n810 & n3326 ;
  assign n6146 = x100 & n814 ;
  assign n6147 = x101 | n6146 ;
  assign n6148 = ( n816 & n6146 ) | ( n816 & n6147 ) | ( n6146 & n6147 ) ;
  assign n6149 = x99 & n885 ;
  assign n6150 = n6148 | n6149 ;
  assign n6151 = ( x17 & n6145 ) | ( x17 & ~n6150 ) | ( n6145 & ~n6150 ) ;
  assign n6152 = ( ~x17 & n6150 ) | ( ~x17 & n6151 ) | ( n6150 & n6151 ) ;
  assign n6153 = ( ~n6145 & n6151 ) | ( ~n6145 & n6152 ) | ( n6151 & n6152 ) ;
  assign n6154 = ( n5930 & n6144 ) | ( n5930 & n6153 ) | ( n6144 & n6153 ) ;
  assign n6155 = ( ~n5930 & n6144 ) | ( ~n5930 & n6153 ) | ( n6144 & n6153 ) ;
  assign n6156 = ( n5930 & ~n6154 ) | ( n5930 & n6155 ) | ( ~n6154 & n6155 ) ;
  assign n6157 = n583 & n3665 ;
  assign n6158 = x103 & n587 ;
  assign n6159 = x104 | n6158 ;
  assign n6160 = ( n589 & n6158 ) | ( n589 & n6159 ) | ( n6158 & n6159 ) ;
  assign n6161 = x102 & n676 ;
  assign n6162 = n6160 | n6161 ;
  assign n6163 = ( x14 & n6157 ) | ( x14 & ~n6162 ) | ( n6157 & ~n6162 ) ;
  assign n6164 = ( ~x14 & n6162 ) | ( ~x14 & n6163 ) | ( n6162 & n6163 ) ;
  assign n6165 = ( ~n6157 & n6163 ) | ( ~n6157 & n6164 ) | ( n6163 & n6164 ) ;
  assign n6166 = ( n5942 & n6156 ) | ( n5942 & n6165 ) | ( n6156 & n6165 ) ;
  assign n6167 = ( ~n5942 & n6156 ) | ( ~n5942 & n6165 ) | ( n6156 & n6165 ) ;
  assign n6168 = ( n5942 & ~n6166 ) | ( n5942 & n6167 ) | ( ~n6166 & n6167 ) ;
  assign n6169 = n407 & n4362 ;
  assign n6170 = x106 & n411 ;
  assign n6171 = x107 | n6170 ;
  assign n6172 = ( n413 & n6170 ) | ( n413 & n6171 ) | ( n6170 & n6171 ) ;
  assign n6173 = x105 & n491 ;
  assign n6174 = n6172 | n6173 ;
  assign n6175 = ( x11 & n6169 ) | ( x11 & ~n6174 ) | ( n6169 & ~n6174 ) ;
  assign n6176 = ( ~x11 & n6174 ) | ( ~x11 & n6175 ) | ( n6174 & n6175 ) ;
  assign n6177 = ( ~n6169 & n6175 ) | ( ~n6169 & n6176 ) | ( n6175 & n6176 ) ;
  assign n6178 = ( n5954 & n6168 ) | ( n5954 & n6177 ) | ( n6168 & n6177 ) ;
  assign n6179 = ( ~n5954 & n6168 ) | ( ~n5954 & n6177 ) | ( n6168 & n6177 ) ;
  assign n6180 = ( n5954 & ~n6178 ) | ( n5954 & n6179 ) | ( ~n6178 & n6179 ) ;
  assign n6181 = ( n5966 & n5995 ) | ( n5966 & n6180 ) | ( n5995 & n6180 ) ;
  assign n6182 = ( ~n5966 & n5995 ) | ( ~n5966 & n6180 ) | ( n5995 & n6180 ) ;
  assign n6183 = ( n5966 & ~n6181 ) | ( n5966 & n6182 ) | ( ~n6181 & n6182 ) ;
  assign n6184 = n186 & n5542 ;
  assign n6185 = x112 & n190 ;
  assign n6186 = x113 | n6185 ;
  assign n6187 = ( n192 & n6185 ) | ( n192 & n6186 ) | ( n6185 & n6186 ) ;
  assign n6188 = x111 & n220 ;
  assign n6189 = n6187 | n6188 ;
  assign n6190 = ( x5 & n6184 ) | ( x5 & ~n6189 ) | ( n6184 & ~n6189 ) ;
  assign n6191 = ( ~x5 & n6189 ) | ( ~x5 & n6190 ) | ( n6189 & n6190 ) ;
  assign n6192 = ( ~n6184 & n6190 ) | ( ~n6184 & n6191 ) | ( n6190 & n6191 ) ;
  assign n6193 = ( n5969 & n6183 ) | ( n5969 & n6192 ) | ( n6183 & n6192 ) ;
  assign n6194 = ( ~n5969 & n6183 ) | ( ~n5969 & n6192 ) | ( n6183 & n6192 ) ;
  assign n6195 = ( n5969 & ~n6193 ) | ( n5969 & n6194 ) | ( ~n6193 & n6194 ) ;
  assign n6196 = ( n5972 & n5986 ) | ( n5972 & n6195 ) | ( n5986 & n6195 ) ;
  assign n6197 = ( ~n5972 & n5986 ) | ( ~n5972 & n6195 ) | ( n5986 & n6195 ) ;
  assign n6198 = ( n5972 & ~n6196 ) | ( n5972 & n6197 ) | ( ~n6196 & n6197 ) ;
  assign n6199 = ( x116 & x117 ) | ( x116 & n5975 ) | ( x117 & n5975 ) ;
  assign n6200 = ( x116 & ~x117 ) | ( x116 & n5975 ) | ( ~x117 & n5975 ) ;
  assign n6201 = ( x117 & ~n6199 ) | ( x117 & n6200 ) | ( ~n6199 & n6200 ) ;
  assign n6202 = n136 & n6201 ;
  assign n6203 = x116 & n138 ;
  assign n6204 = x117 | n6203 ;
  assign n6205 = ( n141 & n6203 ) | ( n141 & n6204 ) | ( n6203 & n6204 ) ;
  assign n6206 = x115 & n154 ;
  assign n6207 = n6205 | n6206 ;
  assign n6208 = ( x2 & n6202 ) | ( x2 & ~n6207 ) | ( n6202 & ~n6207 ) ;
  assign n6209 = ( ~x2 & n6207 ) | ( ~x2 & n6208 ) | ( n6207 & n6208 ) ;
  assign n6210 = ( ~n6202 & n6208 ) | ( ~n6202 & n6209 ) | ( n6208 & n6209 ) ;
  assign n6211 = n291 & n5130 ;
  assign n6212 = x110 & n295 ;
  assign n6213 = x111 | n6212 ;
  assign n6214 = ( n297 & n6212 ) | ( n297 & n6213 ) | ( n6212 & n6213 ) ;
  assign n6215 = x109 & n330 ;
  assign n6216 = n6214 | n6215 ;
  assign n6217 = ( x8 & n6211 ) | ( x8 & ~n6216 ) | ( n6211 & ~n6216 ) ;
  assign n6218 = ( ~x8 & n6216 ) | ( ~x8 & n6217 ) | ( n6216 & n6217 ) ;
  assign n6219 = ( ~n6211 & n6217 ) | ( ~n6211 & n6218 ) | ( n6217 & n6218 ) ;
  assign n6220 = n1297 & n2449 ;
  assign n6221 = x95 & n1301 ;
  assign n6222 = x96 | n6221 ;
  assign n6223 = ( n1303 & n6221 ) | ( n1303 & n6222 ) | ( n6221 & n6222 ) ;
  assign n6224 = x94 & n1426 ;
  assign n6225 = n6223 | n6224 ;
  assign n6226 = ( x23 & n6220 ) | ( x23 & ~n6225 ) | ( n6220 & ~n6225 ) ;
  assign n6227 = ( ~x23 & n6225 ) | ( ~x23 & n6226 ) | ( n6225 & n6226 ) ;
  assign n6228 = ( ~n6220 & n6226 ) | ( ~n6220 & n6227 ) | ( n6226 & n6227 ) ;
  assign n6229 = n1617 & n2057 ;
  assign n6230 = x92 & n1621 ;
  assign n6231 = x93 | n6230 ;
  assign n6232 = ( n1623 & n6230 ) | ( n1623 & n6231 ) | ( n6230 & n6231 ) ;
  assign n6233 = x91 & n1749 ;
  assign n6234 = n6232 | n6233 ;
  assign n6235 = ( x26 & n6229 ) | ( x26 & ~n6234 ) | ( n6229 & ~n6234 ) ;
  assign n6236 = ( ~x26 & n6234 ) | ( ~x26 & n6235 ) | ( n6234 & n6235 ) ;
  assign n6237 = ( ~n6229 & n6235 ) | ( ~n6229 & n6236 ) | ( n6235 & n6236 ) ;
  assign n6238 = n1701 & n1949 ;
  assign n6239 = x89 & n1953 ;
  assign n6240 = x90 | n6239 ;
  assign n6241 = ( n1955 & n6239 ) | ( n1955 & n6240 ) | ( n6239 & n6240 ) ;
  assign n6242 = x88 & n2114 ;
  assign n6243 = n6241 | n6242 ;
  assign n6244 = ( x29 & n6238 ) | ( x29 & ~n6243 ) | ( n6238 & ~n6243 ) ;
  assign n6245 = ( ~x29 & n6243 ) | ( ~x29 & n6244 ) | ( n6243 & n6244 ) ;
  assign n6246 = ( ~n6238 & n6244 ) | ( ~n6238 & n6245 ) | ( n6244 & n6245 ) ;
  assign n6247 = n1466 & n2320 ;
  assign n6248 = x86 & n2324 ;
  assign n6249 = x87 | n6248 ;
  assign n6250 = ( n2326 & n6248 ) | ( n2326 & n6249 ) | ( n6248 & n6249 ) ;
  assign n6251 = x85 & n2497 ;
  assign n6252 = n6250 | n6251 ;
  assign n6253 = ( x32 & n6247 ) | ( x32 & ~n6252 ) | ( n6247 & ~n6252 ) ;
  assign n6254 = ( ~x32 & n6252 ) | ( ~x32 & n6253 ) | ( n6252 & n6253 ) ;
  assign n6255 = ( ~n6247 & n6253 ) | ( ~n6247 & n6254 ) | ( n6253 & n6254 ) ;
  assign n6256 = n1097 & n2766 ;
  assign n6257 = x83 & n2770 ;
  assign n6258 = x84 | n6257 ;
  assign n6259 = ( n2772 & n6257 ) | ( n2772 & n6258 ) | ( n6257 & n6258 ) ;
  assign n6260 = x82 & n2943 ;
  assign n6261 = n6259 | n6260 ;
  assign n6262 = ( x35 & n6256 ) | ( x35 & ~n6261 ) | ( n6256 & ~n6261 ) ;
  assign n6263 = ( ~x35 & n6261 ) | ( ~x35 & n6262 ) | ( n6261 & n6262 ) ;
  assign n6264 = ( ~n6256 & n6262 ) | ( ~n6256 & n6263 ) | ( n6262 & n6263 ) ;
  assign n6265 = n910 & n3224 ;
  assign n6266 = x80 & n3228 ;
  assign n6267 = x81 | n6266 ;
  assign n6268 = ( n3230 & n6266 ) | ( n3230 & n6267 ) | ( n6266 & n6267 ) ;
  assign n6269 = x79 & n3413 ;
  assign n6270 = n6268 | n6269 ;
  assign n6271 = ( x38 & n6265 ) | ( x38 & ~n6270 ) | ( n6265 & ~n6270 ) ;
  assign n6272 = ( ~x38 & n6270 ) | ( ~x38 & n6271 ) | ( n6270 & n6271 ) ;
  assign n6273 = ( ~n6265 & n6271 ) | ( ~n6265 & n6272 ) | ( n6271 & n6272 ) ;
  assign n6274 = n461 & n4227 ;
  assign n6275 = x74 & n4231 ;
  assign n6276 = x75 | n6275 ;
  assign n6277 = ( n4233 & n6275 ) | ( n4233 & n6276 ) | ( n6275 & n6276 ) ;
  assign n6278 = x73 & n4470 ;
  assign n6279 = n6277 | n6278 ;
  assign n6280 = ( x44 & n6274 ) | ( x44 & ~n6279 ) | ( n6274 & ~n6279 ) ;
  assign n6281 = ( ~x44 & n6279 ) | ( ~x44 & n6280 ) | ( n6279 & n6280 ) ;
  assign n6282 = ( ~n6274 & n6280 ) | ( ~n6274 & n6281 ) | ( n6280 & n6281 ) ;
  assign n6283 = n346 & n4787 ;
  assign n6284 = x71 & n4791 ;
  assign n6285 = x72 | n6284 ;
  assign n6286 = ( n4793 & n6284 ) | ( n4793 & n6285 ) | ( n6284 & n6285 ) ;
  assign n6287 = x70 & n5030 ;
  assign n6288 = n6286 | n6287 ;
  assign n6289 = ( x47 & n6283 ) | ( x47 & ~n6288 ) | ( n6283 & ~n6288 ) ;
  assign n6290 = ( ~x47 & n6288 ) | ( ~x47 & n6289 ) | ( n6288 & n6289 ) ;
  assign n6291 = ( ~n6283 & n6289 ) | ( ~n6283 & n6290 ) | ( n6289 & n6290 ) ;
  assign n6292 = n230 & n5374 ;
  assign n6293 = x68 & n5378 ;
  assign n6294 = x69 | n6293 ;
  assign n6295 = ( n5380 & n6293 ) | ( n5380 & n6294 ) | ( n6293 & n6294 ) ;
  assign n6296 = x67 & n5638 ;
  assign n6297 = n6295 | n6296 ;
  assign n6298 = ( ~x50 & n6292 ) | ( ~x50 & n6297 ) | ( n6292 & n6297 ) ;
  assign n6299 = ( n6292 & n6297 ) | ( n6292 & ~n6298 ) | ( n6297 & ~n6298 ) ;
  assign n6300 = ( x50 & n6298 ) | ( x50 & ~n6299 ) | ( n6298 & ~n6299 ) ;
  assign n6301 = ( x53 & n6023 ) | ( x53 & n6037 ) | ( n6023 & n6037 ) ;
  assign n6302 = ( x50 & ~x52 ) | ( x50 & n6026 ) | ( ~x52 & n6026 ) ;
  assign n6303 = ( ~n5839 & n6030 ) | ( ~n5839 & n6302 ) | ( n6030 & n6302 ) ;
  assign n6304 = x64 & n6303 ;
  assign n6305 = x65 & n6031 ;
  assign n6306 = x66 | n6305 ;
  assign n6307 = ( n6033 & n6305 ) | ( n6033 & n6306 ) | ( n6305 & n6306 ) ;
  assign n6308 = ( n151 & n152 ) | ( n151 & n6027 ) | ( n152 & n6027 ) ;
  assign n6309 = ( ~n6304 & n6307 ) | ( ~n6304 & n6308 ) | ( n6307 & n6308 ) ;
  assign n6310 = n6304 | n6309 ;
  assign n6311 = n6301 | n6310 ;
  assign n6312 = ( n6301 & n6310 ) | ( n6301 & ~n6311 ) | ( n6310 & ~n6311 ) ;
  assign n6313 = n6311 & ~n6312 ;
  assign n6314 = ( n6049 & n6300 ) | ( n6049 & n6313 ) | ( n6300 & n6313 ) ;
  assign n6315 = ( ~n6049 & n6300 ) | ( ~n6049 & n6313 ) | ( n6300 & n6313 ) ;
  assign n6316 = ( n6049 & ~n6314 ) | ( n6049 & n6315 ) | ( ~n6314 & n6315 ) ;
  assign n6317 = ( n6061 & n6291 ) | ( n6061 & n6316 ) | ( n6291 & n6316 ) ;
  assign n6318 = ( ~n6061 & n6291 ) | ( ~n6061 & n6316 ) | ( n6291 & n6316 ) ;
  assign n6319 = ( n6061 & ~n6317 ) | ( n6061 & n6318 ) | ( ~n6317 & n6318 ) ;
  assign n6320 = ( n6073 & n6282 ) | ( n6073 & n6319 ) | ( n6282 & n6319 ) ;
  assign n6321 = ( ~n6073 & n6282 ) | ( ~n6073 & n6319 ) | ( n6282 & n6319 ) ;
  assign n6322 = ( n6073 & ~n6320 ) | ( n6073 & n6321 ) | ( ~n6320 & n6321 ) ;
  assign n6323 = n637 & n3715 ;
  assign n6324 = x77 & n3719 ;
  assign n6325 = x78 | n6324 ;
  assign n6326 = ( n3721 & n6324 ) | ( n3721 & n6325 ) | ( n6324 & n6325 ) ;
  assign n6327 = x76 & n3922 ;
  assign n6328 = n6326 | n6327 ;
  assign n6329 = ( x41 & n6323 ) | ( x41 & ~n6328 ) | ( n6323 & ~n6328 ) ;
  assign n6330 = ( ~x41 & n6328 ) | ( ~x41 & n6329 ) | ( n6328 & n6329 ) ;
  assign n6331 = ( ~n6323 & n6329 ) | ( ~n6323 & n6330 ) | ( n6329 & n6330 ) ;
  assign n6332 = ( n6076 & n6322 ) | ( n6076 & n6331 ) | ( n6322 & n6331 ) ;
  assign n6333 = ( ~n6076 & n6322 ) | ( ~n6076 & n6331 ) | ( n6322 & n6331 ) ;
  assign n6334 = ( n6076 & ~n6332 ) | ( n6076 & n6333 ) | ( ~n6332 & n6333 ) ;
  assign n6335 = ( n6088 & n6273 ) | ( n6088 & n6334 ) | ( n6273 & n6334 ) ;
  assign n6336 = ( ~n6088 & n6273 ) | ( ~n6088 & n6334 ) | ( n6273 & n6334 ) ;
  assign n6337 = ( n6088 & ~n6335 ) | ( n6088 & n6336 ) | ( ~n6335 & n6336 ) ;
  assign n6338 = ( n6100 & n6264 ) | ( n6100 & n6337 ) | ( n6264 & n6337 ) ;
  assign n6339 = ( ~n6100 & n6264 ) | ( ~n6100 & n6337 ) | ( n6264 & n6337 ) ;
  assign n6340 = ( n6100 & ~n6338 ) | ( n6100 & n6339 ) | ( ~n6338 & n6339 ) ;
  assign n6341 = ( n6103 & n6255 ) | ( n6103 & n6340 ) | ( n6255 & n6340 ) ;
  assign n6342 = ( ~n6103 & n6255 ) | ( ~n6103 & n6340 ) | ( n6255 & n6340 ) ;
  assign n6343 = ( n6103 & ~n6341 ) | ( n6103 & n6342 ) | ( ~n6341 & n6342 ) ;
  assign n6344 = ( n6115 & n6246 ) | ( n6115 & n6343 ) | ( n6246 & n6343 ) ;
  assign n6345 = ( ~n6115 & n6246 ) | ( ~n6115 & n6343 ) | ( n6246 & n6343 ) ;
  assign n6346 = ( n6115 & ~n6344 ) | ( n6115 & n6345 ) | ( ~n6344 & n6345 ) ;
  assign n6347 = ( n6118 & n6237 ) | ( n6118 & n6346 ) | ( n6237 & n6346 ) ;
  assign n6348 = ( ~n6118 & n6237 ) | ( ~n6118 & n6346 ) | ( n6237 & n6346 ) ;
  assign n6349 = ( n6118 & ~n6347 ) | ( n6118 & n6348 ) | ( ~n6347 & n6348 ) ;
  assign n6350 = ( n6130 & n6228 ) | ( n6130 & n6349 ) | ( n6228 & n6349 ) ;
  assign n6351 = ( ~n6130 & n6228 ) | ( ~n6130 & n6349 ) | ( n6228 & n6349 ) ;
  assign n6352 = ( n6130 & ~n6350 ) | ( n6130 & n6351 ) | ( ~n6350 & n6351 ) ;
  assign n6353 = n1016 & n2877 ;
  assign n6354 = x98 & n1020 ;
  assign n6355 = x99 | n6354 ;
  assign n6356 = ( n1022 & n6354 ) | ( n1022 & n6355 ) | ( n6354 & n6355 ) ;
  assign n6357 = x97 & n1145 ;
  assign n6358 = n6356 | n6357 ;
  assign n6359 = ( x20 & n6353 ) | ( x20 & ~n6358 ) | ( n6353 & ~n6358 ) ;
  assign n6360 = ( ~x20 & n6358 ) | ( ~x20 & n6359 ) | ( n6358 & n6359 ) ;
  assign n6361 = ( ~n6353 & n6359 ) | ( ~n6353 & n6360 ) | ( n6359 & n6360 ) ;
  assign n6362 = ( n6142 & n6352 ) | ( n6142 & n6361 ) | ( n6352 & n6361 ) ;
  assign n6363 = ( ~n6142 & n6352 ) | ( ~n6142 & n6361 ) | ( n6352 & n6361 ) ;
  assign n6364 = ( n6142 & ~n6362 ) | ( n6142 & n6363 ) | ( ~n6362 & n6363 ) ;
  assign n6365 = n810 & n3486 ;
  assign n6366 = x101 & n814 ;
  assign n6367 = x102 | n6366 ;
  assign n6368 = ( n816 & n6366 ) | ( n816 & n6367 ) | ( n6366 & n6367 ) ;
  assign n6369 = x100 & n885 ;
  assign n6370 = n6368 | n6369 ;
  assign n6371 = ( x17 & n6365 ) | ( x17 & ~n6370 ) | ( n6365 & ~n6370 ) ;
  assign n6372 = ( ~x17 & n6370 ) | ( ~x17 & n6371 ) | ( n6370 & n6371 ) ;
  assign n6373 = ( ~n6365 & n6371 ) | ( ~n6365 & n6372 ) | ( n6371 & n6372 ) ;
  assign n6374 = ( n6154 & n6364 ) | ( n6154 & n6373 ) | ( n6364 & n6373 ) ;
  assign n6375 = ( ~n6154 & n6364 ) | ( ~n6154 & n6373 ) | ( n6364 & n6373 ) ;
  assign n6376 = ( n6154 & ~n6374 ) | ( n6154 & n6375 ) | ( ~n6374 & n6375 ) ;
  assign n6377 = n583 & n3998 ;
  assign n6378 = x104 & n587 ;
  assign n6379 = x105 | n6378 ;
  assign n6380 = ( n589 & n6378 ) | ( n589 & n6379 ) | ( n6378 & n6379 ) ;
  assign n6381 = x103 & n676 ;
  assign n6382 = n6380 | n6381 ;
  assign n6383 = ( x14 & n6377 ) | ( x14 & ~n6382 ) | ( n6377 & ~n6382 ) ;
  assign n6384 = ( ~x14 & n6382 ) | ( ~x14 & n6383 ) | ( n6382 & n6383 ) ;
  assign n6385 = ( ~n6377 & n6383 ) | ( ~n6377 & n6384 ) | ( n6383 & n6384 ) ;
  assign n6386 = ( n6166 & n6376 ) | ( n6166 & n6385 ) | ( n6376 & n6385 ) ;
  assign n6387 = ( ~n6166 & n6376 ) | ( ~n6166 & n6385 ) | ( n6376 & n6385 ) ;
  assign n6388 = ( n6166 & ~n6386 ) | ( n6166 & n6387 ) | ( ~n6386 & n6387 ) ;
  assign n6389 = n407 & n4377 ;
  assign n6390 = x107 & n411 ;
  assign n6391 = x108 | n6390 ;
  assign n6392 = ( n413 & n6390 ) | ( n413 & n6391 ) | ( n6390 & n6391 ) ;
  assign n6393 = x106 & n491 ;
  assign n6394 = n6392 | n6393 ;
  assign n6395 = ( x11 & n6389 ) | ( x11 & ~n6394 ) | ( n6389 & ~n6394 ) ;
  assign n6396 = ( ~x11 & n6394 ) | ( ~x11 & n6395 ) | ( n6394 & n6395 ) ;
  assign n6397 = ( ~n6389 & n6395 ) | ( ~n6389 & n6396 ) | ( n6395 & n6396 ) ;
  assign n6398 = ( n6178 & n6388 ) | ( n6178 & n6397 ) | ( n6388 & n6397 ) ;
  assign n6399 = ( ~n6178 & n6388 ) | ( ~n6178 & n6397 ) | ( n6388 & n6397 ) ;
  assign n6400 = ( n6178 & ~n6398 ) | ( n6178 & n6399 ) | ( ~n6398 & n6399 ) ;
  assign n6401 = ( n6181 & n6219 ) | ( n6181 & n6400 ) | ( n6219 & n6400 ) ;
  assign n6402 = ( ~n6181 & n6219 ) | ( ~n6181 & n6400 ) | ( n6219 & n6400 ) ;
  assign n6403 = ( n6181 & ~n6401 ) | ( n6181 & n6402 ) | ( ~n6401 & n6402 ) ;
  assign n6404 = n186 & n5750 ;
  assign n6405 = x113 & n190 ;
  assign n6406 = x114 | n6405 ;
  assign n6407 = ( n192 & n6405 ) | ( n192 & n6406 ) | ( n6405 & n6406 ) ;
  assign n6408 = x112 & n220 ;
  assign n6409 = n6407 | n6408 ;
  assign n6410 = ( x5 & n6404 ) | ( x5 & ~n6409 ) | ( n6404 & ~n6409 ) ;
  assign n6411 = ( ~x5 & n6409 ) | ( ~x5 & n6410 ) | ( n6409 & n6410 ) ;
  assign n6412 = ( ~n6404 & n6410 ) | ( ~n6404 & n6411 ) | ( n6410 & n6411 ) ;
  assign n6413 = ( n6193 & n6403 ) | ( n6193 & n6412 ) | ( n6403 & n6412 ) ;
  assign n6414 = ( ~n6193 & n6403 ) | ( ~n6193 & n6412 ) | ( n6403 & n6412 ) ;
  assign n6415 = ( n6193 & ~n6413 ) | ( n6193 & n6414 ) | ( ~n6413 & n6414 ) ;
  assign n6416 = ( n6196 & n6210 ) | ( n6196 & n6415 ) | ( n6210 & n6415 ) ;
  assign n6417 = ( ~n6196 & n6210 ) | ( ~n6196 & n6415 ) | ( n6210 & n6415 ) ;
  assign n6418 = ( n6196 & ~n6416 ) | ( n6196 & n6417 ) | ( ~n6416 & n6417 ) ;
  assign n6419 = ( x117 & x118 ) | ( x117 & n6199 ) | ( x118 & n6199 ) ;
  assign n6420 = ( x117 & ~x118 ) | ( x117 & n6199 ) | ( ~x118 & n6199 ) ;
  assign n6421 = ( x118 & ~n6419 ) | ( x118 & n6420 ) | ( ~n6419 & n6420 ) ;
  assign n6422 = n136 & n6421 ;
  assign n6423 = x117 & n138 ;
  assign n6424 = x118 | n6423 ;
  assign n6425 = ( n141 & n6423 ) | ( n141 & n6424 ) | ( n6423 & n6424 ) ;
  assign n6426 = x116 & n154 ;
  assign n6427 = n6425 | n6426 ;
  assign n6428 = ( x2 & n6422 ) | ( x2 & ~n6427 ) | ( n6422 & ~n6427 ) ;
  assign n6429 = ( ~x2 & n6427 ) | ( ~x2 & n6428 ) | ( n6427 & n6428 ) ;
  assign n6430 = ( ~n6422 & n6428 ) | ( ~n6422 & n6429 ) | ( n6428 & n6429 ) ;
  assign n6431 = n291 & n5145 ;
  assign n6432 = x111 & n295 ;
  assign n6433 = x112 | n6432 ;
  assign n6434 = ( n297 & n6432 ) | ( n297 & n6433 ) | ( n6432 & n6433 ) ;
  assign n6435 = x110 & n330 ;
  assign n6436 = n6434 | n6435 ;
  assign n6437 = ( x8 & n6431 ) | ( x8 & ~n6436 ) | ( n6431 & ~n6436 ) ;
  assign n6438 = ( ~x8 & n6436 ) | ( ~x8 & n6437 ) | ( n6436 & n6437 ) ;
  assign n6439 = ( ~n6431 & n6437 ) | ( ~n6431 & n6438 ) | ( n6437 & n6438 ) ;
  assign n6440 = n407 & n4734 ;
  assign n6441 = x108 & n411 ;
  assign n6442 = x109 | n6441 ;
  assign n6443 = ( n413 & n6441 ) | ( n413 & n6442 ) | ( n6441 & n6442 ) ;
  assign n6444 = x107 & n491 ;
  assign n6445 = n6443 | n6444 ;
  assign n6446 = ( x11 & n6440 ) | ( x11 & ~n6445 ) | ( n6440 & ~n6445 ) ;
  assign n6447 = ( ~x11 & n6445 ) | ( ~x11 & n6446 ) | ( n6445 & n6446 ) ;
  assign n6448 = ( ~n6440 & n6446 ) | ( ~n6440 & n6447 ) | ( n6446 & n6447 ) ;
  assign n6449 = n1016 & n3162 ;
  assign n6450 = x99 & n1020 ;
  assign n6451 = x100 | n6450 ;
  assign n6452 = ( n1022 & n6450 ) | ( n1022 & n6451 ) | ( n6450 & n6451 ) ;
  assign n6453 = x98 & n1145 ;
  assign n6454 = n6452 | n6453 ;
  assign n6455 = ( x20 & n6449 ) | ( x20 & ~n6454 ) | ( n6449 & ~n6454 ) ;
  assign n6456 = ( ~x20 & n6454 ) | ( ~x20 & n6455 ) | ( n6454 & n6455 ) ;
  assign n6457 = ( ~n6449 & n6455 ) | ( ~n6449 & n6456 ) | ( n6455 & n6456 ) ;
  assign n6458 = n1617 & n2294 ;
  assign n6459 = x93 & n1621 ;
  assign n6460 = x94 | n6459 ;
  assign n6461 = ( n1623 & n6459 ) | ( n1623 & n6460 ) | ( n6459 & n6460 ) ;
  assign n6462 = x92 & n1749 ;
  assign n6463 = n6461 | n6462 ;
  assign n6464 = ( x26 & n6458 ) | ( x26 & ~n6463 ) | ( n6458 & ~n6463 ) ;
  assign n6465 = ( ~x26 & n6463 ) | ( ~x26 & n6464 ) | ( n6463 & n6464 ) ;
  assign n6466 = ( ~n6458 & n6464 ) | ( ~n6458 & n6465 ) | ( n6464 & n6465 ) ;
  assign n6467 = n1914 & n1949 ;
  assign n6468 = x90 & n1953 ;
  assign n6469 = x91 | n6468 ;
  assign n6470 = ( n1955 & n6468 ) | ( n1955 & n6469 ) | ( n6468 & n6469 ) ;
  assign n6471 = x89 & n2114 ;
  assign n6472 = n6470 | n6471 ;
  assign n6473 = ( x29 & n6467 ) | ( x29 & ~n6472 ) | ( n6467 & ~n6472 ) ;
  assign n6474 = ( ~x29 & n6472 ) | ( ~x29 & n6473 ) | ( n6472 & n6473 ) ;
  assign n6475 = ( ~n6467 & n6473 ) | ( ~n6467 & n6474 ) | ( n6473 & n6474 ) ;
  assign n6476 = n1481 & n2320 ;
  assign n6477 = x87 & n2324 ;
  assign n6478 = x88 | n6477 ;
  assign n6479 = ( n2326 & n6477 ) | ( n2326 & n6478 ) | ( n6477 & n6478 ) ;
  assign n6480 = x86 & n2497 ;
  assign n6481 = n6479 | n6480 ;
  assign n6482 = ( x32 & n6476 ) | ( x32 & ~n6481 ) | ( n6476 & ~n6481 ) ;
  assign n6483 = ( ~x32 & n6481 ) | ( ~x32 & n6482 ) | ( n6481 & n6482 ) ;
  assign n6484 = ( ~n6476 & n6482 ) | ( ~n6476 & n6483 ) | ( n6482 & n6483 ) ;
  assign n6485 = n1262 & n2766 ;
  assign n6486 = x84 & n2770 ;
  assign n6487 = x85 | n6486 ;
  assign n6488 = ( n2772 & n6486 ) | ( n2772 & n6487 ) | ( n6486 & n6487 ) ;
  assign n6489 = x83 & n2943 ;
  assign n6490 = n6488 | n6489 ;
  assign n6491 = ( x35 & n6485 ) | ( x35 & ~n6490 ) | ( n6485 & ~n6490 ) ;
  assign n6492 = ( ~x35 & n6490 ) | ( ~x35 & n6491 ) | ( n6490 & n6491 ) ;
  assign n6493 = ( ~n6485 & n6491 ) | ( ~n6485 & n6492 ) | ( n6491 & n6492 ) ;
  assign n6494 = n990 & n3224 ;
  assign n6495 = x81 & n3228 ;
  assign n6496 = x82 | n6495 ;
  assign n6497 = ( n3230 & n6495 ) | ( n3230 & n6496 ) | ( n6495 & n6496 ) ;
  assign n6498 = x80 & n3413 ;
  assign n6499 = n6497 | n6498 ;
  assign n6500 = ( x38 & n6494 ) | ( x38 & ~n6499 ) | ( n6494 & ~n6499 ) ;
  assign n6501 = ( ~x38 & n6499 ) | ( ~x38 & n6500 ) | ( n6499 & n6500 ) ;
  assign n6502 = ( ~n6494 & n6500 ) | ( ~n6494 & n6501 ) | ( n6500 & n6501 ) ;
  assign n6503 = n701 & n3715 ;
  assign n6504 = x78 & n3719 ;
  assign n6505 = x79 | n6504 ;
  assign n6506 = ( n3721 & n6504 ) | ( n3721 & n6505 ) | ( n6504 & n6505 ) ;
  assign n6507 = x77 & n3922 ;
  assign n6508 = n6506 | n6507 ;
  assign n6509 = ( x41 & n6503 ) | ( x41 & ~n6508 ) | ( n6503 & ~n6508 ) ;
  assign n6510 = ( ~x41 & n6508 ) | ( ~x41 & n6509 ) | ( n6508 & n6509 ) ;
  assign n6511 = ( ~n6503 & n6509 ) | ( ~n6503 & n6510 ) | ( n6509 & n6510 ) ;
  assign n6512 = n554 & n4227 ;
  assign n6513 = x75 & n4231 ;
  assign n6514 = x76 | n6513 ;
  assign n6515 = ( n4233 & n6513 ) | ( n4233 & n6514 ) | ( n6513 & n6514 ) ;
  assign n6516 = x74 & n4470 ;
  assign n6517 = n6515 | n6516 ;
  assign n6518 = ( x44 & n6512 ) | ( x44 & ~n6517 ) | ( n6512 & ~n6517 ) ;
  assign n6519 = ( ~x44 & n6517 ) | ( ~x44 & n6518 ) | ( n6517 & n6518 ) ;
  assign n6520 = ( ~n6512 & n6518 ) | ( ~n6512 & n6519 ) | ( n6518 & n6519 ) ;
  assign n6521 = n390 & n4787 ;
  assign n6522 = x72 & n4791 ;
  assign n6523 = x73 | n6522 ;
  assign n6524 = ( n4793 & n6522 ) | ( n4793 & n6523 ) | ( n6522 & n6523 ) ;
  assign n6525 = x71 & n5030 ;
  assign n6526 = n6524 | n6525 ;
  assign n6527 = ( x47 & n6521 ) | ( x47 & ~n6526 ) | ( n6521 & ~n6526 ) ;
  assign n6528 = ( ~x47 & n6526 ) | ( ~x47 & n6527 ) | ( n6526 & n6527 ) ;
  assign n6529 = ( ~n6521 & n6527 ) | ( ~n6521 & n6528 ) | ( n6527 & n6528 ) ;
  assign n6530 = x66 & n6031 ;
  assign n6531 = x67 | n6530 ;
  assign n6532 = ( n6033 & n6530 ) | ( n6033 & n6531 ) | ( n6530 & n6531 ) ;
  assign n6533 = x65 & n6303 ;
  assign n6534 = n6532 | n6533 ;
  assign n6535 = n164 & n6027 ;
  assign n6536 = ( x53 & n6534 ) | ( x53 & ~n6535 ) | ( n6534 & ~n6535 ) ;
  assign n6537 = ( ~x53 & n6535 ) | ( ~x53 & n6536 ) | ( n6535 & n6536 ) ;
  assign n6538 = ( ~n6534 & n6536 ) | ( ~n6534 & n6537 ) | ( n6536 & n6537 ) ;
  assign n6539 = x53 & x54 ;
  assign n6540 = x53 | x54 ;
  assign n6541 = ~n6539 & n6540 ;
  assign n6542 = x64 & n6541 ;
  assign n6543 = x53 & ~n6311 ;
  assign n6544 = ( n6538 & n6542 ) | ( n6538 & n6543 ) | ( n6542 & n6543 ) ;
  assign n6545 = ( ~n6538 & n6542 ) | ( ~n6538 & n6543 ) | ( n6542 & n6543 ) ;
  assign n6546 = ( n6538 & ~n6544 ) | ( n6538 & n6545 ) | ( ~n6544 & n6545 ) ;
  assign n6547 = n245 & n5374 ;
  assign n6548 = x69 & n5378 ;
  assign n6549 = x70 | n6548 ;
  assign n6550 = ( n5380 & n6548 ) | ( n5380 & n6549 ) | ( n6548 & n6549 ) ;
  assign n6551 = x68 & n5638 ;
  assign n6552 = n6550 | n6551 ;
  assign n6553 = ( x50 & n6547 ) | ( x50 & ~n6552 ) | ( n6547 & ~n6552 ) ;
  assign n6554 = ( ~x50 & n6552 ) | ( ~x50 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6555 = ( ~n6547 & n6553 ) | ( ~n6547 & n6554 ) | ( n6553 & n6554 ) ;
  assign n6556 = ( n6314 & n6546 ) | ( n6314 & n6555 ) | ( n6546 & n6555 ) ;
  assign n6557 = ( ~n6314 & n6546 ) | ( ~n6314 & n6555 ) | ( n6546 & n6555 ) ;
  assign n6558 = ( n6314 & ~n6556 ) | ( n6314 & n6557 ) | ( ~n6556 & n6557 ) ;
  assign n6559 = ( n6317 & n6529 ) | ( n6317 & n6558 ) | ( n6529 & n6558 ) ;
  assign n6560 = ( ~n6317 & n6529 ) | ( ~n6317 & n6558 ) | ( n6529 & n6558 ) ;
  assign n6561 = ( n6317 & ~n6559 ) | ( n6317 & n6560 ) | ( ~n6559 & n6560 ) ;
  assign n6562 = ( n6320 & n6520 ) | ( n6320 & n6561 ) | ( n6520 & n6561 ) ;
  assign n6563 = ( ~n6320 & n6520 ) | ( ~n6320 & n6561 ) | ( n6520 & n6561 ) ;
  assign n6564 = ( n6320 & ~n6562 ) | ( n6320 & n6563 ) | ( ~n6562 & n6563 ) ;
  assign n6565 = ( n6332 & n6511 ) | ( n6332 & n6564 ) | ( n6511 & n6564 ) ;
  assign n6566 = ( ~n6332 & n6511 ) | ( ~n6332 & n6564 ) | ( n6511 & n6564 ) ;
  assign n6567 = ( n6332 & ~n6565 ) | ( n6332 & n6566 ) | ( ~n6565 & n6566 ) ;
  assign n6568 = ( n6335 & n6502 ) | ( n6335 & n6567 ) | ( n6502 & n6567 ) ;
  assign n6569 = ( ~n6335 & n6502 ) | ( ~n6335 & n6567 ) | ( n6502 & n6567 ) ;
  assign n6570 = ( n6335 & ~n6568 ) | ( n6335 & n6569 ) | ( ~n6568 & n6569 ) ;
  assign n6571 = ( n6338 & n6493 ) | ( n6338 & n6570 ) | ( n6493 & n6570 ) ;
  assign n6572 = ( ~n6338 & n6493 ) | ( ~n6338 & n6570 ) | ( n6493 & n6570 ) ;
  assign n6573 = ( n6338 & ~n6571 ) | ( n6338 & n6572 ) | ( ~n6571 & n6572 ) ;
  assign n6574 = ( n6341 & n6484 ) | ( n6341 & n6573 ) | ( n6484 & n6573 ) ;
  assign n6575 = ( ~n6341 & n6484 ) | ( ~n6341 & n6573 ) | ( n6484 & n6573 ) ;
  assign n6576 = ( n6341 & ~n6574 ) | ( n6341 & n6575 ) | ( ~n6574 & n6575 ) ;
  assign n6577 = ( n6344 & n6475 ) | ( n6344 & n6576 ) | ( n6475 & n6576 ) ;
  assign n6578 = ( ~n6344 & n6475 ) | ( ~n6344 & n6576 ) | ( n6475 & n6576 ) ;
  assign n6579 = ( n6344 & ~n6577 ) | ( n6344 & n6578 ) | ( ~n6577 & n6578 ) ;
  assign n6580 = ( n6347 & n6466 ) | ( n6347 & n6579 ) | ( n6466 & n6579 ) ;
  assign n6581 = ( ~n6347 & n6466 ) | ( ~n6347 & n6579 ) | ( n6466 & n6579 ) ;
  assign n6582 = ( n6347 & ~n6580 ) | ( n6347 & n6581 ) | ( ~n6580 & n6581 ) ;
  assign n6583 = n1297 & n2585 ;
  assign n6584 = x96 & n1301 ;
  assign n6585 = x97 | n6584 ;
  assign n6586 = ( n1303 & n6584 ) | ( n1303 & n6585 ) | ( n6584 & n6585 ) ;
  assign n6587 = x95 & n1426 ;
  assign n6588 = n6586 | n6587 ;
  assign n6589 = ( x23 & n6583 ) | ( x23 & ~n6588 ) | ( n6583 & ~n6588 ) ;
  assign n6590 = ( ~x23 & n6588 ) | ( ~x23 & n6589 ) | ( n6588 & n6589 ) ;
  assign n6591 = ( ~n6583 & n6589 ) | ( ~n6583 & n6590 ) | ( n6589 & n6590 ) ;
  assign n6592 = ( n6350 & n6582 ) | ( n6350 & n6591 ) | ( n6582 & n6591 ) ;
  assign n6593 = ( ~n6350 & n6582 ) | ( ~n6350 & n6591 ) | ( n6582 & n6591 ) ;
  assign n6594 = ( n6350 & ~n6592 ) | ( n6350 & n6593 ) | ( ~n6592 & n6593 ) ;
  assign n6595 = ( n6362 & n6457 ) | ( n6362 & n6594 ) | ( n6457 & n6594 ) ;
  assign n6596 = ( ~n6362 & n6457 ) | ( ~n6362 & n6594 ) | ( n6457 & n6594 ) ;
  assign n6597 = ( n6362 & ~n6595 ) | ( n6362 & n6596 ) | ( ~n6595 & n6596 ) ;
  assign n6598 = n810 & n3650 ;
  assign n6599 = x102 & n814 ;
  assign n6600 = x103 | n6599 ;
  assign n6601 = ( n816 & n6599 ) | ( n816 & n6600 ) | ( n6599 & n6600 ) ;
  assign n6602 = x101 & n885 ;
  assign n6603 = n6601 | n6602 ;
  assign n6604 = ( x17 & n6598 ) | ( x17 & ~n6603 ) | ( n6598 & ~n6603 ) ;
  assign n6605 = ( ~x17 & n6603 ) | ( ~x17 & n6604 ) | ( n6603 & n6604 ) ;
  assign n6606 = ( ~n6598 & n6604 ) | ( ~n6598 & n6605 ) | ( n6604 & n6605 ) ;
  assign n6607 = ( n6374 & n6597 ) | ( n6374 & n6606 ) | ( n6597 & n6606 ) ;
  assign n6608 = ( ~n6374 & n6597 ) | ( ~n6374 & n6606 ) | ( n6597 & n6606 ) ;
  assign n6609 = ( n6374 & ~n6607 ) | ( n6374 & n6608 ) | ( ~n6607 & n6608 ) ;
  assign n6610 = n583 & n4013 ;
  assign n6611 = x105 & n587 ;
  assign n6612 = x106 | n6611 ;
  assign n6613 = ( n589 & n6611 ) | ( n589 & n6612 ) | ( n6611 & n6612 ) ;
  assign n6614 = x104 & n676 ;
  assign n6615 = n6613 | n6614 ;
  assign n6616 = ( x14 & n6610 ) | ( x14 & ~n6615 ) | ( n6610 & ~n6615 ) ;
  assign n6617 = ( ~x14 & n6615 ) | ( ~x14 & n6616 ) | ( n6615 & n6616 ) ;
  assign n6618 = ( ~n6610 & n6616 ) | ( ~n6610 & n6617 ) | ( n6616 & n6617 ) ;
  assign n6619 = ( n6386 & n6609 ) | ( n6386 & n6618 ) | ( n6609 & n6618 ) ;
  assign n6620 = ( ~n6386 & n6609 ) | ( ~n6386 & n6618 ) | ( n6609 & n6618 ) ;
  assign n6621 = ( n6386 & ~n6619 ) | ( n6386 & n6620 ) | ( ~n6619 & n6620 ) ;
  assign n6622 = ( n6398 & n6448 ) | ( n6398 & n6621 ) | ( n6448 & n6621 ) ;
  assign n6623 = ( ~n6398 & n6448 ) | ( ~n6398 & n6621 ) | ( n6448 & n6621 ) ;
  assign n6624 = ( n6398 & ~n6622 ) | ( n6398 & n6623 ) | ( ~n6622 & n6623 ) ;
  assign n6625 = ( n6401 & n6439 ) | ( n6401 & n6624 ) | ( n6439 & n6624 ) ;
  assign n6626 = ( ~n6401 & n6439 ) | ( ~n6401 & n6624 ) | ( n6439 & n6624 ) ;
  assign n6627 = ( n6401 & ~n6625 ) | ( n6401 & n6626 ) | ( ~n6625 & n6626 ) ;
  assign n6628 = n186 & n5765 ;
  assign n6629 = x114 & n190 ;
  assign n6630 = x115 | n6629 ;
  assign n6631 = ( n192 & n6629 ) | ( n192 & n6630 ) | ( n6629 & n6630 ) ;
  assign n6632 = x113 & n220 ;
  assign n6633 = n6631 | n6632 ;
  assign n6634 = ( x5 & n6628 ) | ( x5 & ~n6633 ) | ( n6628 & ~n6633 ) ;
  assign n6635 = ( ~x5 & n6633 ) | ( ~x5 & n6634 ) | ( n6633 & n6634 ) ;
  assign n6636 = ( ~n6628 & n6634 ) | ( ~n6628 & n6635 ) | ( n6634 & n6635 ) ;
  assign n6637 = ( n6413 & n6627 ) | ( n6413 & n6636 ) | ( n6627 & n6636 ) ;
  assign n6638 = ( ~n6413 & n6627 ) | ( ~n6413 & n6636 ) | ( n6627 & n6636 ) ;
  assign n6639 = ( n6413 & ~n6637 ) | ( n6413 & n6638 ) | ( ~n6637 & n6638 ) ;
  assign n6640 = ( n6416 & n6430 ) | ( n6416 & n6639 ) | ( n6430 & n6639 ) ;
  assign n6641 = ( ~n6416 & n6430 ) | ( ~n6416 & n6639 ) | ( n6430 & n6639 ) ;
  assign n6642 = ( n6416 & ~n6640 ) | ( n6416 & n6641 ) | ( ~n6640 & n6641 ) ;
  assign n6643 = ( x118 & x119 ) | ( x118 & n6419 ) | ( x119 & n6419 ) ;
  assign n6644 = ( x118 & ~x119 ) | ( x118 & n6419 ) | ( ~x119 & n6419 ) ;
  assign n6645 = ( x119 & ~n6643 ) | ( x119 & n6644 ) | ( ~n6643 & n6644 ) ;
  assign n6646 = n136 & n6645 ;
  assign n6647 = x118 & n138 ;
  assign n6648 = x119 | n6647 ;
  assign n6649 = ( n141 & n6647 ) | ( n141 & n6648 ) | ( n6647 & n6648 ) ;
  assign n6650 = x117 & n154 ;
  assign n6651 = n6649 | n6650 ;
  assign n6652 = ( x2 & n6646 ) | ( x2 & ~n6651 ) | ( n6646 & ~n6651 ) ;
  assign n6653 = ( ~x2 & n6651 ) | ( ~x2 & n6652 ) | ( n6651 & n6652 ) ;
  assign n6654 = ( ~n6646 & n6652 ) | ( ~n6646 & n6653 ) | ( n6652 & n6653 ) ;
  assign n6655 = n291 & n5542 ;
  assign n6656 = x112 & n295 ;
  assign n6657 = x113 | n6656 ;
  assign n6658 = ( n297 & n6656 ) | ( n297 & n6657 ) | ( n6656 & n6657 ) ;
  assign n6659 = x111 & n330 ;
  assign n6660 = n6658 | n6659 ;
  assign n6661 = ( x8 & n6655 ) | ( x8 & ~n6660 ) | ( n6655 & ~n6660 ) ;
  assign n6662 = ( ~x8 & n6660 ) | ( ~x8 & n6661 ) | ( n6660 & n6661 ) ;
  assign n6663 = ( ~n6655 & n6661 ) | ( ~n6655 & n6662 ) | ( n6661 & n6662 ) ;
  assign n6664 = n407 & n4934 ;
  assign n6665 = x109 & n411 ;
  assign n6666 = x110 | n6665 ;
  assign n6667 = ( n413 & n6665 ) | ( n413 & n6666 ) | ( n6665 & n6666 ) ;
  assign n6668 = x108 & n491 ;
  assign n6669 = n6667 | n6668 ;
  assign n6670 = ( x11 & n6664 ) | ( x11 & ~n6669 ) | ( n6664 & ~n6669 ) ;
  assign n6671 = ( ~x11 & n6669 ) | ( ~x11 & n6670 ) | ( n6669 & n6670 ) ;
  assign n6672 = ( ~n6664 & n6670 ) | ( ~n6664 & n6671 ) | ( n6670 & n6671 ) ;
  assign n6673 = n1366 & n2766 ;
  assign n6674 = x85 & n2770 ;
  assign n6675 = x86 | n6674 ;
  assign n6676 = ( n2772 & n6674 ) | ( n2772 & n6675 ) | ( n6674 & n6675 ) ;
  assign n6677 = x84 & n2943 ;
  assign n6678 = n6676 | n6677 ;
  assign n6679 = ( x35 & n6673 ) | ( x35 & ~n6678 ) | ( n6673 & ~n6678 ) ;
  assign n6680 = ( ~x35 & n6678 ) | ( ~x35 & n6679 ) | ( n6678 & n6679 ) ;
  assign n6681 = ( ~n6673 & n6679 ) | ( ~n6673 & n6680 ) | ( n6679 & n6680 ) ;
  assign n6682 = n569 & n4227 ;
  assign n6683 = x76 & n4231 ;
  assign n6684 = x77 | n6683 ;
  assign n6685 = ( n4233 & n6683 ) | ( n4233 & n6684 ) | ( n6683 & n6684 ) ;
  assign n6686 = x75 & n4470 ;
  assign n6687 = n6685 | n6686 ;
  assign n6688 = ( x44 & n6682 ) | ( x44 & ~n6687 ) | ( n6682 & ~n6687 ) ;
  assign n6689 = ( ~x44 & n6687 ) | ( ~x44 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6690 = ( ~n6682 & n6688 ) | ( ~n6682 & n6689 ) | ( n6688 & n6689 ) ;
  assign n6691 = n446 & n4787 ;
  assign n6692 = x73 & n4791 ;
  assign n6693 = x74 | n6692 ;
  assign n6694 = ( n4793 & n6692 ) | ( n4793 & n6693 ) | ( n6692 & n6693 ) ;
  assign n6695 = x72 & n5030 ;
  assign n6696 = n6694 | n6695 ;
  assign n6697 = ( x47 & n6691 ) | ( x47 & ~n6696 ) | ( n6691 & ~n6696 ) ;
  assign n6698 = ( ~x47 & n6696 ) | ( ~x47 & n6697 ) | ( n6696 & n6697 ) ;
  assign n6699 = ( ~n6691 & n6697 ) | ( ~n6691 & n6698 ) | ( n6697 & n6698 ) ;
  assign n6700 = n277 & n5374 ;
  assign n6701 = x70 & n5378 ;
  assign n6702 = x71 | n6701 ;
  assign n6703 = ( n5380 & n6701 ) | ( n5380 & n6702 ) | ( n6701 & n6702 ) ;
  assign n6704 = x69 & n5638 ;
  assign n6705 = n6703 | n6704 ;
  assign n6706 = ( x50 & n6700 ) | ( x50 & ~n6705 ) | ( n6700 & ~n6705 ) ;
  assign n6707 = ( ~x50 & n6705 ) | ( ~x50 & n6706 ) | ( n6705 & n6706 ) ;
  assign n6708 = ( ~n6700 & n6706 ) | ( ~n6700 & n6707 ) | ( n6706 & n6707 ) ;
  assign n6709 = x56 & n6542 ;
  assign n6710 = x55 | x56 ;
  assign n6711 = ( x55 & x56 ) | ( x55 & ~n6710 ) | ( x56 & ~n6710 ) ;
  assign n6712 = n6710 & ~n6711 ;
  assign n6713 = n6541 & n6712 ;
  assign n6714 = n133 & n6713 ;
  assign n6715 = ~x53 & x55 ;
  assign n6716 = x54 & x55 ;
  assign n6717 = ( n6539 & n6715 ) | ( n6539 & ~n6716 ) | ( n6715 & ~n6716 ) ;
  assign n6718 = x64 & n6717 ;
  assign n6719 = ( n6541 & ~n6710 ) | ( n6541 & n6711 ) | ( ~n6710 & n6711 ) ;
  assign n6720 = x65 | n6718 ;
  assign n6721 = ( n6718 & n6719 ) | ( n6718 & n6720 ) | ( n6719 & n6720 ) ;
  assign n6722 = ( n6709 & n6714 ) | ( n6709 & n6721 ) | ( n6714 & n6721 ) ;
  assign n6723 = n6714 | n6721 ;
  assign n6724 = ~n6709 & n6723 ;
  assign n6725 = ( n6709 & ~n6722 ) | ( n6709 & n6724 ) | ( ~n6722 & n6724 ) ;
  assign n6726 = x67 & n6031 ;
  assign n6727 = x68 | n6726 ;
  assign n6728 = ( n6033 & n6726 ) | ( n6033 & n6727 ) | ( n6726 & n6727 ) ;
  assign n6729 = x66 & n6303 ;
  assign n6730 = n6728 | n6729 ;
  assign n6731 = n201 & n6027 ;
  assign n6732 = ( x53 & n6730 ) | ( x53 & ~n6731 ) | ( n6730 & ~n6731 ) ;
  assign n6733 = ( ~x53 & n6731 ) | ( ~x53 & n6732 ) | ( n6731 & n6732 ) ;
  assign n6734 = ( ~n6730 & n6732 ) | ( ~n6730 & n6733 ) | ( n6732 & n6733 ) ;
  assign n6735 = ( n6544 & n6725 ) | ( n6544 & n6734 ) | ( n6725 & n6734 ) ;
  assign n6736 = ( ~n6544 & n6725 ) | ( ~n6544 & n6734 ) | ( n6725 & n6734 ) ;
  assign n6737 = ( n6544 & ~n6735 ) | ( n6544 & n6736 ) | ( ~n6735 & n6736 ) ;
  assign n6738 = ( n6556 & n6708 ) | ( n6556 & n6737 ) | ( n6708 & n6737 ) ;
  assign n6739 = ( ~n6556 & n6708 ) | ( ~n6556 & n6737 ) | ( n6708 & n6737 ) ;
  assign n6740 = ( n6556 & ~n6738 ) | ( n6556 & n6739 ) | ( ~n6738 & n6739 ) ;
  assign n6741 = ( n6559 & n6699 ) | ( n6559 & n6740 ) | ( n6699 & n6740 ) ;
  assign n6742 = ( ~n6559 & n6699 ) | ( ~n6559 & n6740 ) | ( n6699 & n6740 ) ;
  assign n6743 = ( n6559 & ~n6741 ) | ( n6559 & n6742 ) | ( ~n6741 & n6742 ) ;
  assign n6744 = ( n6562 & n6690 ) | ( n6562 & n6743 ) | ( n6690 & n6743 ) ;
  assign n6745 = ( ~n6562 & n6690 ) | ( ~n6562 & n6743 ) | ( n6690 & n6743 ) ;
  assign n6746 = ( n6562 & ~n6744 ) | ( n6562 & n6745 ) | ( ~n6744 & n6745 ) ;
  assign n6747 = n769 & n3715 ;
  assign n6748 = x79 & n3719 ;
  assign n6749 = x80 | n6748 ;
  assign n6750 = ( n3721 & n6748 ) | ( n3721 & n6749 ) | ( n6748 & n6749 ) ;
  assign n6751 = x78 & n3922 ;
  assign n6752 = n6750 | n6751 ;
  assign n6753 = ( x41 & n6747 ) | ( x41 & ~n6752 ) | ( n6747 & ~n6752 ) ;
  assign n6754 = ( ~x41 & n6752 ) | ( ~x41 & n6753 ) | ( n6752 & n6753 ) ;
  assign n6755 = ( ~n6747 & n6753 ) | ( ~n6747 & n6754 ) | ( n6753 & n6754 ) ;
  assign n6756 = ( n6565 & n6746 ) | ( n6565 & n6755 ) | ( n6746 & n6755 ) ;
  assign n6757 = ( ~n6565 & n6746 ) | ( ~n6565 & n6755 ) | ( n6746 & n6755 ) ;
  assign n6758 = ( n6565 & ~n6756 ) | ( n6565 & n6757 ) | ( ~n6756 & n6757 ) ;
  assign n6759 = n1082 & n3224 ;
  assign n6760 = x82 & n3228 ;
  assign n6761 = x83 | n6760 ;
  assign n6762 = ( n3230 & n6760 ) | ( n3230 & n6761 ) | ( n6760 & n6761 ) ;
  assign n6763 = x81 & n3413 ;
  assign n6764 = n6762 | n6763 ;
  assign n6765 = ( x38 & n6759 ) | ( x38 & ~n6764 ) | ( n6759 & ~n6764 ) ;
  assign n6766 = ( ~x38 & n6764 ) | ( ~x38 & n6765 ) | ( n6764 & n6765 ) ;
  assign n6767 = ( ~n6759 & n6765 ) | ( ~n6759 & n6766 ) | ( n6765 & n6766 ) ;
  assign n6768 = ( n6568 & n6758 ) | ( n6568 & n6767 ) | ( n6758 & n6767 ) ;
  assign n6769 = ( ~n6568 & n6758 ) | ( ~n6568 & n6767 ) | ( n6758 & n6767 ) ;
  assign n6770 = ( n6568 & ~n6768 ) | ( n6568 & n6769 ) | ( ~n6768 & n6769 ) ;
  assign n6771 = ( n6571 & n6681 ) | ( n6571 & n6770 ) | ( n6681 & n6770 ) ;
  assign n6772 = ( ~n6571 & n6681 ) | ( ~n6571 & n6770 ) | ( n6681 & n6770 ) ;
  assign n6773 = ( n6571 & ~n6771 ) | ( n6571 & n6772 ) | ( ~n6771 & n6772 ) ;
  assign n6774 = n1585 & n2320 ;
  assign n6775 = x88 & n2324 ;
  assign n6776 = x89 | n6775 ;
  assign n6777 = ( n2326 & n6775 ) | ( n2326 & n6776 ) | ( n6775 & n6776 ) ;
  assign n6778 = x87 & n2497 ;
  assign n6779 = n6777 | n6778 ;
  assign n6780 = ( x32 & n6774 ) | ( x32 & ~n6779 ) | ( n6774 & ~n6779 ) ;
  assign n6781 = ( ~x32 & n6779 ) | ( ~x32 & n6780 ) | ( n6779 & n6780 ) ;
  assign n6782 = ( ~n6774 & n6780 ) | ( ~n6774 & n6781 ) | ( n6780 & n6781 ) ;
  assign n6783 = ( n6574 & n6773 ) | ( n6574 & n6782 ) | ( n6773 & n6782 ) ;
  assign n6784 = ( ~n6574 & n6773 ) | ( ~n6574 & n6782 ) | ( n6773 & n6782 ) ;
  assign n6785 = ( n6574 & ~n6783 ) | ( n6574 & n6784 ) | ( ~n6783 & n6784 ) ;
  assign n6786 = n1949 & n2042 ;
  assign n6787 = x91 & n1953 ;
  assign n6788 = x92 | n6787 ;
  assign n6789 = ( n1955 & n6787 ) | ( n1955 & n6788 ) | ( n6787 & n6788 ) ;
  assign n6790 = x90 & n2114 ;
  assign n6791 = n6789 | n6790 ;
  assign n6792 = ( x29 & n6786 ) | ( x29 & ~n6791 ) | ( n6786 & ~n6791 ) ;
  assign n6793 = ( ~x29 & n6791 ) | ( ~x29 & n6792 ) | ( n6791 & n6792 ) ;
  assign n6794 = ( ~n6786 & n6792 ) | ( ~n6786 & n6793 ) | ( n6792 & n6793 ) ;
  assign n6795 = ( n6577 & n6785 ) | ( n6577 & n6794 ) | ( n6785 & n6794 ) ;
  assign n6796 = ( ~n6577 & n6785 ) | ( ~n6577 & n6794 ) | ( n6785 & n6794 ) ;
  assign n6797 = ( n6577 & ~n6795 ) | ( n6577 & n6796 ) | ( ~n6795 & n6796 ) ;
  assign n6798 = n1617 & n2434 ;
  assign n6799 = x94 & n1621 ;
  assign n6800 = x95 | n6799 ;
  assign n6801 = ( n1623 & n6799 ) | ( n1623 & n6800 ) | ( n6799 & n6800 ) ;
  assign n6802 = x93 & n1749 ;
  assign n6803 = n6801 | n6802 ;
  assign n6804 = ( x26 & n6798 ) | ( x26 & ~n6803 ) | ( n6798 & ~n6803 ) ;
  assign n6805 = ( ~x26 & n6803 ) | ( ~x26 & n6804 ) | ( n6803 & n6804 ) ;
  assign n6806 = ( ~n6798 & n6804 ) | ( ~n6798 & n6805 ) | ( n6804 & n6805 ) ;
  assign n6807 = ( n6580 & n6797 ) | ( n6580 & n6806 ) | ( n6797 & n6806 ) ;
  assign n6808 = ( ~n6580 & n6797 ) | ( ~n6580 & n6806 ) | ( n6797 & n6806 ) ;
  assign n6809 = ( n6580 & ~n6807 ) | ( n6580 & n6808 ) | ( ~n6807 & n6808 ) ;
  assign n6810 = n1297 & n2725 ;
  assign n6811 = x97 & n1301 ;
  assign n6812 = x98 | n6811 ;
  assign n6813 = ( n1303 & n6811 ) | ( n1303 & n6812 ) | ( n6811 & n6812 ) ;
  assign n6814 = x96 & n1426 ;
  assign n6815 = n6813 | n6814 ;
  assign n6816 = ( x23 & n6810 ) | ( x23 & ~n6815 ) | ( n6810 & ~n6815 ) ;
  assign n6817 = ( ~x23 & n6815 ) | ( ~x23 & n6816 ) | ( n6815 & n6816 ) ;
  assign n6818 = ( ~n6810 & n6816 ) | ( ~n6810 & n6817 ) | ( n6816 & n6817 ) ;
  assign n6819 = ( n6592 & n6809 ) | ( n6592 & n6818 ) | ( n6809 & n6818 ) ;
  assign n6820 = ( ~n6592 & n6809 ) | ( ~n6592 & n6818 ) | ( n6809 & n6818 ) ;
  assign n6821 = ( n6592 & ~n6819 ) | ( n6592 & n6820 ) | ( ~n6819 & n6820 ) ;
  assign n6822 = n1016 & n3326 ;
  assign n6823 = x100 & n1020 ;
  assign n6824 = x101 | n6823 ;
  assign n6825 = ( n1022 & n6823 ) | ( n1022 & n6824 ) | ( n6823 & n6824 ) ;
  assign n6826 = x99 & n1145 ;
  assign n6827 = n6825 | n6826 ;
  assign n6828 = ( x20 & n6822 ) | ( x20 & ~n6827 ) | ( n6822 & ~n6827 ) ;
  assign n6829 = ( ~x20 & n6827 ) | ( ~x20 & n6828 ) | ( n6827 & n6828 ) ;
  assign n6830 = ( ~n6822 & n6828 ) | ( ~n6822 & n6829 ) | ( n6828 & n6829 ) ;
  assign n6831 = ( n6595 & n6821 ) | ( n6595 & n6830 ) | ( n6821 & n6830 ) ;
  assign n6832 = ( ~n6595 & n6821 ) | ( ~n6595 & n6830 ) | ( n6821 & n6830 ) ;
  assign n6833 = ( n6595 & ~n6831 ) | ( n6595 & n6832 ) | ( ~n6831 & n6832 ) ;
  assign n6834 = n810 & n3665 ;
  assign n6835 = x103 & n814 ;
  assign n6836 = x104 | n6835 ;
  assign n6837 = ( n816 & n6835 ) | ( n816 & n6836 ) | ( n6835 & n6836 ) ;
  assign n6838 = x102 & n885 ;
  assign n6839 = n6837 | n6838 ;
  assign n6840 = ( x17 & n6834 ) | ( x17 & ~n6839 ) | ( n6834 & ~n6839 ) ;
  assign n6841 = ( ~x17 & n6839 ) | ( ~x17 & n6840 ) | ( n6839 & n6840 ) ;
  assign n6842 = ( ~n6834 & n6840 ) | ( ~n6834 & n6841 ) | ( n6840 & n6841 ) ;
  assign n6843 = ( n6607 & n6833 ) | ( n6607 & n6842 ) | ( n6833 & n6842 ) ;
  assign n6844 = ( ~n6607 & n6833 ) | ( ~n6607 & n6842 ) | ( n6833 & n6842 ) ;
  assign n6845 = ( n6607 & ~n6843 ) | ( n6607 & n6844 ) | ( ~n6843 & n6844 ) ;
  assign n6846 = n583 & n4362 ;
  assign n6847 = x106 & n587 ;
  assign n6848 = x107 | n6847 ;
  assign n6849 = ( n589 & n6847 ) | ( n589 & n6848 ) | ( n6847 & n6848 ) ;
  assign n6850 = x105 & n676 ;
  assign n6851 = n6849 | n6850 ;
  assign n6852 = ( x14 & n6846 ) | ( x14 & ~n6851 ) | ( n6846 & ~n6851 ) ;
  assign n6853 = ( ~x14 & n6851 ) | ( ~x14 & n6852 ) | ( n6851 & n6852 ) ;
  assign n6854 = ( ~n6846 & n6852 ) | ( ~n6846 & n6853 ) | ( n6852 & n6853 ) ;
  assign n6855 = ( n6619 & n6845 ) | ( n6619 & n6854 ) | ( n6845 & n6854 ) ;
  assign n6856 = ( ~n6619 & n6845 ) | ( ~n6619 & n6854 ) | ( n6845 & n6854 ) ;
  assign n6857 = ( n6619 & ~n6855 ) | ( n6619 & n6856 ) | ( ~n6855 & n6856 ) ;
  assign n6858 = ( n6622 & n6672 ) | ( n6622 & n6857 ) | ( n6672 & n6857 ) ;
  assign n6859 = ( ~n6622 & n6672 ) | ( ~n6622 & n6857 ) | ( n6672 & n6857 ) ;
  assign n6860 = ( n6622 & ~n6858 ) | ( n6622 & n6859 ) | ( ~n6858 & n6859 ) ;
  assign n6861 = ( n6625 & n6663 ) | ( n6625 & n6860 ) | ( n6663 & n6860 ) ;
  assign n6862 = ( ~n6625 & n6663 ) | ( ~n6625 & n6860 ) | ( n6663 & n6860 ) ;
  assign n6863 = ( n6625 & ~n6861 ) | ( n6625 & n6862 ) | ( ~n6861 & n6862 ) ;
  assign n6864 = n186 & n5977 ;
  assign n6865 = x115 & n190 ;
  assign n6866 = x116 | n6865 ;
  assign n6867 = ( n192 & n6865 ) | ( n192 & n6866 ) | ( n6865 & n6866 ) ;
  assign n6868 = x114 & n220 ;
  assign n6869 = n6867 | n6868 ;
  assign n6870 = ( x5 & n6864 ) | ( x5 & ~n6869 ) | ( n6864 & ~n6869 ) ;
  assign n6871 = ( ~x5 & n6869 ) | ( ~x5 & n6870 ) | ( n6869 & n6870 ) ;
  assign n6872 = ( ~n6864 & n6870 ) | ( ~n6864 & n6871 ) | ( n6870 & n6871 ) ;
  assign n6873 = ( n6637 & n6863 ) | ( n6637 & n6872 ) | ( n6863 & n6872 ) ;
  assign n6874 = ( ~n6637 & n6863 ) | ( ~n6637 & n6872 ) | ( n6863 & n6872 ) ;
  assign n6875 = ( n6637 & ~n6873 ) | ( n6637 & n6874 ) | ( ~n6873 & n6874 ) ;
  assign n6876 = ( n6640 & n6654 ) | ( n6640 & n6875 ) | ( n6654 & n6875 ) ;
  assign n6877 = ( ~n6640 & n6654 ) | ( ~n6640 & n6875 ) | ( n6654 & n6875 ) ;
  assign n6878 = ( n6640 & ~n6876 ) | ( n6640 & n6877 ) | ( ~n6876 & n6877 ) ;
  assign n6879 = n186 & n6201 ;
  assign n6880 = x116 & n190 ;
  assign n6881 = x117 | n6880 ;
  assign n6882 = ( n192 & n6880 ) | ( n192 & n6881 ) | ( n6880 & n6881 ) ;
  assign n6883 = x115 & n220 ;
  assign n6884 = n6882 | n6883 ;
  assign n6885 = ( x5 & n6879 ) | ( x5 & ~n6884 ) | ( n6879 & ~n6884 ) ;
  assign n6886 = ( ~x5 & n6884 ) | ( ~x5 & n6885 ) | ( n6884 & n6885 ) ;
  assign n6887 = ( ~n6879 & n6885 ) | ( ~n6879 & n6886 ) | ( n6885 & n6886 ) ;
  assign n6888 = n291 & n5750 ;
  assign n6889 = x113 & n295 ;
  assign n6890 = x114 | n6889 ;
  assign n6891 = ( n297 & n6889 ) | ( n297 & n6890 ) | ( n6889 & n6890 ) ;
  assign n6892 = x112 & n330 ;
  assign n6893 = n6891 | n6892 ;
  assign n6894 = ( x8 & n6888 ) | ( x8 & ~n6893 ) | ( n6888 & ~n6893 ) ;
  assign n6895 = ( ~x8 & n6893 ) | ( ~x8 & n6894 ) | ( n6893 & n6894 ) ;
  assign n6896 = ( ~n6888 & n6894 ) | ( ~n6888 & n6895 ) | ( n6894 & n6895 ) ;
  assign n6897 = n407 & n5130 ;
  assign n6898 = x110 & n411 ;
  assign n6899 = x111 | n6898 ;
  assign n6900 = ( n413 & n6898 ) | ( n413 & n6899 ) | ( n6898 & n6899 ) ;
  assign n6901 = x109 & n491 ;
  assign n6902 = n6900 | n6901 ;
  assign n6903 = ( x11 & n6897 ) | ( x11 & ~n6902 ) | ( n6897 & ~n6902 ) ;
  assign n6904 = ( ~x11 & n6902 ) | ( ~x11 & n6903 ) | ( n6902 & n6903 ) ;
  assign n6905 = ( ~n6897 & n6903 ) | ( ~n6897 & n6904 ) | ( n6903 & n6904 ) ;
  assign n6906 = n1617 & n2449 ;
  assign n6907 = x95 & n1621 ;
  assign n6908 = x96 | n6907 ;
  assign n6909 = ( n1623 & n6907 ) | ( n1623 & n6908 ) | ( n6907 & n6908 ) ;
  assign n6910 = x94 & n1749 ;
  assign n6911 = n6909 | n6910 ;
  assign n6912 = ( x26 & n6906 ) | ( x26 & ~n6911 ) | ( n6906 & ~n6911 ) ;
  assign n6913 = ( ~x26 & n6911 ) | ( ~x26 & n6912 ) | ( n6911 & n6912 ) ;
  assign n6914 = ( ~n6906 & n6912 ) | ( ~n6906 & n6913 ) | ( n6912 & n6913 ) ;
  assign n6915 = n1949 & n2057 ;
  assign n6916 = x92 & n1953 ;
  assign n6917 = x93 | n6916 ;
  assign n6918 = ( n1955 & n6916 ) | ( n1955 & n6917 ) | ( n6916 & n6917 ) ;
  assign n6919 = x91 & n2114 ;
  assign n6920 = n6918 | n6919 ;
  assign n6921 = ( x29 & n6915 ) | ( x29 & ~n6920 ) | ( n6915 & ~n6920 ) ;
  assign n6922 = ( ~x29 & n6920 ) | ( ~x29 & n6921 ) | ( n6920 & n6921 ) ;
  assign n6923 = ( ~n6915 & n6921 ) | ( ~n6915 & n6922 ) | ( n6921 & n6922 ) ;
  assign n6924 = n1466 & n2766 ;
  assign n6925 = x86 & n2770 ;
  assign n6926 = x87 | n6925 ;
  assign n6927 = ( n2772 & n6925 ) | ( n2772 & n6926 ) | ( n6925 & n6926 ) ;
  assign n6928 = x85 & n2943 ;
  assign n6929 = n6927 | n6928 ;
  assign n6930 = ( x35 & n6924 ) | ( x35 & ~n6929 ) | ( n6924 & ~n6929 ) ;
  assign n6931 = ( ~x35 & n6929 ) | ( ~x35 & n6930 ) | ( n6929 & n6930 ) ;
  assign n6932 = ( ~n6924 & n6930 ) | ( ~n6924 & n6931 ) | ( n6930 & n6931 ) ;
  assign n6933 = n1097 & n3224 ;
  assign n6934 = x83 & n3228 ;
  assign n6935 = x84 | n6934 ;
  assign n6936 = ( n3230 & n6934 ) | ( n3230 & n6935 ) | ( n6934 & n6935 ) ;
  assign n6937 = x82 & n3413 ;
  assign n6938 = n6936 | n6937 ;
  assign n6939 = ( x38 & n6933 ) | ( x38 & ~n6938 ) | ( n6933 & ~n6938 ) ;
  assign n6940 = ( ~x38 & n6938 ) | ( ~x38 & n6939 ) | ( n6938 & n6939 ) ;
  assign n6941 = ( ~n6933 & n6939 ) | ( ~n6933 & n6940 ) | ( n6939 & n6940 ) ;
  assign n6942 = n910 & n3715 ;
  assign n6943 = x80 & n3719 ;
  assign n6944 = x81 | n6943 ;
  assign n6945 = ( n3721 & n6943 ) | ( n3721 & n6944 ) | ( n6943 & n6944 ) ;
  assign n6946 = x79 & n3922 ;
  assign n6947 = n6945 | n6946 ;
  assign n6948 = ( x41 & n6942 ) | ( x41 & ~n6947 ) | ( n6942 & ~n6947 ) ;
  assign n6949 = ( ~x41 & n6947 ) | ( ~x41 & n6948 ) | ( n6947 & n6948 ) ;
  assign n6950 = ( ~n6942 & n6948 ) | ( ~n6942 & n6949 ) | ( n6948 & n6949 ) ;
  assign n6951 = n461 & n4787 ;
  assign n6952 = x74 & n4791 ;
  assign n6953 = x75 | n6952 ;
  assign n6954 = ( n4793 & n6952 ) | ( n4793 & n6953 ) | ( n6952 & n6953 ) ;
  assign n6955 = x73 & n5030 ;
  assign n6956 = n6954 | n6955 ;
  assign n6957 = ( x47 & n6951 ) | ( x47 & ~n6956 ) | ( n6951 & ~n6956 ) ;
  assign n6958 = ( ~x47 & n6956 ) | ( ~x47 & n6957 ) | ( n6956 & n6957 ) ;
  assign n6959 = ( ~n6951 & n6957 ) | ( ~n6951 & n6958 ) | ( n6957 & n6958 ) ;
  assign n6960 = n346 & n5374 ;
  assign n6961 = x71 & n5378 ;
  assign n6962 = x72 | n6961 ;
  assign n6963 = ( n5380 & n6961 ) | ( n5380 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6964 = x70 & n5638 ;
  assign n6965 = n6963 | n6964 ;
  assign n6966 = ( x50 & n6960 ) | ( x50 & ~n6965 ) | ( n6960 & ~n6965 ) ;
  assign n6967 = ( ~x50 & n6965 ) | ( ~x50 & n6966 ) | ( n6965 & n6966 ) ;
  assign n6968 = ( ~n6960 & n6966 ) | ( ~n6960 & n6967 ) | ( n6966 & n6967 ) ;
  assign n6969 = n230 & n6027 ;
  assign n6970 = x68 & n6031 ;
  assign n6971 = x69 | n6970 ;
  assign n6972 = ( n6033 & n6970 ) | ( n6033 & n6971 ) | ( n6970 & n6971 ) ;
  assign n6973 = x67 & n6303 ;
  assign n6974 = n6972 | n6973 ;
  assign n6975 = ( ~x53 & n6969 ) | ( ~x53 & n6974 ) | ( n6969 & n6974 ) ;
  assign n6976 = ( n6969 & n6974 ) | ( n6969 & ~n6975 ) | ( n6974 & ~n6975 ) ;
  assign n6977 = ( x53 & n6975 ) | ( x53 & ~n6976 ) | ( n6975 & ~n6976 ) ;
  assign n6978 = ( x56 & n6709 ) | ( x56 & n6723 ) | ( n6709 & n6723 ) ;
  assign n6979 = ( x53 & ~x55 ) | ( x53 & n6712 ) | ( ~x55 & n6712 ) ;
  assign n6980 = ( ~n6540 & n6716 ) | ( ~n6540 & n6979 ) | ( n6716 & n6979 ) ;
  assign n6981 = x64 & n6980 ;
  assign n6982 = x65 & n6717 ;
  assign n6983 = x66 | n6982 ;
  assign n6984 = ( n6719 & n6982 ) | ( n6719 & n6983 ) | ( n6982 & n6983 ) ;
  assign n6985 = ( n151 & n152 ) | ( n151 & n6713 ) | ( n152 & n6713 ) ;
  assign n6986 = ( ~n6981 & n6984 ) | ( ~n6981 & n6985 ) | ( n6984 & n6985 ) ;
  assign n6987 = n6981 | n6986 ;
  assign n6988 = n6978 | n6987 ;
  assign n6989 = ( n6978 & n6987 ) | ( n6978 & ~n6988 ) | ( n6987 & ~n6988 ) ;
  assign n6990 = n6988 & ~n6989 ;
  assign n6991 = ( n6735 & n6977 ) | ( n6735 & n6990 ) | ( n6977 & n6990 ) ;
  assign n6992 = ( ~n6735 & n6977 ) | ( ~n6735 & n6990 ) | ( n6977 & n6990 ) ;
  assign n6993 = ( n6735 & ~n6991 ) | ( n6735 & n6992 ) | ( ~n6991 & n6992 ) ;
  assign n6994 = ( n6738 & n6968 ) | ( n6738 & n6993 ) | ( n6968 & n6993 ) ;
  assign n6995 = ( ~n6738 & n6968 ) | ( ~n6738 & n6993 ) | ( n6968 & n6993 ) ;
  assign n6996 = ( n6738 & ~n6994 ) | ( n6738 & n6995 ) | ( ~n6994 & n6995 ) ;
  assign n6997 = ( n6741 & n6959 ) | ( n6741 & n6996 ) | ( n6959 & n6996 ) ;
  assign n6998 = ( ~n6741 & n6959 ) | ( ~n6741 & n6996 ) | ( n6959 & n6996 ) ;
  assign n6999 = ( n6741 & ~n6997 ) | ( n6741 & n6998 ) | ( ~n6997 & n6998 ) ;
  assign n7000 = n637 & n4227 ;
  assign n7001 = x77 & n4231 ;
  assign n7002 = x78 | n7001 ;
  assign n7003 = ( n4233 & n7001 ) | ( n4233 & n7002 ) | ( n7001 & n7002 ) ;
  assign n7004 = x76 & n4470 ;
  assign n7005 = n7003 | n7004 ;
  assign n7006 = ( x44 & n7000 ) | ( x44 & ~n7005 ) | ( n7000 & ~n7005 ) ;
  assign n7007 = ( ~x44 & n7005 ) | ( ~x44 & n7006 ) | ( n7005 & n7006 ) ;
  assign n7008 = ( ~n7000 & n7006 ) | ( ~n7000 & n7007 ) | ( n7006 & n7007 ) ;
  assign n7009 = ( n6744 & n6999 ) | ( n6744 & n7008 ) | ( n6999 & n7008 ) ;
  assign n7010 = ( ~n6744 & n6999 ) | ( ~n6744 & n7008 ) | ( n6999 & n7008 ) ;
  assign n7011 = ( n6744 & ~n7009 ) | ( n6744 & n7010 ) | ( ~n7009 & n7010 ) ;
  assign n7012 = ( n6756 & n6950 ) | ( n6756 & n7011 ) | ( n6950 & n7011 ) ;
  assign n7013 = ( ~n6756 & n6950 ) | ( ~n6756 & n7011 ) | ( n6950 & n7011 ) ;
  assign n7014 = ( n6756 & ~n7012 ) | ( n6756 & n7013 ) | ( ~n7012 & n7013 ) ;
  assign n7015 = ( n6768 & n6941 ) | ( n6768 & n7014 ) | ( n6941 & n7014 ) ;
  assign n7016 = ( ~n6768 & n6941 ) | ( ~n6768 & n7014 ) | ( n6941 & n7014 ) ;
  assign n7017 = ( n6768 & ~n7015 ) | ( n6768 & n7016 ) | ( ~n7015 & n7016 ) ;
  assign n7018 = ( n6771 & n6932 ) | ( n6771 & n7017 ) | ( n6932 & n7017 ) ;
  assign n7019 = ( ~n6771 & n6932 ) | ( ~n6771 & n7017 ) | ( n6932 & n7017 ) ;
  assign n7020 = ( n6771 & ~n7018 ) | ( n6771 & n7019 ) | ( ~n7018 & n7019 ) ;
  assign n7021 = n1701 & n2320 ;
  assign n7022 = x89 & n2324 ;
  assign n7023 = x90 | n7022 ;
  assign n7024 = ( n2326 & n7022 ) | ( n2326 & n7023 ) | ( n7022 & n7023 ) ;
  assign n7025 = x88 & n2497 ;
  assign n7026 = n7024 | n7025 ;
  assign n7027 = ( x32 & n7021 ) | ( x32 & ~n7026 ) | ( n7021 & ~n7026 ) ;
  assign n7028 = ( ~x32 & n7026 ) | ( ~x32 & n7027 ) | ( n7026 & n7027 ) ;
  assign n7029 = ( ~n7021 & n7027 ) | ( ~n7021 & n7028 ) | ( n7027 & n7028 ) ;
  assign n7030 = ( n6783 & n7020 ) | ( n6783 & n7029 ) | ( n7020 & n7029 ) ;
  assign n7031 = ( ~n6783 & n7020 ) | ( ~n6783 & n7029 ) | ( n7020 & n7029 ) ;
  assign n7032 = ( n6783 & ~n7030 ) | ( n6783 & n7031 ) | ( ~n7030 & n7031 ) ;
  assign n7033 = ( n6795 & n6923 ) | ( n6795 & n7032 ) | ( n6923 & n7032 ) ;
  assign n7034 = ( ~n6795 & n6923 ) | ( ~n6795 & n7032 ) | ( n6923 & n7032 ) ;
  assign n7035 = ( n6795 & ~n7033 ) | ( n6795 & n7034 ) | ( ~n7033 & n7034 ) ;
  assign n7036 = ( n6807 & n6914 ) | ( n6807 & n7035 ) | ( n6914 & n7035 ) ;
  assign n7037 = ( ~n6807 & n6914 ) | ( ~n6807 & n7035 ) | ( n6914 & n7035 ) ;
  assign n7038 = ( n6807 & ~n7036 ) | ( n6807 & n7037 ) | ( ~n7036 & n7037 ) ;
  assign n7039 = n1297 & n2877 ;
  assign n7040 = x98 & n1301 ;
  assign n7041 = x99 | n7040 ;
  assign n7042 = ( n1303 & n7040 ) | ( n1303 & n7041 ) | ( n7040 & n7041 ) ;
  assign n7043 = x97 & n1426 ;
  assign n7044 = n7042 | n7043 ;
  assign n7045 = ( x23 & n7039 ) | ( x23 & ~n7044 ) | ( n7039 & ~n7044 ) ;
  assign n7046 = ( ~x23 & n7044 ) | ( ~x23 & n7045 ) | ( n7044 & n7045 ) ;
  assign n7047 = ( ~n7039 & n7045 ) | ( ~n7039 & n7046 ) | ( n7045 & n7046 ) ;
  assign n7048 = ( n6819 & n7038 ) | ( n6819 & n7047 ) | ( n7038 & n7047 ) ;
  assign n7049 = ( ~n6819 & n7038 ) | ( ~n6819 & n7047 ) | ( n7038 & n7047 ) ;
  assign n7050 = ( n6819 & ~n7048 ) | ( n6819 & n7049 ) | ( ~n7048 & n7049 ) ;
  assign n7051 = n1016 & n3486 ;
  assign n7052 = x101 & n1020 ;
  assign n7053 = x102 | n7052 ;
  assign n7054 = ( n1022 & n7052 ) | ( n1022 & n7053 ) | ( n7052 & n7053 ) ;
  assign n7055 = x100 & n1145 ;
  assign n7056 = n7054 | n7055 ;
  assign n7057 = ( x20 & n7051 ) | ( x20 & ~n7056 ) | ( n7051 & ~n7056 ) ;
  assign n7058 = ( ~x20 & n7056 ) | ( ~x20 & n7057 ) | ( n7056 & n7057 ) ;
  assign n7059 = ( ~n7051 & n7057 ) | ( ~n7051 & n7058 ) | ( n7057 & n7058 ) ;
  assign n7060 = ( n6831 & n7050 ) | ( n6831 & n7059 ) | ( n7050 & n7059 ) ;
  assign n7061 = ( ~n6831 & n7050 ) | ( ~n6831 & n7059 ) | ( n7050 & n7059 ) ;
  assign n7062 = ( n6831 & ~n7060 ) | ( n6831 & n7061 ) | ( ~n7060 & n7061 ) ;
  assign n7063 = n810 & n3998 ;
  assign n7064 = x104 & n814 ;
  assign n7065 = x105 | n7064 ;
  assign n7066 = ( n816 & n7064 ) | ( n816 & n7065 ) | ( n7064 & n7065 ) ;
  assign n7067 = x103 & n885 ;
  assign n7068 = n7066 | n7067 ;
  assign n7069 = ( x17 & n7063 ) | ( x17 & ~n7068 ) | ( n7063 & ~n7068 ) ;
  assign n7070 = ( ~x17 & n7068 ) | ( ~x17 & n7069 ) | ( n7068 & n7069 ) ;
  assign n7071 = ( ~n7063 & n7069 ) | ( ~n7063 & n7070 ) | ( n7069 & n7070 ) ;
  assign n7072 = ( n6843 & n7062 ) | ( n6843 & n7071 ) | ( n7062 & n7071 ) ;
  assign n7073 = ( ~n6843 & n7062 ) | ( ~n6843 & n7071 ) | ( n7062 & n7071 ) ;
  assign n7074 = ( n6843 & ~n7072 ) | ( n6843 & n7073 ) | ( ~n7072 & n7073 ) ;
  assign n7075 = n583 & n4377 ;
  assign n7076 = x107 & n587 ;
  assign n7077 = x108 | n7076 ;
  assign n7078 = ( n589 & n7076 ) | ( n589 & n7077 ) | ( n7076 & n7077 ) ;
  assign n7079 = x106 & n676 ;
  assign n7080 = n7078 | n7079 ;
  assign n7081 = ( x14 & n7075 ) | ( x14 & ~n7080 ) | ( n7075 & ~n7080 ) ;
  assign n7082 = ( ~x14 & n7080 ) | ( ~x14 & n7081 ) | ( n7080 & n7081 ) ;
  assign n7083 = ( ~n7075 & n7081 ) | ( ~n7075 & n7082 ) | ( n7081 & n7082 ) ;
  assign n7084 = ( n6855 & n7074 ) | ( n6855 & n7083 ) | ( n7074 & n7083 ) ;
  assign n7085 = ( ~n6855 & n7074 ) | ( ~n6855 & n7083 ) | ( n7074 & n7083 ) ;
  assign n7086 = ( n6855 & ~n7084 ) | ( n6855 & n7085 ) | ( ~n7084 & n7085 ) ;
  assign n7087 = ( n6858 & n6905 ) | ( n6858 & n7086 ) | ( n6905 & n7086 ) ;
  assign n7088 = ( ~n6858 & n6905 ) | ( ~n6858 & n7086 ) | ( n6905 & n7086 ) ;
  assign n7089 = ( n6858 & ~n7087 ) | ( n6858 & n7088 ) | ( ~n7087 & n7088 ) ;
  assign n7090 = ( n6861 & n6896 ) | ( n6861 & n7089 ) | ( n6896 & n7089 ) ;
  assign n7091 = ( ~n6861 & n6896 ) | ( ~n6861 & n7089 ) | ( n6896 & n7089 ) ;
  assign n7092 = ( n6861 & ~n7090 ) | ( n6861 & n7091 ) | ( ~n7090 & n7091 ) ;
  assign n7093 = ( n6873 & n6887 ) | ( n6873 & n7092 ) | ( n6887 & n7092 ) ;
  assign n7094 = ( ~n6873 & n6887 ) | ( ~n6873 & n7092 ) | ( n6887 & n7092 ) ;
  assign n7095 = ( n6873 & ~n7093 ) | ( n6873 & n7094 ) | ( ~n7093 & n7094 ) ;
  assign n7096 = ( x119 & x120 ) | ( x119 & n6643 ) | ( x120 & n6643 ) ;
  assign n7097 = ( x119 & ~x120 ) | ( x119 & n6643 ) | ( ~x120 & n6643 ) ;
  assign n7098 = ( x120 & ~n7096 ) | ( x120 & n7097 ) | ( ~n7096 & n7097 ) ;
  assign n7099 = n136 & n7098 ;
  assign n7100 = x119 & n138 ;
  assign n7101 = x120 | n7100 ;
  assign n7102 = ( n141 & n7100 ) | ( n141 & n7101 ) | ( n7100 & n7101 ) ;
  assign n7103 = x118 & n154 ;
  assign n7104 = n7102 | n7103 ;
  assign n7105 = ( x2 & n7099 ) | ( x2 & ~n7104 ) | ( n7099 & ~n7104 ) ;
  assign n7106 = ( ~x2 & n7104 ) | ( ~x2 & n7105 ) | ( n7104 & n7105 ) ;
  assign n7107 = ( ~n7099 & n7105 ) | ( ~n7099 & n7106 ) | ( n7105 & n7106 ) ;
  assign n7108 = ( n6876 & n7095 ) | ( n6876 & n7107 ) | ( n7095 & n7107 ) ;
  assign n7109 = ( ~n6876 & n7095 ) | ( ~n6876 & n7107 ) | ( n7095 & n7107 ) ;
  assign n7110 = ( n6876 & ~n7108 ) | ( n6876 & n7109 ) | ( ~n7108 & n7109 ) ;
  assign n7111 = ( x120 & x121 ) | ( x120 & n7096 ) | ( x121 & n7096 ) ;
  assign n7112 = ( x120 & ~x121 ) | ( x120 & n7096 ) | ( ~x121 & n7096 ) ;
  assign n7113 = ( x121 & ~n7111 ) | ( x121 & n7112 ) | ( ~n7111 & n7112 ) ;
  assign n7114 = n136 & n7113 ;
  assign n7115 = x120 & n138 ;
  assign n7116 = x121 | n7115 ;
  assign n7117 = ( n141 & n7115 ) | ( n141 & n7116 ) | ( n7115 & n7116 ) ;
  assign n7118 = x119 & n154 ;
  assign n7119 = n7117 | n7118 ;
  assign n7120 = ( x2 & n7114 ) | ( x2 & ~n7119 ) | ( n7114 & ~n7119 ) ;
  assign n7121 = ( ~x2 & n7119 ) | ( ~x2 & n7120 ) | ( n7119 & n7120 ) ;
  assign n7122 = ( ~n7114 & n7120 ) | ( ~n7114 & n7121 ) | ( n7120 & n7121 ) ;
  assign n7123 = n186 & n6421 ;
  assign n7124 = x117 & n190 ;
  assign n7125 = x118 | n7124 ;
  assign n7126 = ( n192 & n7124 ) | ( n192 & n7125 ) | ( n7124 & n7125 ) ;
  assign n7127 = x116 & n220 ;
  assign n7128 = n7126 | n7127 ;
  assign n7129 = ( x5 & n7123 ) | ( x5 & ~n7128 ) | ( n7123 & ~n7128 ) ;
  assign n7130 = ( ~x5 & n7128 ) | ( ~x5 & n7129 ) | ( n7128 & n7129 ) ;
  assign n7131 = ( ~n7123 & n7129 ) | ( ~n7123 & n7130 ) | ( n7129 & n7130 ) ;
  assign n7132 = n291 & n5765 ;
  assign n7133 = x114 & n295 ;
  assign n7134 = x115 | n7133 ;
  assign n7135 = ( n297 & n7133 ) | ( n297 & n7134 ) | ( n7133 & n7134 ) ;
  assign n7136 = x113 & n330 ;
  assign n7137 = n7135 | n7136 ;
  assign n7138 = ( x8 & n7132 ) | ( x8 & ~n7137 ) | ( n7132 & ~n7137 ) ;
  assign n7139 = ( ~x8 & n7137 ) | ( ~x8 & n7138 ) | ( n7137 & n7138 ) ;
  assign n7140 = ( ~n7132 & n7138 ) | ( ~n7132 & n7139 ) | ( n7138 & n7139 ) ;
  assign n7141 = n407 & n5145 ;
  assign n7142 = x111 & n411 ;
  assign n7143 = x112 | n7142 ;
  assign n7144 = ( n413 & n7142 ) | ( n413 & n7143 ) | ( n7142 & n7143 ) ;
  assign n7145 = x110 & n491 ;
  assign n7146 = n7144 | n7145 ;
  assign n7147 = ( x11 & n7141 ) | ( x11 & ~n7146 ) | ( n7141 & ~n7146 ) ;
  assign n7148 = ( ~x11 & n7146 ) | ( ~x11 & n7147 ) | ( n7146 & n7147 ) ;
  assign n7149 = ( ~n7141 & n7147 ) | ( ~n7141 & n7148 ) | ( n7147 & n7148 ) ;
  assign n7150 = n583 & n4734 ;
  assign n7151 = x108 & n587 ;
  assign n7152 = x109 | n7151 ;
  assign n7153 = ( n589 & n7151 ) | ( n589 & n7152 ) | ( n7151 & n7152 ) ;
  assign n7154 = x107 & n676 ;
  assign n7155 = n7153 | n7154 ;
  assign n7156 = ( x14 & n7150 ) | ( x14 & ~n7155 ) | ( n7150 & ~n7155 ) ;
  assign n7157 = ( ~x14 & n7155 ) | ( ~x14 & n7156 ) | ( n7155 & n7156 ) ;
  assign n7158 = ( ~n7150 & n7156 ) | ( ~n7150 & n7157 ) | ( n7156 & n7157 ) ;
  assign n7159 = n1297 & n3162 ;
  assign n7160 = x99 & n1301 ;
  assign n7161 = x100 | n7160 ;
  assign n7162 = ( n1303 & n7160 ) | ( n1303 & n7161 ) | ( n7160 & n7161 ) ;
  assign n7163 = x98 & n1426 ;
  assign n7164 = n7162 | n7163 ;
  assign n7165 = ( x23 & n7159 ) | ( x23 & ~n7164 ) | ( n7159 & ~n7164 ) ;
  assign n7166 = ( ~x23 & n7164 ) | ( ~x23 & n7165 ) | ( n7164 & n7165 ) ;
  assign n7167 = ( ~n7159 & n7165 ) | ( ~n7159 & n7166 ) | ( n7165 & n7166 ) ;
  assign n7168 = n1949 & n2294 ;
  assign n7169 = x93 & n1953 ;
  assign n7170 = x94 | n7169 ;
  assign n7171 = ( n1955 & n7169 ) | ( n1955 & n7170 ) | ( n7169 & n7170 ) ;
  assign n7172 = x92 & n2114 ;
  assign n7173 = n7171 | n7172 ;
  assign n7174 = ( x29 & n7168 ) | ( x29 & ~n7173 ) | ( n7168 & ~n7173 ) ;
  assign n7175 = ( ~x29 & n7173 ) | ( ~x29 & n7174 ) | ( n7173 & n7174 ) ;
  assign n7176 = ( ~n7168 & n7174 ) | ( ~n7168 & n7175 ) | ( n7174 & n7175 ) ;
  assign n7177 = n1262 & n3224 ;
  assign n7178 = x84 & n3228 ;
  assign n7179 = x85 | n7178 ;
  assign n7180 = ( n3230 & n7178 ) | ( n3230 & n7179 ) | ( n7178 & n7179 ) ;
  assign n7181 = x83 & n3413 ;
  assign n7182 = n7180 | n7181 ;
  assign n7183 = ( x38 & n7177 ) | ( x38 & ~n7182 ) | ( n7177 & ~n7182 ) ;
  assign n7184 = ( ~x38 & n7182 ) | ( ~x38 & n7183 ) | ( n7182 & n7183 ) ;
  assign n7185 = ( ~n7177 & n7183 ) | ( ~n7177 & n7184 ) | ( n7183 & n7184 ) ;
  assign n7186 = n990 & n3715 ;
  assign n7187 = x81 & n3719 ;
  assign n7188 = x82 | n7187 ;
  assign n7189 = ( n3721 & n7187 ) | ( n3721 & n7188 ) | ( n7187 & n7188 ) ;
  assign n7190 = x80 & n3922 ;
  assign n7191 = n7189 | n7190 ;
  assign n7192 = ( x41 & n7186 ) | ( x41 & ~n7191 ) | ( n7186 & ~n7191 ) ;
  assign n7193 = ( ~x41 & n7191 ) | ( ~x41 & n7192 ) | ( n7191 & n7192 ) ;
  assign n7194 = ( ~n7186 & n7192 ) | ( ~n7186 & n7193 ) | ( n7192 & n7193 ) ;
  assign n7195 = n701 & n4227 ;
  assign n7196 = x78 & n4231 ;
  assign n7197 = x79 | n7196 ;
  assign n7198 = ( n4233 & n7196 ) | ( n4233 & n7197 ) | ( n7196 & n7197 ) ;
  assign n7199 = x77 & n4470 ;
  assign n7200 = n7198 | n7199 ;
  assign n7201 = ( x44 & n7195 ) | ( x44 & ~n7200 ) | ( n7195 & ~n7200 ) ;
  assign n7202 = ( ~x44 & n7200 ) | ( ~x44 & n7201 ) | ( n7200 & n7201 ) ;
  assign n7203 = ( ~n7195 & n7201 ) | ( ~n7195 & n7202 ) | ( n7201 & n7202 ) ;
  assign n7204 = n554 & n4787 ;
  assign n7205 = x75 & n4791 ;
  assign n7206 = x76 | n7205 ;
  assign n7207 = ( n4793 & n7205 ) | ( n4793 & n7206 ) | ( n7205 & n7206 ) ;
  assign n7208 = x74 & n5030 ;
  assign n7209 = n7207 | n7208 ;
  assign n7210 = ( x47 & n7204 ) | ( x47 & ~n7209 ) | ( n7204 & ~n7209 ) ;
  assign n7211 = ( ~x47 & n7209 ) | ( ~x47 & n7210 ) | ( n7209 & n7210 ) ;
  assign n7212 = ( ~n7204 & n7210 ) | ( ~n7204 & n7211 ) | ( n7210 & n7211 ) ;
  assign n7213 = n390 & n5374 ;
  assign n7214 = x72 & n5378 ;
  assign n7215 = x73 | n7214 ;
  assign n7216 = ( n5380 & n7214 ) | ( n5380 & n7215 ) | ( n7214 & n7215 ) ;
  assign n7217 = x71 & n5638 ;
  assign n7218 = n7216 | n7217 ;
  assign n7219 = ( x50 & n7213 ) | ( x50 & ~n7218 ) | ( n7213 & ~n7218 ) ;
  assign n7220 = ( ~x50 & n7218 ) | ( ~x50 & n7219 ) | ( n7218 & n7219 ) ;
  assign n7221 = ( ~n7213 & n7219 ) | ( ~n7213 & n7220 ) | ( n7219 & n7220 ) ;
  assign n7222 = x66 & n6717 ;
  assign n7223 = x67 | n7222 ;
  assign n7224 = ( n6719 & n7222 ) | ( n6719 & n7223 ) | ( n7222 & n7223 ) ;
  assign n7225 = x65 & n6980 ;
  assign n7226 = n7224 | n7225 ;
  assign n7227 = n164 & n6713 ;
  assign n7228 = ( x56 & n7226 ) | ( x56 & ~n7227 ) | ( n7226 & ~n7227 ) ;
  assign n7229 = ( ~x56 & n7227 ) | ( ~x56 & n7228 ) | ( n7227 & n7228 ) ;
  assign n7230 = ( ~n7226 & n7228 ) | ( ~n7226 & n7229 ) | ( n7228 & n7229 ) ;
  assign n7231 = x56 & x57 ;
  assign n7232 = x56 | x57 ;
  assign n7233 = ~n7231 & n7232 ;
  assign n7234 = x64 & n7233 ;
  assign n7235 = x56 & ~n6988 ;
  assign n7236 = ( n7230 & n7234 ) | ( n7230 & n7235 ) | ( n7234 & n7235 ) ;
  assign n7237 = ( ~n7230 & n7234 ) | ( ~n7230 & n7235 ) | ( n7234 & n7235 ) ;
  assign n7238 = ( n7230 & ~n7236 ) | ( n7230 & n7237 ) | ( ~n7236 & n7237 ) ;
  assign n7239 = n245 & n6027 ;
  assign n7240 = x69 & n6031 ;
  assign n7241 = x70 | n7240 ;
  assign n7242 = ( n6033 & n7240 ) | ( n6033 & n7241 ) | ( n7240 & n7241 ) ;
  assign n7243 = x68 & n6303 ;
  assign n7244 = n7242 | n7243 ;
  assign n7245 = ( x53 & n7239 ) | ( x53 & ~n7244 ) | ( n7239 & ~n7244 ) ;
  assign n7246 = ( ~x53 & n7244 ) | ( ~x53 & n7245 ) | ( n7244 & n7245 ) ;
  assign n7247 = ( ~n7239 & n7245 ) | ( ~n7239 & n7246 ) | ( n7245 & n7246 ) ;
  assign n7248 = ( n6991 & n7238 ) | ( n6991 & n7247 ) | ( n7238 & n7247 ) ;
  assign n7249 = ( ~n6991 & n7238 ) | ( ~n6991 & n7247 ) | ( n7238 & n7247 ) ;
  assign n7250 = ( n6991 & ~n7248 ) | ( n6991 & n7249 ) | ( ~n7248 & n7249 ) ;
  assign n7251 = ( n6994 & n7221 ) | ( n6994 & n7250 ) | ( n7221 & n7250 ) ;
  assign n7252 = ( ~n6994 & n7221 ) | ( ~n6994 & n7250 ) | ( n7221 & n7250 ) ;
  assign n7253 = ( n6994 & ~n7251 ) | ( n6994 & n7252 ) | ( ~n7251 & n7252 ) ;
  assign n7254 = ( n6997 & n7212 ) | ( n6997 & n7253 ) | ( n7212 & n7253 ) ;
  assign n7255 = ( ~n6997 & n7212 ) | ( ~n6997 & n7253 ) | ( n7212 & n7253 ) ;
  assign n7256 = ( n6997 & ~n7254 ) | ( n6997 & n7255 ) | ( ~n7254 & n7255 ) ;
  assign n7257 = ( n7009 & n7203 ) | ( n7009 & n7256 ) | ( n7203 & n7256 ) ;
  assign n7258 = ( ~n7009 & n7203 ) | ( ~n7009 & n7256 ) | ( n7203 & n7256 ) ;
  assign n7259 = ( n7009 & ~n7257 ) | ( n7009 & n7258 ) | ( ~n7257 & n7258 ) ;
  assign n7260 = ( n7012 & n7194 ) | ( n7012 & n7259 ) | ( n7194 & n7259 ) ;
  assign n7261 = ( ~n7012 & n7194 ) | ( ~n7012 & n7259 ) | ( n7194 & n7259 ) ;
  assign n7262 = ( n7012 & ~n7260 ) | ( n7012 & n7261 ) | ( ~n7260 & n7261 ) ;
  assign n7263 = ( n7015 & n7185 ) | ( n7015 & n7262 ) | ( n7185 & n7262 ) ;
  assign n7264 = ( ~n7015 & n7185 ) | ( ~n7015 & n7262 ) | ( n7185 & n7262 ) ;
  assign n7265 = ( n7015 & ~n7263 ) | ( n7015 & n7264 ) | ( ~n7263 & n7264 ) ;
  assign n7266 = n1481 & n2766 ;
  assign n7267 = x87 & n2770 ;
  assign n7268 = x88 | n7267 ;
  assign n7269 = ( n2772 & n7267 ) | ( n2772 & n7268 ) | ( n7267 & n7268 ) ;
  assign n7270 = x86 & n2943 ;
  assign n7271 = n7269 | n7270 ;
  assign n7272 = ( x35 & n7266 ) | ( x35 & ~n7271 ) | ( n7266 & ~n7271 ) ;
  assign n7273 = ( ~x35 & n7271 ) | ( ~x35 & n7272 ) | ( n7271 & n7272 ) ;
  assign n7274 = ( ~n7266 & n7272 ) | ( ~n7266 & n7273 ) | ( n7272 & n7273 ) ;
  assign n7275 = ( n7018 & n7265 ) | ( n7018 & n7274 ) | ( n7265 & n7274 ) ;
  assign n7276 = ( ~n7018 & n7265 ) | ( ~n7018 & n7274 ) | ( n7265 & n7274 ) ;
  assign n7277 = ( n7018 & ~n7275 ) | ( n7018 & n7276 ) | ( ~n7275 & n7276 ) ;
  assign n7278 = n1914 & n2320 ;
  assign n7279 = x90 & n2324 ;
  assign n7280 = x91 | n7279 ;
  assign n7281 = ( n2326 & n7279 ) | ( n2326 & n7280 ) | ( n7279 & n7280 ) ;
  assign n7282 = x89 & n2497 ;
  assign n7283 = n7281 | n7282 ;
  assign n7284 = ( x32 & n7278 ) | ( x32 & ~n7283 ) | ( n7278 & ~n7283 ) ;
  assign n7285 = ( ~x32 & n7283 ) | ( ~x32 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7286 = ( ~n7278 & n7284 ) | ( ~n7278 & n7285 ) | ( n7284 & n7285 ) ;
  assign n7287 = ( n7030 & n7277 ) | ( n7030 & n7286 ) | ( n7277 & n7286 ) ;
  assign n7288 = ( ~n7030 & n7277 ) | ( ~n7030 & n7286 ) | ( n7277 & n7286 ) ;
  assign n7289 = ( n7030 & ~n7287 ) | ( n7030 & n7288 ) | ( ~n7287 & n7288 ) ;
  assign n7290 = ( n7033 & n7176 ) | ( n7033 & n7289 ) | ( n7176 & n7289 ) ;
  assign n7291 = ( ~n7033 & n7176 ) | ( ~n7033 & n7289 ) | ( n7176 & n7289 ) ;
  assign n7292 = ( n7033 & ~n7290 ) | ( n7033 & n7291 ) | ( ~n7290 & n7291 ) ;
  assign n7293 = n1617 & n2585 ;
  assign n7294 = x96 & n1621 ;
  assign n7295 = x97 | n7294 ;
  assign n7296 = ( n1623 & n7294 ) | ( n1623 & n7295 ) | ( n7294 & n7295 ) ;
  assign n7297 = x95 & n1749 ;
  assign n7298 = n7296 | n7297 ;
  assign n7299 = ( x26 & n7293 ) | ( x26 & ~n7298 ) | ( n7293 & ~n7298 ) ;
  assign n7300 = ( ~x26 & n7298 ) | ( ~x26 & n7299 ) | ( n7298 & n7299 ) ;
  assign n7301 = ( ~n7293 & n7299 ) | ( ~n7293 & n7300 ) | ( n7299 & n7300 ) ;
  assign n7302 = ( n7036 & n7292 ) | ( n7036 & n7301 ) | ( n7292 & n7301 ) ;
  assign n7303 = ( ~n7036 & n7292 ) | ( ~n7036 & n7301 ) | ( n7292 & n7301 ) ;
  assign n7304 = ( n7036 & ~n7302 ) | ( n7036 & n7303 ) | ( ~n7302 & n7303 ) ;
  assign n7305 = ( n7048 & n7167 ) | ( n7048 & n7304 ) | ( n7167 & n7304 ) ;
  assign n7306 = ( ~n7048 & n7167 ) | ( ~n7048 & n7304 ) | ( n7167 & n7304 ) ;
  assign n7307 = ( n7048 & ~n7305 ) | ( n7048 & n7306 ) | ( ~n7305 & n7306 ) ;
  assign n7308 = n1016 & n3650 ;
  assign n7309 = x102 & n1020 ;
  assign n7310 = x103 | n7309 ;
  assign n7311 = ( n1022 & n7309 ) | ( n1022 & n7310 ) | ( n7309 & n7310 ) ;
  assign n7312 = x101 & n1145 ;
  assign n7313 = n7311 | n7312 ;
  assign n7314 = ( x20 & n7308 ) | ( x20 & ~n7313 ) | ( n7308 & ~n7313 ) ;
  assign n7315 = ( ~x20 & n7313 ) | ( ~x20 & n7314 ) | ( n7313 & n7314 ) ;
  assign n7316 = ( ~n7308 & n7314 ) | ( ~n7308 & n7315 ) | ( n7314 & n7315 ) ;
  assign n7317 = ( n7060 & n7307 ) | ( n7060 & n7316 ) | ( n7307 & n7316 ) ;
  assign n7318 = ( ~n7060 & n7307 ) | ( ~n7060 & n7316 ) | ( n7307 & n7316 ) ;
  assign n7319 = ( n7060 & ~n7317 ) | ( n7060 & n7318 ) | ( ~n7317 & n7318 ) ;
  assign n7320 = n810 & n4013 ;
  assign n7321 = x105 & n814 ;
  assign n7322 = x106 | n7321 ;
  assign n7323 = ( n816 & n7321 ) | ( n816 & n7322 ) | ( n7321 & n7322 ) ;
  assign n7324 = x104 & n885 ;
  assign n7325 = n7323 | n7324 ;
  assign n7326 = ( x17 & n7320 ) | ( x17 & ~n7325 ) | ( n7320 & ~n7325 ) ;
  assign n7327 = ( ~x17 & n7325 ) | ( ~x17 & n7326 ) | ( n7325 & n7326 ) ;
  assign n7328 = ( ~n7320 & n7326 ) | ( ~n7320 & n7327 ) | ( n7326 & n7327 ) ;
  assign n7329 = ( n7072 & n7319 ) | ( n7072 & n7328 ) | ( n7319 & n7328 ) ;
  assign n7330 = ( ~n7072 & n7319 ) | ( ~n7072 & n7328 ) | ( n7319 & n7328 ) ;
  assign n7331 = ( n7072 & ~n7329 ) | ( n7072 & n7330 ) | ( ~n7329 & n7330 ) ;
  assign n7332 = ( n7084 & n7158 ) | ( n7084 & n7331 ) | ( n7158 & n7331 ) ;
  assign n7333 = ( ~n7084 & n7158 ) | ( ~n7084 & n7331 ) | ( n7158 & n7331 ) ;
  assign n7334 = ( n7084 & ~n7332 ) | ( n7084 & n7333 ) | ( ~n7332 & n7333 ) ;
  assign n7335 = ( n7087 & n7149 ) | ( n7087 & n7334 ) | ( n7149 & n7334 ) ;
  assign n7336 = ( ~n7087 & n7149 ) | ( ~n7087 & n7334 ) | ( n7149 & n7334 ) ;
  assign n7337 = ( n7087 & ~n7335 ) | ( n7087 & n7336 ) | ( ~n7335 & n7336 ) ;
  assign n7338 = ( n7090 & n7140 ) | ( n7090 & n7337 ) | ( n7140 & n7337 ) ;
  assign n7339 = ( ~n7090 & n7140 ) | ( ~n7090 & n7337 ) | ( n7140 & n7337 ) ;
  assign n7340 = ( n7090 & ~n7338 ) | ( n7090 & n7339 ) | ( ~n7338 & n7339 ) ;
  assign n7341 = ( n7093 & n7131 ) | ( n7093 & n7340 ) | ( n7131 & n7340 ) ;
  assign n7342 = ( ~n7093 & n7131 ) | ( ~n7093 & n7340 ) | ( n7131 & n7340 ) ;
  assign n7343 = ( n7093 & ~n7341 ) | ( n7093 & n7342 ) | ( ~n7341 & n7342 ) ;
  assign n7344 = ( n7108 & n7122 ) | ( n7108 & n7343 ) | ( n7122 & n7343 ) ;
  assign n7345 = ( ~n7108 & n7122 ) | ( ~n7108 & n7343 ) | ( n7122 & n7343 ) ;
  assign n7346 = ( n7108 & ~n7344 ) | ( n7108 & n7345 ) | ( ~n7344 & n7345 ) ;
  assign n7347 = n186 & n6645 ;
  assign n7348 = x118 & n190 ;
  assign n7349 = x119 | n7348 ;
  assign n7350 = ( n192 & n7348 ) | ( n192 & n7349 ) | ( n7348 & n7349 ) ;
  assign n7351 = x117 & n220 ;
  assign n7352 = n7350 | n7351 ;
  assign n7353 = ( x5 & n7347 ) | ( x5 & ~n7352 ) | ( n7347 & ~n7352 ) ;
  assign n7354 = ( ~x5 & n7352 ) | ( ~x5 & n7353 ) | ( n7352 & n7353 ) ;
  assign n7355 = ( ~n7347 & n7353 ) | ( ~n7347 & n7354 ) | ( n7353 & n7354 ) ;
  assign n7356 = n291 & n5977 ;
  assign n7357 = x115 & n295 ;
  assign n7358 = x116 | n7357 ;
  assign n7359 = ( n297 & n7357 ) | ( n297 & n7358 ) | ( n7357 & n7358 ) ;
  assign n7360 = x114 & n330 ;
  assign n7361 = n7359 | n7360 ;
  assign n7362 = ( x8 & n7356 ) | ( x8 & ~n7361 ) | ( n7356 & ~n7361 ) ;
  assign n7363 = ( ~x8 & n7361 ) | ( ~x8 & n7362 ) | ( n7361 & n7362 ) ;
  assign n7364 = ( ~n7356 & n7362 ) | ( ~n7356 & n7363 ) | ( n7362 & n7363 ) ;
  assign n7365 = n407 & n5542 ;
  assign n7366 = x112 & n411 ;
  assign n7367 = x113 | n7366 ;
  assign n7368 = ( n413 & n7366 ) | ( n413 & n7367 ) | ( n7366 & n7367 ) ;
  assign n7369 = x111 & n491 ;
  assign n7370 = n7368 | n7369 ;
  assign n7371 = ( x11 & n7365 ) | ( x11 & ~n7370 ) | ( n7365 & ~n7370 ) ;
  assign n7372 = ( ~x11 & n7370 ) | ( ~x11 & n7371 ) | ( n7370 & n7371 ) ;
  assign n7373 = ( ~n7365 & n7371 ) | ( ~n7365 & n7372 ) | ( n7371 & n7372 ) ;
  assign n7374 = n583 & n4934 ;
  assign n7375 = x109 & n587 ;
  assign n7376 = x110 | n7375 ;
  assign n7377 = ( n589 & n7375 ) | ( n589 & n7376 ) | ( n7375 & n7376 ) ;
  assign n7378 = x108 & n676 ;
  assign n7379 = n7377 | n7378 ;
  assign n7380 = ( x14 & n7374 ) | ( x14 & ~n7379 ) | ( n7374 & ~n7379 ) ;
  assign n7381 = ( ~x14 & n7379 ) | ( ~x14 & n7380 ) | ( n7379 & n7380 ) ;
  assign n7382 = ( ~n7374 & n7380 ) | ( ~n7374 & n7381 ) | ( n7380 & n7381 ) ;
  assign n7383 = n1949 & n2434 ;
  assign n7384 = x94 & n1953 ;
  assign n7385 = x95 | n7384 ;
  assign n7386 = ( n1955 & n7384 ) | ( n1955 & n7385 ) | ( n7384 & n7385 ) ;
  assign n7387 = x93 & n2114 ;
  assign n7388 = n7386 | n7387 ;
  assign n7389 = ( x29 & n7383 ) | ( x29 & ~n7388 ) | ( n7383 & ~n7388 ) ;
  assign n7390 = ( ~x29 & n7388 ) | ( ~x29 & n7389 ) | ( n7388 & n7389 ) ;
  assign n7391 = ( ~n7383 & n7389 ) | ( ~n7383 & n7390 ) | ( n7389 & n7390 ) ;
  assign n7392 = n1366 & n3224 ;
  assign n7393 = x85 & n3228 ;
  assign n7394 = x86 | n7393 ;
  assign n7395 = ( n3230 & n7393 ) | ( n3230 & n7394 ) | ( n7393 & n7394 ) ;
  assign n7396 = x84 & n3413 ;
  assign n7397 = n7395 | n7396 ;
  assign n7398 = ( x38 & n7392 ) | ( x38 & ~n7397 ) | ( n7392 & ~n7397 ) ;
  assign n7399 = ( ~x38 & n7397 ) | ( ~x38 & n7398 ) | ( n7397 & n7398 ) ;
  assign n7400 = ( ~n7392 & n7398 ) | ( ~n7392 & n7399 ) | ( n7398 & n7399 ) ;
  assign n7401 = n769 & n4227 ;
  assign n7402 = x79 & n4231 ;
  assign n7403 = x80 | n7402 ;
  assign n7404 = ( n4233 & n7402 ) | ( n4233 & n7403 ) | ( n7402 & n7403 ) ;
  assign n7405 = x78 & n4470 ;
  assign n7406 = n7404 | n7405 ;
  assign n7407 = ( x44 & n7401 ) | ( x44 & ~n7406 ) | ( n7401 & ~n7406 ) ;
  assign n7408 = ( ~x44 & n7406 ) | ( ~x44 & n7407 ) | ( n7406 & n7407 ) ;
  assign n7409 = ( ~n7401 & n7407 ) | ( ~n7401 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7410 = n277 & n6027 ;
  assign n7411 = x70 & n6031 ;
  assign n7412 = x71 | n7411 ;
  assign n7413 = ( n6033 & n7411 ) | ( n6033 & n7412 ) | ( n7411 & n7412 ) ;
  assign n7414 = x69 & n6303 ;
  assign n7415 = n7413 | n7414 ;
  assign n7416 = ( x53 & n7410 ) | ( x53 & ~n7415 ) | ( n7410 & ~n7415 ) ;
  assign n7417 = ( ~x53 & n7415 ) | ( ~x53 & n7416 ) | ( n7415 & n7416 ) ;
  assign n7418 = ( ~n7410 & n7416 ) | ( ~n7410 & n7417 ) | ( n7416 & n7417 ) ;
  assign n7419 = x59 & n7234 ;
  assign n7420 = x58 | x59 ;
  assign n7421 = ( x58 & x59 ) | ( x58 & ~n7420 ) | ( x59 & ~n7420 ) ;
  assign n7422 = n7420 & ~n7421 ;
  assign n7423 = n7233 & n7422 ;
  assign n7424 = n133 & n7423 ;
  assign n7425 = ~x56 & x58 ;
  assign n7426 = x57 & x58 ;
  assign n7427 = ( n7231 & n7425 ) | ( n7231 & ~n7426 ) | ( n7425 & ~n7426 ) ;
  assign n7428 = x64 & n7427 ;
  assign n7429 = ( n7233 & ~n7420 ) | ( n7233 & n7421 ) | ( ~n7420 & n7421 ) ;
  assign n7430 = x65 | n7428 ;
  assign n7431 = ( n7428 & n7429 ) | ( n7428 & n7430 ) | ( n7429 & n7430 ) ;
  assign n7432 = ( n7419 & n7424 ) | ( n7419 & n7431 ) | ( n7424 & n7431 ) ;
  assign n7433 = n7424 | n7431 ;
  assign n7434 = ~n7419 & n7433 ;
  assign n7435 = ( n7419 & ~n7432 ) | ( n7419 & n7434 ) | ( ~n7432 & n7434 ) ;
  assign n7436 = x67 & n6717 ;
  assign n7437 = x68 | n7436 ;
  assign n7438 = ( n6719 & n7436 ) | ( n6719 & n7437 ) | ( n7436 & n7437 ) ;
  assign n7439 = x66 & n6980 ;
  assign n7440 = n7438 | n7439 ;
  assign n7441 = n201 & n6713 ;
  assign n7442 = ( x56 & n7440 ) | ( x56 & ~n7441 ) | ( n7440 & ~n7441 ) ;
  assign n7443 = ( ~x56 & n7441 ) | ( ~x56 & n7442 ) | ( n7441 & n7442 ) ;
  assign n7444 = ( ~n7440 & n7442 ) | ( ~n7440 & n7443 ) | ( n7442 & n7443 ) ;
  assign n7445 = ( n7236 & n7435 ) | ( n7236 & n7444 ) | ( n7435 & n7444 ) ;
  assign n7446 = ( ~n7236 & n7435 ) | ( ~n7236 & n7444 ) | ( n7435 & n7444 ) ;
  assign n7447 = ( n7236 & ~n7445 ) | ( n7236 & n7446 ) | ( ~n7445 & n7446 ) ;
  assign n7448 = ( n7248 & n7418 ) | ( n7248 & n7447 ) | ( n7418 & n7447 ) ;
  assign n7449 = ( ~n7248 & n7418 ) | ( ~n7248 & n7447 ) | ( n7418 & n7447 ) ;
  assign n7450 = ( n7248 & ~n7448 ) | ( n7248 & n7449 ) | ( ~n7448 & n7449 ) ;
  assign n7451 = n446 & n5374 ;
  assign n7452 = x73 & n5378 ;
  assign n7453 = x74 | n7452 ;
  assign n7454 = ( n5380 & n7452 ) | ( n5380 & n7453 ) | ( n7452 & n7453 ) ;
  assign n7455 = x72 & n5638 ;
  assign n7456 = n7454 | n7455 ;
  assign n7457 = ( x50 & n7451 ) | ( x50 & ~n7456 ) | ( n7451 & ~n7456 ) ;
  assign n7458 = ( ~x50 & n7456 ) | ( ~x50 & n7457 ) | ( n7456 & n7457 ) ;
  assign n7459 = ( ~n7451 & n7457 ) | ( ~n7451 & n7458 ) | ( n7457 & n7458 ) ;
  assign n7460 = ( n7251 & n7450 ) | ( n7251 & n7459 ) | ( n7450 & n7459 ) ;
  assign n7461 = ( ~n7251 & n7450 ) | ( ~n7251 & n7459 ) | ( n7450 & n7459 ) ;
  assign n7462 = ( n7251 & ~n7460 ) | ( n7251 & n7461 ) | ( ~n7460 & n7461 ) ;
  assign n7463 = n569 & n4787 ;
  assign n7464 = x76 & n4791 ;
  assign n7465 = x77 | n7464 ;
  assign n7466 = ( n4793 & n7464 ) | ( n4793 & n7465 ) | ( n7464 & n7465 ) ;
  assign n7467 = x75 & n5030 ;
  assign n7468 = n7466 | n7467 ;
  assign n7469 = ( x47 & n7463 ) | ( x47 & ~n7468 ) | ( n7463 & ~n7468 ) ;
  assign n7470 = ( ~x47 & n7468 ) | ( ~x47 & n7469 ) | ( n7468 & n7469 ) ;
  assign n7471 = ( ~n7463 & n7469 ) | ( ~n7463 & n7470 ) | ( n7469 & n7470 ) ;
  assign n7472 = ( n7254 & n7462 ) | ( n7254 & n7471 ) | ( n7462 & n7471 ) ;
  assign n7473 = ( ~n7254 & n7462 ) | ( ~n7254 & n7471 ) | ( n7462 & n7471 ) ;
  assign n7474 = ( n7254 & ~n7472 ) | ( n7254 & n7473 ) | ( ~n7472 & n7473 ) ;
  assign n7475 = ( n7257 & n7409 ) | ( n7257 & n7474 ) | ( n7409 & n7474 ) ;
  assign n7476 = ( ~n7257 & n7409 ) | ( ~n7257 & n7474 ) | ( n7409 & n7474 ) ;
  assign n7477 = ( n7257 & ~n7475 ) | ( n7257 & n7476 ) | ( ~n7475 & n7476 ) ;
  assign n7478 = n1082 & n3715 ;
  assign n7479 = x82 & n3719 ;
  assign n7480 = x83 | n7479 ;
  assign n7481 = ( n3721 & n7479 ) | ( n3721 & n7480 ) | ( n7479 & n7480 ) ;
  assign n7482 = x81 & n3922 ;
  assign n7483 = n7481 | n7482 ;
  assign n7484 = ( x41 & n7478 ) | ( x41 & ~n7483 ) | ( n7478 & ~n7483 ) ;
  assign n7485 = ( ~x41 & n7483 ) | ( ~x41 & n7484 ) | ( n7483 & n7484 ) ;
  assign n7486 = ( ~n7478 & n7484 ) | ( ~n7478 & n7485 ) | ( n7484 & n7485 ) ;
  assign n7487 = ( n7260 & n7477 ) | ( n7260 & n7486 ) | ( n7477 & n7486 ) ;
  assign n7488 = ( ~n7260 & n7477 ) | ( ~n7260 & n7486 ) | ( n7477 & n7486 ) ;
  assign n7489 = ( n7260 & ~n7487 ) | ( n7260 & n7488 ) | ( ~n7487 & n7488 ) ;
  assign n7490 = ( n7263 & n7400 ) | ( n7263 & n7489 ) | ( n7400 & n7489 ) ;
  assign n7491 = ( ~n7263 & n7400 ) | ( ~n7263 & n7489 ) | ( n7400 & n7489 ) ;
  assign n7492 = ( n7263 & ~n7490 ) | ( n7263 & n7491 ) | ( ~n7490 & n7491 ) ;
  assign n7493 = n1585 & n2766 ;
  assign n7494 = x88 & n2770 ;
  assign n7495 = x89 | n7494 ;
  assign n7496 = ( n2772 & n7494 ) | ( n2772 & n7495 ) | ( n7494 & n7495 ) ;
  assign n7497 = x87 & n2943 ;
  assign n7498 = n7496 | n7497 ;
  assign n7499 = ( x35 & n7493 ) | ( x35 & ~n7498 ) | ( n7493 & ~n7498 ) ;
  assign n7500 = ( ~x35 & n7498 ) | ( ~x35 & n7499 ) | ( n7498 & n7499 ) ;
  assign n7501 = ( ~n7493 & n7499 ) | ( ~n7493 & n7500 ) | ( n7499 & n7500 ) ;
  assign n7502 = ( n7275 & n7492 ) | ( n7275 & n7501 ) | ( n7492 & n7501 ) ;
  assign n7503 = ( ~n7275 & n7492 ) | ( ~n7275 & n7501 ) | ( n7492 & n7501 ) ;
  assign n7504 = ( n7275 & ~n7502 ) | ( n7275 & n7503 ) | ( ~n7502 & n7503 ) ;
  assign n7505 = n2042 & n2320 ;
  assign n7506 = x91 & n2324 ;
  assign n7507 = x92 | n7506 ;
  assign n7508 = ( n2326 & n7506 ) | ( n2326 & n7507 ) | ( n7506 & n7507 ) ;
  assign n7509 = x90 & n2497 ;
  assign n7510 = n7508 | n7509 ;
  assign n7511 = ( x32 & n7505 ) | ( x32 & ~n7510 ) | ( n7505 & ~n7510 ) ;
  assign n7512 = ( ~x32 & n7510 ) | ( ~x32 & n7511 ) | ( n7510 & n7511 ) ;
  assign n7513 = ( ~n7505 & n7511 ) | ( ~n7505 & n7512 ) | ( n7511 & n7512 ) ;
  assign n7514 = ( n7287 & n7504 ) | ( n7287 & n7513 ) | ( n7504 & n7513 ) ;
  assign n7515 = ( ~n7287 & n7504 ) | ( ~n7287 & n7513 ) | ( n7504 & n7513 ) ;
  assign n7516 = ( n7287 & ~n7514 ) | ( n7287 & n7515 ) | ( ~n7514 & n7515 ) ;
  assign n7517 = ( n7290 & n7391 ) | ( n7290 & n7516 ) | ( n7391 & n7516 ) ;
  assign n7518 = ( ~n7290 & n7391 ) | ( ~n7290 & n7516 ) | ( n7391 & n7516 ) ;
  assign n7519 = ( n7290 & ~n7517 ) | ( n7290 & n7518 ) | ( ~n7517 & n7518 ) ;
  assign n7520 = n1617 & n2725 ;
  assign n7521 = x97 & n1621 ;
  assign n7522 = x98 | n7521 ;
  assign n7523 = ( n1623 & n7521 ) | ( n1623 & n7522 ) | ( n7521 & n7522 ) ;
  assign n7524 = x96 & n1749 ;
  assign n7525 = n7523 | n7524 ;
  assign n7526 = ( x26 & n7520 ) | ( x26 & ~n7525 ) | ( n7520 & ~n7525 ) ;
  assign n7527 = ( ~x26 & n7525 ) | ( ~x26 & n7526 ) | ( n7525 & n7526 ) ;
  assign n7528 = ( ~n7520 & n7526 ) | ( ~n7520 & n7527 ) | ( n7526 & n7527 ) ;
  assign n7529 = ( n7302 & n7519 ) | ( n7302 & n7528 ) | ( n7519 & n7528 ) ;
  assign n7530 = ( ~n7302 & n7519 ) | ( ~n7302 & n7528 ) | ( n7519 & n7528 ) ;
  assign n7531 = ( n7302 & ~n7529 ) | ( n7302 & n7530 ) | ( ~n7529 & n7530 ) ;
  assign n7532 = n1297 & n3326 ;
  assign n7533 = x100 & n1301 ;
  assign n7534 = x101 | n7533 ;
  assign n7535 = ( n1303 & n7533 ) | ( n1303 & n7534 ) | ( n7533 & n7534 ) ;
  assign n7536 = x99 & n1426 ;
  assign n7537 = n7535 | n7536 ;
  assign n7538 = ( x23 & n7532 ) | ( x23 & ~n7537 ) | ( n7532 & ~n7537 ) ;
  assign n7539 = ( ~x23 & n7537 ) | ( ~x23 & n7538 ) | ( n7537 & n7538 ) ;
  assign n7540 = ( ~n7532 & n7538 ) | ( ~n7532 & n7539 ) | ( n7538 & n7539 ) ;
  assign n7541 = ( n7305 & n7531 ) | ( n7305 & n7540 ) | ( n7531 & n7540 ) ;
  assign n7542 = ( ~n7305 & n7531 ) | ( ~n7305 & n7540 ) | ( n7531 & n7540 ) ;
  assign n7543 = ( n7305 & ~n7541 ) | ( n7305 & n7542 ) | ( ~n7541 & n7542 ) ;
  assign n7544 = n1016 & n3665 ;
  assign n7545 = x103 & n1020 ;
  assign n7546 = x104 | n7545 ;
  assign n7547 = ( n1022 & n7545 ) | ( n1022 & n7546 ) | ( n7545 & n7546 ) ;
  assign n7548 = x102 & n1145 ;
  assign n7549 = n7547 | n7548 ;
  assign n7550 = ( x20 & n7544 ) | ( x20 & ~n7549 ) | ( n7544 & ~n7549 ) ;
  assign n7551 = ( ~x20 & n7549 ) | ( ~x20 & n7550 ) | ( n7549 & n7550 ) ;
  assign n7552 = ( ~n7544 & n7550 ) | ( ~n7544 & n7551 ) | ( n7550 & n7551 ) ;
  assign n7553 = ( n7317 & n7543 ) | ( n7317 & n7552 ) | ( n7543 & n7552 ) ;
  assign n7554 = ( ~n7317 & n7543 ) | ( ~n7317 & n7552 ) | ( n7543 & n7552 ) ;
  assign n7555 = ( n7317 & ~n7553 ) | ( n7317 & n7554 ) | ( ~n7553 & n7554 ) ;
  assign n7556 = n810 & n4362 ;
  assign n7557 = x106 & n814 ;
  assign n7558 = x107 | n7557 ;
  assign n7559 = ( n816 & n7557 ) | ( n816 & n7558 ) | ( n7557 & n7558 ) ;
  assign n7560 = x105 & n885 ;
  assign n7561 = n7559 | n7560 ;
  assign n7562 = ( x17 & n7556 ) | ( x17 & ~n7561 ) | ( n7556 & ~n7561 ) ;
  assign n7563 = ( ~x17 & n7561 ) | ( ~x17 & n7562 ) | ( n7561 & n7562 ) ;
  assign n7564 = ( ~n7556 & n7562 ) | ( ~n7556 & n7563 ) | ( n7562 & n7563 ) ;
  assign n7565 = ( n7329 & n7555 ) | ( n7329 & n7564 ) | ( n7555 & n7564 ) ;
  assign n7566 = ( ~n7329 & n7555 ) | ( ~n7329 & n7564 ) | ( n7555 & n7564 ) ;
  assign n7567 = ( n7329 & ~n7565 ) | ( n7329 & n7566 ) | ( ~n7565 & n7566 ) ;
  assign n7568 = ( n7332 & n7382 ) | ( n7332 & n7567 ) | ( n7382 & n7567 ) ;
  assign n7569 = ( ~n7332 & n7382 ) | ( ~n7332 & n7567 ) | ( n7382 & n7567 ) ;
  assign n7570 = ( n7332 & ~n7568 ) | ( n7332 & n7569 ) | ( ~n7568 & n7569 ) ;
  assign n7571 = ( n7335 & n7373 ) | ( n7335 & n7570 ) | ( n7373 & n7570 ) ;
  assign n7572 = ( ~n7335 & n7373 ) | ( ~n7335 & n7570 ) | ( n7373 & n7570 ) ;
  assign n7573 = ( n7335 & ~n7571 ) | ( n7335 & n7572 ) | ( ~n7571 & n7572 ) ;
  assign n7574 = ( n7338 & n7364 ) | ( n7338 & n7573 ) | ( n7364 & n7573 ) ;
  assign n7575 = ( ~n7338 & n7364 ) | ( ~n7338 & n7573 ) | ( n7364 & n7573 ) ;
  assign n7576 = ( n7338 & ~n7574 ) | ( n7338 & n7575 ) | ( ~n7574 & n7575 ) ;
  assign n7577 = ( n7341 & n7355 ) | ( n7341 & n7576 ) | ( n7355 & n7576 ) ;
  assign n7578 = ( ~n7341 & n7355 ) | ( ~n7341 & n7576 ) | ( n7355 & n7576 ) ;
  assign n7579 = ( n7341 & ~n7577 ) | ( n7341 & n7578 ) | ( ~n7577 & n7578 ) ;
  assign n7580 = ( x121 & x122 ) | ( x121 & n7111 ) | ( x122 & n7111 ) ;
  assign n7581 = ( x121 & ~x122 ) | ( x121 & n7111 ) | ( ~x122 & n7111 ) ;
  assign n7582 = ( x122 & ~n7580 ) | ( x122 & n7581 ) | ( ~n7580 & n7581 ) ;
  assign n7583 = n136 & n7582 ;
  assign n7584 = x121 & n138 ;
  assign n7585 = x122 | n7584 ;
  assign n7586 = ( n141 & n7584 ) | ( n141 & n7585 ) | ( n7584 & n7585 ) ;
  assign n7587 = x120 & n154 ;
  assign n7588 = n7586 | n7587 ;
  assign n7589 = ( x2 & n7583 ) | ( x2 & ~n7588 ) | ( n7583 & ~n7588 ) ;
  assign n7590 = ( ~x2 & n7588 ) | ( ~x2 & n7589 ) | ( n7588 & n7589 ) ;
  assign n7591 = ( ~n7583 & n7589 ) | ( ~n7583 & n7590 ) | ( n7589 & n7590 ) ;
  assign n7592 = ( n7344 & n7579 ) | ( n7344 & n7591 ) | ( n7579 & n7591 ) ;
  assign n7593 = ( ~n7344 & n7579 ) | ( ~n7344 & n7591 ) | ( n7579 & n7591 ) ;
  assign n7594 = ( n7344 & ~n7592 ) | ( n7344 & n7593 ) | ( ~n7592 & n7593 ) ;
  assign n7595 = ( x122 & x123 ) | ( x122 & n7580 ) | ( x123 & n7580 ) ;
  assign n7596 = ( x122 & ~x123 ) | ( x122 & n7580 ) | ( ~x123 & n7580 ) ;
  assign n7597 = ( x123 & ~n7595 ) | ( x123 & n7596 ) | ( ~n7595 & n7596 ) ;
  assign n7598 = n136 & n7597 ;
  assign n7599 = x122 & n138 ;
  assign n7600 = x123 | n7599 ;
  assign n7601 = ( n141 & n7599 ) | ( n141 & n7600 ) | ( n7599 & n7600 ) ;
  assign n7602 = x121 & n154 ;
  assign n7603 = n7601 | n7602 ;
  assign n7604 = ( x2 & n7598 ) | ( x2 & ~n7603 ) | ( n7598 & ~n7603 ) ;
  assign n7605 = ( ~x2 & n7603 ) | ( ~x2 & n7604 ) | ( n7603 & n7604 ) ;
  assign n7606 = ( ~n7598 & n7604 ) | ( ~n7598 & n7605 ) | ( n7604 & n7605 ) ;
  assign n7607 = n186 & n7098 ;
  assign n7608 = x119 & n190 ;
  assign n7609 = x120 | n7608 ;
  assign n7610 = ( n192 & n7608 ) | ( n192 & n7609 ) | ( n7608 & n7609 ) ;
  assign n7611 = x118 & n220 ;
  assign n7612 = n7610 | n7611 ;
  assign n7613 = ( x5 & n7607 ) | ( x5 & ~n7612 ) | ( n7607 & ~n7612 ) ;
  assign n7614 = ( ~x5 & n7612 ) | ( ~x5 & n7613 ) | ( n7612 & n7613 ) ;
  assign n7615 = ( ~n7607 & n7613 ) | ( ~n7607 & n7614 ) | ( n7613 & n7614 ) ;
  assign n7616 = n291 & n6201 ;
  assign n7617 = x116 & n295 ;
  assign n7618 = x117 | n7617 ;
  assign n7619 = ( n297 & n7617 ) | ( n297 & n7618 ) | ( n7617 & n7618 ) ;
  assign n7620 = x115 & n330 ;
  assign n7621 = n7619 | n7620 ;
  assign n7622 = ( x8 & n7616 ) | ( x8 & ~n7621 ) | ( n7616 & ~n7621 ) ;
  assign n7623 = ( ~x8 & n7621 ) | ( ~x8 & n7622 ) | ( n7621 & n7622 ) ;
  assign n7624 = ( ~n7616 & n7622 ) | ( ~n7616 & n7623 ) | ( n7622 & n7623 ) ;
  assign n7625 = n583 & n5130 ;
  assign n7626 = x110 & n587 ;
  assign n7627 = x111 | n7626 ;
  assign n7628 = ( n589 & n7626 ) | ( n589 & n7627 ) | ( n7626 & n7627 ) ;
  assign n7629 = x109 & n676 ;
  assign n7630 = n7628 | n7629 ;
  assign n7631 = ( x14 & n7625 ) | ( x14 & ~n7630 ) | ( n7625 & ~n7630 ) ;
  assign n7632 = ( ~x14 & n7630 ) | ( ~x14 & n7631 ) | ( n7630 & n7631 ) ;
  assign n7633 = ( ~n7625 & n7631 ) | ( ~n7625 & n7632 ) | ( n7631 & n7632 ) ;
  assign n7634 = n810 & n4377 ;
  assign n7635 = x107 & n814 ;
  assign n7636 = x108 | n7635 ;
  assign n7637 = ( n816 & n7635 ) | ( n816 & n7636 ) | ( n7635 & n7636 ) ;
  assign n7638 = x106 & n885 ;
  assign n7639 = n7637 | n7638 ;
  assign n7640 = ( x17 & n7634 ) | ( x17 & ~n7639 ) | ( n7634 & ~n7639 ) ;
  assign n7641 = ( ~x17 & n7639 ) | ( ~x17 & n7640 ) | ( n7639 & n7640 ) ;
  assign n7642 = ( ~n7634 & n7640 ) | ( ~n7634 & n7641 ) | ( n7640 & n7641 ) ;
  assign n7643 = n1949 & n2449 ;
  assign n7644 = x95 & n1953 ;
  assign n7645 = x96 | n7644 ;
  assign n7646 = ( n1955 & n7644 ) | ( n1955 & n7645 ) | ( n7644 & n7645 ) ;
  assign n7647 = x94 & n2114 ;
  assign n7648 = n7646 | n7647 ;
  assign n7649 = ( x29 & n7643 ) | ( x29 & ~n7648 ) | ( n7643 & ~n7648 ) ;
  assign n7650 = ( ~x29 & n7648 ) | ( ~x29 & n7649 ) | ( n7648 & n7649 ) ;
  assign n7651 = ( ~n7643 & n7649 ) | ( ~n7643 & n7650 ) | ( n7649 & n7650 ) ;
  assign n7652 = n1466 & n3224 ;
  assign n7653 = x86 & n3228 ;
  assign n7654 = x87 | n7653 ;
  assign n7655 = ( n3230 & n7653 ) | ( n3230 & n7654 ) | ( n7653 & n7654 ) ;
  assign n7656 = x85 & n3413 ;
  assign n7657 = n7655 | n7656 ;
  assign n7658 = ( x38 & n7652 ) | ( x38 & ~n7657 ) | ( n7652 & ~n7657 ) ;
  assign n7659 = ( ~x38 & n7657 ) | ( ~x38 & n7658 ) | ( n7657 & n7658 ) ;
  assign n7660 = ( ~n7652 & n7658 ) | ( ~n7652 & n7659 ) | ( n7658 & n7659 ) ;
  assign n7661 = n1097 & n3715 ;
  assign n7662 = x83 & n3719 ;
  assign n7663 = x84 | n7662 ;
  assign n7664 = ( n3721 & n7662 ) | ( n3721 & n7663 ) | ( n7662 & n7663 ) ;
  assign n7665 = x82 & n3922 ;
  assign n7666 = n7664 | n7665 ;
  assign n7667 = ( x41 & n7661 ) | ( x41 & ~n7666 ) | ( n7661 & ~n7666 ) ;
  assign n7668 = ( ~x41 & n7666 ) | ( ~x41 & n7667 ) | ( n7666 & n7667 ) ;
  assign n7669 = ( ~n7661 & n7667 ) | ( ~n7661 & n7668 ) | ( n7667 & n7668 ) ;
  assign n7670 = n910 & n4227 ;
  assign n7671 = x80 & n4231 ;
  assign n7672 = x81 | n7671 ;
  assign n7673 = ( n4233 & n7671 ) | ( n4233 & n7672 ) | ( n7671 & n7672 ) ;
  assign n7674 = x79 & n4470 ;
  assign n7675 = n7673 | n7674 ;
  assign n7676 = ( x44 & n7670 ) | ( x44 & ~n7675 ) | ( n7670 & ~n7675 ) ;
  assign n7677 = ( ~x44 & n7675 ) | ( ~x44 & n7676 ) | ( n7675 & n7676 ) ;
  assign n7678 = ( ~n7670 & n7676 ) | ( ~n7670 & n7677 ) | ( n7676 & n7677 ) ;
  assign n7679 = n461 & n5374 ;
  assign n7680 = x74 & n5378 ;
  assign n7681 = x75 | n7680 ;
  assign n7682 = ( n5380 & n7680 ) | ( n5380 & n7681 ) | ( n7680 & n7681 ) ;
  assign n7683 = x73 & n5638 ;
  assign n7684 = n7682 | n7683 ;
  assign n7685 = ( x50 & n7679 ) | ( x50 & ~n7684 ) | ( n7679 & ~n7684 ) ;
  assign n7686 = ( ~x50 & n7684 ) | ( ~x50 & n7685 ) | ( n7684 & n7685 ) ;
  assign n7687 = ( ~n7679 & n7685 ) | ( ~n7679 & n7686 ) | ( n7685 & n7686 ) ;
  assign n7688 = n346 & n6027 ;
  assign n7689 = x71 & n6031 ;
  assign n7690 = x72 | n7689 ;
  assign n7691 = ( n6033 & n7689 ) | ( n6033 & n7690 ) | ( n7689 & n7690 ) ;
  assign n7692 = x70 & n6303 ;
  assign n7693 = n7691 | n7692 ;
  assign n7694 = ( x53 & n7688 ) | ( x53 & ~n7693 ) | ( n7688 & ~n7693 ) ;
  assign n7695 = ( ~x53 & n7693 ) | ( ~x53 & n7694 ) | ( n7693 & n7694 ) ;
  assign n7696 = ( ~n7688 & n7694 ) | ( ~n7688 & n7695 ) | ( n7694 & n7695 ) ;
  assign n7697 = n230 & n6713 ;
  assign n7698 = x68 & n6717 ;
  assign n7699 = x69 | n7698 ;
  assign n7700 = ( n6719 & n7698 ) | ( n6719 & n7699 ) | ( n7698 & n7699 ) ;
  assign n7701 = x67 & n6980 ;
  assign n7702 = n7700 | n7701 ;
  assign n7703 = ( ~x56 & n7697 ) | ( ~x56 & n7702 ) | ( n7697 & n7702 ) ;
  assign n7704 = ( n7697 & n7702 ) | ( n7697 & ~n7703 ) | ( n7702 & ~n7703 ) ;
  assign n7705 = ( x56 & n7703 ) | ( x56 & ~n7704 ) | ( n7703 & ~n7704 ) ;
  assign n7706 = ( x59 & n7419 ) | ( x59 & n7433 ) | ( n7419 & n7433 ) ;
  assign n7707 = ( x56 & ~x58 ) | ( x56 & n7422 ) | ( ~x58 & n7422 ) ;
  assign n7708 = ( ~n7232 & n7426 ) | ( ~n7232 & n7707 ) | ( n7426 & n7707 ) ;
  assign n7709 = x64 & n7708 ;
  assign n7710 = x65 & n7427 ;
  assign n7711 = x66 | n7710 ;
  assign n7712 = ( n7429 & n7710 ) | ( n7429 & n7711 ) | ( n7710 & n7711 ) ;
  assign n7713 = ( n151 & n152 ) | ( n151 & n7423 ) | ( n152 & n7423 ) ;
  assign n7714 = ( ~n7709 & n7712 ) | ( ~n7709 & n7713 ) | ( n7712 & n7713 ) ;
  assign n7715 = n7709 | n7714 ;
  assign n7716 = n7706 | n7715 ;
  assign n7717 = ( n7706 & n7715 ) | ( n7706 & ~n7716 ) | ( n7715 & ~n7716 ) ;
  assign n7718 = n7716 & ~n7717 ;
  assign n7719 = ( n7445 & n7705 ) | ( n7445 & n7718 ) | ( n7705 & n7718 ) ;
  assign n7720 = ( ~n7445 & n7705 ) | ( ~n7445 & n7718 ) | ( n7705 & n7718 ) ;
  assign n7721 = ( n7445 & ~n7719 ) | ( n7445 & n7720 ) | ( ~n7719 & n7720 ) ;
  assign n7722 = ( n7448 & n7696 ) | ( n7448 & n7721 ) | ( n7696 & n7721 ) ;
  assign n7723 = ( ~n7448 & n7696 ) | ( ~n7448 & n7721 ) | ( n7696 & n7721 ) ;
  assign n7724 = ( n7448 & ~n7722 ) | ( n7448 & n7723 ) | ( ~n7722 & n7723 ) ;
  assign n7725 = ( n7460 & n7687 ) | ( n7460 & n7724 ) | ( n7687 & n7724 ) ;
  assign n7726 = ( ~n7460 & n7687 ) | ( ~n7460 & n7724 ) | ( n7687 & n7724 ) ;
  assign n7727 = ( n7460 & ~n7725 ) | ( n7460 & n7726 ) | ( ~n7725 & n7726 ) ;
  assign n7728 = n637 & n4787 ;
  assign n7729 = x77 & n4791 ;
  assign n7730 = x78 | n7729 ;
  assign n7731 = ( n4793 & n7729 ) | ( n4793 & n7730 ) | ( n7729 & n7730 ) ;
  assign n7732 = x76 & n5030 ;
  assign n7733 = n7731 | n7732 ;
  assign n7734 = ( x47 & n7728 ) | ( x47 & ~n7733 ) | ( n7728 & ~n7733 ) ;
  assign n7735 = ( ~x47 & n7733 ) | ( ~x47 & n7734 ) | ( n7733 & n7734 ) ;
  assign n7736 = ( ~n7728 & n7734 ) | ( ~n7728 & n7735 ) | ( n7734 & n7735 ) ;
  assign n7737 = ( n7472 & n7727 ) | ( n7472 & n7736 ) | ( n7727 & n7736 ) ;
  assign n7738 = ( ~n7472 & n7727 ) | ( ~n7472 & n7736 ) | ( n7727 & n7736 ) ;
  assign n7739 = ( n7472 & ~n7737 ) | ( n7472 & n7738 ) | ( ~n7737 & n7738 ) ;
  assign n7740 = ( n7475 & n7678 ) | ( n7475 & n7739 ) | ( n7678 & n7739 ) ;
  assign n7741 = ( ~n7475 & n7678 ) | ( ~n7475 & n7739 ) | ( n7678 & n7739 ) ;
  assign n7742 = ( n7475 & ~n7740 ) | ( n7475 & n7741 ) | ( ~n7740 & n7741 ) ;
  assign n7743 = ( n7487 & n7669 ) | ( n7487 & n7742 ) | ( n7669 & n7742 ) ;
  assign n7744 = ( ~n7487 & n7669 ) | ( ~n7487 & n7742 ) | ( n7669 & n7742 ) ;
  assign n7745 = ( n7487 & ~n7743 ) | ( n7487 & n7744 ) | ( ~n7743 & n7744 ) ;
  assign n7746 = ( n7490 & n7660 ) | ( n7490 & n7745 ) | ( n7660 & n7745 ) ;
  assign n7747 = ( ~n7490 & n7660 ) | ( ~n7490 & n7745 ) | ( n7660 & n7745 ) ;
  assign n7748 = ( n7490 & ~n7746 ) | ( n7490 & n7747 ) | ( ~n7746 & n7747 ) ;
  assign n7749 = n1701 & n2766 ;
  assign n7750 = x89 & n2770 ;
  assign n7751 = x90 | n7750 ;
  assign n7752 = ( n2772 & n7750 ) | ( n2772 & n7751 ) | ( n7750 & n7751 ) ;
  assign n7753 = x88 & n2943 ;
  assign n7754 = n7752 | n7753 ;
  assign n7755 = ( x35 & n7749 ) | ( x35 & ~n7754 ) | ( n7749 & ~n7754 ) ;
  assign n7756 = ( ~x35 & n7754 ) | ( ~x35 & n7755 ) | ( n7754 & n7755 ) ;
  assign n7757 = ( ~n7749 & n7755 ) | ( ~n7749 & n7756 ) | ( n7755 & n7756 ) ;
  assign n7758 = ( n7502 & n7748 ) | ( n7502 & n7757 ) | ( n7748 & n7757 ) ;
  assign n7759 = ( ~n7502 & n7748 ) | ( ~n7502 & n7757 ) | ( n7748 & n7757 ) ;
  assign n7760 = ( n7502 & ~n7758 ) | ( n7502 & n7759 ) | ( ~n7758 & n7759 ) ;
  assign n7761 = n2057 & n2320 ;
  assign n7762 = x92 & n2324 ;
  assign n7763 = x93 | n7762 ;
  assign n7764 = ( n2326 & n7762 ) | ( n2326 & n7763 ) | ( n7762 & n7763 ) ;
  assign n7765 = x91 & n2497 ;
  assign n7766 = n7764 | n7765 ;
  assign n7767 = ( x32 & n7761 ) | ( x32 & ~n7766 ) | ( n7761 & ~n7766 ) ;
  assign n7768 = ( ~x32 & n7766 ) | ( ~x32 & n7767 ) | ( n7766 & n7767 ) ;
  assign n7769 = ( ~n7761 & n7767 ) | ( ~n7761 & n7768 ) | ( n7767 & n7768 ) ;
  assign n7770 = ( n7514 & n7760 ) | ( n7514 & n7769 ) | ( n7760 & n7769 ) ;
  assign n7771 = ( ~n7514 & n7760 ) | ( ~n7514 & n7769 ) | ( n7760 & n7769 ) ;
  assign n7772 = ( n7514 & ~n7770 ) | ( n7514 & n7771 ) | ( ~n7770 & n7771 ) ;
  assign n7773 = ( n7517 & n7651 ) | ( n7517 & n7772 ) | ( n7651 & n7772 ) ;
  assign n7774 = ( ~n7517 & n7651 ) | ( ~n7517 & n7772 ) | ( n7651 & n7772 ) ;
  assign n7775 = ( n7517 & ~n7773 ) | ( n7517 & n7774 ) | ( ~n7773 & n7774 ) ;
  assign n7776 = n1617 & n2877 ;
  assign n7777 = x98 & n1621 ;
  assign n7778 = x99 | n7777 ;
  assign n7779 = ( n1623 & n7777 ) | ( n1623 & n7778 ) | ( n7777 & n7778 ) ;
  assign n7780 = x97 & n1749 ;
  assign n7781 = n7779 | n7780 ;
  assign n7782 = ( x26 & n7776 ) | ( x26 & ~n7781 ) | ( n7776 & ~n7781 ) ;
  assign n7783 = ( ~x26 & n7781 ) | ( ~x26 & n7782 ) | ( n7781 & n7782 ) ;
  assign n7784 = ( ~n7776 & n7782 ) | ( ~n7776 & n7783 ) | ( n7782 & n7783 ) ;
  assign n7785 = ( n7529 & n7775 ) | ( n7529 & n7784 ) | ( n7775 & n7784 ) ;
  assign n7786 = ( ~n7529 & n7775 ) | ( ~n7529 & n7784 ) | ( n7775 & n7784 ) ;
  assign n7787 = ( n7529 & ~n7785 ) | ( n7529 & n7786 ) | ( ~n7785 & n7786 ) ;
  assign n7788 = n1297 & n3486 ;
  assign n7789 = x101 & n1301 ;
  assign n7790 = x102 | n7789 ;
  assign n7791 = ( n1303 & n7789 ) | ( n1303 & n7790 ) | ( n7789 & n7790 ) ;
  assign n7792 = x100 & n1426 ;
  assign n7793 = n7791 | n7792 ;
  assign n7794 = ( x23 & n7788 ) | ( x23 & ~n7793 ) | ( n7788 & ~n7793 ) ;
  assign n7795 = ( ~x23 & n7793 ) | ( ~x23 & n7794 ) | ( n7793 & n7794 ) ;
  assign n7796 = ( ~n7788 & n7794 ) | ( ~n7788 & n7795 ) | ( n7794 & n7795 ) ;
  assign n7797 = ( n7541 & n7787 ) | ( n7541 & n7796 ) | ( n7787 & n7796 ) ;
  assign n7798 = ( ~n7541 & n7787 ) | ( ~n7541 & n7796 ) | ( n7787 & n7796 ) ;
  assign n7799 = ( n7541 & ~n7797 ) | ( n7541 & n7798 ) | ( ~n7797 & n7798 ) ;
  assign n7800 = n1016 & n3998 ;
  assign n7801 = x104 & n1020 ;
  assign n7802 = x105 | n7801 ;
  assign n7803 = ( n1022 & n7801 ) | ( n1022 & n7802 ) | ( n7801 & n7802 ) ;
  assign n7804 = x103 & n1145 ;
  assign n7805 = n7803 | n7804 ;
  assign n7806 = ( x20 & n7800 ) | ( x20 & ~n7805 ) | ( n7800 & ~n7805 ) ;
  assign n7807 = ( ~x20 & n7805 ) | ( ~x20 & n7806 ) | ( n7805 & n7806 ) ;
  assign n7808 = ( ~n7800 & n7806 ) | ( ~n7800 & n7807 ) | ( n7806 & n7807 ) ;
  assign n7809 = ( n7553 & n7799 ) | ( n7553 & n7808 ) | ( n7799 & n7808 ) ;
  assign n7810 = ( ~n7553 & n7799 ) | ( ~n7553 & n7808 ) | ( n7799 & n7808 ) ;
  assign n7811 = ( n7553 & ~n7809 ) | ( n7553 & n7810 ) | ( ~n7809 & n7810 ) ;
  assign n7812 = ( n7565 & n7642 ) | ( n7565 & n7811 ) | ( n7642 & n7811 ) ;
  assign n7813 = ( ~n7565 & n7642 ) | ( ~n7565 & n7811 ) | ( n7642 & n7811 ) ;
  assign n7814 = ( n7565 & ~n7812 ) | ( n7565 & n7813 ) | ( ~n7812 & n7813 ) ;
  assign n7815 = ( n7568 & n7633 ) | ( n7568 & n7814 ) | ( n7633 & n7814 ) ;
  assign n7816 = ( ~n7568 & n7633 ) | ( ~n7568 & n7814 ) | ( n7633 & n7814 ) ;
  assign n7817 = ( n7568 & ~n7815 ) | ( n7568 & n7816 ) | ( ~n7815 & n7816 ) ;
  assign n7818 = n407 & n5750 ;
  assign n7819 = x113 & n411 ;
  assign n7820 = x114 | n7819 ;
  assign n7821 = ( n413 & n7819 ) | ( n413 & n7820 ) | ( n7819 & n7820 ) ;
  assign n7822 = x112 & n491 ;
  assign n7823 = n7821 | n7822 ;
  assign n7824 = ( x11 & n7818 ) | ( x11 & ~n7823 ) | ( n7818 & ~n7823 ) ;
  assign n7825 = ( ~x11 & n7823 ) | ( ~x11 & n7824 ) | ( n7823 & n7824 ) ;
  assign n7826 = ( ~n7818 & n7824 ) | ( ~n7818 & n7825 ) | ( n7824 & n7825 ) ;
  assign n7827 = ( n7571 & n7817 ) | ( n7571 & n7826 ) | ( n7817 & n7826 ) ;
  assign n7828 = ( ~n7571 & n7817 ) | ( ~n7571 & n7826 ) | ( n7817 & n7826 ) ;
  assign n7829 = ( n7571 & ~n7827 ) | ( n7571 & n7828 ) | ( ~n7827 & n7828 ) ;
  assign n7830 = ( n7574 & n7624 ) | ( n7574 & n7829 ) | ( n7624 & n7829 ) ;
  assign n7831 = ( ~n7574 & n7624 ) | ( ~n7574 & n7829 ) | ( n7624 & n7829 ) ;
  assign n7832 = ( n7574 & ~n7830 ) | ( n7574 & n7831 ) | ( ~n7830 & n7831 ) ;
  assign n7833 = ( n7606 & n7615 ) | ( n7606 & n7832 ) | ( n7615 & n7832 ) ;
  assign n7834 = ( ~n7606 & n7615 ) | ( ~n7606 & n7832 ) | ( n7615 & n7832 ) ;
  assign n7835 = ( n7606 & ~n7833 ) | ( n7606 & n7834 ) | ( ~n7833 & n7834 ) ;
  assign n7836 = ( n7577 & n7592 ) | ( n7577 & n7835 ) | ( n7592 & n7835 ) ;
  assign n7837 = ( n7577 & ~n7592 ) | ( n7577 & n7835 ) | ( ~n7592 & n7835 ) ;
  assign n7838 = ( n7592 & ~n7836 ) | ( n7592 & n7837 ) | ( ~n7836 & n7837 ) ;
  assign n7839 = ( x123 & x124 ) | ( x123 & n7595 ) | ( x124 & n7595 ) ;
  assign n7840 = ( x123 & ~x124 ) | ( x123 & n7595 ) | ( ~x124 & n7595 ) ;
  assign n7841 = ( x124 & ~n7839 ) | ( x124 & n7840 ) | ( ~n7839 & n7840 ) ;
  assign n7842 = n136 & n7841 ;
  assign n7843 = x123 & n138 ;
  assign n7844 = x124 | n7843 ;
  assign n7845 = ( n141 & n7843 ) | ( n141 & n7844 ) | ( n7843 & n7844 ) ;
  assign n7846 = x122 & n154 ;
  assign n7847 = n7845 | n7846 ;
  assign n7848 = ( x2 & n7842 ) | ( x2 & ~n7847 ) | ( n7842 & ~n7847 ) ;
  assign n7849 = ( ~x2 & n7847 ) | ( ~x2 & n7848 ) | ( n7847 & n7848 ) ;
  assign n7850 = ( ~n7842 & n7848 ) | ( ~n7842 & n7849 ) | ( n7848 & n7849 ) ;
  assign n7851 = n186 & n7113 ;
  assign n7852 = x120 & n190 ;
  assign n7853 = x121 | n7852 ;
  assign n7854 = ( n192 & n7852 ) | ( n192 & n7853 ) | ( n7852 & n7853 ) ;
  assign n7855 = x119 & n220 ;
  assign n7856 = n7854 | n7855 ;
  assign n7857 = ( x5 & n7851 ) | ( x5 & ~n7856 ) | ( n7851 & ~n7856 ) ;
  assign n7858 = ( ~x5 & n7856 ) | ( ~x5 & n7857 ) | ( n7856 & n7857 ) ;
  assign n7859 = ( ~n7851 & n7857 ) | ( ~n7851 & n7858 ) | ( n7857 & n7858 ) ;
  assign n7860 = n291 & n6421 ;
  assign n7861 = x117 & n295 ;
  assign n7862 = x118 | n7861 ;
  assign n7863 = ( n297 & n7861 ) | ( n297 & n7862 ) | ( n7861 & n7862 ) ;
  assign n7864 = x116 & n330 ;
  assign n7865 = n7863 | n7864 ;
  assign n7866 = ( x8 & n7860 ) | ( x8 & ~n7865 ) | ( n7860 & ~n7865 ) ;
  assign n7867 = ( ~x8 & n7865 ) | ( ~x8 & n7866 ) | ( n7865 & n7866 ) ;
  assign n7868 = ( ~n7860 & n7866 ) | ( ~n7860 & n7867 ) | ( n7866 & n7867 ) ;
  assign n7869 = n407 & n5765 ;
  assign n7870 = x114 & n411 ;
  assign n7871 = x115 | n7870 ;
  assign n7872 = ( n413 & n7870 ) | ( n413 & n7871 ) | ( n7870 & n7871 ) ;
  assign n7873 = x113 & n491 ;
  assign n7874 = n7872 | n7873 ;
  assign n7875 = ( x11 & n7869 ) | ( x11 & ~n7874 ) | ( n7869 & ~n7874 ) ;
  assign n7876 = ( ~x11 & n7874 ) | ( ~x11 & n7875 ) | ( n7874 & n7875 ) ;
  assign n7877 = ( ~n7869 & n7875 ) | ( ~n7869 & n7876 ) | ( n7875 & n7876 ) ;
  assign n7878 = n583 & n5145 ;
  assign n7879 = x111 & n587 ;
  assign n7880 = x112 | n7879 ;
  assign n7881 = ( n589 & n7879 ) | ( n589 & n7880 ) | ( n7879 & n7880 ) ;
  assign n7882 = x110 & n676 ;
  assign n7883 = n7881 | n7882 ;
  assign n7884 = ( x14 & n7878 ) | ( x14 & ~n7883 ) | ( n7878 & ~n7883 ) ;
  assign n7885 = ( ~x14 & n7883 ) | ( ~x14 & n7884 ) | ( n7883 & n7884 ) ;
  assign n7886 = ( ~n7878 & n7884 ) | ( ~n7878 & n7885 ) | ( n7884 & n7885 ) ;
  assign n7887 = n810 & n4734 ;
  assign n7888 = x108 & n814 ;
  assign n7889 = x109 | n7888 ;
  assign n7890 = ( n816 & n7888 ) | ( n816 & n7889 ) | ( n7888 & n7889 ) ;
  assign n7891 = x107 & n885 ;
  assign n7892 = n7890 | n7891 ;
  assign n7893 = ( x17 & n7887 ) | ( x17 & ~n7892 ) | ( n7887 & ~n7892 ) ;
  assign n7894 = ( ~x17 & n7892 ) | ( ~x17 & n7893 ) | ( n7892 & n7893 ) ;
  assign n7895 = ( ~n7887 & n7893 ) | ( ~n7887 & n7894 ) | ( n7893 & n7894 ) ;
  assign n7896 = n1617 & n3162 ;
  assign n7897 = x99 & n1621 ;
  assign n7898 = x100 | n7897 ;
  assign n7899 = ( n1623 & n7897 ) | ( n1623 & n7898 ) | ( n7897 & n7898 ) ;
  assign n7900 = x98 & n1749 ;
  assign n7901 = n7899 | n7900 ;
  assign n7902 = ( x26 & n7896 ) | ( x26 & ~n7901 ) | ( n7896 & ~n7901 ) ;
  assign n7903 = ( ~x26 & n7901 ) | ( ~x26 & n7902 ) | ( n7901 & n7902 ) ;
  assign n7904 = ( ~n7896 & n7902 ) | ( ~n7896 & n7903 ) | ( n7902 & n7903 ) ;
  assign n7905 = n1262 & n3715 ;
  assign n7906 = x84 & n3719 ;
  assign n7907 = x85 | n7906 ;
  assign n7908 = ( n3721 & n7906 ) | ( n3721 & n7907 ) | ( n7906 & n7907 ) ;
  assign n7909 = x83 & n3922 ;
  assign n7910 = n7908 | n7909 ;
  assign n7911 = ( x41 & n7905 ) | ( x41 & ~n7910 ) | ( n7905 & ~n7910 ) ;
  assign n7912 = ( ~x41 & n7910 ) | ( ~x41 & n7911 ) | ( n7910 & n7911 ) ;
  assign n7913 = ( ~n7905 & n7911 ) | ( ~n7905 & n7912 ) | ( n7911 & n7912 ) ;
  assign n7914 = n990 & n4227 ;
  assign n7915 = x81 & n4231 ;
  assign n7916 = x82 | n7915 ;
  assign n7917 = ( n4233 & n7915 ) | ( n4233 & n7916 ) | ( n7915 & n7916 ) ;
  assign n7918 = x80 & n4470 ;
  assign n7919 = n7917 | n7918 ;
  assign n7920 = ( x44 & n7914 ) | ( x44 & ~n7919 ) | ( n7914 & ~n7919 ) ;
  assign n7921 = ( ~x44 & n7919 ) | ( ~x44 & n7920 ) | ( n7919 & n7920 ) ;
  assign n7922 = ( ~n7914 & n7920 ) | ( ~n7914 & n7921 ) | ( n7920 & n7921 ) ;
  assign n7923 = n701 & n4787 ;
  assign n7924 = x78 & n4791 ;
  assign n7925 = x79 | n7924 ;
  assign n7926 = ( n4793 & n7924 ) | ( n4793 & n7925 ) | ( n7924 & n7925 ) ;
  assign n7927 = x77 & n5030 ;
  assign n7928 = n7926 | n7927 ;
  assign n7929 = ( x47 & n7923 ) | ( x47 & ~n7928 ) | ( n7923 & ~n7928 ) ;
  assign n7930 = ( ~x47 & n7928 ) | ( ~x47 & n7929 ) | ( n7928 & n7929 ) ;
  assign n7931 = ( ~n7923 & n7929 ) | ( ~n7923 & n7930 ) | ( n7929 & n7930 ) ;
  assign n7932 = n554 & n5374 ;
  assign n7933 = x75 & n5378 ;
  assign n7934 = x76 | n7933 ;
  assign n7935 = ( n5380 & n7933 ) | ( n5380 & n7934 ) | ( n7933 & n7934 ) ;
  assign n7936 = x74 & n5638 ;
  assign n7937 = n7935 | n7936 ;
  assign n7938 = ( x50 & n7932 ) | ( x50 & ~n7937 ) | ( n7932 & ~n7937 ) ;
  assign n7939 = ( ~x50 & n7937 ) | ( ~x50 & n7938 ) | ( n7937 & n7938 ) ;
  assign n7940 = ( ~n7932 & n7938 ) | ( ~n7932 & n7939 ) | ( n7938 & n7939 ) ;
  assign n7941 = n390 & n6027 ;
  assign n7942 = x72 & n6031 ;
  assign n7943 = x73 | n7942 ;
  assign n7944 = ( n6033 & n7942 ) | ( n6033 & n7943 ) | ( n7942 & n7943 ) ;
  assign n7945 = x71 & n6303 ;
  assign n7946 = n7944 | n7945 ;
  assign n7947 = ( x53 & n7941 ) | ( x53 & ~n7946 ) | ( n7941 & ~n7946 ) ;
  assign n7948 = ( ~x53 & n7946 ) | ( ~x53 & n7947 ) | ( n7946 & n7947 ) ;
  assign n7949 = ( ~n7941 & n7947 ) | ( ~n7941 & n7948 ) | ( n7947 & n7948 ) ;
  assign n7950 = x66 & n7427 ;
  assign n7951 = x67 | n7950 ;
  assign n7952 = ( n7429 & n7950 ) | ( n7429 & n7951 ) | ( n7950 & n7951 ) ;
  assign n7953 = x65 & n7708 ;
  assign n7954 = n7952 | n7953 ;
  assign n7955 = n164 & n7423 ;
  assign n7956 = ( x59 & n7954 ) | ( x59 & ~n7955 ) | ( n7954 & ~n7955 ) ;
  assign n7957 = ( ~x59 & n7955 ) | ( ~x59 & n7956 ) | ( n7955 & n7956 ) ;
  assign n7958 = ( ~n7954 & n7956 ) | ( ~n7954 & n7957 ) | ( n7956 & n7957 ) ;
  assign n7959 = x59 & x60 ;
  assign n7960 = x59 | x60 ;
  assign n7961 = ~n7959 & n7960 ;
  assign n7962 = x64 & n7961 ;
  assign n7963 = x59 & ~n7716 ;
  assign n7964 = ( n7958 & n7962 ) | ( n7958 & n7963 ) | ( n7962 & n7963 ) ;
  assign n7965 = ( ~n7958 & n7962 ) | ( ~n7958 & n7963 ) | ( n7962 & n7963 ) ;
  assign n7966 = ( n7958 & ~n7964 ) | ( n7958 & n7965 ) | ( ~n7964 & n7965 ) ;
  assign n7967 = n245 & n6713 ;
  assign n7968 = x69 & n6717 ;
  assign n7969 = x70 | n7968 ;
  assign n7970 = ( n6719 & n7968 ) | ( n6719 & n7969 ) | ( n7968 & n7969 ) ;
  assign n7971 = x68 & n6980 ;
  assign n7972 = n7970 | n7971 ;
  assign n7973 = ( x56 & n7967 ) | ( x56 & ~n7972 ) | ( n7967 & ~n7972 ) ;
  assign n7974 = ( ~x56 & n7972 ) | ( ~x56 & n7973 ) | ( n7972 & n7973 ) ;
  assign n7975 = ( ~n7967 & n7973 ) | ( ~n7967 & n7974 ) | ( n7973 & n7974 ) ;
  assign n7976 = ( n7719 & n7966 ) | ( n7719 & n7975 ) | ( n7966 & n7975 ) ;
  assign n7977 = ( ~n7719 & n7966 ) | ( ~n7719 & n7975 ) | ( n7966 & n7975 ) ;
  assign n7978 = ( n7719 & ~n7976 ) | ( n7719 & n7977 ) | ( ~n7976 & n7977 ) ;
  assign n7979 = ( n7722 & n7949 ) | ( n7722 & n7978 ) | ( n7949 & n7978 ) ;
  assign n7980 = ( ~n7722 & n7949 ) | ( ~n7722 & n7978 ) | ( n7949 & n7978 ) ;
  assign n7981 = ( n7722 & ~n7979 ) | ( n7722 & n7980 ) | ( ~n7979 & n7980 ) ;
  assign n7982 = ( n7725 & n7940 ) | ( n7725 & n7981 ) | ( n7940 & n7981 ) ;
  assign n7983 = ( ~n7725 & n7940 ) | ( ~n7725 & n7981 ) | ( n7940 & n7981 ) ;
  assign n7984 = ( n7725 & ~n7982 ) | ( n7725 & n7983 ) | ( ~n7982 & n7983 ) ;
  assign n7985 = ( n7737 & n7931 ) | ( n7737 & n7984 ) | ( n7931 & n7984 ) ;
  assign n7986 = ( ~n7737 & n7931 ) | ( ~n7737 & n7984 ) | ( n7931 & n7984 ) ;
  assign n7987 = ( n7737 & ~n7985 ) | ( n7737 & n7986 ) | ( ~n7985 & n7986 ) ;
  assign n7988 = ( n7740 & n7922 ) | ( n7740 & n7987 ) | ( n7922 & n7987 ) ;
  assign n7989 = ( ~n7740 & n7922 ) | ( ~n7740 & n7987 ) | ( n7922 & n7987 ) ;
  assign n7990 = ( n7740 & ~n7988 ) | ( n7740 & n7989 ) | ( ~n7988 & n7989 ) ;
  assign n7991 = ( n7743 & n7913 ) | ( n7743 & n7990 ) | ( n7913 & n7990 ) ;
  assign n7992 = ( ~n7743 & n7913 ) | ( ~n7743 & n7990 ) | ( n7913 & n7990 ) ;
  assign n7993 = ( n7743 & ~n7991 ) | ( n7743 & n7992 ) | ( ~n7991 & n7992 ) ;
  assign n7994 = n1481 & n3224 ;
  assign n7995 = x87 & n3228 ;
  assign n7996 = x88 | n7995 ;
  assign n7997 = ( n3230 & n7995 ) | ( n3230 & n7996 ) | ( n7995 & n7996 ) ;
  assign n7998 = x86 & n3413 ;
  assign n7999 = n7997 | n7998 ;
  assign n8000 = ( x38 & n7994 ) | ( x38 & ~n7999 ) | ( n7994 & ~n7999 ) ;
  assign n8001 = ( ~x38 & n7999 ) | ( ~x38 & n8000 ) | ( n7999 & n8000 ) ;
  assign n8002 = ( ~n7994 & n8000 ) | ( ~n7994 & n8001 ) | ( n8000 & n8001 ) ;
  assign n8003 = ( n7746 & n7993 ) | ( n7746 & n8002 ) | ( n7993 & n8002 ) ;
  assign n8004 = ( ~n7746 & n7993 ) | ( ~n7746 & n8002 ) | ( n7993 & n8002 ) ;
  assign n8005 = ( n7746 & ~n8003 ) | ( n7746 & n8004 ) | ( ~n8003 & n8004 ) ;
  assign n8006 = n1914 & n2766 ;
  assign n8007 = x90 & n2770 ;
  assign n8008 = x91 | n8007 ;
  assign n8009 = ( n2772 & n8007 ) | ( n2772 & n8008 ) | ( n8007 & n8008 ) ;
  assign n8010 = x89 & n2943 ;
  assign n8011 = n8009 | n8010 ;
  assign n8012 = ( x35 & n8006 ) | ( x35 & ~n8011 ) | ( n8006 & ~n8011 ) ;
  assign n8013 = ( ~x35 & n8011 ) | ( ~x35 & n8012 ) | ( n8011 & n8012 ) ;
  assign n8014 = ( ~n8006 & n8012 ) | ( ~n8006 & n8013 ) | ( n8012 & n8013 ) ;
  assign n8015 = ( n7758 & n8005 ) | ( n7758 & n8014 ) | ( n8005 & n8014 ) ;
  assign n8016 = ( ~n7758 & n8005 ) | ( ~n7758 & n8014 ) | ( n8005 & n8014 ) ;
  assign n8017 = ( n7758 & ~n8015 ) | ( n7758 & n8016 ) | ( ~n8015 & n8016 ) ;
  assign n8018 = n2294 & n2320 ;
  assign n8019 = x93 & n2324 ;
  assign n8020 = x94 | n8019 ;
  assign n8021 = ( n2326 & n8019 ) | ( n2326 & n8020 ) | ( n8019 & n8020 ) ;
  assign n8022 = x92 & n2497 ;
  assign n8023 = n8021 | n8022 ;
  assign n8024 = ( x32 & n8018 ) | ( x32 & ~n8023 ) | ( n8018 & ~n8023 ) ;
  assign n8025 = ( ~x32 & n8023 ) | ( ~x32 & n8024 ) | ( n8023 & n8024 ) ;
  assign n8026 = ( ~n8018 & n8024 ) | ( ~n8018 & n8025 ) | ( n8024 & n8025 ) ;
  assign n8027 = ( n7770 & n8017 ) | ( n7770 & n8026 ) | ( n8017 & n8026 ) ;
  assign n8028 = ( ~n7770 & n8017 ) | ( ~n7770 & n8026 ) | ( n8017 & n8026 ) ;
  assign n8029 = ( n7770 & ~n8027 ) | ( n7770 & n8028 ) | ( ~n8027 & n8028 ) ;
  assign n8030 = n1949 & n2585 ;
  assign n8031 = x96 & n1953 ;
  assign n8032 = x97 | n8031 ;
  assign n8033 = ( n1955 & n8031 ) | ( n1955 & n8032 ) | ( n8031 & n8032 ) ;
  assign n8034 = x95 & n2114 ;
  assign n8035 = n8033 | n8034 ;
  assign n8036 = ( x29 & n8030 ) | ( x29 & ~n8035 ) | ( n8030 & ~n8035 ) ;
  assign n8037 = ( ~x29 & n8035 ) | ( ~x29 & n8036 ) | ( n8035 & n8036 ) ;
  assign n8038 = ( ~n8030 & n8036 ) | ( ~n8030 & n8037 ) | ( n8036 & n8037 ) ;
  assign n8039 = ( n7773 & n8029 ) | ( n7773 & n8038 ) | ( n8029 & n8038 ) ;
  assign n8040 = ( ~n7773 & n8029 ) | ( ~n7773 & n8038 ) | ( n8029 & n8038 ) ;
  assign n8041 = ( n7773 & ~n8039 ) | ( n7773 & n8040 ) | ( ~n8039 & n8040 ) ;
  assign n8042 = ( n7785 & n7904 ) | ( n7785 & n8041 ) | ( n7904 & n8041 ) ;
  assign n8043 = ( ~n7785 & n7904 ) | ( ~n7785 & n8041 ) | ( n7904 & n8041 ) ;
  assign n8044 = ( n7785 & ~n8042 ) | ( n7785 & n8043 ) | ( ~n8042 & n8043 ) ;
  assign n8045 = n1297 & n3650 ;
  assign n8046 = x102 & n1301 ;
  assign n8047 = x103 | n8046 ;
  assign n8048 = ( n1303 & n8046 ) | ( n1303 & n8047 ) | ( n8046 & n8047 ) ;
  assign n8049 = x101 & n1426 ;
  assign n8050 = n8048 | n8049 ;
  assign n8051 = ( x23 & n8045 ) | ( x23 & ~n8050 ) | ( n8045 & ~n8050 ) ;
  assign n8052 = ( ~x23 & n8050 ) | ( ~x23 & n8051 ) | ( n8050 & n8051 ) ;
  assign n8053 = ( ~n8045 & n8051 ) | ( ~n8045 & n8052 ) | ( n8051 & n8052 ) ;
  assign n8054 = ( n7797 & n8044 ) | ( n7797 & n8053 ) | ( n8044 & n8053 ) ;
  assign n8055 = ( ~n7797 & n8044 ) | ( ~n7797 & n8053 ) | ( n8044 & n8053 ) ;
  assign n8056 = ( n7797 & ~n8054 ) | ( n7797 & n8055 ) | ( ~n8054 & n8055 ) ;
  assign n8057 = n1016 & n4013 ;
  assign n8058 = x105 & n1020 ;
  assign n8059 = x106 | n8058 ;
  assign n8060 = ( n1022 & n8058 ) | ( n1022 & n8059 ) | ( n8058 & n8059 ) ;
  assign n8061 = x104 & n1145 ;
  assign n8062 = n8060 | n8061 ;
  assign n8063 = ( x20 & n8057 ) | ( x20 & ~n8062 ) | ( n8057 & ~n8062 ) ;
  assign n8064 = ( ~x20 & n8062 ) | ( ~x20 & n8063 ) | ( n8062 & n8063 ) ;
  assign n8065 = ( ~n8057 & n8063 ) | ( ~n8057 & n8064 ) | ( n8063 & n8064 ) ;
  assign n8066 = ( n7809 & n8056 ) | ( n7809 & n8065 ) | ( n8056 & n8065 ) ;
  assign n8067 = ( ~n7809 & n8056 ) | ( ~n7809 & n8065 ) | ( n8056 & n8065 ) ;
  assign n8068 = ( n7809 & ~n8066 ) | ( n7809 & n8067 ) | ( ~n8066 & n8067 ) ;
  assign n8069 = ( n7812 & n7895 ) | ( n7812 & n8068 ) | ( n7895 & n8068 ) ;
  assign n8070 = ( ~n7812 & n7895 ) | ( ~n7812 & n8068 ) | ( n7895 & n8068 ) ;
  assign n8071 = ( n7812 & ~n8069 ) | ( n7812 & n8070 ) | ( ~n8069 & n8070 ) ;
  assign n8072 = ( n7815 & n7886 ) | ( n7815 & n8071 ) | ( n7886 & n8071 ) ;
  assign n8073 = ( ~n7815 & n7886 ) | ( ~n7815 & n8071 ) | ( n7886 & n8071 ) ;
  assign n8074 = ( n7815 & ~n8072 ) | ( n7815 & n8073 ) | ( ~n8072 & n8073 ) ;
  assign n8075 = ( n7827 & n7877 ) | ( n7827 & n8074 ) | ( n7877 & n8074 ) ;
  assign n8076 = ( ~n7827 & n7877 ) | ( ~n7827 & n8074 ) | ( n7877 & n8074 ) ;
  assign n8077 = ( n7827 & ~n8075 ) | ( n7827 & n8076 ) | ( ~n8075 & n8076 ) ;
  assign n8078 = ( n7830 & n7868 ) | ( n7830 & n8077 ) | ( n7868 & n8077 ) ;
  assign n8079 = ( ~n7830 & n7868 ) | ( ~n7830 & n8077 ) | ( n7868 & n8077 ) ;
  assign n8080 = ( n7830 & ~n8078 ) | ( n7830 & n8079 ) | ( ~n8078 & n8079 ) ;
  assign n8081 = ( n7850 & n7859 ) | ( n7850 & n8080 ) | ( n7859 & n8080 ) ;
  assign n8082 = ( ~n7850 & n7859 ) | ( ~n7850 & n8080 ) | ( n7859 & n8080 ) ;
  assign n8083 = ( n7850 & ~n8081 ) | ( n7850 & n8082 ) | ( ~n8081 & n8082 ) ;
  assign n8084 = ( n7833 & n7836 ) | ( n7833 & n8083 ) | ( n7836 & n8083 ) ;
  assign n8085 = ( n7833 & ~n7836 ) | ( n7833 & n8083 ) | ( ~n7836 & n8083 ) ;
  assign n8086 = ( n7836 & ~n8084 ) | ( n7836 & n8085 ) | ( ~n8084 & n8085 ) ;
  assign n8087 = n407 & n5977 ;
  assign n8088 = x115 & n411 ;
  assign n8089 = x116 | n8088 ;
  assign n8090 = ( n413 & n8088 ) | ( n413 & n8089 ) | ( n8088 & n8089 ) ;
  assign n8091 = x114 & n491 ;
  assign n8092 = n8090 | n8091 ;
  assign n8093 = ( x11 & n8087 ) | ( x11 & ~n8092 ) | ( n8087 & ~n8092 ) ;
  assign n8094 = ( ~x11 & n8092 ) | ( ~x11 & n8093 ) | ( n8092 & n8093 ) ;
  assign n8095 = ( ~n8087 & n8093 ) | ( ~n8087 & n8094 ) | ( n8093 & n8094 ) ;
  assign n8096 = n583 & n5542 ;
  assign n8097 = x112 & n587 ;
  assign n8098 = x113 | n8097 ;
  assign n8099 = ( n589 & n8097 ) | ( n589 & n8098 ) | ( n8097 & n8098 ) ;
  assign n8100 = x111 & n676 ;
  assign n8101 = n8099 | n8100 ;
  assign n8102 = ( x14 & n8096 ) | ( x14 & ~n8101 ) | ( n8096 & ~n8101 ) ;
  assign n8103 = ( ~x14 & n8101 ) | ( ~x14 & n8102 ) | ( n8101 & n8102 ) ;
  assign n8104 = ( ~n8096 & n8102 ) | ( ~n8096 & n8103 ) | ( n8102 & n8103 ) ;
  assign n8105 = n810 & n4934 ;
  assign n8106 = x109 & n814 ;
  assign n8107 = x110 | n8106 ;
  assign n8108 = ( n816 & n8106 ) | ( n816 & n8107 ) | ( n8106 & n8107 ) ;
  assign n8109 = x108 & n885 ;
  assign n8110 = n8108 | n8109 ;
  assign n8111 = ( x17 & n8105 ) | ( x17 & ~n8110 ) | ( n8105 & ~n8110 ) ;
  assign n8112 = ( ~x17 & n8110 ) | ( ~x17 & n8111 ) | ( n8110 & n8111 ) ;
  assign n8113 = ( ~n8105 & n8111 ) | ( ~n8105 & n8112 ) | ( n8111 & n8112 ) ;
  assign n8114 = n1949 & n2725 ;
  assign n8115 = x97 & n1953 ;
  assign n8116 = x98 | n8115 ;
  assign n8117 = ( n1955 & n8115 ) | ( n1955 & n8116 ) | ( n8115 & n8116 ) ;
  assign n8118 = x96 & n2114 ;
  assign n8119 = n8117 | n8118 ;
  assign n8120 = ( x29 & n8114 ) | ( x29 & ~n8119 ) | ( n8114 & ~n8119 ) ;
  assign n8121 = ( ~x29 & n8119 ) | ( ~x29 & n8120 ) | ( n8119 & n8120 ) ;
  assign n8122 = ( ~n8114 & n8120 ) | ( ~n8114 & n8121 ) | ( n8120 & n8121 ) ;
  assign n8123 = n1366 & n3715 ;
  assign n8124 = x85 & n3719 ;
  assign n8125 = x86 | n8124 ;
  assign n8126 = ( n3721 & n8124 ) | ( n3721 & n8125 ) | ( n8124 & n8125 ) ;
  assign n8127 = x84 & n3922 ;
  assign n8128 = n8126 | n8127 ;
  assign n8129 = ( x41 & n8123 ) | ( x41 & ~n8128 ) | ( n8123 & ~n8128 ) ;
  assign n8130 = ( ~x41 & n8128 ) | ( ~x41 & n8129 ) | ( n8128 & n8129 ) ;
  assign n8131 = ( ~n8123 & n8129 ) | ( ~n8123 & n8130 ) | ( n8129 & n8130 ) ;
  assign n8132 = n769 & n4787 ;
  assign n8133 = x79 & n4791 ;
  assign n8134 = x80 | n8133 ;
  assign n8135 = ( n4793 & n8133 ) | ( n4793 & n8134 ) | ( n8133 & n8134 ) ;
  assign n8136 = x78 & n5030 ;
  assign n8137 = n8135 | n8136 ;
  assign n8138 = ( x47 & n8132 ) | ( x47 & ~n8137 ) | ( n8132 & ~n8137 ) ;
  assign n8139 = ( ~x47 & n8137 ) | ( ~x47 & n8138 ) | ( n8137 & n8138 ) ;
  assign n8140 = ( ~n8132 & n8138 ) | ( ~n8132 & n8139 ) | ( n8138 & n8139 ) ;
  assign n8141 = n277 & n6713 ;
  assign n8142 = x70 & n6717 ;
  assign n8143 = x71 | n8142 ;
  assign n8144 = ( n6719 & n8142 ) | ( n6719 & n8143 ) | ( n8142 & n8143 ) ;
  assign n8145 = x69 & n6980 ;
  assign n8146 = n8144 | n8145 ;
  assign n8147 = ( x56 & n8141 ) | ( x56 & ~n8146 ) | ( n8141 & ~n8146 ) ;
  assign n8148 = ( ~x56 & n8146 ) | ( ~x56 & n8147 ) | ( n8146 & n8147 ) ;
  assign n8149 = ( ~n8141 & n8147 ) | ( ~n8141 & n8148 ) | ( n8147 & n8148 ) ;
  assign n8150 = x62 & n7962 ;
  assign n8151 = x61 | x62 ;
  assign n8152 = ( x61 & x62 ) | ( x61 & ~n8151 ) | ( x62 & ~n8151 ) ;
  assign n8153 = n8151 & ~n8152 ;
  assign n8154 = n7961 & n8153 ;
  assign n8155 = n133 & n8154 ;
  assign n8156 = ~x59 & x61 ;
  assign n8157 = x60 & x61 ;
  assign n8158 = ( n7959 & n8156 ) | ( n7959 & ~n8157 ) | ( n8156 & ~n8157 ) ;
  assign n8159 = x64 & n8158 ;
  assign n8160 = ( n7961 & ~n8151 ) | ( n7961 & n8152 ) | ( ~n8151 & n8152 ) ;
  assign n8161 = x65 | n8159 ;
  assign n8162 = ( n8159 & n8160 ) | ( n8159 & n8161 ) | ( n8160 & n8161 ) ;
  assign n8163 = ( n8150 & n8155 ) | ( n8150 & n8162 ) | ( n8155 & n8162 ) ;
  assign n8164 = n8155 | n8162 ;
  assign n8165 = ~n8150 & n8164 ;
  assign n8166 = ( n8150 & ~n8163 ) | ( n8150 & n8165 ) | ( ~n8163 & n8165 ) ;
  assign n8167 = x67 & n7427 ;
  assign n8168 = x68 | n8167 ;
  assign n8169 = ( n7429 & n8167 ) | ( n7429 & n8168 ) | ( n8167 & n8168 ) ;
  assign n8170 = x66 & n7708 ;
  assign n8171 = n8169 | n8170 ;
  assign n8172 = n201 & n7423 ;
  assign n8173 = ( x59 & n8171 ) | ( x59 & ~n8172 ) | ( n8171 & ~n8172 ) ;
  assign n8174 = ( ~x59 & n8172 ) | ( ~x59 & n8173 ) | ( n8172 & n8173 ) ;
  assign n8175 = ( ~n8171 & n8173 ) | ( ~n8171 & n8174 ) | ( n8173 & n8174 ) ;
  assign n8176 = ( n7964 & n8166 ) | ( n7964 & n8175 ) | ( n8166 & n8175 ) ;
  assign n8177 = ( ~n7964 & n8166 ) | ( ~n7964 & n8175 ) | ( n8166 & n8175 ) ;
  assign n8178 = ( n7964 & ~n8176 ) | ( n7964 & n8177 ) | ( ~n8176 & n8177 ) ;
  assign n8179 = ( n7976 & n8149 ) | ( n7976 & n8178 ) | ( n8149 & n8178 ) ;
  assign n8180 = ( ~n7976 & n8149 ) | ( ~n7976 & n8178 ) | ( n8149 & n8178 ) ;
  assign n8181 = ( n7976 & ~n8179 ) | ( n7976 & n8180 ) | ( ~n8179 & n8180 ) ;
  assign n8182 = n446 & n6027 ;
  assign n8183 = x73 & n6031 ;
  assign n8184 = x74 | n8183 ;
  assign n8185 = ( n6033 & n8183 ) | ( n6033 & n8184 ) | ( n8183 & n8184 ) ;
  assign n8186 = x72 & n6303 ;
  assign n8187 = n8185 | n8186 ;
  assign n8188 = ( x53 & n8182 ) | ( x53 & ~n8187 ) | ( n8182 & ~n8187 ) ;
  assign n8189 = ( ~x53 & n8187 ) | ( ~x53 & n8188 ) | ( n8187 & n8188 ) ;
  assign n8190 = ( ~n8182 & n8188 ) | ( ~n8182 & n8189 ) | ( n8188 & n8189 ) ;
  assign n8191 = ( n7979 & n8181 ) | ( n7979 & n8190 ) | ( n8181 & n8190 ) ;
  assign n8192 = ( ~n7979 & n8181 ) | ( ~n7979 & n8190 ) | ( n8181 & n8190 ) ;
  assign n8193 = ( n7979 & ~n8191 ) | ( n7979 & n8192 ) | ( ~n8191 & n8192 ) ;
  assign n8194 = n569 & n5374 ;
  assign n8195 = x76 & n5378 ;
  assign n8196 = x77 | n8195 ;
  assign n8197 = ( n5380 & n8195 ) | ( n5380 & n8196 ) | ( n8195 & n8196 ) ;
  assign n8198 = x75 & n5638 ;
  assign n8199 = n8197 | n8198 ;
  assign n8200 = ( x50 & n8194 ) | ( x50 & ~n8199 ) | ( n8194 & ~n8199 ) ;
  assign n8201 = ( ~x50 & n8199 ) | ( ~x50 & n8200 ) | ( n8199 & n8200 ) ;
  assign n8202 = ( ~n8194 & n8200 ) | ( ~n8194 & n8201 ) | ( n8200 & n8201 ) ;
  assign n8203 = ( n7982 & n8193 ) | ( n7982 & n8202 ) | ( n8193 & n8202 ) ;
  assign n8204 = ( ~n7982 & n8193 ) | ( ~n7982 & n8202 ) | ( n8193 & n8202 ) ;
  assign n8205 = ( n7982 & ~n8203 ) | ( n7982 & n8204 ) | ( ~n8203 & n8204 ) ;
  assign n8206 = ( n7985 & n8140 ) | ( n7985 & n8205 ) | ( n8140 & n8205 ) ;
  assign n8207 = ( ~n7985 & n8140 ) | ( ~n7985 & n8205 ) | ( n8140 & n8205 ) ;
  assign n8208 = ( n7985 & ~n8206 ) | ( n7985 & n8207 ) | ( ~n8206 & n8207 ) ;
  assign n8209 = n1082 & n4227 ;
  assign n8210 = x82 & n4231 ;
  assign n8211 = x83 | n8210 ;
  assign n8212 = ( n4233 & n8210 ) | ( n4233 & n8211 ) | ( n8210 & n8211 ) ;
  assign n8213 = x81 & n4470 ;
  assign n8214 = n8212 | n8213 ;
  assign n8215 = ( x44 & n8209 ) | ( x44 & ~n8214 ) | ( n8209 & ~n8214 ) ;
  assign n8216 = ( ~x44 & n8214 ) | ( ~x44 & n8215 ) | ( n8214 & n8215 ) ;
  assign n8217 = ( ~n8209 & n8215 ) | ( ~n8209 & n8216 ) | ( n8215 & n8216 ) ;
  assign n8218 = ( n7988 & n8208 ) | ( n7988 & n8217 ) | ( n8208 & n8217 ) ;
  assign n8219 = ( ~n7988 & n8208 ) | ( ~n7988 & n8217 ) | ( n8208 & n8217 ) ;
  assign n8220 = ( n7988 & ~n8218 ) | ( n7988 & n8219 ) | ( ~n8218 & n8219 ) ;
  assign n8221 = ( n7991 & n8131 ) | ( n7991 & n8220 ) | ( n8131 & n8220 ) ;
  assign n8222 = ( ~n7991 & n8131 ) | ( ~n7991 & n8220 ) | ( n8131 & n8220 ) ;
  assign n8223 = ( n7991 & ~n8221 ) | ( n7991 & n8222 ) | ( ~n8221 & n8222 ) ;
  assign n8224 = n1585 & n3224 ;
  assign n8225 = x88 & n3228 ;
  assign n8226 = x89 | n8225 ;
  assign n8227 = ( n3230 & n8225 ) | ( n3230 & n8226 ) | ( n8225 & n8226 ) ;
  assign n8228 = x87 & n3413 ;
  assign n8229 = n8227 | n8228 ;
  assign n8230 = ( x38 & n8224 ) | ( x38 & ~n8229 ) | ( n8224 & ~n8229 ) ;
  assign n8231 = ( ~x38 & n8229 ) | ( ~x38 & n8230 ) | ( n8229 & n8230 ) ;
  assign n8232 = ( ~n8224 & n8230 ) | ( ~n8224 & n8231 ) | ( n8230 & n8231 ) ;
  assign n8233 = ( n8003 & n8223 ) | ( n8003 & n8232 ) | ( n8223 & n8232 ) ;
  assign n8234 = ( ~n8003 & n8223 ) | ( ~n8003 & n8232 ) | ( n8223 & n8232 ) ;
  assign n8235 = ( n8003 & ~n8233 ) | ( n8003 & n8234 ) | ( ~n8233 & n8234 ) ;
  assign n8236 = n2042 & n2766 ;
  assign n8237 = x91 & n2770 ;
  assign n8238 = x92 | n8237 ;
  assign n8239 = ( n2772 & n8237 ) | ( n2772 & n8238 ) | ( n8237 & n8238 ) ;
  assign n8240 = x90 & n2943 ;
  assign n8241 = n8239 | n8240 ;
  assign n8242 = ( x35 & n8236 ) | ( x35 & ~n8241 ) | ( n8236 & ~n8241 ) ;
  assign n8243 = ( ~x35 & n8241 ) | ( ~x35 & n8242 ) | ( n8241 & n8242 ) ;
  assign n8244 = ( ~n8236 & n8242 ) | ( ~n8236 & n8243 ) | ( n8242 & n8243 ) ;
  assign n8245 = ( n8015 & n8235 ) | ( n8015 & n8244 ) | ( n8235 & n8244 ) ;
  assign n8246 = ( ~n8015 & n8235 ) | ( ~n8015 & n8244 ) | ( n8235 & n8244 ) ;
  assign n8247 = ( n8015 & ~n8245 ) | ( n8015 & n8246 ) | ( ~n8245 & n8246 ) ;
  assign n8248 = n2320 & n2434 ;
  assign n8249 = x94 & n2324 ;
  assign n8250 = x95 | n8249 ;
  assign n8251 = ( n2326 & n8249 ) | ( n2326 & n8250 ) | ( n8249 & n8250 ) ;
  assign n8252 = x93 & n2497 ;
  assign n8253 = n8251 | n8252 ;
  assign n8254 = ( x32 & n8248 ) | ( x32 & ~n8253 ) | ( n8248 & ~n8253 ) ;
  assign n8255 = ( ~x32 & n8253 ) | ( ~x32 & n8254 ) | ( n8253 & n8254 ) ;
  assign n8256 = ( ~n8248 & n8254 ) | ( ~n8248 & n8255 ) | ( n8254 & n8255 ) ;
  assign n8257 = ( n8027 & n8247 ) | ( n8027 & n8256 ) | ( n8247 & n8256 ) ;
  assign n8258 = ( ~n8027 & n8247 ) | ( ~n8027 & n8256 ) | ( n8247 & n8256 ) ;
  assign n8259 = ( n8027 & ~n8257 ) | ( n8027 & n8258 ) | ( ~n8257 & n8258 ) ;
  assign n8260 = ( n8039 & n8122 ) | ( n8039 & n8259 ) | ( n8122 & n8259 ) ;
  assign n8261 = ( ~n8039 & n8122 ) | ( ~n8039 & n8259 ) | ( n8122 & n8259 ) ;
  assign n8262 = ( n8039 & ~n8260 ) | ( n8039 & n8261 ) | ( ~n8260 & n8261 ) ;
  assign n8263 = n1617 & n3326 ;
  assign n8264 = x100 & n1621 ;
  assign n8265 = x101 | n8264 ;
  assign n8266 = ( n1623 & n8264 ) | ( n1623 & n8265 ) | ( n8264 & n8265 ) ;
  assign n8267 = x99 & n1749 ;
  assign n8268 = n8266 | n8267 ;
  assign n8269 = ( x26 & n8263 ) | ( x26 & ~n8268 ) | ( n8263 & ~n8268 ) ;
  assign n8270 = ( ~x26 & n8268 ) | ( ~x26 & n8269 ) | ( n8268 & n8269 ) ;
  assign n8271 = ( ~n8263 & n8269 ) | ( ~n8263 & n8270 ) | ( n8269 & n8270 ) ;
  assign n8272 = ( n8042 & n8262 ) | ( n8042 & n8271 ) | ( n8262 & n8271 ) ;
  assign n8273 = ( ~n8042 & n8262 ) | ( ~n8042 & n8271 ) | ( n8262 & n8271 ) ;
  assign n8274 = ( n8042 & ~n8272 ) | ( n8042 & n8273 ) | ( ~n8272 & n8273 ) ;
  assign n8275 = n1297 & n3665 ;
  assign n8276 = x103 & n1301 ;
  assign n8277 = x104 | n8276 ;
  assign n8278 = ( n1303 & n8276 ) | ( n1303 & n8277 ) | ( n8276 & n8277 ) ;
  assign n8279 = x102 & n1426 ;
  assign n8280 = n8278 | n8279 ;
  assign n8281 = ( x23 & n8275 ) | ( x23 & ~n8280 ) | ( n8275 & ~n8280 ) ;
  assign n8282 = ( ~x23 & n8280 ) | ( ~x23 & n8281 ) | ( n8280 & n8281 ) ;
  assign n8283 = ( ~n8275 & n8281 ) | ( ~n8275 & n8282 ) | ( n8281 & n8282 ) ;
  assign n8284 = ( n8054 & n8274 ) | ( n8054 & n8283 ) | ( n8274 & n8283 ) ;
  assign n8285 = ( ~n8054 & n8274 ) | ( ~n8054 & n8283 ) | ( n8274 & n8283 ) ;
  assign n8286 = ( n8054 & ~n8284 ) | ( n8054 & n8285 ) | ( ~n8284 & n8285 ) ;
  assign n8287 = n1016 & n4362 ;
  assign n8288 = x106 & n1020 ;
  assign n8289 = x107 | n8288 ;
  assign n8290 = ( n1022 & n8288 ) | ( n1022 & n8289 ) | ( n8288 & n8289 ) ;
  assign n8291 = x105 & n1145 ;
  assign n8292 = n8290 | n8291 ;
  assign n8293 = ( x20 & n8287 ) | ( x20 & ~n8292 ) | ( n8287 & ~n8292 ) ;
  assign n8294 = ( ~x20 & n8292 ) | ( ~x20 & n8293 ) | ( n8292 & n8293 ) ;
  assign n8295 = ( ~n8287 & n8293 ) | ( ~n8287 & n8294 ) | ( n8293 & n8294 ) ;
  assign n8296 = ( n8066 & n8286 ) | ( n8066 & n8295 ) | ( n8286 & n8295 ) ;
  assign n8297 = ( ~n8066 & n8286 ) | ( ~n8066 & n8295 ) | ( n8286 & n8295 ) ;
  assign n8298 = ( n8066 & ~n8296 ) | ( n8066 & n8297 ) | ( ~n8296 & n8297 ) ;
  assign n8299 = ( n8069 & n8113 ) | ( n8069 & n8298 ) | ( n8113 & n8298 ) ;
  assign n8300 = ( ~n8069 & n8113 ) | ( ~n8069 & n8298 ) | ( n8113 & n8298 ) ;
  assign n8301 = ( n8069 & ~n8299 ) | ( n8069 & n8300 ) | ( ~n8299 & n8300 ) ;
  assign n8302 = ( n8072 & n8104 ) | ( n8072 & n8301 ) | ( n8104 & n8301 ) ;
  assign n8303 = ( ~n8072 & n8104 ) | ( ~n8072 & n8301 ) | ( n8104 & n8301 ) ;
  assign n8304 = ( n8072 & ~n8302 ) | ( n8072 & n8303 ) | ( ~n8302 & n8303 ) ;
  assign n8305 = ( n8075 & n8095 ) | ( n8075 & n8304 ) | ( n8095 & n8304 ) ;
  assign n8306 = ( ~n8075 & n8095 ) | ( ~n8075 & n8304 ) | ( n8095 & n8304 ) ;
  assign n8307 = ( n8075 & ~n8305 ) | ( n8075 & n8306 ) | ( ~n8305 & n8306 ) ;
  assign n8308 = n291 & n6645 ;
  assign n8309 = x118 & n295 ;
  assign n8310 = x119 | n8309 ;
  assign n8311 = ( n297 & n8309 ) | ( n297 & n8310 ) | ( n8309 & n8310 ) ;
  assign n8312 = x117 & n330 ;
  assign n8313 = n8311 | n8312 ;
  assign n8314 = ( x8 & n8308 ) | ( x8 & ~n8313 ) | ( n8308 & ~n8313 ) ;
  assign n8315 = ( ~x8 & n8313 ) | ( ~x8 & n8314 ) | ( n8313 & n8314 ) ;
  assign n8316 = ( ~n8308 & n8314 ) | ( ~n8308 & n8315 ) | ( n8314 & n8315 ) ;
  assign n8317 = ( n8078 & n8307 ) | ( n8078 & n8316 ) | ( n8307 & n8316 ) ;
  assign n8318 = ( ~n8078 & n8307 ) | ( ~n8078 & n8316 ) | ( n8307 & n8316 ) ;
  assign n8319 = ( n8078 & ~n8317 ) | ( n8078 & n8318 ) | ( ~n8317 & n8318 ) ;
  assign n8320 = n186 & n7582 ;
  assign n8321 = x121 & n190 ;
  assign n8322 = x122 | n8321 ;
  assign n8323 = ( n192 & n8321 ) | ( n192 & n8322 ) | ( n8321 & n8322 ) ;
  assign n8324 = x120 & n220 ;
  assign n8325 = n8323 | n8324 ;
  assign n8326 = ( x5 & n8320 ) | ( x5 & ~n8325 ) | ( n8320 & ~n8325 ) ;
  assign n8327 = ( ~x5 & n8325 ) | ( ~x5 & n8326 ) | ( n8325 & n8326 ) ;
  assign n8328 = ( ~n8320 & n8326 ) | ( ~n8320 & n8327 ) | ( n8326 & n8327 ) ;
  assign n8329 = ( x124 & x125 ) | ( x124 & n7839 ) | ( x125 & n7839 ) ;
  assign n8330 = ( x124 & ~x125 ) | ( x124 & n7839 ) | ( ~x125 & n7839 ) ;
  assign n8331 = ( x125 & ~n8329 ) | ( x125 & n8330 ) | ( ~n8329 & n8330 ) ;
  assign n8332 = n136 & n8331 ;
  assign n8333 = x124 & n138 ;
  assign n8334 = x125 | n8333 ;
  assign n8335 = ( n141 & n8333 ) | ( n141 & n8334 ) | ( n8333 & n8334 ) ;
  assign n8336 = x123 & n154 ;
  assign n8337 = n8335 | n8336 ;
  assign n8338 = ( x2 & n8332 ) | ( x2 & ~n8337 ) | ( n8332 & ~n8337 ) ;
  assign n8339 = ( ~x2 & n8337 ) | ( ~x2 & n8338 ) | ( n8337 & n8338 ) ;
  assign n8340 = ( ~n8332 & n8338 ) | ( ~n8332 & n8339 ) | ( n8338 & n8339 ) ;
  assign n8341 = ( n8319 & n8328 ) | ( n8319 & n8340 ) | ( n8328 & n8340 ) ;
  assign n8342 = ( ~n8319 & n8328 ) | ( ~n8319 & n8340 ) | ( n8328 & n8340 ) ;
  assign n8343 = ( n8319 & ~n8341 ) | ( n8319 & n8342 ) | ( ~n8341 & n8342 ) ;
  assign n8344 = ( n8081 & n8084 ) | ( n8081 & n8343 ) | ( n8084 & n8343 ) ;
  assign n8345 = ( ~n8081 & n8084 ) | ( ~n8081 & n8343 ) | ( n8084 & n8343 ) ;
  assign n8346 = ( n8081 & ~n8344 ) | ( n8081 & n8345 ) | ( ~n8344 & n8345 ) ;
  assign n8347 = n407 & n6201 ;
  assign n8348 = x116 & n411 ;
  assign n8349 = x117 | n8348 ;
  assign n8350 = ( n413 & n8348 ) | ( n413 & n8349 ) | ( n8348 & n8349 ) ;
  assign n8351 = x115 & n491 ;
  assign n8352 = n8350 | n8351 ;
  assign n8353 = ( x11 & n8347 ) | ( x11 & ~n8352 ) | ( n8347 & ~n8352 ) ;
  assign n8354 = ( ~x11 & n8352 ) | ( ~x11 & n8353 ) | ( n8352 & n8353 ) ;
  assign n8355 = ( ~n8347 & n8353 ) | ( ~n8347 & n8354 ) | ( n8353 & n8354 ) ;
  assign n8356 = n810 & n5130 ;
  assign n8357 = x110 & n814 ;
  assign n8358 = x111 | n8357 ;
  assign n8359 = ( n816 & n8357 ) | ( n816 & n8358 ) | ( n8357 & n8358 ) ;
  assign n8360 = x109 & n885 ;
  assign n8361 = n8359 | n8360 ;
  assign n8362 = ( x17 & n8356 ) | ( x17 & ~n8361 ) | ( n8356 & ~n8361 ) ;
  assign n8363 = ( ~x17 & n8361 ) | ( ~x17 & n8362 ) | ( n8361 & n8362 ) ;
  assign n8364 = ( ~n8356 & n8362 ) | ( ~n8356 & n8363 ) | ( n8362 & n8363 ) ;
  assign n8365 = n1016 & n4377 ;
  assign n8366 = x107 & n1020 ;
  assign n8367 = x108 | n8366 ;
  assign n8368 = ( n1022 & n8366 ) | ( n1022 & n8367 ) | ( n8366 & n8367 ) ;
  assign n8369 = x106 & n1145 ;
  assign n8370 = n8368 | n8369 ;
  assign n8371 = ( x20 & n8365 ) | ( x20 & ~n8370 ) | ( n8365 & ~n8370 ) ;
  assign n8372 = ( ~x20 & n8370 ) | ( ~x20 & n8371 ) | ( n8370 & n8371 ) ;
  assign n8373 = ( ~n8365 & n8371 ) | ( ~n8365 & n8372 ) | ( n8371 & n8372 ) ;
  assign n8374 = n1949 & n2877 ;
  assign n8375 = x98 & n1953 ;
  assign n8376 = x99 | n8375 ;
  assign n8377 = ( n1955 & n8375 ) | ( n1955 & n8376 ) | ( n8375 & n8376 ) ;
  assign n8378 = x97 & n2114 ;
  assign n8379 = n8377 | n8378 ;
  assign n8380 = ( x29 & n8374 ) | ( x29 & ~n8379 ) | ( n8374 & ~n8379 ) ;
  assign n8381 = ( ~x29 & n8379 ) | ( ~x29 & n8380 ) | ( n8379 & n8380 ) ;
  assign n8382 = ( ~n8374 & n8380 ) | ( ~n8374 & n8381 ) | ( n8380 & n8381 ) ;
  assign n8383 = n1466 & n3715 ;
  assign n8384 = x86 & n3719 ;
  assign n8385 = x87 | n8384 ;
  assign n8386 = ( n3721 & n8384 ) | ( n3721 & n8385 ) | ( n8384 & n8385 ) ;
  assign n8387 = x85 & n3922 ;
  assign n8388 = n8386 | n8387 ;
  assign n8389 = ( x41 & n8383 ) | ( x41 & ~n8388 ) | ( n8383 & ~n8388 ) ;
  assign n8390 = ( ~x41 & n8388 ) | ( ~x41 & n8389 ) | ( n8388 & n8389 ) ;
  assign n8391 = ( ~n8383 & n8389 ) | ( ~n8383 & n8390 ) | ( n8389 & n8390 ) ;
  assign n8392 = n1097 & n4227 ;
  assign n8393 = x83 & n4231 ;
  assign n8394 = x84 | n8393 ;
  assign n8395 = ( n4233 & n8393 ) | ( n4233 & n8394 ) | ( n8393 & n8394 ) ;
  assign n8396 = x82 & n4470 ;
  assign n8397 = n8395 | n8396 ;
  assign n8398 = ( x44 & n8392 ) | ( x44 & ~n8397 ) | ( n8392 & ~n8397 ) ;
  assign n8399 = ( ~x44 & n8397 ) | ( ~x44 & n8398 ) | ( n8397 & n8398 ) ;
  assign n8400 = ( ~n8392 & n8398 ) | ( ~n8392 & n8399 ) | ( n8398 & n8399 ) ;
  assign n8401 = n910 & n4787 ;
  assign n8402 = x80 & n4791 ;
  assign n8403 = x81 | n8402 ;
  assign n8404 = ( n4793 & n8402 ) | ( n4793 & n8403 ) | ( n8402 & n8403 ) ;
  assign n8405 = x79 & n5030 ;
  assign n8406 = n8404 | n8405 ;
  assign n8407 = ( x47 & n8401 ) | ( x47 & ~n8406 ) | ( n8401 & ~n8406 ) ;
  assign n8408 = ( ~x47 & n8406 ) | ( ~x47 & n8407 ) | ( n8406 & n8407 ) ;
  assign n8409 = ( ~n8401 & n8407 ) | ( ~n8401 & n8408 ) | ( n8407 & n8408 ) ;
  assign n8410 = n461 & n6027 ;
  assign n8411 = x74 & n6031 ;
  assign n8412 = x75 | n8411 ;
  assign n8413 = ( n6033 & n8411 ) | ( n6033 & n8412 ) | ( n8411 & n8412 ) ;
  assign n8414 = x73 & n6303 ;
  assign n8415 = n8413 | n8414 ;
  assign n8416 = ( x53 & n8410 ) | ( x53 & ~n8415 ) | ( n8410 & ~n8415 ) ;
  assign n8417 = ( ~x53 & n8415 ) | ( ~x53 & n8416 ) | ( n8415 & n8416 ) ;
  assign n8418 = ( ~n8410 & n8416 ) | ( ~n8410 & n8417 ) | ( n8416 & n8417 ) ;
  assign n8419 = n346 & n6713 ;
  assign n8420 = x71 & n6717 ;
  assign n8421 = x72 | n8420 ;
  assign n8422 = ( n6719 & n8420 ) | ( n6719 & n8421 ) | ( n8420 & n8421 ) ;
  assign n8423 = x70 & n6980 ;
  assign n8424 = n8422 | n8423 ;
  assign n8425 = ( x56 & n8419 ) | ( x56 & ~n8424 ) | ( n8419 & ~n8424 ) ;
  assign n8426 = ( ~x56 & n8424 ) | ( ~x56 & n8425 ) | ( n8424 & n8425 ) ;
  assign n8427 = ( ~n8419 & n8425 ) | ( ~n8419 & n8426 ) | ( n8425 & n8426 ) ;
  assign n8428 = n230 & n7423 ;
  assign n8429 = x68 & n7427 ;
  assign n8430 = x69 | n8429 ;
  assign n8431 = ( n7429 & n8429 ) | ( n7429 & n8430 ) | ( n8429 & n8430 ) ;
  assign n8432 = x67 & n7708 ;
  assign n8433 = n8431 | n8432 ;
  assign n8434 = ( ~x59 & n8428 ) | ( ~x59 & n8433 ) | ( n8428 & n8433 ) ;
  assign n8435 = ( n8428 & n8433 ) | ( n8428 & ~n8434 ) | ( n8433 & ~n8434 ) ;
  assign n8436 = ( x59 & n8434 ) | ( x59 & ~n8435 ) | ( n8434 & ~n8435 ) ;
  assign n8437 = ( x62 & n8150 ) | ( x62 & n8164 ) | ( n8150 & n8164 ) ;
  assign n8438 = ( x59 & ~x61 ) | ( x59 & n8153 ) | ( ~x61 & n8153 ) ;
  assign n8439 = ( ~n7960 & n8157 ) | ( ~n7960 & n8438 ) | ( n8157 & n8438 ) ;
  assign n8440 = x64 & n8439 ;
  assign n8441 = x65 & n8158 ;
  assign n8442 = x66 | n8441 ;
  assign n8443 = ( n8160 & n8441 ) | ( n8160 & n8442 ) | ( n8441 & n8442 ) ;
  assign n8444 = ( n151 & n152 ) | ( n151 & n8154 ) | ( n152 & n8154 ) ;
  assign n8445 = ( ~n8440 & n8443 ) | ( ~n8440 & n8444 ) | ( n8443 & n8444 ) ;
  assign n8446 = n8440 | n8445 ;
  assign n8447 = n8437 | n8446 ;
  assign n8448 = ( n8437 & n8446 ) | ( n8437 & ~n8447 ) | ( n8446 & ~n8447 ) ;
  assign n8449 = n8447 & ~n8448 ;
  assign n8450 = ( n8176 & n8436 ) | ( n8176 & n8449 ) | ( n8436 & n8449 ) ;
  assign n8451 = ( ~n8176 & n8436 ) | ( ~n8176 & n8449 ) | ( n8436 & n8449 ) ;
  assign n8452 = ( n8176 & ~n8450 ) | ( n8176 & n8451 ) | ( ~n8450 & n8451 ) ;
  assign n8453 = ( n8179 & n8427 ) | ( n8179 & n8452 ) | ( n8427 & n8452 ) ;
  assign n8454 = ( ~n8179 & n8427 ) | ( ~n8179 & n8452 ) | ( n8427 & n8452 ) ;
  assign n8455 = ( n8179 & ~n8453 ) | ( n8179 & n8454 ) | ( ~n8453 & n8454 ) ;
  assign n8456 = ( n8191 & n8418 ) | ( n8191 & n8455 ) | ( n8418 & n8455 ) ;
  assign n8457 = ( ~n8191 & n8418 ) | ( ~n8191 & n8455 ) | ( n8418 & n8455 ) ;
  assign n8458 = ( n8191 & ~n8456 ) | ( n8191 & n8457 ) | ( ~n8456 & n8457 ) ;
  assign n8459 = n637 & n5374 ;
  assign n8460 = x77 & n5378 ;
  assign n8461 = x78 | n8460 ;
  assign n8462 = ( n5380 & n8460 ) | ( n5380 & n8461 ) | ( n8460 & n8461 ) ;
  assign n8463 = x76 & n5638 ;
  assign n8464 = n8462 | n8463 ;
  assign n8465 = ( x50 & n8459 ) | ( x50 & ~n8464 ) | ( n8459 & ~n8464 ) ;
  assign n8466 = ( ~x50 & n8464 ) | ( ~x50 & n8465 ) | ( n8464 & n8465 ) ;
  assign n8467 = ( ~n8459 & n8465 ) | ( ~n8459 & n8466 ) | ( n8465 & n8466 ) ;
  assign n8468 = ( n8203 & n8458 ) | ( n8203 & n8467 ) | ( n8458 & n8467 ) ;
  assign n8469 = ( ~n8203 & n8458 ) | ( ~n8203 & n8467 ) | ( n8458 & n8467 ) ;
  assign n8470 = ( n8203 & ~n8468 ) | ( n8203 & n8469 ) | ( ~n8468 & n8469 ) ;
  assign n8471 = ( n8206 & n8409 ) | ( n8206 & n8470 ) | ( n8409 & n8470 ) ;
  assign n8472 = ( ~n8206 & n8409 ) | ( ~n8206 & n8470 ) | ( n8409 & n8470 ) ;
  assign n8473 = ( n8206 & ~n8471 ) | ( n8206 & n8472 ) | ( ~n8471 & n8472 ) ;
  assign n8474 = ( n8218 & n8400 ) | ( n8218 & n8473 ) | ( n8400 & n8473 ) ;
  assign n8475 = ( ~n8218 & n8400 ) | ( ~n8218 & n8473 ) | ( n8400 & n8473 ) ;
  assign n8476 = ( n8218 & ~n8474 ) | ( n8218 & n8475 ) | ( ~n8474 & n8475 ) ;
  assign n8477 = ( n8221 & n8391 ) | ( n8221 & n8476 ) | ( n8391 & n8476 ) ;
  assign n8478 = ( ~n8221 & n8391 ) | ( ~n8221 & n8476 ) | ( n8391 & n8476 ) ;
  assign n8479 = ( n8221 & ~n8477 ) | ( n8221 & n8478 ) | ( ~n8477 & n8478 ) ;
  assign n8480 = n1701 & n3224 ;
  assign n8481 = x89 & n3228 ;
  assign n8482 = x90 | n8481 ;
  assign n8483 = ( n3230 & n8481 ) | ( n3230 & n8482 ) | ( n8481 & n8482 ) ;
  assign n8484 = x88 & n3413 ;
  assign n8485 = n8483 | n8484 ;
  assign n8486 = ( x38 & n8480 ) | ( x38 & ~n8485 ) | ( n8480 & ~n8485 ) ;
  assign n8487 = ( ~x38 & n8485 ) | ( ~x38 & n8486 ) | ( n8485 & n8486 ) ;
  assign n8488 = ( ~n8480 & n8486 ) | ( ~n8480 & n8487 ) | ( n8486 & n8487 ) ;
  assign n8489 = ( n8233 & n8479 ) | ( n8233 & n8488 ) | ( n8479 & n8488 ) ;
  assign n8490 = ( ~n8233 & n8479 ) | ( ~n8233 & n8488 ) | ( n8479 & n8488 ) ;
  assign n8491 = ( n8233 & ~n8489 ) | ( n8233 & n8490 ) | ( ~n8489 & n8490 ) ;
  assign n8492 = n2057 & n2766 ;
  assign n8493 = x92 & n2770 ;
  assign n8494 = x93 | n8493 ;
  assign n8495 = ( n2772 & n8493 ) | ( n2772 & n8494 ) | ( n8493 & n8494 ) ;
  assign n8496 = x91 & n2943 ;
  assign n8497 = n8495 | n8496 ;
  assign n8498 = ( x35 & n8492 ) | ( x35 & ~n8497 ) | ( n8492 & ~n8497 ) ;
  assign n8499 = ( ~x35 & n8497 ) | ( ~x35 & n8498 ) | ( n8497 & n8498 ) ;
  assign n8500 = ( ~n8492 & n8498 ) | ( ~n8492 & n8499 ) | ( n8498 & n8499 ) ;
  assign n8501 = ( n8245 & n8491 ) | ( n8245 & n8500 ) | ( n8491 & n8500 ) ;
  assign n8502 = ( ~n8245 & n8491 ) | ( ~n8245 & n8500 ) | ( n8491 & n8500 ) ;
  assign n8503 = ( n8245 & ~n8501 ) | ( n8245 & n8502 ) | ( ~n8501 & n8502 ) ;
  assign n8504 = n2320 & n2449 ;
  assign n8505 = x95 & n2324 ;
  assign n8506 = x96 | n8505 ;
  assign n8507 = ( n2326 & n8505 ) | ( n2326 & n8506 ) | ( n8505 & n8506 ) ;
  assign n8508 = x94 & n2497 ;
  assign n8509 = n8507 | n8508 ;
  assign n8510 = ( x32 & n8504 ) | ( x32 & ~n8509 ) | ( n8504 & ~n8509 ) ;
  assign n8511 = ( ~x32 & n8509 ) | ( ~x32 & n8510 ) | ( n8509 & n8510 ) ;
  assign n8512 = ( ~n8504 & n8510 ) | ( ~n8504 & n8511 ) | ( n8510 & n8511 ) ;
  assign n8513 = ( n8257 & n8503 ) | ( n8257 & n8512 ) | ( n8503 & n8512 ) ;
  assign n8514 = ( ~n8257 & n8503 ) | ( ~n8257 & n8512 ) | ( n8503 & n8512 ) ;
  assign n8515 = ( n8257 & ~n8513 ) | ( n8257 & n8514 ) | ( ~n8513 & n8514 ) ;
  assign n8516 = ( n8260 & n8382 ) | ( n8260 & n8515 ) | ( n8382 & n8515 ) ;
  assign n8517 = ( ~n8260 & n8382 ) | ( ~n8260 & n8515 ) | ( n8382 & n8515 ) ;
  assign n8518 = ( n8260 & ~n8516 ) | ( n8260 & n8517 ) | ( ~n8516 & n8517 ) ;
  assign n8519 = n1617 & n3486 ;
  assign n8520 = x101 & n1621 ;
  assign n8521 = x102 | n8520 ;
  assign n8522 = ( n1623 & n8520 ) | ( n1623 & n8521 ) | ( n8520 & n8521 ) ;
  assign n8523 = x100 & n1749 ;
  assign n8524 = n8522 | n8523 ;
  assign n8525 = ( x26 & n8519 ) | ( x26 & ~n8524 ) | ( n8519 & ~n8524 ) ;
  assign n8526 = ( ~x26 & n8524 ) | ( ~x26 & n8525 ) | ( n8524 & n8525 ) ;
  assign n8527 = ( ~n8519 & n8525 ) | ( ~n8519 & n8526 ) | ( n8525 & n8526 ) ;
  assign n8528 = ( n8272 & n8518 ) | ( n8272 & n8527 ) | ( n8518 & n8527 ) ;
  assign n8529 = ( ~n8272 & n8518 ) | ( ~n8272 & n8527 ) | ( n8518 & n8527 ) ;
  assign n8530 = ( n8272 & ~n8528 ) | ( n8272 & n8529 ) | ( ~n8528 & n8529 ) ;
  assign n8531 = n1297 & n3998 ;
  assign n8532 = x104 & n1301 ;
  assign n8533 = x105 | n8532 ;
  assign n8534 = ( n1303 & n8532 ) | ( n1303 & n8533 ) | ( n8532 & n8533 ) ;
  assign n8535 = x103 & n1426 ;
  assign n8536 = n8534 | n8535 ;
  assign n8537 = ( x23 & n8531 ) | ( x23 & ~n8536 ) | ( n8531 & ~n8536 ) ;
  assign n8538 = ( ~x23 & n8536 ) | ( ~x23 & n8537 ) | ( n8536 & n8537 ) ;
  assign n8539 = ( ~n8531 & n8537 ) | ( ~n8531 & n8538 ) | ( n8537 & n8538 ) ;
  assign n8540 = ( n8284 & n8530 ) | ( n8284 & n8539 ) | ( n8530 & n8539 ) ;
  assign n8541 = ( ~n8284 & n8530 ) | ( ~n8284 & n8539 ) | ( n8530 & n8539 ) ;
  assign n8542 = ( n8284 & ~n8540 ) | ( n8284 & n8541 ) | ( ~n8540 & n8541 ) ;
  assign n8543 = ( n8296 & n8373 ) | ( n8296 & n8542 ) | ( n8373 & n8542 ) ;
  assign n8544 = ( ~n8296 & n8373 ) | ( ~n8296 & n8542 ) | ( n8373 & n8542 ) ;
  assign n8545 = ( n8296 & ~n8543 ) | ( n8296 & n8544 ) | ( ~n8543 & n8544 ) ;
  assign n8546 = ( n8299 & n8364 ) | ( n8299 & n8545 ) | ( n8364 & n8545 ) ;
  assign n8547 = ( ~n8299 & n8364 ) | ( ~n8299 & n8545 ) | ( n8364 & n8545 ) ;
  assign n8548 = ( n8299 & ~n8546 ) | ( n8299 & n8547 ) | ( ~n8546 & n8547 ) ;
  assign n8549 = n583 & n5750 ;
  assign n8550 = x113 & n587 ;
  assign n8551 = x114 | n8550 ;
  assign n8552 = ( n589 & n8550 ) | ( n589 & n8551 ) | ( n8550 & n8551 ) ;
  assign n8553 = x112 & n676 ;
  assign n8554 = n8552 | n8553 ;
  assign n8555 = ( x14 & n8549 ) | ( x14 & ~n8554 ) | ( n8549 & ~n8554 ) ;
  assign n8556 = ( ~x14 & n8554 ) | ( ~x14 & n8555 ) | ( n8554 & n8555 ) ;
  assign n8557 = ( ~n8549 & n8555 ) | ( ~n8549 & n8556 ) | ( n8555 & n8556 ) ;
  assign n8558 = ( n8302 & n8548 ) | ( n8302 & n8557 ) | ( n8548 & n8557 ) ;
  assign n8559 = ( ~n8302 & n8548 ) | ( ~n8302 & n8557 ) | ( n8548 & n8557 ) ;
  assign n8560 = ( n8302 & ~n8558 ) | ( n8302 & n8559 ) | ( ~n8558 & n8559 ) ;
  assign n8561 = ( n8305 & n8355 ) | ( n8305 & n8560 ) | ( n8355 & n8560 ) ;
  assign n8562 = ( ~n8305 & n8355 ) | ( ~n8305 & n8560 ) | ( n8355 & n8560 ) ;
  assign n8563 = ( n8305 & ~n8561 ) | ( n8305 & n8562 ) | ( ~n8561 & n8562 ) ;
  assign n8564 = n291 & n7098 ;
  assign n8565 = x119 & n295 ;
  assign n8566 = x120 | n8565 ;
  assign n8567 = ( n297 & n8565 ) | ( n297 & n8566 ) | ( n8565 & n8566 ) ;
  assign n8568 = x118 & n330 ;
  assign n8569 = n8567 | n8568 ;
  assign n8570 = ( x8 & n8564 ) | ( x8 & ~n8569 ) | ( n8564 & ~n8569 ) ;
  assign n8571 = ( ~x8 & n8569 ) | ( ~x8 & n8570 ) | ( n8569 & n8570 ) ;
  assign n8572 = ( ~n8564 & n8570 ) | ( ~n8564 & n8571 ) | ( n8570 & n8571 ) ;
  assign n8573 = n186 & n7597 ;
  assign n8574 = x122 & n190 ;
  assign n8575 = x123 | n8574 ;
  assign n8576 = ( n192 & n8574 ) | ( n192 & n8575 ) | ( n8574 & n8575 ) ;
  assign n8577 = x121 & n220 ;
  assign n8578 = n8576 | n8577 ;
  assign n8579 = ( x5 & n8573 ) | ( x5 & ~n8578 ) | ( n8573 & ~n8578 ) ;
  assign n8580 = ( ~x5 & n8578 ) | ( ~x5 & n8579 ) | ( n8578 & n8579 ) ;
  assign n8581 = ( ~n8573 & n8579 ) | ( ~n8573 & n8580 ) | ( n8579 & n8580 ) ;
  assign n8582 = ( n8563 & n8572 ) | ( n8563 & n8581 ) | ( n8572 & n8581 ) ;
  assign n8583 = ( ~n8563 & n8572 ) | ( ~n8563 & n8581 ) | ( n8572 & n8581 ) ;
  assign n8584 = ( n8563 & ~n8582 ) | ( n8563 & n8583 ) | ( ~n8582 & n8583 ) ;
  assign n8585 = ( x125 & x126 ) | ( x125 & n8329 ) | ( x126 & n8329 ) ;
  assign n8586 = ( x125 & ~x126 ) | ( x125 & n8329 ) | ( ~x126 & n8329 ) ;
  assign n8587 = ( x126 & ~n8585 ) | ( x126 & n8586 ) | ( ~n8585 & n8586 ) ;
  assign n8588 = n136 & n8587 ;
  assign n8589 = x125 & n138 ;
  assign n8590 = x126 | n8589 ;
  assign n8591 = ( n141 & n8589 ) | ( n141 & n8590 ) | ( n8589 & n8590 ) ;
  assign n8592 = x124 & n154 ;
  assign n8593 = n8591 | n8592 ;
  assign n8594 = ( x2 & n8588 ) | ( x2 & ~n8593 ) | ( n8588 & ~n8593 ) ;
  assign n8595 = ( ~x2 & n8593 ) | ( ~x2 & n8594 ) | ( n8593 & n8594 ) ;
  assign n8596 = ( ~n8588 & n8594 ) | ( ~n8588 & n8595 ) | ( n8594 & n8595 ) ;
  assign n8597 = ( n8317 & n8584 ) | ( n8317 & n8596 ) | ( n8584 & n8596 ) ;
  assign n8598 = ( ~n8317 & n8584 ) | ( ~n8317 & n8596 ) | ( n8584 & n8596 ) ;
  assign n8599 = ( n8317 & ~n8597 ) | ( n8317 & n8598 ) | ( ~n8597 & n8598 ) ;
  assign n8600 = ( n8341 & n8344 ) | ( n8341 & n8599 ) | ( n8344 & n8599 ) ;
  assign n8601 = ( n8341 & ~n8344 ) | ( n8341 & n8599 ) | ( ~n8344 & n8599 ) ;
  assign n8602 = ( n8344 & ~n8600 ) | ( n8344 & n8601 ) | ( ~n8600 & n8601 ) ;
  assign n8603 = n186 & n7841 ;
  assign n8604 = x123 & n190 ;
  assign n8605 = x124 | n8604 ;
  assign n8606 = ( n192 & n8604 ) | ( n192 & n8605 ) | ( n8604 & n8605 ) ;
  assign n8607 = x122 & n220 ;
  assign n8608 = n8606 | n8607 ;
  assign n8609 = ( x5 & n8603 ) | ( x5 & ~n8608 ) | ( n8603 & ~n8608 ) ;
  assign n8610 = ( ~x5 & n8608 ) | ( ~x5 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8611 = ( ~n8603 & n8609 ) | ( ~n8603 & n8610 ) | ( n8609 & n8610 ) ;
  assign n8612 = n583 & n5765 ;
  assign n8613 = x114 & n587 ;
  assign n8614 = x115 | n8613 ;
  assign n8615 = ( n589 & n8613 ) | ( n589 & n8614 ) | ( n8613 & n8614 ) ;
  assign n8616 = x113 & n676 ;
  assign n8617 = n8615 | n8616 ;
  assign n8618 = ( x14 & n8612 ) | ( x14 & ~n8617 ) | ( n8612 & ~n8617 ) ;
  assign n8619 = ( ~x14 & n8617 ) | ( ~x14 & n8618 ) | ( n8617 & n8618 ) ;
  assign n8620 = ( ~n8612 & n8618 ) | ( ~n8612 & n8619 ) | ( n8618 & n8619 ) ;
  assign n8621 = n810 & n5145 ;
  assign n8622 = x111 & n814 ;
  assign n8623 = x112 | n8622 ;
  assign n8624 = ( n816 & n8622 ) | ( n816 & n8623 ) | ( n8622 & n8623 ) ;
  assign n8625 = x110 & n885 ;
  assign n8626 = n8624 | n8625 ;
  assign n8627 = ( x17 & n8621 ) | ( x17 & ~n8626 ) | ( n8621 & ~n8626 ) ;
  assign n8628 = ( ~x17 & n8626 ) | ( ~x17 & n8627 ) | ( n8626 & n8627 ) ;
  assign n8629 = ( ~n8621 & n8627 ) | ( ~n8621 & n8628 ) | ( n8627 & n8628 ) ;
  assign n8630 = n1016 & n4734 ;
  assign n8631 = x108 & n1020 ;
  assign n8632 = x109 | n8631 ;
  assign n8633 = ( n1022 & n8631 ) | ( n1022 & n8632 ) | ( n8631 & n8632 ) ;
  assign n8634 = x107 & n1145 ;
  assign n8635 = n8633 | n8634 ;
  assign n8636 = ( x20 & n8630 ) | ( x20 & ~n8635 ) | ( n8630 & ~n8635 ) ;
  assign n8637 = ( ~x20 & n8635 ) | ( ~x20 & n8636 ) | ( n8635 & n8636 ) ;
  assign n8638 = ( ~n8630 & n8636 ) | ( ~n8630 & n8637 ) | ( n8636 & n8637 ) ;
  assign n8639 = n1297 & n4013 ;
  assign n8640 = x105 & n1301 ;
  assign n8641 = x106 | n8640 ;
  assign n8642 = ( n1303 & n8640 ) | ( n1303 & n8641 ) | ( n8640 & n8641 ) ;
  assign n8643 = x104 & n1426 ;
  assign n8644 = n8642 | n8643 ;
  assign n8645 = ( x23 & n8639 ) | ( x23 & ~n8644 ) | ( n8639 & ~n8644 ) ;
  assign n8646 = ( ~x23 & n8644 ) | ( ~x23 & n8645 ) | ( n8644 & n8645 ) ;
  assign n8647 = ( ~n8639 & n8645 ) | ( ~n8639 & n8646 ) | ( n8645 & n8646 ) ;
  assign n8648 = n1949 & n3162 ;
  assign n8649 = x99 & n1953 ;
  assign n8650 = x100 | n8649 ;
  assign n8651 = ( n1955 & n8649 ) | ( n1955 & n8650 ) | ( n8649 & n8650 ) ;
  assign n8652 = x98 & n2114 ;
  assign n8653 = n8651 | n8652 ;
  assign n8654 = ( x29 & n8648 ) | ( x29 & ~n8653 ) | ( n8648 & ~n8653 ) ;
  assign n8655 = ( ~x29 & n8653 ) | ( ~x29 & n8654 ) | ( n8653 & n8654 ) ;
  assign n8656 = ( ~n8648 & n8654 ) | ( ~n8648 & n8655 ) | ( n8654 & n8655 ) ;
  assign n8657 = n1262 & n4227 ;
  assign n8658 = x84 & n4231 ;
  assign n8659 = x85 | n8658 ;
  assign n8660 = ( n4233 & n8658 ) | ( n4233 & n8659 ) | ( n8658 & n8659 ) ;
  assign n8661 = x83 & n4470 ;
  assign n8662 = n8660 | n8661 ;
  assign n8663 = ( x44 & n8657 ) | ( x44 & ~n8662 ) | ( n8657 & ~n8662 ) ;
  assign n8664 = ( ~x44 & n8662 ) | ( ~x44 & n8663 ) | ( n8662 & n8663 ) ;
  assign n8665 = ( ~n8657 & n8663 ) | ( ~n8657 & n8664 ) | ( n8663 & n8664 ) ;
  assign n8666 = n554 & n6027 ;
  assign n8667 = x75 & n6031 ;
  assign n8668 = x76 | n8667 ;
  assign n8669 = ( n6033 & n8667 ) | ( n6033 & n8668 ) | ( n8667 & n8668 ) ;
  assign n8670 = x74 & n6303 ;
  assign n8671 = n8669 | n8670 ;
  assign n8672 = ( x53 & n8666 ) | ( x53 & ~n8671 ) | ( n8666 & ~n8671 ) ;
  assign n8673 = ( ~x53 & n8671 ) | ( ~x53 & n8672 ) | ( n8671 & n8672 ) ;
  assign n8674 = ( ~n8666 & n8672 ) | ( ~n8666 & n8673 ) | ( n8672 & n8673 ) ;
  assign n8675 = n245 & n7423 ;
  assign n8676 = x69 & n7427 ;
  assign n8677 = x70 | n8676 ;
  assign n8678 = ( n7429 & n8676 ) | ( n7429 & n8677 ) | ( n8676 & n8677 ) ;
  assign n8679 = x68 & n7708 ;
  assign n8680 = n8678 | n8679 ;
  assign n8681 = ( x59 & n8675 ) | ( x59 & ~n8680 ) | ( n8675 & ~n8680 ) ;
  assign n8682 = ( ~x59 & n8680 ) | ( ~x59 & n8681 ) | ( n8680 & n8681 ) ;
  assign n8683 = ( ~n8675 & n8681 ) | ( ~n8675 & n8682 ) | ( n8681 & n8682 ) ;
  assign n8684 = x66 & n8158 ;
  assign n8685 = x67 | n8684 ;
  assign n8686 = ( n8160 & n8684 ) | ( n8160 & n8685 ) | ( n8684 & n8685 ) ;
  assign n8687 = x65 & n8439 ;
  assign n8688 = n8686 | n8687 ;
  assign n8689 = n164 & n8154 ;
  assign n8690 = ( x62 & n8688 ) | ( x62 & ~n8689 ) | ( n8688 & ~n8689 ) ;
  assign n8691 = ( ~x62 & n8689 ) | ( ~x62 & n8690 ) | ( n8689 & n8690 ) ;
  assign n8692 = ( ~n8688 & n8690 ) | ( ~n8688 & n8691 ) | ( n8690 & n8691 ) ;
  assign n8693 = x62 | x63 ;
  assign n8694 = ( x62 & x63 ) | ( x62 & ~x64 ) | ( x63 & ~x64 ) ;
  assign n8695 = n8693 & ~n8694 ;
  assign n8696 = x62 & ~n8447 ;
  assign n8697 = ( n8692 & n8695 ) | ( n8692 & n8696 ) | ( n8695 & n8696 ) ;
  assign n8698 = ( ~n8692 & n8695 ) | ( ~n8692 & n8696 ) | ( n8695 & n8696 ) ;
  assign n8699 = ( n8692 & ~n8697 ) | ( n8692 & n8698 ) | ( ~n8697 & n8698 ) ;
  assign n8700 = ( n8450 & n8683 ) | ( n8450 & n8699 ) | ( n8683 & n8699 ) ;
  assign n8701 = ( ~n8450 & n8683 ) | ( ~n8450 & n8699 ) | ( n8683 & n8699 ) ;
  assign n8702 = ( n8450 & ~n8700 ) | ( n8450 & n8701 ) | ( ~n8700 & n8701 ) ;
  assign n8703 = n390 & n6713 ;
  assign n8704 = x72 & n6717 ;
  assign n8705 = x73 | n8704 ;
  assign n8706 = ( n6719 & n8704 ) | ( n6719 & n8705 ) | ( n8704 & n8705 ) ;
  assign n8707 = x71 & n6980 ;
  assign n8708 = n8706 | n8707 ;
  assign n8709 = ( x56 & n8703 ) | ( x56 & ~n8708 ) | ( n8703 & ~n8708 ) ;
  assign n8710 = ( ~x56 & n8708 ) | ( ~x56 & n8709 ) | ( n8708 & n8709 ) ;
  assign n8711 = ( ~n8703 & n8709 ) | ( ~n8703 & n8710 ) | ( n8709 & n8710 ) ;
  assign n8712 = ( n8453 & n8702 ) | ( n8453 & n8711 ) | ( n8702 & n8711 ) ;
  assign n8713 = ( ~n8453 & n8702 ) | ( ~n8453 & n8711 ) | ( n8702 & n8711 ) ;
  assign n8714 = ( n8453 & ~n8712 ) | ( n8453 & n8713 ) | ( ~n8712 & n8713 ) ;
  assign n8715 = ( n8456 & n8674 ) | ( n8456 & n8714 ) | ( n8674 & n8714 ) ;
  assign n8716 = ( ~n8456 & n8674 ) | ( ~n8456 & n8714 ) | ( n8674 & n8714 ) ;
  assign n8717 = ( n8456 & ~n8715 ) | ( n8456 & n8716 ) | ( ~n8715 & n8716 ) ;
  assign n8718 = n701 & n5374 ;
  assign n8719 = x78 & n5378 ;
  assign n8720 = x79 | n8719 ;
  assign n8721 = ( n5380 & n8719 ) | ( n5380 & n8720 ) | ( n8719 & n8720 ) ;
  assign n8722 = x77 & n5638 ;
  assign n8723 = n8721 | n8722 ;
  assign n8724 = ( x50 & n8718 ) | ( x50 & ~n8723 ) | ( n8718 & ~n8723 ) ;
  assign n8725 = ( ~x50 & n8723 ) | ( ~x50 & n8724 ) | ( n8723 & n8724 ) ;
  assign n8726 = ( ~n8718 & n8724 ) | ( ~n8718 & n8725 ) | ( n8724 & n8725 ) ;
  assign n8727 = ( n8468 & n8717 ) | ( n8468 & n8726 ) | ( n8717 & n8726 ) ;
  assign n8728 = ( ~n8468 & n8717 ) | ( ~n8468 & n8726 ) | ( n8717 & n8726 ) ;
  assign n8729 = ( n8468 & ~n8727 ) | ( n8468 & n8728 ) | ( ~n8727 & n8728 ) ;
  assign n8730 = n990 & n4787 ;
  assign n8731 = x81 & n4791 ;
  assign n8732 = x82 | n8731 ;
  assign n8733 = ( n4793 & n8731 ) | ( n4793 & n8732 ) | ( n8731 & n8732 ) ;
  assign n8734 = x80 & n5030 ;
  assign n8735 = n8733 | n8734 ;
  assign n8736 = ( x47 & n8730 ) | ( x47 & ~n8735 ) | ( n8730 & ~n8735 ) ;
  assign n8737 = ( ~x47 & n8735 ) | ( ~x47 & n8736 ) | ( n8735 & n8736 ) ;
  assign n8738 = ( ~n8730 & n8736 ) | ( ~n8730 & n8737 ) | ( n8736 & n8737 ) ;
  assign n8739 = ( n8471 & n8729 ) | ( n8471 & n8738 ) | ( n8729 & n8738 ) ;
  assign n8740 = ( ~n8471 & n8729 ) | ( ~n8471 & n8738 ) | ( n8729 & n8738 ) ;
  assign n8741 = ( n8471 & ~n8739 ) | ( n8471 & n8740 ) | ( ~n8739 & n8740 ) ;
  assign n8742 = ( n8474 & n8665 ) | ( n8474 & n8741 ) | ( n8665 & n8741 ) ;
  assign n8743 = ( ~n8474 & n8665 ) | ( ~n8474 & n8741 ) | ( n8665 & n8741 ) ;
  assign n8744 = ( n8474 & ~n8742 ) | ( n8474 & n8743 ) | ( ~n8742 & n8743 ) ;
  assign n8745 = n1481 & n3715 ;
  assign n8746 = x87 & n3719 ;
  assign n8747 = x88 | n8746 ;
  assign n8748 = ( n3721 & n8746 ) | ( n3721 & n8747 ) | ( n8746 & n8747 ) ;
  assign n8749 = x86 & n3922 ;
  assign n8750 = n8748 | n8749 ;
  assign n8751 = ( x41 & n8745 ) | ( x41 & ~n8750 ) | ( n8745 & ~n8750 ) ;
  assign n8752 = ( ~x41 & n8750 ) | ( ~x41 & n8751 ) | ( n8750 & n8751 ) ;
  assign n8753 = ( ~n8745 & n8751 ) | ( ~n8745 & n8752 ) | ( n8751 & n8752 ) ;
  assign n8754 = ( n8477 & n8744 ) | ( n8477 & n8753 ) | ( n8744 & n8753 ) ;
  assign n8755 = ( ~n8477 & n8744 ) | ( ~n8477 & n8753 ) | ( n8744 & n8753 ) ;
  assign n8756 = ( n8477 & ~n8754 ) | ( n8477 & n8755 ) | ( ~n8754 & n8755 ) ;
  assign n8757 = n1914 & n3224 ;
  assign n8758 = x90 & n3228 ;
  assign n8759 = x91 | n8758 ;
  assign n8760 = ( n3230 & n8758 ) | ( n3230 & n8759 ) | ( n8758 & n8759 ) ;
  assign n8761 = x89 & n3413 ;
  assign n8762 = n8760 | n8761 ;
  assign n8763 = ( x38 & n8757 ) | ( x38 & ~n8762 ) | ( n8757 & ~n8762 ) ;
  assign n8764 = ( ~x38 & n8762 ) | ( ~x38 & n8763 ) | ( n8762 & n8763 ) ;
  assign n8765 = ( ~n8757 & n8763 ) | ( ~n8757 & n8764 ) | ( n8763 & n8764 ) ;
  assign n8766 = ( n8489 & n8756 ) | ( n8489 & n8765 ) | ( n8756 & n8765 ) ;
  assign n8767 = ( ~n8489 & n8756 ) | ( ~n8489 & n8765 ) | ( n8756 & n8765 ) ;
  assign n8768 = ( n8489 & ~n8766 ) | ( n8489 & n8767 ) | ( ~n8766 & n8767 ) ;
  assign n8769 = n2294 & n2766 ;
  assign n8770 = x93 & n2770 ;
  assign n8771 = x94 | n8770 ;
  assign n8772 = ( n2772 & n8770 ) | ( n2772 & n8771 ) | ( n8770 & n8771 ) ;
  assign n8773 = x92 & n2943 ;
  assign n8774 = n8772 | n8773 ;
  assign n8775 = ( x35 & n8769 ) | ( x35 & ~n8774 ) | ( n8769 & ~n8774 ) ;
  assign n8776 = ( ~x35 & n8774 ) | ( ~x35 & n8775 ) | ( n8774 & n8775 ) ;
  assign n8777 = ( ~n8769 & n8775 ) | ( ~n8769 & n8776 ) | ( n8775 & n8776 ) ;
  assign n8778 = ( n8501 & n8768 ) | ( n8501 & n8777 ) | ( n8768 & n8777 ) ;
  assign n8779 = ( n8501 & ~n8768 ) | ( n8501 & n8777 ) | ( ~n8768 & n8777 ) ;
  assign n8780 = ( n8768 & ~n8778 ) | ( n8768 & n8779 ) | ( ~n8778 & n8779 ) ;
  assign n8781 = n2320 & n2585 ;
  assign n8782 = x96 & n2324 ;
  assign n8783 = x97 | n8782 ;
  assign n8784 = ( n2326 & n8782 ) | ( n2326 & n8783 ) | ( n8782 & n8783 ) ;
  assign n8785 = x95 & n2497 ;
  assign n8786 = n8784 | n8785 ;
  assign n8787 = ( x32 & n8781 ) | ( x32 & ~n8786 ) | ( n8781 & ~n8786 ) ;
  assign n8788 = ( ~x32 & n8786 ) | ( ~x32 & n8787 ) | ( n8786 & n8787 ) ;
  assign n8789 = ( ~n8781 & n8787 ) | ( ~n8781 & n8788 ) | ( n8787 & n8788 ) ;
  assign n8790 = ( n8513 & n8780 ) | ( n8513 & n8789 ) | ( n8780 & n8789 ) ;
  assign n8791 = ( ~n8513 & n8780 ) | ( ~n8513 & n8789 ) | ( n8780 & n8789 ) ;
  assign n8792 = ( n8513 & ~n8790 ) | ( n8513 & n8791 ) | ( ~n8790 & n8791 ) ;
  assign n8793 = ( n8516 & n8656 ) | ( n8516 & n8792 ) | ( n8656 & n8792 ) ;
  assign n8794 = ( ~n8516 & n8656 ) | ( ~n8516 & n8792 ) | ( n8656 & n8792 ) ;
  assign n8795 = ( n8516 & ~n8793 ) | ( n8516 & n8794 ) | ( ~n8793 & n8794 ) ;
  assign n8796 = n1617 & n3650 ;
  assign n8797 = x102 & n1621 ;
  assign n8798 = x103 | n8797 ;
  assign n8799 = ( n1623 & n8797 ) | ( n1623 & n8798 ) | ( n8797 & n8798 ) ;
  assign n8800 = x101 & n1749 ;
  assign n8801 = n8799 | n8800 ;
  assign n8802 = ( x26 & n8796 ) | ( x26 & ~n8801 ) | ( n8796 & ~n8801 ) ;
  assign n8803 = ( ~x26 & n8801 ) | ( ~x26 & n8802 ) | ( n8801 & n8802 ) ;
  assign n8804 = ( ~n8796 & n8802 ) | ( ~n8796 & n8803 ) | ( n8802 & n8803 ) ;
  assign n8805 = ( n8528 & n8795 ) | ( n8528 & n8804 ) | ( n8795 & n8804 ) ;
  assign n8806 = ( ~n8528 & n8795 ) | ( ~n8528 & n8804 ) | ( n8795 & n8804 ) ;
  assign n8807 = ( n8528 & ~n8805 ) | ( n8528 & n8806 ) | ( ~n8805 & n8806 ) ;
  assign n8808 = ( n8540 & n8647 ) | ( n8540 & n8807 ) | ( n8647 & n8807 ) ;
  assign n8809 = ( ~n8540 & n8647 ) | ( ~n8540 & n8807 ) | ( n8647 & n8807 ) ;
  assign n8810 = ( n8540 & ~n8808 ) | ( n8540 & n8809 ) | ( ~n8808 & n8809 ) ;
  assign n8811 = ( n8543 & n8638 ) | ( n8543 & n8810 ) | ( n8638 & n8810 ) ;
  assign n8812 = ( ~n8543 & n8638 ) | ( ~n8543 & n8810 ) | ( n8638 & n8810 ) ;
  assign n8813 = ( n8543 & ~n8811 ) | ( n8543 & n8812 ) | ( ~n8811 & n8812 ) ;
  assign n8814 = ( n8546 & n8629 ) | ( n8546 & n8813 ) | ( n8629 & n8813 ) ;
  assign n8815 = ( ~n8546 & n8629 ) | ( ~n8546 & n8813 ) | ( n8629 & n8813 ) ;
  assign n8816 = ( n8546 & ~n8814 ) | ( n8546 & n8815 ) | ( ~n8814 & n8815 ) ;
  assign n8817 = ( n8558 & n8620 ) | ( n8558 & n8816 ) | ( n8620 & n8816 ) ;
  assign n8818 = ( ~n8558 & n8620 ) | ( ~n8558 & n8816 ) | ( n8620 & n8816 ) ;
  assign n8819 = ( n8558 & ~n8817 ) | ( n8558 & n8818 ) | ( ~n8817 & n8818 ) ;
  assign n8820 = n407 & n6421 ;
  assign n8821 = x117 & n411 ;
  assign n8822 = x118 | n8821 ;
  assign n8823 = ( n413 & n8821 ) | ( n413 & n8822 ) | ( n8821 & n8822 ) ;
  assign n8824 = x116 & n491 ;
  assign n8825 = n8823 | n8824 ;
  assign n8826 = ( x11 & n8820 ) | ( x11 & ~n8825 ) | ( n8820 & ~n8825 ) ;
  assign n8827 = ( ~x11 & n8825 ) | ( ~x11 & n8826 ) | ( n8825 & n8826 ) ;
  assign n8828 = ( ~n8820 & n8826 ) | ( ~n8820 & n8827 ) | ( n8826 & n8827 ) ;
  assign n8829 = ( n8561 & n8819 ) | ( n8561 & n8828 ) | ( n8819 & n8828 ) ;
  assign n8830 = ( ~n8561 & n8819 ) | ( ~n8561 & n8828 ) | ( n8819 & n8828 ) ;
  assign n8831 = ( n8561 & ~n8829 ) | ( n8561 & n8830 ) | ( ~n8829 & n8830 ) ;
  assign n8832 = n291 & n7113 ;
  assign n8833 = x120 & n295 ;
  assign n8834 = x121 | n8833 ;
  assign n8835 = ( n297 & n8833 ) | ( n297 & n8834 ) | ( n8833 & n8834 ) ;
  assign n8836 = x119 & n330 ;
  assign n8837 = n8835 | n8836 ;
  assign n8838 = ( x8 & n8832 ) | ( x8 & ~n8837 ) | ( n8832 & ~n8837 ) ;
  assign n8839 = ( ~x8 & n8837 ) | ( ~x8 & n8838 ) | ( n8837 & n8838 ) ;
  assign n8840 = ( ~n8832 & n8838 ) | ( ~n8832 & n8839 ) | ( n8838 & n8839 ) ;
  assign n8841 = ( n8611 & n8831 ) | ( n8611 & n8840 ) | ( n8831 & n8840 ) ;
  assign n8842 = ( ~n8611 & n8831 ) | ( ~n8611 & n8840 ) | ( n8831 & n8840 ) ;
  assign n8843 = ( n8611 & ~n8841 ) | ( n8611 & n8842 ) | ( ~n8841 & n8842 ) ;
  assign n8844 = ( x126 & x127 ) | ( x126 & n8585 ) | ( x127 & n8585 ) ;
  assign n8845 = ( ~x126 & x127 ) | ( ~x126 & n8585 ) | ( x127 & n8585 ) ;
  assign n8846 = ( x126 & ~n8844 ) | ( x126 & n8845 ) | ( ~n8844 & n8845 ) ;
  assign n8847 = n136 & n8846 ;
  assign n8848 = x125 & n154 ;
  assign n8849 = ( x0 & x126 ) | ( x0 & ~n134 ) | ( x126 & ~n134 ) ;
  assign n8850 = x127 & n141 ;
  assign n8851 = ( n138 & n8849 ) | ( n138 & n8850 ) | ( n8849 & n8850 ) ;
  assign n8852 = n8848 | n8851 ;
  assign n8853 = ( x2 & n8847 ) | ( x2 & ~n8852 ) | ( n8847 & ~n8852 ) ;
  assign n8854 = ( ~x2 & n8852 ) | ( ~x2 & n8853 ) | ( n8852 & n8853 ) ;
  assign n8855 = ( ~n8847 & n8853 ) | ( ~n8847 & n8854 ) | ( n8853 & n8854 ) ;
  assign n8856 = ( n8582 & n8843 ) | ( n8582 & n8855 ) | ( n8843 & n8855 ) ;
  assign n8857 = ( ~n8582 & n8843 ) | ( ~n8582 & n8855 ) | ( n8843 & n8855 ) ;
  assign n8858 = ( n8582 & ~n8856 ) | ( n8582 & n8857 ) | ( ~n8856 & n8857 ) ;
  assign n8859 = ( n8597 & n8600 ) | ( n8597 & n8858 ) | ( n8600 & n8858 ) ;
  assign n8860 = ( n8597 & ~n8600 ) | ( n8597 & n8858 ) | ( ~n8600 & n8858 ) ;
  assign n8861 = ( n8600 & ~n8859 ) | ( n8600 & n8860 ) | ( ~n8859 & n8860 ) ;
  assign n8862 = x126 | n8585 ;
  assign n8863 = x126 & ~x127 ;
  assign n8864 = x127 | n8585 ;
  assign n8865 = ( ~n8862 & n8863 ) | ( ~n8862 & n8864 ) | ( n8863 & n8864 ) ;
  assign n8866 = n136 & n8865 ;
  assign n8867 = x127 & n138 ;
  assign n8868 = ( x126 & ~n8849 ) | ( x126 & n8867 ) | ( ~n8849 & n8867 ) ;
  assign n8869 = ( x2 & n8866 ) | ( x2 & ~n8868 ) | ( n8866 & ~n8868 ) ;
  assign n8870 = ( ~x2 & n8868 ) | ( ~x2 & n8869 ) | ( n8868 & n8869 ) ;
  assign n8871 = ( ~n8866 & n8869 ) | ( ~n8866 & n8870 ) | ( n8869 & n8870 ) ;
  assign n8872 = n186 & n8331 ;
  assign n8873 = x124 & n190 ;
  assign n8874 = x125 | n8873 ;
  assign n8875 = ( n192 & n8873 ) | ( n192 & n8874 ) | ( n8873 & n8874 ) ;
  assign n8876 = x123 & n220 ;
  assign n8877 = n8875 | n8876 ;
  assign n8878 = ( x5 & n8872 ) | ( x5 & ~n8877 ) | ( n8872 & ~n8877 ) ;
  assign n8879 = ( ~x5 & n8877 ) | ( ~x5 & n8878 ) | ( n8877 & n8878 ) ;
  assign n8880 = ( ~n8872 & n8878 ) | ( ~n8872 & n8879 ) | ( n8878 & n8879 ) ;
  assign n8881 = n407 & n6645 ;
  assign n8882 = x118 & n411 ;
  assign n8883 = x119 | n8882 ;
  assign n8884 = ( n413 & n8882 ) | ( n413 & n8883 ) | ( n8882 & n8883 ) ;
  assign n8885 = x117 & n491 ;
  assign n8886 = n8884 | n8885 ;
  assign n8887 = ( x11 & n8881 ) | ( x11 & ~n8886 ) | ( n8881 & ~n8886 ) ;
  assign n8888 = ( ~x11 & n8886 ) | ( ~x11 & n8887 ) | ( n8886 & n8887 ) ;
  assign n8889 = ( ~n8881 & n8887 ) | ( ~n8881 & n8888 ) | ( n8887 & n8888 ) ;
  assign n8890 = n583 & n5977 ;
  assign n8891 = x115 & n587 ;
  assign n8892 = x116 | n8891 ;
  assign n8893 = ( n589 & n8891 ) | ( n589 & n8892 ) | ( n8891 & n8892 ) ;
  assign n8894 = x114 & n676 ;
  assign n8895 = n8893 | n8894 ;
  assign n8896 = ( x14 & n8890 ) | ( x14 & ~n8895 ) | ( n8890 & ~n8895 ) ;
  assign n8897 = ( ~x14 & n8895 ) | ( ~x14 & n8896 ) | ( n8895 & n8896 ) ;
  assign n8898 = ( ~n8890 & n8896 ) | ( ~n8890 & n8897 ) | ( n8896 & n8897 ) ;
  assign n8899 = n810 & n5542 ;
  assign n8900 = x112 & n814 ;
  assign n8901 = x113 | n8900 ;
  assign n8902 = ( n816 & n8900 ) | ( n816 & n8901 ) | ( n8900 & n8901 ) ;
  assign n8903 = x111 & n885 ;
  assign n8904 = n8902 | n8903 ;
  assign n8905 = ( x17 & n8899 ) | ( x17 & ~n8904 ) | ( n8899 & ~n8904 ) ;
  assign n8906 = ( ~x17 & n8904 ) | ( ~x17 & n8905 ) | ( n8904 & n8905 ) ;
  assign n8907 = ( ~n8899 & n8905 ) | ( ~n8899 & n8906 ) | ( n8905 & n8906 ) ;
  assign n8908 = n1016 & n4934 ;
  assign n8909 = x109 & n1020 ;
  assign n8910 = x110 | n8909 ;
  assign n8911 = ( n1022 & n8909 ) | ( n1022 & n8910 ) | ( n8909 & n8910 ) ;
  assign n8912 = x108 & n1145 ;
  assign n8913 = n8911 | n8912 ;
  assign n8914 = ( x20 & n8908 ) | ( x20 & ~n8913 ) | ( n8908 & ~n8913 ) ;
  assign n8915 = ( ~x20 & n8913 ) | ( ~x20 & n8914 ) | ( n8913 & n8914 ) ;
  assign n8916 = ( ~n8908 & n8914 ) | ( ~n8908 & n8915 ) | ( n8914 & n8915 ) ;
  assign n8917 = n1297 & n4362 ;
  assign n8918 = x106 & n1301 ;
  assign n8919 = x107 | n8918 ;
  assign n8920 = ( n1303 & n8918 ) | ( n1303 & n8919 ) | ( n8918 & n8919 ) ;
  assign n8921 = x105 & n1426 ;
  assign n8922 = n8920 | n8921 ;
  assign n8923 = ( x23 & n8917 ) | ( x23 & ~n8922 ) | ( n8917 & ~n8922 ) ;
  assign n8924 = ( ~x23 & n8922 ) | ( ~x23 & n8923 ) | ( n8922 & n8923 ) ;
  assign n8925 = ( ~n8917 & n8923 ) | ( ~n8917 & n8924 ) | ( n8923 & n8924 ) ;
  assign n8926 = ( x62 & x63 ) | ( x62 & x65 ) | ( x63 & x65 ) ;
  assign n8927 = x62 & x63 ;
  assign n8928 = x64 | n8927 ;
  assign n8929 = ( x64 & n8926 ) | ( x64 & ~n8928 ) | ( n8926 & ~n8928 ) ;
  assign n8930 = x67 & n8158 ;
  assign n8931 = x68 | n8930 ;
  assign n8932 = ( n8160 & n8930 ) | ( n8160 & n8931 ) | ( n8930 & n8931 ) ;
  assign n8933 = x66 & n8439 ;
  assign n8934 = n8932 | n8933 ;
  assign n8935 = n201 & n8154 ;
  assign n8936 = ( x62 & n8934 ) | ( x62 & ~n8935 ) | ( n8934 & ~n8935 ) ;
  assign n8937 = ( ~x62 & n8935 ) | ( ~x62 & n8936 ) | ( n8935 & n8936 ) ;
  assign n8938 = ( ~n8934 & n8936 ) | ( ~n8934 & n8937 ) | ( n8936 & n8937 ) ;
  assign n8939 = ( n8697 & n8929 ) | ( n8697 & n8938 ) | ( n8929 & n8938 ) ;
  assign n8940 = ( ~n8697 & n8929 ) | ( ~n8697 & n8938 ) | ( n8929 & n8938 ) ;
  assign n8941 = ( n8697 & ~n8939 ) | ( n8697 & n8940 ) | ( ~n8939 & n8940 ) ;
  assign n8942 = n277 & n7423 ;
  assign n8943 = x70 & n7427 ;
  assign n8944 = x71 | n8943 ;
  assign n8945 = ( n7429 & n8943 ) | ( n7429 & n8944 ) | ( n8943 & n8944 ) ;
  assign n8946 = x69 & n7708 ;
  assign n8947 = n8945 | n8946 ;
  assign n8948 = ( x59 & n8942 ) | ( x59 & ~n8947 ) | ( n8942 & ~n8947 ) ;
  assign n8949 = ( ~x59 & n8947 ) | ( ~x59 & n8948 ) | ( n8947 & n8948 ) ;
  assign n8950 = ( ~n8942 & n8948 ) | ( ~n8942 & n8949 ) | ( n8948 & n8949 ) ;
  assign n8951 = ( n8700 & n8941 ) | ( n8700 & n8950 ) | ( n8941 & n8950 ) ;
  assign n8952 = ( ~n8700 & n8941 ) | ( ~n8700 & n8950 ) | ( n8941 & n8950 ) ;
  assign n8953 = ( n8700 & ~n8951 ) | ( n8700 & n8952 ) | ( ~n8951 & n8952 ) ;
  assign n8954 = n446 & n6713 ;
  assign n8955 = x73 & n6717 ;
  assign n8956 = x74 | n8955 ;
  assign n8957 = ( n6719 & n8955 ) | ( n6719 & n8956 ) | ( n8955 & n8956 ) ;
  assign n8958 = x72 & n6980 ;
  assign n8959 = n8957 | n8958 ;
  assign n8960 = ( x56 & n8954 ) | ( x56 & ~n8959 ) | ( n8954 & ~n8959 ) ;
  assign n8961 = ( ~x56 & n8959 ) | ( ~x56 & n8960 ) | ( n8959 & n8960 ) ;
  assign n8962 = ( ~n8954 & n8960 ) | ( ~n8954 & n8961 ) | ( n8960 & n8961 ) ;
  assign n8963 = ( n8712 & n8953 ) | ( n8712 & n8962 ) | ( n8953 & n8962 ) ;
  assign n8964 = ( ~n8712 & n8953 ) | ( ~n8712 & n8962 ) | ( n8953 & n8962 ) ;
  assign n8965 = ( n8712 & ~n8963 ) | ( n8712 & n8964 ) | ( ~n8963 & n8964 ) ;
  assign n8966 = n569 & n6027 ;
  assign n8967 = x76 & n6031 ;
  assign n8968 = x77 | n8967 ;
  assign n8969 = ( n6033 & n8967 ) | ( n6033 & n8968 ) | ( n8967 & n8968 ) ;
  assign n8970 = x75 & n6303 ;
  assign n8971 = n8969 | n8970 ;
  assign n8972 = ( x53 & n8966 ) | ( x53 & ~n8971 ) | ( n8966 & ~n8971 ) ;
  assign n8973 = ( ~x53 & n8971 ) | ( ~x53 & n8972 ) | ( n8971 & n8972 ) ;
  assign n8974 = ( ~n8966 & n8972 ) | ( ~n8966 & n8973 ) | ( n8972 & n8973 ) ;
  assign n8975 = ( n8715 & n8965 ) | ( n8715 & n8974 ) | ( n8965 & n8974 ) ;
  assign n8976 = ( n8715 & ~n8965 ) | ( n8715 & n8974 ) | ( ~n8965 & n8974 ) ;
  assign n8977 = ( n8965 & ~n8975 ) | ( n8965 & n8976 ) | ( ~n8975 & n8976 ) ;
  assign n8978 = n769 & n5374 ;
  assign n8979 = x79 & n5378 ;
  assign n8980 = x80 | n8979 ;
  assign n8981 = ( n5380 & n8979 ) | ( n5380 & n8980 ) | ( n8979 & n8980 ) ;
  assign n8982 = x78 & n5638 ;
  assign n8983 = n8981 | n8982 ;
  assign n8984 = ( x50 & n8978 ) | ( x50 & ~n8983 ) | ( n8978 & ~n8983 ) ;
  assign n8985 = ( ~x50 & n8983 ) | ( ~x50 & n8984 ) | ( n8983 & n8984 ) ;
  assign n8986 = ( ~n8978 & n8984 ) | ( ~n8978 & n8985 ) | ( n8984 & n8985 ) ;
  assign n8987 = ( n8727 & n8977 ) | ( n8727 & n8986 ) | ( n8977 & n8986 ) ;
  assign n8988 = ( ~n8727 & n8977 ) | ( ~n8727 & n8986 ) | ( n8977 & n8986 ) ;
  assign n8989 = ( n8727 & ~n8987 ) | ( n8727 & n8988 ) | ( ~n8987 & n8988 ) ;
  assign n8990 = n1082 & n4787 ;
  assign n8991 = x82 & n4791 ;
  assign n8992 = x83 | n8991 ;
  assign n8993 = ( n4793 & n8991 ) | ( n4793 & n8992 ) | ( n8991 & n8992 ) ;
  assign n8994 = x81 & n5030 ;
  assign n8995 = n8993 | n8994 ;
  assign n8996 = ( x47 & n8990 ) | ( x47 & ~n8995 ) | ( n8990 & ~n8995 ) ;
  assign n8997 = ( ~x47 & n8995 ) | ( ~x47 & n8996 ) | ( n8995 & n8996 ) ;
  assign n8998 = ( ~n8990 & n8996 ) | ( ~n8990 & n8997 ) | ( n8996 & n8997 ) ;
  assign n8999 = ( n8739 & n8989 ) | ( n8739 & n8998 ) | ( n8989 & n8998 ) ;
  assign n9000 = ( n8739 & ~n8989 ) | ( n8739 & n8998 ) | ( ~n8989 & n8998 ) ;
  assign n9001 = ( n8989 & ~n8999 ) | ( n8989 & n9000 ) | ( ~n8999 & n9000 ) ;
  assign n9002 = n1366 & n4227 ;
  assign n9003 = x85 & n4231 ;
  assign n9004 = x86 | n9003 ;
  assign n9005 = ( n4233 & n9003 ) | ( n4233 & n9004 ) | ( n9003 & n9004 ) ;
  assign n9006 = x84 & n4470 ;
  assign n9007 = n9005 | n9006 ;
  assign n9008 = ( x44 & n9002 ) | ( x44 & ~n9007 ) | ( n9002 & ~n9007 ) ;
  assign n9009 = ( ~x44 & n9007 ) | ( ~x44 & n9008 ) | ( n9007 & n9008 ) ;
  assign n9010 = ( ~n9002 & n9008 ) | ( ~n9002 & n9009 ) | ( n9008 & n9009 ) ;
  assign n9011 = ( n8742 & n9001 ) | ( n8742 & n9010 ) | ( n9001 & n9010 ) ;
  assign n9012 = ( ~n8742 & n9001 ) | ( ~n8742 & n9010 ) | ( n9001 & n9010 ) ;
  assign n9013 = ( n8742 & ~n9011 ) | ( n8742 & n9012 ) | ( ~n9011 & n9012 ) ;
  assign n9014 = n1585 & n3715 ;
  assign n9015 = x88 & n3719 ;
  assign n9016 = x89 | n9015 ;
  assign n9017 = ( n3721 & n9015 ) | ( n3721 & n9016 ) | ( n9015 & n9016 ) ;
  assign n9018 = x87 & n3922 ;
  assign n9019 = n9017 | n9018 ;
  assign n9020 = ( x41 & n9014 ) | ( x41 & ~n9019 ) | ( n9014 & ~n9019 ) ;
  assign n9021 = ( ~x41 & n9019 ) | ( ~x41 & n9020 ) | ( n9019 & n9020 ) ;
  assign n9022 = ( ~n9014 & n9020 ) | ( ~n9014 & n9021 ) | ( n9020 & n9021 ) ;
  assign n9023 = ( n8754 & n9013 ) | ( n8754 & n9022 ) | ( n9013 & n9022 ) ;
  assign n9024 = ( ~n8754 & n9013 ) | ( ~n8754 & n9022 ) | ( n9013 & n9022 ) ;
  assign n9025 = ( n8754 & ~n9023 ) | ( n8754 & n9024 ) | ( ~n9023 & n9024 ) ;
  assign n9026 = n2042 & n3224 ;
  assign n9027 = x91 & n3228 ;
  assign n9028 = x92 | n9027 ;
  assign n9029 = ( n3230 & n9027 ) | ( n3230 & n9028 ) | ( n9027 & n9028 ) ;
  assign n9030 = x90 & n3413 ;
  assign n9031 = n9029 | n9030 ;
  assign n9032 = ( x38 & n9026 ) | ( x38 & ~n9031 ) | ( n9026 & ~n9031 ) ;
  assign n9033 = ( ~x38 & n9031 ) | ( ~x38 & n9032 ) | ( n9031 & n9032 ) ;
  assign n9034 = ( ~n9026 & n9032 ) | ( ~n9026 & n9033 ) | ( n9032 & n9033 ) ;
  assign n9035 = ( n8766 & n9025 ) | ( n8766 & n9034 ) | ( n9025 & n9034 ) ;
  assign n9036 = ( ~n8766 & n9025 ) | ( ~n8766 & n9034 ) | ( n9025 & n9034 ) ;
  assign n9037 = ( n8766 & ~n9035 ) | ( n8766 & n9036 ) | ( ~n9035 & n9036 ) ;
  assign n9038 = n2434 & n2766 ;
  assign n9039 = x94 & n2770 ;
  assign n9040 = x95 | n9039 ;
  assign n9041 = ( n2772 & n9039 ) | ( n2772 & n9040 ) | ( n9039 & n9040 ) ;
  assign n9042 = x93 & n2943 ;
  assign n9043 = n9041 | n9042 ;
  assign n9044 = ( x35 & n9038 ) | ( x35 & ~n9043 ) | ( n9038 & ~n9043 ) ;
  assign n9045 = ( ~x35 & n9043 ) | ( ~x35 & n9044 ) | ( n9043 & n9044 ) ;
  assign n9046 = ( ~n9038 & n9044 ) | ( ~n9038 & n9045 ) | ( n9044 & n9045 ) ;
  assign n9047 = ( n8778 & n9037 ) | ( n8778 & n9046 ) | ( n9037 & n9046 ) ;
  assign n9048 = ( n8778 & ~n9037 ) | ( n8778 & n9046 ) | ( ~n9037 & n9046 ) ;
  assign n9049 = ( n9037 & ~n9047 ) | ( n9037 & n9048 ) | ( ~n9047 & n9048 ) ;
  assign n9050 = n2320 & n2725 ;
  assign n9051 = x97 & n2324 ;
  assign n9052 = x98 | n9051 ;
  assign n9053 = ( n2326 & n9051 ) | ( n2326 & n9052 ) | ( n9051 & n9052 ) ;
  assign n9054 = x96 & n2497 ;
  assign n9055 = n9053 | n9054 ;
  assign n9056 = ( x32 & n9050 ) | ( x32 & ~n9055 ) | ( n9050 & ~n9055 ) ;
  assign n9057 = ( ~x32 & n9055 ) | ( ~x32 & n9056 ) | ( n9055 & n9056 ) ;
  assign n9058 = ( ~n9050 & n9056 ) | ( ~n9050 & n9057 ) | ( n9056 & n9057 ) ;
  assign n9059 = ( n8790 & n9049 ) | ( n8790 & n9058 ) | ( n9049 & n9058 ) ;
  assign n9060 = ( ~n8790 & n9049 ) | ( ~n8790 & n9058 ) | ( n9049 & n9058 ) ;
  assign n9061 = ( n8790 & ~n9059 ) | ( n8790 & n9060 ) | ( ~n9059 & n9060 ) ;
  assign n9062 = n1949 & n3326 ;
  assign n9063 = x100 & n1953 ;
  assign n9064 = x101 | n9063 ;
  assign n9065 = ( n1955 & n9063 ) | ( n1955 & n9064 ) | ( n9063 & n9064 ) ;
  assign n9066 = x99 & n2114 ;
  assign n9067 = n9065 | n9066 ;
  assign n9068 = ( x29 & n9062 ) | ( x29 & ~n9067 ) | ( n9062 & ~n9067 ) ;
  assign n9069 = ( ~x29 & n9067 ) | ( ~x29 & n9068 ) | ( n9067 & n9068 ) ;
  assign n9070 = ( ~n9062 & n9068 ) | ( ~n9062 & n9069 ) | ( n9068 & n9069 ) ;
  assign n9071 = ( n8793 & n9061 ) | ( n8793 & n9070 ) | ( n9061 & n9070 ) ;
  assign n9072 = ( ~n8793 & n9061 ) | ( ~n8793 & n9070 ) | ( n9061 & n9070 ) ;
  assign n9073 = ( n8793 & ~n9071 ) | ( n8793 & n9072 ) | ( ~n9071 & n9072 ) ;
  assign n9074 = n1617 & n3665 ;
  assign n9075 = x103 & n1621 ;
  assign n9076 = x104 | n9075 ;
  assign n9077 = ( n1623 & n9075 ) | ( n1623 & n9076 ) | ( n9075 & n9076 ) ;
  assign n9078 = x102 & n1749 ;
  assign n9079 = n9077 | n9078 ;
  assign n9080 = ( x26 & n9074 ) | ( x26 & ~n9079 ) | ( n9074 & ~n9079 ) ;
  assign n9081 = ( ~x26 & n9079 ) | ( ~x26 & n9080 ) | ( n9079 & n9080 ) ;
  assign n9082 = ( ~n9074 & n9080 ) | ( ~n9074 & n9081 ) | ( n9080 & n9081 ) ;
  assign n9083 = ( n8805 & n9073 ) | ( n8805 & n9082 ) | ( n9073 & n9082 ) ;
  assign n9084 = ( ~n8805 & n9073 ) | ( ~n8805 & n9082 ) | ( n9073 & n9082 ) ;
  assign n9085 = ( n8805 & ~n9083 ) | ( n8805 & n9084 ) | ( ~n9083 & n9084 ) ;
  assign n9086 = ( n8808 & n8925 ) | ( n8808 & n9085 ) | ( n8925 & n9085 ) ;
  assign n9087 = ( ~n8808 & n8925 ) | ( ~n8808 & n9085 ) | ( n8925 & n9085 ) ;
  assign n9088 = ( n8808 & ~n9086 ) | ( n8808 & n9087 ) | ( ~n9086 & n9087 ) ;
  assign n9089 = ( n8811 & n8916 ) | ( n8811 & n9088 ) | ( n8916 & n9088 ) ;
  assign n9090 = ( ~n8811 & n8916 ) | ( ~n8811 & n9088 ) | ( n8916 & n9088 ) ;
  assign n9091 = ( n8811 & ~n9089 ) | ( n8811 & n9090 ) | ( ~n9089 & n9090 ) ;
  assign n9092 = ( n8814 & n8907 ) | ( n8814 & n9091 ) | ( n8907 & n9091 ) ;
  assign n9093 = ( ~n8814 & n8907 ) | ( ~n8814 & n9091 ) | ( n8907 & n9091 ) ;
  assign n9094 = ( n8814 & ~n9092 ) | ( n8814 & n9093 ) | ( ~n9092 & n9093 ) ;
  assign n9095 = ( n8817 & n8898 ) | ( n8817 & n9094 ) | ( n8898 & n9094 ) ;
  assign n9096 = ( ~n8817 & n8898 ) | ( ~n8817 & n9094 ) | ( n8898 & n9094 ) ;
  assign n9097 = ( n8817 & ~n9095 ) | ( n8817 & n9096 ) | ( ~n9095 & n9096 ) ;
  assign n9098 = ( n8829 & n8889 ) | ( n8829 & n9097 ) | ( n8889 & n9097 ) ;
  assign n9099 = ( ~n8829 & n8889 ) | ( ~n8829 & n9097 ) | ( n8889 & n9097 ) ;
  assign n9100 = ( n8829 & ~n9098 ) | ( n8829 & n9099 ) | ( ~n9098 & n9099 ) ;
  assign n9101 = n291 & n7582 ;
  assign n9102 = x121 & n295 ;
  assign n9103 = x122 | n9102 ;
  assign n9104 = ( n297 & n9102 ) | ( n297 & n9103 ) | ( n9102 & n9103 ) ;
  assign n9105 = x120 & n330 ;
  assign n9106 = n9104 | n9105 ;
  assign n9107 = ( x8 & n9101 ) | ( x8 & ~n9106 ) | ( n9101 & ~n9106 ) ;
  assign n9108 = ( ~x8 & n9106 ) | ( ~x8 & n9107 ) | ( n9106 & n9107 ) ;
  assign n9109 = ( ~n9101 & n9107 ) | ( ~n9101 & n9108 ) | ( n9107 & n9108 ) ;
  assign n9110 = ( n8880 & n9100 ) | ( n8880 & n9109 ) | ( n9100 & n9109 ) ;
  assign n9111 = ( ~n8880 & n9100 ) | ( ~n8880 & n9109 ) | ( n9100 & n9109 ) ;
  assign n9112 = ( n8880 & ~n9110 ) | ( n8880 & n9111 ) | ( ~n9110 & n9111 ) ;
  assign n9113 = ( n8841 & n8871 ) | ( n8841 & n9112 ) | ( n8871 & n9112 ) ;
  assign n9114 = ( n8841 & ~n8871 ) | ( n8841 & n9112 ) | ( ~n8871 & n9112 ) ;
  assign n9115 = ( n8871 & ~n9113 ) | ( n8871 & n9114 ) | ( ~n9113 & n9114 ) ;
  assign n9116 = ( n8856 & n8859 ) | ( n8856 & n9115 ) | ( n8859 & n9115 ) ;
  assign n9117 = ( n8856 & ~n8859 ) | ( n8856 & n9115 ) | ( ~n8859 & n9115 ) ;
  assign n9118 = ( n8859 & ~n9116 ) | ( n8859 & n9117 ) | ( ~n9116 & n9117 ) ;
  assign n9119 = x127 & n136 ;
  assign n9120 = n8862 & n9119 ;
  assign n9121 = x2 | n9120 ;
  assign n9122 = x127 & n154 ;
  assign n9123 = ( x2 & n9120 ) | ( x2 & n9122 ) | ( n9120 & n9122 ) ;
  assign n9124 = n9121 & ~n9123 ;
  assign n9125 = n810 & n5750 ;
  assign n9126 = x113 & n814 ;
  assign n9127 = x114 | n9126 ;
  assign n9128 = ( n816 & n9126 ) | ( n816 & n9127 ) | ( n9126 & n9127 ) ;
  assign n9129 = x112 & n885 ;
  assign n9130 = n9128 | n9129 ;
  assign n9131 = ( x17 & n9125 ) | ( x17 & ~n9130 ) | ( n9125 & ~n9130 ) ;
  assign n9132 = ( ~x17 & n9130 ) | ( ~x17 & n9131 ) | ( n9130 & n9131 ) ;
  assign n9133 = ( ~n9125 & n9131 ) | ( ~n9125 & n9132 ) | ( n9131 & n9132 ) ;
  assign n9134 = n1016 & n5130 ;
  assign n9135 = x110 & n1020 ;
  assign n9136 = x111 | n9135 ;
  assign n9137 = ( n1022 & n9135 ) | ( n1022 & n9136 ) | ( n9135 & n9136 ) ;
  assign n9138 = x109 & n1145 ;
  assign n9139 = n9137 | n9138 ;
  assign n9140 = ( x20 & n9134 ) | ( x20 & ~n9139 ) | ( n9134 & ~n9139 ) ;
  assign n9141 = ( ~x20 & n9139 ) | ( ~x20 & n9140 ) | ( n9139 & n9140 ) ;
  assign n9142 = ( ~n9134 & n9140 ) | ( ~n9134 & n9141 ) | ( n9140 & n9141 ) ;
  assign n9143 = n1297 & n4377 ;
  assign n9144 = x107 & n1301 ;
  assign n9145 = x108 | n9144 ;
  assign n9146 = ( n1303 & n9144 ) | ( n1303 & n9145 ) | ( n9144 & n9145 ) ;
  assign n9147 = x106 & n1426 ;
  assign n9148 = n9146 | n9147 ;
  assign n9149 = ( x23 & n9143 ) | ( x23 & ~n9148 ) | ( n9143 & ~n9148 ) ;
  assign n9150 = ( ~x23 & n9148 ) | ( ~x23 & n9149 ) | ( n9148 & n9149 ) ;
  assign n9151 = ( ~n9143 & n9149 ) | ( ~n9143 & n9150 ) | ( n9149 & n9150 ) ;
  assign n9152 = n2320 & n2877 ;
  assign n9153 = x98 & n2324 ;
  assign n9154 = x99 | n9153 ;
  assign n9155 = ( n2326 & n9153 ) | ( n2326 & n9154 ) | ( n9153 & n9154 ) ;
  assign n9156 = x97 & n2497 ;
  assign n9157 = n9155 | n9156 ;
  assign n9158 = ( x32 & n9152 ) | ( x32 & ~n9157 ) | ( n9152 & ~n9157 ) ;
  assign n9159 = ( ~x32 & n9157 ) | ( ~x32 & n9158 ) | ( n9157 & n9158 ) ;
  assign n9160 = ( ~n9152 & n9158 ) | ( ~n9152 & n9159 ) | ( n9158 & n9159 ) ;
  assign n9161 = n1466 & n4227 ;
  assign n9162 = x86 & n4231 ;
  assign n9163 = x87 | n9162 ;
  assign n9164 = ( n4233 & n9162 ) | ( n4233 & n9163 ) | ( n9162 & n9163 ) ;
  assign n9165 = x85 & n4470 ;
  assign n9166 = n9164 | n9165 ;
  assign n9167 = ( x44 & n9161 ) | ( x44 & ~n9166 ) | ( n9161 & ~n9166 ) ;
  assign n9168 = ( ~x44 & n9166 ) | ( ~x44 & n9167 ) | ( n9166 & n9167 ) ;
  assign n9169 = ( ~n9161 & n9167 ) | ( ~n9161 & n9168 ) | ( n9167 & n9168 ) ;
  assign n9170 = n910 & n5374 ;
  assign n9171 = x80 & n5378 ;
  assign n9172 = x81 | n9171 ;
  assign n9173 = ( n5380 & n9171 ) | ( n5380 & n9172 ) | ( n9171 & n9172 ) ;
  assign n9174 = x79 & n5638 ;
  assign n9175 = n9173 | n9174 ;
  assign n9176 = ( x50 & n9170 ) | ( x50 & ~n9175 ) | ( n9170 & ~n9175 ) ;
  assign n9177 = ( ~x50 & n9175 ) | ( ~x50 & n9176 ) | ( n9175 & n9176 ) ;
  assign n9178 = ( ~n9170 & n9176 ) | ( ~n9170 & n9177 ) | ( n9176 & n9177 ) ;
  assign n9179 = n461 & n6713 ;
  assign n9180 = x74 & n6717 ;
  assign n9181 = x75 | n9180 ;
  assign n9182 = ( n6719 & n9180 ) | ( n6719 & n9181 ) | ( n9180 & n9181 ) ;
  assign n9183 = x73 & n6980 ;
  assign n9184 = n9182 | n9183 ;
  assign n9185 = ( x56 & n9179 ) | ( x56 & ~n9184 ) | ( n9179 & ~n9184 ) ;
  assign n9186 = ( ~x56 & n9184 ) | ( ~x56 & n9185 ) | ( n9184 & n9185 ) ;
  assign n9187 = ( ~n9179 & n9185 ) | ( ~n9179 & n9186 ) | ( n9185 & n9186 ) ;
  assign n9188 = x65 & n8927 ;
  assign n9189 = ( ~x66 & n8693 ) | ( ~x66 & n8927 ) | ( n8693 & n8927 ) ;
  assign n9190 = ( n8693 & n9188 ) | ( n8693 & ~n9189 ) | ( n9188 & ~n9189 ) ;
  assign n9191 = n230 & n8154 ;
  assign n9192 = x68 & n8158 ;
  assign n9193 = x69 | n9192 ;
  assign n9194 = ( n8160 & n9192 ) | ( n8160 & n9193 ) | ( n9192 & n9193 ) ;
  assign n9195 = x67 & n8439 ;
  assign n9196 = n9194 | n9195 ;
  assign n9197 = ( ~x62 & n9191 ) | ( ~x62 & n9196 ) | ( n9191 & n9196 ) ;
  assign n9198 = ( n9191 & n9196 ) | ( n9191 & ~n9197 ) | ( n9196 & ~n9197 ) ;
  assign n9199 = ( x62 & n9197 ) | ( x62 & ~n9198 ) | ( n9197 & ~n9198 ) ;
  assign n9200 = ( n8939 & n9190 ) | ( n8939 & n9199 ) | ( n9190 & n9199 ) ;
  assign n9201 = ( ~n8939 & n9190 ) | ( ~n8939 & n9199 ) | ( n9190 & n9199 ) ;
  assign n9202 = ( n8939 & ~n9200 ) | ( n8939 & n9201 ) | ( ~n9200 & n9201 ) ;
  assign n9203 = n346 & n7423 ;
  assign n9204 = x71 & n7427 ;
  assign n9205 = x72 | n9204 ;
  assign n9206 = ( n7429 & n9204 ) | ( n7429 & n9205 ) | ( n9204 & n9205 ) ;
  assign n9207 = x70 & n7708 ;
  assign n9208 = n9206 | n9207 ;
  assign n9209 = ( x59 & n9203 ) | ( x59 & ~n9208 ) | ( n9203 & ~n9208 ) ;
  assign n9210 = ( ~x59 & n9208 ) | ( ~x59 & n9209 ) | ( n9208 & n9209 ) ;
  assign n9211 = ( ~n9203 & n9209 ) | ( ~n9203 & n9210 ) | ( n9209 & n9210 ) ;
  assign n9212 = ( n8951 & n9202 ) | ( n8951 & n9211 ) | ( n9202 & n9211 ) ;
  assign n9213 = ( ~n8951 & n9202 ) | ( ~n8951 & n9211 ) | ( n9202 & n9211 ) ;
  assign n9214 = ( n8951 & ~n9212 ) | ( n8951 & n9213 ) | ( ~n9212 & n9213 ) ;
  assign n9215 = ( n8963 & n9187 ) | ( n8963 & n9214 ) | ( n9187 & n9214 ) ;
  assign n9216 = ( ~n8963 & n9187 ) | ( ~n8963 & n9214 ) | ( n9187 & n9214 ) ;
  assign n9217 = ( n8963 & ~n9215 ) | ( n8963 & n9216 ) | ( ~n9215 & n9216 ) ;
  assign n9218 = n637 & n6027 ;
  assign n9219 = x77 & n6031 ;
  assign n9220 = x78 | n9219 ;
  assign n9221 = ( n6033 & n9219 ) | ( n6033 & n9220 ) | ( n9219 & n9220 ) ;
  assign n9222 = x76 & n6303 ;
  assign n9223 = n9221 | n9222 ;
  assign n9224 = ( x53 & n9218 ) | ( x53 & ~n9223 ) | ( n9218 & ~n9223 ) ;
  assign n9225 = ( ~x53 & n9223 ) | ( ~x53 & n9224 ) | ( n9223 & n9224 ) ;
  assign n9226 = ( ~n9218 & n9224 ) | ( ~n9218 & n9225 ) | ( n9224 & n9225 ) ;
  assign n9227 = ( n8975 & n9217 ) | ( n8975 & n9226 ) | ( n9217 & n9226 ) ;
  assign n9228 = ( ~n8975 & n9217 ) | ( ~n8975 & n9226 ) | ( n9217 & n9226 ) ;
  assign n9229 = ( n8975 & ~n9227 ) | ( n8975 & n9228 ) | ( ~n9227 & n9228 ) ;
  assign n9230 = ( n8987 & n9178 ) | ( n8987 & n9229 ) | ( n9178 & n9229 ) ;
  assign n9231 = ( ~n8987 & n9178 ) | ( ~n8987 & n9229 ) | ( n9178 & n9229 ) ;
  assign n9232 = ( n8987 & ~n9230 ) | ( n8987 & n9231 ) | ( ~n9230 & n9231 ) ;
  assign n9233 = n1097 & n4787 ;
  assign n9234 = x83 & n4791 ;
  assign n9235 = x84 | n9234 ;
  assign n9236 = ( n4793 & n9234 ) | ( n4793 & n9235 ) | ( n9234 & n9235 ) ;
  assign n9237 = x82 & n5030 ;
  assign n9238 = n9236 | n9237 ;
  assign n9239 = ( x47 & n9233 ) | ( x47 & ~n9238 ) | ( n9233 & ~n9238 ) ;
  assign n9240 = ( ~x47 & n9238 ) | ( ~x47 & n9239 ) | ( n9238 & n9239 ) ;
  assign n9241 = ( ~n9233 & n9239 ) | ( ~n9233 & n9240 ) | ( n9239 & n9240 ) ;
  assign n9242 = ( n8999 & n9232 ) | ( n8999 & n9241 ) | ( n9232 & n9241 ) ;
  assign n9243 = ( ~n8999 & n9232 ) | ( ~n8999 & n9241 ) | ( n9232 & n9241 ) ;
  assign n9244 = ( n8999 & ~n9242 ) | ( n8999 & n9243 ) | ( ~n9242 & n9243 ) ;
  assign n9245 = ( n9011 & n9169 ) | ( n9011 & n9244 ) | ( n9169 & n9244 ) ;
  assign n9246 = ( ~n9011 & n9169 ) | ( ~n9011 & n9244 ) | ( n9169 & n9244 ) ;
  assign n9247 = ( n9011 & ~n9245 ) | ( n9011 & n9246 ) | ( ~n9245 & n9246 ) ;
  assign n9248 = n1701 & n3715 ;
  assign n9249 = x89 & n3719 ;
  assign n9250 = x90 | n9249 ;
  assign n9251 = ( n3721 & n9249 ) | ( n3721 & n9250 ) | ( n9249 & n9250 ) ;
  assign n9252 = x88 & n3922 ;
  assign n9253 = n9251 | n9252 ;
  assign n9254 = ( x41 & n9248 ) | ( x41 & ~n9253 ) | ( n9248 & ~n9253 ) ;
  assign n9255 = ( ~x41 & n9253 ) | ( ~x41 & n9254 ) | ( n9253 & n9254 ) ;
  assign n9256 = ( ~n9248 & n9254 ) | ( ~n9248 & n9255 ) | ( n9254 & n9255 ) ;
  assign n9257 = ( n9023 & n9247 ) | ( n9023 & n9256 ) | ( n9247 & n9256 ) ;
  assign n9258 = ( ~n9023 & n9247 ) | ( ~n9023 & n9256 ) | ( n9247 & n9256 ) ;
  assign n9259 = ( n9023 & ~n9257 ) | ( n9023 & n9258 ) | ( ~n9257 & n9258 ) ;
  assign n9260 = n2057 & n3224 ;
  assign n9261 = x92 & n3228 ;
  assign n9262 = x93 | n9261 ;
  assign n9263 = ( n3230 & n9261 ) | ( n3230 & n9262 ) | ( n9261 & n9262 ) ;
  assign n9264 = x91 & n3413 ;
  assign n9265 = n9263 | n9264 ;
  assign n9266 = ( x38 & n9260 ) | ( x38 & ~n9265 ) | ( n9260 & ~n9265 ) ;
  assign n9267 = ( ~x38 & n9265 ) | ( ~x38 & n9266 ) | ( n9265 & n9266 ) ;
  assign n9268 = ( ~n9260 & n9266 ) | ( ~n9260 & n9267 ) | ( n9266 & n9267 ) ;
  assign n9269 = ( n9035 & n9259 ) | ( n9035 & n9268 ) | ( n9259 & n9268 ) ;
  assign n9270 = ( ~n9035 & n9259 ) | ( ~n9035 & n9268 ) | ( n9259 & n9268 ) ;
  assign n9271 = ( n9035 & ~n9269 ) | ( n9035 & n9270 ) | ( ~n9269 & n9270 ) ;
  assign n9272 = n2449 & n2766 ;
  assign n9273 = x95 & n2770 ;
  assign n9274 = x96 | n9273 ;
  assign n9275 = ( n2772 & n9273 ) | ( n2772 & n9274 ) | ( n9273 & n9274 ) ;
  assign n9276 = x94 & n2943 ;
  assign n9277 = n9275 | n9276 ;
  assign n9278 = ( x35 & n9272 ) | ( x35 & ~n9277 ) | ( n9272 & ~n9277 ) ;
  assign n9279 = ( ~x35 & n9277 ) | ( ~x35 & n9278 ) | ( n9277 & n9278 ) ;
  assign n9280 = ( ~n9272 & n9278 ) | ( ~n9272 & n9279 ) | ( n9278 & n9279 ) ;
  assign n9281 = ( n9047 & n9271 ) | ( n9047 & n9280 ) | ( n9271 & n9280 ) ;
  assign n9282 = ( ~n9047 & n9271 ) | ( ~n9047 & n9280 ) | ( n9271 & n9280 ) ;
  assign n9283 = ( n9047 & ~n9281 ) | ( n9047 & n9282 ) | ( ~n9281 & n9282 ) ;
  assign n9284 = ( n9059 & n9160 ) | ( n9059 & n9283 ) | ( n9160 & n9283 ) ;
  assign n9285 = ( ~n9059 & n9160 ) | ( ~n9059 & n9283 ) | ( n9160 & n9283 ) ;
  assign n9286 = ( n9059 & ~n9284 ) | ( n9059 & n9285 ) | ( ~n9284 & n9285 ) ;
  assign n9287 = n1949 & n3486 ;
  assign n9288 = x101 & n1953 ;
  assign n9289 = x102 | n9288 ;
  assign n9290 = ( n1955 & n9288 ) | ( n1955 & n9289 ) | ( n9288 & n9289 ) ;
  assign n9291 = x100 & n2114 ;
  assign n9292 = n9290 | n9291 ;
  assign n9293 = ( x29 & n9287 ) | ( x29 & ~n9292 ) | ( n9287 & ~n9292 ) ;
  assign n9294 = ( ~x29 & n9292 ) | ( ~x29 & n9293 ) | ( n9292 & n9293 ) ;
  assign n9295 = ( ~n9287 & n9293 ) | ( ~n9287 & n9294 ) | ( n9293 & n9294 ) ;
  assign n9296 = ( n9071 & n9286 ) | ( n9071 & n9295 ) | ( n9286 & n9295 ) ;
  assign n9297 = ( ~n9071 & n9286 ) | ( ~n9071 & n9295 ) | ( n9286 & n9295 ) ;
  assign n9298 = ( n9071 & ~n9296 ) | ( n9071 & n9297 ) | ( ~n9296 & n9297 ) ;
  assign n9299 = n1617 & n3998 ;
  assign n9300 = x104 & n1621 ;
  assign n9301 = x105 | n9300 ;
  assign n9302 = ( n1623 & n9300 ) | ( n1623 & n9301 ) | ( n9300 & n9301 ) ;
  assign n9303 = x103 & n1749 ;
  assign n9304 = n9302 | n9303 ;
  assign n9305 = ( x26 & n9299 ) | ( x26 & ~n9304 ) | ( n9299 & ~n9304 ) ;
  assign n9306 = ( ~x26 & n9304 ) | ( ~x26 & n9305 ) | ( n9304 & n9305 ) ;
  assign n9307 = ( ~n9299 & n9305 ) | ( ~n9299 & n9306 ) | ( n9305 & n9306 ) ;
  assign n9308 = ( n9083 & n9298 ) | ( n9083 & n9307 ) | ( n9298 & n9307 ) ;
  assign n9309 = ( ~n9083 & n9298 ) | ( ~n9083 & n9307 ) | ( n9298 & n9307 ) ;
  assign n9310 = ( n9083 & ~n9308 ) | ( n9083 & n9309 ) | ( ~n9308 & n9309 ) ;
  assign n9311 = ( n9086 & n9151 ) | ( n9086 & n9310 ) | ( n9151 & n9310 ) ;
  assign n9312 = ( ~n9086 & n9151 ) | ( ~n9086 & n9310 ) | ( n9151 & n9310 ) ;
  assign n9313 = ( n9086 & ~n9311 ) | ( n9086 & n9312 ) | ( ~n9311 & n9312 ) ;
  assign n9314 = ( n9089 & n9142 ) | ( n9089 & n9313 ) | ( n9142 & n9313 ) ;
  assign n9315 = ( ~n9089 & n9142 ) | ( ~n9089 & n9313 ) | ( n9142 & n9313 ) ;
  assign n9316 = ( n9089 & ~n9314 ) | ( n9089 & n9315 ) | ( ~n9314 & n9315 ) ;
  assign n9317 = ( n9092 & n9133 ) | ( n9092 & n9316 ) | ( n9133 & n9316 ) ;
  assign n9318 = ( ~n9092 & n9133 ) | ( ~n9092 & n9316 ) | ( n9133 & n9316 ) ;
  assign n9319 = ( n9092 & ~n9317 ) | ( n9092 & n9318 ) | ( ~n9317 & n9318 ) ;
  assign n9320 = n583 & n6201 ;
  assign n9321 = x116 & n587 ;
  assign n9322 = x117 | n9321 ;
  assign n9323 = ( n589 & n9321 ) | ( n589 & n9322 ) | ( n9321 & n9322 ) ;
  assign n9324 = x115 & n676 ;
  assign n9325 = n9323 | n9324 ;
  assign n9326 = ( x14 & n9320 ) | ( x14 & ~n9325 ) | ( n9320 & ~n9325 ) ;
  assign n9327 = ( ~x14 & n9325 ) | ( ~x14 & n9326 ) | ( n9325 & n9326 ) ;
  assign n9328 = ( ~n9320 & n9326 ) | ( ~n9320 & n9327 ) | ( n9326 & n9327 ) ;
  assign n9329 = ( n9095 & n9319 ) | ( n9095 & n9328 ) | ( n9319 & n9328 ) ;
  assign n9330 = ( ~n9095 & n9319 ) | ( ~n9095 & n9328 ) | ( n9319 & n9328 ) ;
  assign n9331 = ( n9095 & ~n9329 ) | ( n9095 & n9330 ) | ( ~n9329 & n9330 ) ;
  assign n9332 = n407 & n7098 ;
  assign n9333 = x119 & n411 ;
  assign n9334 = x120 | n9333 ;
  assign n9335 = ( n413 & n9333 ) | ( n413 & n9334 ) | ( n9333 & n9334 ) ;
  assign n9336 = x118 & n491 ;
  assign n9337 = n9335 | n9336 ;
  assign n9338 = ( x11 & n9332 ) | ( x11 & ~n9337 ) | ( n9332 & ~n9337 ) ;
  assign n9339 = ( ~x11 & n9337 ) | ( ~x11 & n9338 ) | ( n9337 & n9338 ) ;
  assign n9340 = ( ~n9332 & n9338 ) | ( ~n9332 & n9339 ) | ( n9338 & n9339 ) ;
  assign n9341 = n291 & n7597 ;
  assign n9342 = x122 & n295 ;
  assign n9343 = x123 | n9342 ;
  assign n9344 = ( n297 & n9342 ) | ( n297 & n9343 ) | ( n9342 & n9343 ) ;
  assign n9345 = x121 & n330 ;
  assign n9346 = n9344 | n9345 ;
  assign n9347 = ( x8 & n9341 ) | ( x8 & ~n9346 ) | ( n9341 & ~n9346 ) ;
  assign n9348 = ( ~x8 & n9346 ) | ( ~x8 & n9347 ) | ( n9346 & n9347 ) ;
  assign n9349 = ( ~n9341 & n9347 ) | ( ~n9341 & n9348 ) | ( n9347 & n9348 ) ;
  assign n9350 = ( n9331 & n9340 ) | ( n9331 & n9349 ) | ( n9340 & n9349 ) ;
  assign n9351 = ( ~n9331 & n9340 ) | ( ~n9331 & n9349 ) | ( n9340 & n9349 ) ;
  assign n9352 = ( n9331 & ~n9350 ) | ( n9331 & n9351 ) | ( ~n9350 & n9351 ) ;
  assign n9353 = n186 & n8587 ;
  assign n9354 = x125 & n190 ;
  assign n9355 = x126 | n9354 ;
  assign n9356 = ( n192 & n9354 ) | ( n192 & n9355 ) | ( n9354 & n9355 ) ;
  assign n9357 = x124 & n220 ;
  assign n9358 = n9356 | n9357 ;
  assign n9359 = ( x5 & n9353 ) | ( x5 & ~n9358 ) | ( n9353 & ~n9358 ) ;
  assign n9360 = ( ~x5 & n9358 ) | ( ~x5 & n9359 ) | ( n9358 & n9359 ) ;
  assign n9361 = ( ~n9353 & n9359 ) | ( ~n9353 & n9360 ) | ( n9359 & n9360 ) ;
  assign n9362 = ( n9098 & n9352 ) | ( n9098 & n9361 ) | ( n9352 & n9361 ) ;
  assign n9363 = ( ~n9098 & n9352 ) | ( ~n9098 & n9361 ) | ( n9352 & n9361 ) ;
  assign n9364 = ( n9098 & ~n9362 ) | ( n9098 & n9363 ) | ( ~n9362 & n9363 ) ;
  assign n9365 = ( n9110 & n9124 ) | ( n9110 & n9364 ) | ( n9124 & n9364 ) ;
  assign n9366 = ( ~n9110 & n9124 ) | ( ~n9110 & n9364 ) | ( n9124 & n9364 ) ;
  assign n9367 = ( n9110 & ~n9365 ) | ( n9110 & n9366 ) | ( ~n9365 & n9366 ) ;
  assign n9368 = ( n9113 & n9116 ) | ( n9113 & n9367 ) | ( n9116 & n9367 ) ;
  assign n9369 = ( ~n9113 & n9116 ) | ( ~n9113 & n9367 ) | ( n9116 & n9367 ) ;
  assign n9370 = ( n9113 & ~n9368 ) | ( n9113 & n9369 ) | ( ~n9368 & n9369 ) ;
  assign n9371 = n407 & n7113 ;
  assign n9372 = x120 & n411 ;
  assign n9373 = x121 | n9372 ;
  assign n9374 = ( n413 & n9372 ) | ( n413 & n9373 ) | ( n9372 & n9373 ) ;
  assign n9375 = x119 & n491 ;
  assign n9376 = n9374 | n9375 ;
  assign n9377 = ( x11 & n9371 ) | ( x11 & ~n9376 ) | ( n9371 & ~n9376 ) ;
  assign n9378 = ( ~x11 & n9376 ) | ( ~x11 & n9377 ) | ( n9376 & n9377 ) ;
  assign n9379 = ( ~n9371 & n9377 ) | ( ~n9371 & n9378 ) | ( n9377 & n9378 ) ;
  assign n9380 = n810 & n5765 ;
  assign n9381 = x114 & n814 ;
  assign n9382 = x115 | n9381 ;
  assign n9383 = ( n816 & n9381 ) | ( n816 & n9382 ) | ( n9381 & n9382 ) ;
  assign n9384 = x113 & n885 ;
  assign n9385 = n9383 | n9384 ;
  assign n9386 = ( x17 & n9380 ) | ( x17 & ~n9385 ) | ( n9380 & ~n9385 ) ;
  assign n9387 = ( ~x17 & n9385 ) | ( ~x17 & n9386 ) | ( n9385 & n9386 ) ;
  assign n9388 = ( ~n9380 & n9386 ) | ( ~n9380 & n9387 ) | ( n9386 & n9387 ) ;
  assign n9389 = n1016 & n5145 ;
  assign n9390 = x111 & n1020 ;
  assign n9391 = x112 | n9390 ;
  assign n9392 = ( n1022 & n9390 ) | ( n1022 & n9391 ) | ( n9390 & n9391 ) ;
  assign n9393 = x110 & n1145 ;
  assign n9394 = n9392 | n9393 ;
  assign n9395 = ( x20 & n9389 ) | ( x20 & ~n9394 ) | ( n9389 & ~n9394 ) ;
  assign n9396 = ( ~x20 & n9394 ) | ( ~x20 & n9395 ) | ( n9394 & n9395 ) ;
  assign n9397 = ( ~n9389 & n9395 ) | ( ~n9389 & n9396 ) | ( n9395 & n9396 ) ;
  assign n9398 = n1617 & n4013 ;
  assign n9399 = x105 & n1621 ;
  assign n9400 = x106 | n9399 ;
  assign n9401 = ( n1623 & n9399 ) | ( n1623 & n9400 ) | ( n9399 & n9400 ) ;
  assign n9402 = x104 & n1749 ;
  assign n9403 = n9401 | n9402 ;
  assign n9404 = ( x26 & n9398 ) | ( x26 & ~n9403 ) | ( n9398 & ~n9403 ) ;
  assign n9405 = ( ~x26 & n9403 ) | ( ~x26 & n9404 ) | ( n9403 & n9404 ) ;
  assign n9406 = ( ~n9398 & n9404 ) | ( ~n9398 & n9405 ) | ( n9404 & n9405 ) ;
  assign n9407 = n1949 & n3650 ;
  assign n9408 = x102 & n1953 ;
  assign n9409 = x103 | n9408 ;
  assign n9410 = ( n1955 & n9408 ) | ( n1955 & n9409 ) | ( n9408 & n9409 ) ;
  assign n9411 = x101 & n2114 ;
  assign n9412 = n9410 | n9411 ;
  assign n9413 = ( x29 & n9407 ) | ( x29 & ~n9412 ) | ( n9407 & ~n9412 ) ;
  assign n9414 = ( ~x29 & n9412 ) | ( ~x29 & n9413 ) | ( n9412 & n9413 ) ;
  assign n9415 = ( ~n9407 & n9413 ) | ( ~n9407 & n9414 ) | ( n9413 & n9414 ) ;
  assign n9416 = n554 & n6713 ;
  assign n9417 = x75 & n6717 ;
  assign n9418 = x76 | n9417 ;
  assign n9419 = ( n6719 & n9417 ) | ( n6719 & n9418 ) | ( n9417 & n9418 ) ;
  assign n9420 = x74 & n6980 ;
  assign n9421 = n9419 | n9420 ;
  assign n9422 = ( x56 & n9416 ) | ( x56 & ~n9421 ) | ( n9416 & ~n9421 ) ;
  assign n9423 = ( ~x56 & n9421 ) | ( ~x56 & n9422 ) | ( n9421 & n9422 ) ;
  assign n9424 = ( ~n9416 & n9422 ) | ( ~n9416 & n9423 ) | ( n9422 & n9423 ) ;
  assign n9425 = x66 & n8927 ;
  assign n9426 = ( ~x67 & n8693 ) | ( ~x67 & n8927 ) | ( n8693 & n8927 ) ;
  assign n9427 = ( n8693 & n9425 ) | ( n8693 & ~n9426 ) | ( n9425 & ~n9426 ) ;
  assign n9428 = n245 & n8154 ;
  assign n9429 = x69 & n8158 ;
  assign n9430 = x70 | n9429 ;
  assign n9431 = ( n8160 & n9429 ) | ( n8160 & n9430 ) | ( n9429 & n9430 ) ;
  assign n9432 = x68 & n8439 ;
  assign n9433 = n9431 | n9432 ;
  assign n9434 = ( x62 & n9428 ) | ( x62 & ~n9433 ) | ( n9428 & ~n9433 ) ;
  assign n9435 = ( ~x62 & n9433 ) | ( ~x62 & n9434 ) | ( n9433 & n9434 ) ;
  assign n9436 = ( ~n9428 & n9434 ) | ( ~n9428 & n9435 ) | ( n9434 & n9435 ) ;
  assign n9437 = ( x2 & n9427 ) | ( x2 & n9436 ) | ( n9427 & n9436 ) ;
  assign n9438 = ( ~x2 & n9427 ) | ( ~x2 & n9436 ) | ( n9427 & n9436 ) ;
  assign n9439 = ( x2 & ~n9437 ) | ( x2 & n9438 ) | ( ~n9437 & n9438 ) ;
  assign n9440 = n390 & n7423 ;
  assign n9441 = x72 & n7427 ;
  assign n9442 = x73 | n9441 ;
  assign n9443 = ( n7429 & n9441 ) | ( n7429 & n9442 ) | ( n9441 & n9442 ) ;
  assign n9444 = x71 & n7708 ;
  assign n9445 = n9443 | n9444 ;
  assign n9446 = ( x59 & n9440 ) | ( x59 & ~n9445 ) | ( n9440 & ~n9445 ) ;
  assign n9447 = ( ~x59 & n9445 ) | ( ~x59 & n9446 ) | ( n9445 & n9446 ) ;
  assign n9448 = ( ~n9440 & n9446 ) | ( ~n9440 & n9447 ) | ( n9446 & n9447 ) ;
  assign n9449 = ( n9200 & n9439 ) | ( n9200 & n9448 ) | ( n9439 & n9448 ) ;
  assign n9450 = ( ~n9200 & n9439 ) | ( ~n9200 & n9448 ) | ( n9439 & n9448 ) ;
  assign n9451 = ( n9200 & ~n9449 ) | ( n9200 & n9450 ) | ( ~n9449 & n9450 ) ;
  assign n9452 = ( n9212 & n9424 ) | ( n9212 & n9451 ) | ( n9424 & n9451 ) ;
  assign n9453 = ( n9212 & ~n9424 ) | ( n9212 & n9451 ) | ( ~n9424 & n9451 ) ;
  assign n9454 = ( n9424 & ~n9452 ) | ( n9424 & n9453 ) | ( ~n9452 & n9453 ) ;
  assign n9455 = n701 & n6027 ;
  assign n9456 = x78 & n6031 ;
  assign n9457 = x79 | n9456 ;
  assign n9458 = ( n6033 & n9456 ) | ( n6033 & n9457 ) | ( n9456 & n9457 ) ;
  assign n9459 = x77 & n6303 ;
  assign n9460 = n9458 | n9459 ;
  assign n9461 = ( x53 & n9455 ) | ( x53 & ~n9460 ) | ( n9455 & ~n9460 ) ;
  assign n9462 = ( ~x53 & n9460 ) | ( ~x53 & n9461 ) | ( n9460 & n9461 ) ;
  assign n9463 = ( ~n9455 & n9461 ) | ( ~n9455 & n9462 ) | ( n9461 & n9462 ) ;
  assign n9464 = ( n9215 & n9454 ) | ( n9215 & n9463 ) | ( n9454 & n9463 ) ;
  assign n9465 = ( ~n9215 & n9454 ) | ( ~n9215 & n9463 ) | ( n9454 & n9463 ) ;
  assign n9466 = ( n9215 & ~n9464 ) | ( n9215 & n9465 ) | ( ~n9464 & n9465 ) ;
  assign n9467 = n990 & n5374 ;
  assign n9468 = x81 & n5378 ;
  assign n9469 = x82 | n9468 ;
  assign n9470 = ( n5380 & n9468 ) | ( n5380 & n9469 ) | ( n9468 & n9469 ) ;
  assign n9471 = x80 & n5638 ;
  assign n9472 = n9470 | n9471 ;
  assign n9473 = ( x50 & n9467 ) | ( x50 & ~n9472 ) | ( n9467 & ~n9472 ) ;
  assign n9474 = ( ~x50 & n9472 ) | ( ~x50 & n9473 ) | ( n9472 & n9473 ) ;
  assign n9475 = ( ~n9467 & n9473 ) | ( ~n9467 & n9474 ) | ( n9473 & n9474 ) ;
  assign n9476 = ( n9227 & n9466 ) | ( n9227 & n9475 ) | ( n9466 & n9475 ) ;
  assign n9477 = ( ~n9227 & n9466 ) | ( ~n9227 & n9475 ) | ( n9466 & n9475 ) ;
  assign n9478 = ( n9227 & ~n9476 ) | ( n9227 & n9477 ) | ( ~n9476 & n9477 ) ;
  assign n9479 = n1262 & n4787 ;
  assign n9480 = x84 & n4791 ;
  assign n9481 = x85 | n9480 ;
  assign n9482 = ( n4793 & n9480 ) | ( n4793 & n9481 ) | ( n9480 & n9481 ) ;
  assign n9483 = x83 & n5030 ;
  assign n9484 = n9482 | n9483 ;
  assign n9485 = ( x47 & n9479 ) | ( x47 & ~n9484 ) | ( n9479 & ~n9484 ) ;
  assign n9486 = ( ~x47 & n9484 ) | ( ~x47 & n9485 ) | ( n9484 & n9485 ) ;
  assign n9487 = ( ~n9479 & n9485 ) | ( ~n9479 & n9486 ) | ( n9485 & n9486 ) ;
  assign n9488 = ( n9230 & n9478 ) | ( n9230 & n9487 ) | ( n9478 & n9487 ) ;
  assign n9489 = ( ~n9230 & n9478 ) | ( ~n9230 & n9487 ) | ( n9478 & n9487 ) ;
  assign n9490 = ( n9230 & ~n9488 ) | ( n9230 & n9489 ) | ( ~n9488 & n9489 ) ;
  assign n9491 = n1481 & n4227 ;
  assign n9492 = x87 & n4231 ;
  assign n9493 = x88 | n9492 ;
  assign n9494 = ( n4233 & n9492 ) | ( n4233 & n9493 ) | ( n9492 & n9493 ) ;
  assign n9495 = x86 & n4470 ;
  assign n9496 = n9494 | n9495 ;
  assign n9497 = ( x44 & n9491 ) | ( x44 & ~n9496 ) | ( n9491 & ~n9496 ) ;
  assign n9498 = ( ~x44 & n9496 ) | ( ~x44 & n9497 ) | ( n9496 & n9497 ) ;
  assign n9499 = ( ~n9491 & n9497 ) | ( ~n9491 & n9498 ) | ( n9497 & n9498 ) ;
  assign n9500 = ( n9242 & n9490 ) | ( n9242 & n9499 ) | ( n9490 & n9499 ) ;
  assign n9501 = ( n9242 & ~n9490 ) | ( n9242 & n9499 ) | ( ~n9490 & n9499 ) ;
  assign n9502 = ( n9490 & ~n9500 ) | ( n9490 & n9501 ) | ( ~n9500 & n9501 ) ;
  assign n9503 = n1914 & n3715 ;
  assign n9504 = x90 & n3719 ;
  assign n9505 = x91 | n9504 ;
  assign n9506 = ( n3721 & n9504 ) | ( n3721 & n9505 ) | ( n9504 & n9505 ) ;
  assign n9507 = x89 & n3922 ;
  assign n9508 = n9506 | n9507 ;
  assign n9509 = ( x41 & n9503 ) | ( x41 & ~n9508 ) | ( n9503 & ~n9508 ) ;
  assign n9510 = ( ~x41 & n9508 ) | ( ~x41 & n9509 ) | ( n9508 & n9509 ) ;
  assign n9511 = ( ~n9503 & n9509 ) | ( ~n9503 & n9510 ) | ( n9509 & n9510 ) ;
  assign n9512 = ( n9245 & n9502 ) | ( n9245 & n9511 ) | ( n9502 & n9511 ) ;
  assign n9513 = ( ~n9245 & n9502 ) | ( ~n9245 & n9511 ) | ( n9502 & n9511 ) ;
  assign n9514 = ( n9245 & ~n9512 ) | ( n9245 & n9513 ) | ( ~n9512 & n9513 ) ;
  assign n9515 = n2294 & n3224 ;
  assign n9516 = x93 & n3228 ;
  assign n9517 = x94 | n9516 ;
  assign n9518 = ( n3230 & n9516 ) | ( n3230 & n9517 ) | ( n9516 & n9517 ) ;
  assign n9519 = x92 & n3413 ;
  assign n9520 = n9518 | n9519 ;
  assign n9521 = ( x38 & n9515 ) | ( x38 & ~n9520 ) | ( n9515 & ~n9520 ) ;
  assign n9522 = ( ~x38 & n9520 ) | ( ~x38 & n9521 ) | ( n9520 & n9521 ) ;
  assign n9523 = ( ~n9515 & n9521 ) | ( ~n9515 & n9522 ) | ( n9521 & n9522 ) ;
  assign n9524 = ( n9257 & n9514 ) | ( n9257 & n9523 ) | ( n9514 & n9523 ) ;
  assign n9525 = ( ~n9257 & n9514 ) | ( ~n9257 & n9523 ) | ( n9514 & n9523 ) ;
  assign n9526 = ( n9257 & ~n9524 ) | ( n9257 & n9525 ) | ( ~n9524 & n9525 ) ;
  assign n9527 = n2585 & n2766 ;
  assign n9528 = x96 & n2770 ;
  assign n9529 = x97 | n9528 ;
  assign n9530 = ( n2772 & n9528 ) | ( n2772 & n9529 ) | ( n9528 & n9529 ) ;
  assign n9531 = x95 & n2943 ;
  assign n9532 = n9530 | n9531 ;
  assign n9533 = ( x35 & n9527 ) | ( x35 & ~n9532 ) | ( n9527 & ~n9532 ) ;
  assign n9534 = ( ~x35 & n9532 ) | ( ~x35 & n9533 ) | ( n9532 & n9533 ) ;
  assign n9535 = ( ~n9527 & n9533 ) | ( ~n9527 & n9534 ) | ( n9533 & n9534 ) ;
  assign n9536 = ( n9269 & n9526 ) | ( n9269 & n9535 ) | ( n9526 & n9535 ) ;
  assign n9537 = ( n9269 & ~n9526 ) | ( n9269 & n9535 ) | ( ~n9526 & n9535 ) ;
  assign n9538 = ( n9526 & ~n9536 ) | ( n9526 & n9537 ) | ( ~n9536 & n9537 ) ;
  assign n9539 = n2320 & n3162 ;
  assign n9540 = x99 & n2324 ;
  assign n9541 = x100 | n9540 ;
  assign n9542 = ( n2326 & n9540 ) | ( n2326 & n9541 ) | ( n9540 & n9541 ) ;
  assign n9543 = x98 & n2497 ;
  assign n9544 = n9542 | n9543 ;
  assign n9545 = ( x32 & n9539 ) | ( x32 & ~n9544 ) | ( n9539 & ~n9544 ) ;
  assign n9546 = ( ~x32 & n9544 ) | ( ~x32 & n9545 ) | ( n9544 & n9545 ) ;
  assign n9547 = ( ~n9539 & n9545 ) | ( ~n9539 & n9546 ) | ( n9545 & n9546 ) ;
  assign n9548 = ( n9281 & n9538 ) | ( n9281 & n9547 ) | ( n9538 & n9547 ) ;
  assign n9549 = ( n9281 & ~n9538 ) | ( n9281 & n9547 ) | ( ~n9538 & n9547 ) ;
  assign n9550 = ( n9538 & ~n9548 ) | ( n9538 & n9549 ) | ( ~n9548 & n9549 ) ;
  assign n9551 = ( n9284 & n9415 ) | ( n9284 & n9550 ) | ( n9415 & n9550 ) ;
  assign n9552 = ( ~n9284 & n9415 ) | ( ~n9284 & n9550 ) | ( n9415 & n9550 ) ;
  assign n9553 = ( n9284 & ~n9551 ) | ( n9284 & n9552 ) | ( ~n9551 & n9552 ) ;
  assign n9554 = ( n9296 & n9406 ) | ( n9296 & n9553 ) | ( n9406 & n9553 ) ;
  assign n9555 = ( n9296 & ~n9406 ) | ( n9296 & n9553 ) | ( ~n9406 & n9553 ) ;
  assign n9556 = ( n9406 & ~n9554 ) | ( n9406 & n9555 ) | ( ~n9554 & n9555 ) ;
  assign n9557 = n1297 & n4734 ;
  assign n9558 = x108 & n1301 ;
  assign n9559 = x109 | n9558 ;
  assign n9560 = ( n1303 & n9558 ) | ( n1303 & n9559 ) | ( n9558 & n9559 ) ;
  assign n9561 = x107 & n1426 ;
  assign n9562 = n9560 | n9561 ;
  assign n9563 = ( x23 & n9557 ) | ( x23 & ~n9562 ) | ( n9557 & ~n9562 ) ;
  assign n9564 = ( ~x23 & n9562 ) | ( ~x23 & n9563 ) | ( n9562 & n9563 ) ;
  assign n9565 = ( ~n9557 & n9563 ) | ( ~n9557 & n9564 ) | ( n9563 & n9564 ) ;
  assign n9566 = ( n9308 & n9556 ) | ( n9308 & n9565 ) | ( n9556 & n9565 ) ;
  assign n9567 = ( n9308 & ~n9556 ) | ( n9308 & n9565 ) | ( ~n9556 & n9565 ) ;
  assign n9568 = ( n9556 & ~n9566 ) | ( n9556 & n9567 ) | ( ~n9566 & n9567 ) ;
  assign n9569 = ( n9311 & n9397 ) | ( n9311 & n9568 ) | ( n9397 & n9568 ) ;
  assign n9570 = ( n9311 & ~n9397 ) | ( n9311 & n9568 ) | ( ~n9397 & n9568 ) ;
  assign n9571 = ( n9397 & ~n9569 ) | ( n9397 & n9570 ) | ( ~n9569 & n9570 ) ;
  assign n9572 = ( n9314 & n9388 ) | ( n9314 & n9571 ) | ( n9388 & n9571 ) ;
  assign n9573 = ( n9314 & ~n9388 ) | ( n9314 & n9571 ) | ( ~n9388 & n9571 ) ;
  assign n9574 = ( n9388 & ~n9572 ) | ( n9388 & n9573 ) | ( ~n9572 & n9573 ) ;
  assign n9575 = n583 & n6421 ;
  assign n9576 = x117 & n587 ;
  assign n9577 = x118 | n9576 ;
  assign n9578 = ( n589 & n9576 ) | ( n589 & n9577 ) | ( n9576 & n9577 ) ;
  assign n9579 = x116 & n676 ;
  assign n9580 = n9578 | n9579 ;
  assign n9581 = ( x14 & n9575 ) | ( x14 & ~n9580 ) | ( n9575 & ~n9580 ) ;
  assign n9582 = ( ~x14 & n9580 ) | ( ~x14 & n9581 ) | ( n9580 & n9581 ) ;
  assign n9583 = ( ~n9575 & n9581 ) | ( ~n9575 & n9582 ) | ( n9581 & n9582 ) ;
  assign n9584 = ( n9317 & n9574 ) | ( n9317 & n9583 ) | ( n9574 & n9583 ) ;
  assign n9585 = ( n9317 & ~n9574 ) | ( n9317 & n9583 ) | ( ~n9574 & n9583 ) ;
  assign n9586 = ( n9574 & ~n9584 ) | ( n9574 & n9585 ) | ( ~n9584 & n9585 ) ;
  assign n9587 = ( n9329 & n9379 ) | ( n9329 & n9586 ) | ( n9379 & n9586 ) ;
  assign n9588 = ( n9329 & ~n9379 ) | ( n9329 & n9586 ) | ( ~n9379 & n9586 ) ;
  assign n9589 = ( n9379 & ~n9587 ) | ( n9379 & n9588 ) | ( ~n9587 & n9588 ) ;
  assign n9590 = n291 & n7841 ;
  assign n9591 = x123 & n295 ;
  assign n9592 = x124 | n9591 ;
  assign n9593 = ( n297 & n9591 ) | ( n297 & n9592 ) | ( n9591 & n9592 ) ;
  assign n9594 = x122 & n330 ;
  assign n9595 = n9593 | n9594 ;
  assign n9596 = ( x8 & n9590 ) | ( x8 & ~n9595 ) | ( n9590 & ~n9595 ) ;
  assign n9597 = ( ~x8 & n9595 ) | ( ~x8 & n9596 ) | ( n9595 & n9596 ) ;
  assign n9598 = ( ~n9590 & n9596 ) | ( ~n9590 & n9597 ) | ( n9596 & n9597 ) ;
  assign n9599 = ( n9350 & n9589 ) | ( n9350 & n9598 ) | ( n9589 & n9598 ) ;
  assign n9600 = ( n9350 & ~n9589 ) | ( n9350 & n9598 ) | ( ~n9589 & n9598 ) ;
  assign n9601 = ( n9589 & ~n9599 ) | ( n9589 & n9600 ) | ( ~n9599 & n9600 ) ;
  assign n9602 = n186 & n8846 ;
  assign n9603 = x126 & n190 ;
  assign n9604 = x127 | n9603 ;
  assign n9605 = ( n192 & n9603 ) | ( n192 & n9604 ) | ( n9603 & n9604 ) ;
  assign n9606 = x125 & n220 ;
  assign n9607 = n9605 | n9606 ;
  assign n9608 = ( x5 & n9602 ) | ( x5 & ~n9607 ) | ( n9602 & ~n9607 ) ;
  assign n9609 = ( ~x5 & n9607 ) | ( ~x5 & n9608 ) | ( n9607 & n9608 ) ;
  assign n9610 = ( ~n9602 & n9608 ) | ( ~n9602 & n9609 ) | ( n9608 & n9609 ) ;
  assign n9611 = ( n9362 & n9601 ) | ( n9362 & n9610 ) | ( n9601 & n9610 ) ;
  assign n9612 = ( n9362 & ~n9601 ) | ( n9362 & n9610 ) | ( ~n9601 & n9610 ) ;
  assign n9613 = ( n9601 & ~n9611 ) | ( n9601 & n9612 ) | ( ~n9611 & n9612 ) ;
  assign n9614 = ( n9365 & n9368 ) | ( n9365 & n9613 ) | ( n9368 & n9613 ) ;
  assign n9615 = ( ~n9365 & n9368 ) | ( ~n9365 & n9613 ) | ( n9368 & n9613 ) ;
  assign n9616 = ( n9365 & ~n9614 ) | ( n9365 & n9615 ) | ( ~n9614 & n9615 ) ;
  assign n9617 = n583 & n6645 ;
  assign n9618 = x118 & n587 ;
  assign n9619 = x119 | n9618 ;
  assign n9620 = ( n589 & n9618 ) | ( n589 & n9619 ) | ( n9618 & n9619 ) ;
  assign n9621 = x117 & n676 ;
  assign n9622 = n9620 | n9621 ;
  assign n9623 = ( x14 & n9617 ) | ( x14 & ~n9622 ) | ( n9617 & ~n9622 ) ;
  assign n9624 = ( ~x14 & n9622 ) | ( ~x14 & n9623 ) | ( n9622 & n9623 ) ;
  assign n9625 = ( ~n9617 & n9623 ) | ( ~n9617 & n9624 ) | ( n9623 & n9624 ) ;
  assign n9626 = n1016 & n5542 ;
  assign n9627 = x112 & n1020 ;
  assign n9628 = x113 | n9627 ;
  assign n9629 = ( n1022 & n9627 ) | ( n1022 & n9628 ) | ( n9627 & n9628 ) ;
  assign n9630 = x111 & n1145 ;
  assign n9631 = n9629 | n9630 ;
  assign n9632 = ( x20 & n9626 ) | ( x20 & ~n9631 ) | ( n9626 & ~n9631 ) ;
  assign n9633 = ( ~x20 & n9631 ) | ( ~x20 & n9632 ) | ( n9631 & n9632 ) ;
  assign n9634 = ( ~n9626 & n9632 ) | ( ~n9626 & n9633 ) | ( n9632 & n9633 ) ;
  assign n9635 = n1617 & n4362 ;
  assign n9636 = x106 & n1621 ;
  assign n9637 = x107 | n9636 ;
  assign n9638 = ( n1623 & n9636 ) | ( n1623 & n9637 ) | ( n9636 & n9637 ) ;
  assign n9639 = x105 & n1749 ;
  assign n9640 = n9638 | n9639 ;
  assign n9641 = ( x26 & n9635 ) | ( x26 & ~n9640 ) | ( n9635 & ~n9640 ) ;
  assign n9642 = ( ~x26 & n9640 ) | ( ~x26 & n9641 ) | ( n9640 & n9641 ) ;
  assign n9643 = ( ~n9635 & n9641 ) | ( ~n9635 & n9642 ) | ( n9641 & n9642 ) ;
  assign n9644 = n2320 & n3326 ;
  assign n9645 = x100 & n2324 ;
  assign n9646 = x101 | n9645 ;
  assign n9647 = ( n2326 & n9645 ) | ( n2326 & n9646 ) | ( n9645 & n9646 ) ;
  assign n9648 = x99 & n2497 ;
  assign n9649 = n9647 | n9648 ;
  assign n9650 = ( x32 & n9644 ) | ( x32 & ~n9649 ) | ( n9644 & ~n9649 ) ;
  assign n9651 = ( ~x32 & n9649 ) | ( ~x32 & n9650 ) | ( n9649 & n9650 ) ;
  assign n9652 = ( ~n9644 & n9650 ) | ( ~n9644 & n9651 ) | ( n9650 & n9651 ) ;
  assign n9653 = n2725 & n2766 ;
  assign n9654 = x97 & n2770 ;
  assign n9655 = x98 | n9654 ;
  assign n9656 = ( n2772 & n9654 ) | ( n2772 & n9655 ) | ( n9654 & n9655 ) ;
  assign n9657 = x96 & n2943 ;
  assign n9658 = n9656 | n9657 ;
  assign n9659 = ( x35 & n9653 ) | ( x35 & ~n9658 ) | ( n9653 & ~n9658 ) ;
  assign n9660 = ( ~x35 & n9658 ) | ( ~x35 & n9659 ) | ( n9658 & n9659 ) ;
  assign n9661 = ( ~n9653 & n9659 ) | ( ~n9653 & n9660 ) | ( n9659 & n9660 ) ;
  assign n9662 = n277 & n8154 ;
  assign n9663 = x70 & n8158 ;
  assign n9664 = x71 | n9663 ;
  assign n9665 = ( n8160 & n9663 ) | ( n8160 & n9664 ) | ( n9663 & n9664 ) ;
  assign n9666 = x69 & n8439 ;
  assign n9667 = n9665 | n9666 ;
  assign n9668 = ( x62 & n9662 ) | ( x62 & ~n9667 ) | ( n9662 & ~n9667 ) ;
  assign n9669 = ( ~x62 & n9667 ) | ( ~x62 & n9668 ) | ( n9667 & n9668 ) ;
  assign n9670 = ( ~n9662 & n9668 ) | ( ~n9662 & n9669 ) | ( n9668 & n9669 ) ;
  assign n9671 = x67 & n8927 ;
  assign n9672 = ( ~x68 & n8693 ) | ( ~x68 & n8927 ) | ( n8693 & n8927 ) ;
  assign n9673 = ( n8693 & n9671 ) | ( n8693 & ~n9672 ) | ( n9671 & ~n9672 ) ;
  assign n9674 = ( x2 & n9670 ) | ( x2 & n9673 ) | ( n9670 & n9673 ) ;
  assign n9675 = ( ~x2 & n9670 ) | ( ~x2 & n9673 ) | ( n9670 & n9673 ) ;
  assign n9676 = ( x2 & ~n9674 ) | ( x2 & n9675 ) | ( ~n9674 & n9675 ) ;
  assign n9677 = n446 & n7423 ;
  assign n9678 = x73 & n7427 ;
  assign n9679 = x74 | n9678 ;
  assign n9680 = ( n7429 & n9678 ) | ( n7429 & n9679 ) | ( n9678 & n9679 ) ;
  assign n9681 = x72 & n7708 ;
  assign n9682 = n9680 | n9681 ;
  assign n9683 = ( x59 & n9677 ) | ( x59 & ~n9682 ) | ( n9677 & ~n9682 ) ;
  assign n9684 = ( ~x59 & n9682 ) | ( ~x59 & n9683 ) | ( n9682 & n9683 ) ;
  assign n9685 = ( ~n9677 & n9683 ) | ( ~n9677 & n9684 ) | ( n9683 & n9684 ) ;
  assign n9686 = ( n9437 & n9676 ) | ( n9437 & n9685 ) | ( n9676 & n9685 ) ;
  assign n9687 = ( ~n9437 & n9676 ) | ( ~n9437 & n9685 ) | ( n9676 & n9685 ) ;
  assign n9688 = ( n9437 & ~n9686 ) | ( n9437 & n9687 ) | ( ~n9686 & n9687 ) ;
  assign n9689 = n569 & n6713 ;
  assign n9690 = x76 & n6717 ;
  assign n9691 = x77 | n9690 ;
  assign n9692 = ( n6719 & n9690 ) | ( n6719 & n9691 ) | ( n9690 & n9691 ) ;
  assign n9693 = x75 & n6980 ;
  assign n9694 = n9692 | n9693 ;
  assign n9695 = ( x56 & n9689 ) | ( x56 & ~n9694 ) | ( n9689 & ~n9694 ) ;
  assign n9696 = ( ~x56 & n9694 ) | ( ~x56 & n9695 ) | ( n9694 & n9695 ) ;
  assign n9697 = ( ~n9689 & n9695 ) | ( ~n9689 & n9696 ) | ( n9695 & n9696 ) ;
  assign n9698 = ( n9449 & n9688 ) | ( n9449 & n9697 ) | ( n9688 & n9697 ) ;
  assign n9699 = ( ~n9449 & n9688 ) | ( ~n9449 & n9697 ) | ( n9688 & n9697 ) ;
  assign n9700 = ( n9449 & ~n9698 ) | ( n9449 & n9699 ) | ( ~n9698 & n9699 ) ;
  assign n9701 = n769 & n6027 ;
  assign n9702 = x79 & n6031 ;
  assign n9703 = x80 | n9702 ;
  assign n9704 = ( n6033 & n9702 ) | ( n6033 & n9703 ) | ( n9702 & n9703 ) ;
  assign n9705 = x78 & n6303 ;
  assign n9706 = n9704 | n9705 ;
  assign n9707 = ( x53 & n9701 ) | ( x53 & ~n9706 ) | ( n9701 & ~n9706 ) ;
  assign n9708 = ( ~x53 & n9706 ) | ( ~x53 & n9707 ) | ( n9706 & n9707 ) ;
  assign n9709 = ( ~n9701 & n9707 ) | ( ~n9701 & n9708 ) | ( n9707 & n9708 ) ;
  assign n9710 = ( n9452 & n9700 ) | ( n9452 & n9709 ) | ( n9700 & n9709 ) ;
  assign n9711 = ( n9452 & ~n9700 ) | ( n9452 & n9709 ) | ( ~n9700 & n9709 ) ;
  assign n9712 = ( n9700 & ~n9710 ) | ( n9700 & n9711 ) | ( ~n9710 & n9711 ) ;
  assign n9713 = n1082 & n5374 ;
  assign n9714 = x82 & n5378 ;
  assign n9715 = x83 | n9714 ;
  assign n9716 = ( n5380 & n9714 ) | ( n5380 & n9715 ) | ( n9714 & n9715 ) ;
  assign n9717 = x81 & n5638 ;
  assign n9718 = n9716 | n9717 ;
  assign n9719 = ( x50 & n9713 ) | ( x50 & ~n9718 ) | ( n9713 & ~n9718 ) ;
  assign n9720 = ( ~x50 & n9718 ) | ( ~x50 & n9719 ) | ( n9718 & n9719 ) ;
  assign n9721 = ( ~n9713 & n9719 ) | ( ~n9713 & n9720 ) | ( n9719 & n9720 ) ;
  assign n9722 = ( n9464 & n9712 ) | ( n9464 & n9721 ) | ( n9712 & n9721 ) ;
  assign n9723 = ( ~n9464 & n9712 ) | ( ~n9464 & n9721 ) | ( n9712 & n9721 ) ;
  assign n9724 = ( n9464 & ~n9722 ) | ( n9464 & n9723 ) | ( ~n9722 & n9723 ) ;
  assign n9725 = n1366 & n4787 ;
  assign n9726 = x85 & n4791 ;
  assign n9727 = x86 | n9726 ;
  assign n9728 = ( n4793 & n9726 ) | ( n4793 & n9727 ) | ( n9726 & n9727 ) ;
  assign n9729 = x84 & n5030 ;
  assign n9730 = n9728 | n9729 ;
  assign n9731 = ( x47 & n9725 ) | ( x47 & ~n9730 ) | ( n9725 & ~n9730 ) ;
  assign n9732 = ( ~x47 & n9730 ) | ( ~x47 & n9731 ) | ( n9730 & n9731 ) ;
  assign n9733 = ( ~n9725 & n9731 ) | ( ~n9725 & n9732 ) | ( n9731 & n9732 ) ;
  assign n9734 = ( n9476 & n9724 ) | ( n9476 & n9733 ) | ( n9724 & n9733 ) ;
  assign n9735 = ( ~n9476 & n9724 ) | ( ~n9476 & n9733 ) | ( n9724 & n9733 ) ;
  assign n9736 = ( n9476 & ~n9734 ) | ( n9476 & n9735 ) | ( ~n9734 & n9735 ) ;
  assign n9737 = n1585 & n4227 ;
  assign n9738 = x88 & n4231 ;
  assign n9739 = x89 | n9738 ;
  assign n9740 = ( n4233 & n9738 ) | ( n4233 & n9739 ) | ( n9738 & n9739 ) ;
  assign n9741 = x87 & n4470 ;
  assign n9742 = n9740 | n9741 ;
  assign n9743 = ( x44 & n9737 ) | ( x44 & ~n9742 ) | ( n9737 & ~n9742 ) ;
  assign n9744 = ( ~x44 & n9742 ) | ( ~x44 & n9743 ) | ( n9742 & n9743 ) ;
  assign n9745 = ( ~n9737 & n9743 ) | ( ~n9737 & n9744 ) | ( n9743 & n9744 ) ;
  assign n9746 = ( n9488 & n9736 ) | ( n9488 & n9745 ) | ( n9736 & n9745 ) ;
  assign n9747 = ( ~n9488 & n9736 ) | ( ~n9488 & n9745 ) | ( n9736 & n9745 ) ;
  assign n9748 = ( n9488 & ~n9746 ) | ( n9488 & n9747 ) | ( ~n9746 & n9747 ) ;
  assign n9749 = n2042 & n3715 ;
  assign n9750 = x91 & n3719 ;
  assign n9751 = x92 | n9750 ;
  assign n9752 = ( n3721 & n9750 ) | ( n3721 & n9751 ) | ( n9750 & n9751 ) ;
  assign n9753 = x90 & n3922 ;
  assign n9754 = n9752 | n9753 ;
  assign n9755 = ( x41 & n9749 ) | ( x41 & ~n9754 ) | ( n9749 & ~n9754 ) ;
  assign n9756 = ( ~x41 & n9754 ) | ( ~x41 & n9755 ) | ( n9754 & n9755 ) ;
  assign n9757 = ( ~n9749 & n9755 ) | ( ~n9749 & n9756 ) | ( n9755 & n9756 ) ;
  assign n9758 = ( n9500 & n9748 ) | ( n9500 & n9757 ) | ( n9748 & n9757 ) ;
  assign n9759 = ( ~n9500 & n9748 ) | ( ~n9500 & n9757 ) | ( n9748 & n9757 ) ;
  assign n9760 = ( n9500 & ~n9758 ) | ( n9500 & n9759 ) | ( ~n9758 & n9759 ) ;
  assign n9761 = n2434 & n3224 ;
  assign n9762 = x94 & n3228 ;
  assign n9763 = x95 | n9762 ;
  assign n9764 = ( n3230 & n9762 ) | ( n3230 & n9763 ) | ( n9762 & n9763 ) ;
  assign n9765 = x93 & n3413 ;
  assign n9766 = n9764 | n9765 ;
  assign n9767 = ( x38 & n9761 ) | ( x38 & ~n9766 ) | ( n9761 & ~n9766 ) ;
  assign n9768 = ( ~x38 & n9766 ) | ( ~x38 & n9767 ) | ( n9766 & n9767 ) ;
  assign n9769 = ( ~n9761 & n9767 ) | ( ~n9761 & n9768 ) | ( n9767 & n9768 ) ;
  assign n9770 = ( n9512 & n9760 ) | ( n9512 & n9769 ) | ( n9760 & n9769 ) ;
  assign n9771 = ( ~n9512 & n9760 ) | ( ~n9512 & n9769 ) | ( n9760 & n9769 ) ;
  assign n9772 = ( n9512 & ~n9770 ) | ( n9512 & n9771 ) | ( ~n9770 & n9771 ) ;
  assign n9773 = ( n9524 & n9661 ) | ( n9524 & n9772 ) | ( n9661 & n9772 ) ;
  assign n9774 = ( n9524 & ~n9661 ) | ( n9524 & n9772 ) | ( ~n9661 & n9772 ) ;
  assign n9775 = ( n9661 & ~n9773 ) | ( n9661 & n9774 ) | ( ~n9773 & n9774 ) ;
  assign n9776 = ( n9536 & n9652 ) | ( n9536 & n9775 ) | ( n9652 & n9775 ) ;
  assign n9777 = ( ~n9536 & n9652 ) | ( ~n9536 & n9775 ) | ( n9652 & n9775 ) ;
  assign n9778 = ( n9536 & ~n9776 ) | ( n9536 & n9777 ) | ( ~n9776 & n9777 ) ;
  assign n9779 = n1949 & n3665 ;
  assign n9780 = x103 & n1953 ;
  assign n9781 = x104 | n9780 ;
  assign n9782 = ( n1955 & n9780 ) | ( n1955 & n9781 ) | ( n9780 & n9781 ) ;
  assign n9783 = x102 & n2114 ;
  assign n9784 = n9782 | n9783 ;
  assign n9785 = ( x29 & n9779 ) | ( x29 & ~n9784 ) | ( n9779 & ~n9784 ) ;
  assign n9786 = ( ~x29 & n9784 ) | ( ~x29 & n9785 ) | ( n9784 & n9785 ) ;
  assign n9787 = ( ~n9779 & n9785 ) | ( ~n9779 & n9786 ) | ( n9785 & n9786 ) ;
  assign n9788 = ( n9548 & n9778 ) | ( n9548 & n9787 ) | ( n9778 & n9787 ) ;
  assign n9789 = ( n9548 & ~n9778 ) | ( n9548 & n9787 ) | ( ~n9778 & n9787 ) ;
  assign n9790 = ( n9778 & ~n9788 ) | ( n9778 & n9789 ) | ( ~n9788 & n9789 ) ;
  assign n9791 = ( n9551 & n9643 ) | ( n9551 & n9790 ) | ( n9643 & n9790 ) ;
  assign n9792 = ( n9551 & ~n9643 ) | ( n9551 & n9790 ) | ( ~n9643 & n9790 ) ;
  assign n9793 = ( n9643 & ~n9791 ) | ( n9643 & n9792 ) | ( ~n9791 & n9792 ) ;
  assign n9794 = n1297 & n4934 ;
  assign n9795 = x109 & n1301 ;
  assign n9796 = x110 | n9795 ;
  assign n9797 = ( n1303 & n9795 ) | ( n1303 & n9796 ) | ( n9795 & n9796 ) ;
  assign n9798 = x108 & n1426 ;
  assign n9799 = n9797 | n9798 ;
  assign n9800 = ( x23 & n9794 ) | ( x23 & ~n9799 ) | ( n9794 & ~n9799 ) ;
  assign n9801 = ( ~x23 & n9799 ) | ( ~x23 & n9800 ) | ( n9799 & n9800 ) ;
  assign n9802 = ( ~n9794 & n9800 ) | ( ~n9794 & n9801 ) | ( n9800 & n9801 ) ;
  assign n9803 = ( n9554 & n9793 ) | ( n9554 & n9802 ) | ( n9793 & n9802 ) ;
  assign n9804 = ( n9554 & ~n9793 ) | ( n9554 & n9802 ) | ( ~n9793 & n9802 ) ;
  assign n9805 = ( n9793 & ~n9803 ) | ( n9793 & n9804 ) | ( ~n9803 & n9804 ) ;
  assign n9806 = ( n9566 & n9634 ) | ( n9566 & n9805 ) | ( n9634 & n9805 ) ;
  assign n9807 = ( n9566 & ~n9634 ) | ( n9566 & n9805 ) | ( ~n9634 & n9805 ) ;
  assign n9808 = ( n9634 & ~n9806 ) | ( n9634 & n9807 ) | ( ~n9806 & n9807 ) ;
  assign n9809 = n810 & n5977 ;
  assign n9810 = x115 & n814 ;
  assign n9811 = x116 | n9810 ;
  assign n9812 = ( n816 & n9810 ) | ( n816 & n9811 ) | ( n9810 & n9811 ) ;
  assign n9813 = x114 & n885 ;
  assign n9814 = n9812 | n9813 ;
  assign n9815 = ( x17 & n9809 ) | ( x17 & ~n9814 ) | ( n9809 & ~n9814 ) ;
  assign n9816 = ( ~x17 & n9814 ) | ( ~x17 & n9815 ) | ( n9814 & n9815 ) ;
  assign n9817 = ( ~n9809 & n9815 ) | ( ~n9809 & n9816 ) | ( n9815 & n9816 ) ;
  assign n9818 = ( n9569 & n9808 ) | ( n9569 & n9817 ) | ( n9808 & n9817 ) ;
  assign n9819 = ( n9569 & ~n9808 ) | ( n9569 & n9817 ) | ( ~n9808 & n9817 ) ;
  assign n9820 = ( n9808 & ~n9818 ) | ( n9808 & n9819 ) | ( ~n9818 & n9819 ) ;
  assign n9821 = ( n9572 & n9625 ) | ( n9572 & n9820 ) | ( n9625 & n9820 ) ;
  assign n9822 = ( n9572 & ~n9625 ) | ( n9572 & n9820 ) | ( ~n9625 & n9820 ) ;
  assign n9823 = ( n9625 & ~n9821 ) | ( n9625 & n9822 ) | ( ~n9821 & n9822 ) ;
  assign n9824 = n407 & n7582 ;
  assign n9825 = x121 & n411 ;
  assign n9826 = x122 | n9825 ;
  assign n9827 = ( n413 & n9825 ) | ( n413 & n9826 ) | ( n9825 & n9826 ) ;
  assign n9828 = x120 & n491 ;
  assign n9829 = n9827 | n9828 ;
  assign n9830 = ( x11 & n9824 ) | ( x11 & ~n9829 ) | ( n9824 & ~n9829 ) ;
  assign n9831 = ( ~x11 & n9829 ) | ( ~x11 & n9830 ) | ( n9829 & n9830 ) ;
  assign n9832 = ( ~n9824 & n9830 ) | ( ~n9824 & n9831 ) | ( n9830 & n9831 ) ;
  assign n9833 = ( n9584 & n9823 ) | ( n9584 & n9832 ) | ( n9823 & n9832 ) ;
  assign n9834 = ( n9584 & ~n9823 ) | ( n9584 & n9832 ) | ( ~n9823 & n9832 ) ;
  assign n9835 = ( n9823 & ~n9833 ) | ( n9823 & n9834 ) | ( ~n9833 & n9834 ) ;
  assign n9836 = n291 & n8331 ;
  assign n9837 = x124 & n295 ;
  assign n9838 = x125 | n9837 ;
  assign n9839 = ( n297 & n9837 ) | ( n297 & n9838 ) | ( n9837 & n9838 ) ;
  assign n9840 = x123 & n330 ;
  assign n9841 = n9839 | n9840 ;
  assign n9842 = ( x8 & n9836 ) | ( x8 & ~n9841 ) | ( n9836 & ~n9841 ) ;
  assign n9843 = ( ~x8 & n9841 ) | ( ~x8 & n9842 ) | ( n9841 & n9842 ) ;
  assign n9844 = ( ~n9836 & n9842 ) | ( ~n9836 & n9843 ) | ( n9842 & n9843 ) ;
  assign n9845 = ( n9587 & n9835 ) | ( n9587 & n9844 ) | ( n9835 & n9844 ) ;
  assign n9846 = ( n9587 & ~n9835 ) | ( n9587 & n9844 ) | ( ~n9835 & n9844 ) ;
  assign n9847 = ( n9835 & ~n9845 ) | ( n9835 & n9846 ) | ( ~n9845 & n9846 ) ;
  assign n9848 = n186 & n8865 ;
  assign n9849 = x127 & n190 ;
  assign n9850 = x126 | n9849 ;
  assign n9851 = ( n220 & n9849 ) | ( n220 & n9850 ) | ( n9849 & n9850 ) ;
  assign n9852 = ( x5 & n9848 ) | ( x5 & ~n9851 ) | ( n9848 & ~n9851 ) ;
  assign n9853 = ( ~x5 & n9851 ) | ( ~x5 & n9852 ) | ( n9851 & n9852 ) ;
  assign n9854 = ( ~n9848 & n9852 ) | ( ~n9848 & n9853 ) | ( n9852 & n9853 ) ;
  assign n9855 = ( n9599 & n9847 ) | ( n9599 & n9854 ) | ( n9847 & n9854 ) ;
  assign n9856 = ( n9599 & ~n9847 ) | ( n9599 & n9854 ) | ( ~n9847 & n9854 ) ;
  assign n9857 = ( n9847 & ~n9855 ) | ( n9847 & n9856 ) | ( ~n9855 & n9856 ) ;
  assign n9858 = ( n9611 & n9614 ) | ( n9611 & n9857 ) | ( n9614 & n9857 ) ;
  assign n9859 = ( n9611 & ~n9614 ) | ( n9611 & n9857 ) | ( ~n9614 & n9857 ) ;
  assign n9860 = ( n9614 & ~n9858 ) | ( n9614 & n9859 ) | ( ~n9858 & n9859 ) ;
  assign n9861 = n407 & n7597 ;
  assign n9862 = x122 & n411 ;
  assign n9863 = x123 | n9862 ;
  assign n9864 = ( n413 & n9862 ) | ( n413 & n9863 ) | ( n9862 & n9863 ) ;
  assign n9865 = x121 & n491 ;
  assign n9866 = n9864 | n9865 ;
  assign n9867 = ( x11 & n9861 ) | ( x11 & ~n9866 ) | ( n9861 & ~n9866 ) ;
  assign n9868 = ( ~x11 & n9866 ) | ( ~x11 & n9867 ) | ( n9866 & n9867 ) ;
  assign n9869 = ( ~n9861 & n9867 ) | ( ~n9861 & n9868 ) | ( n9867 & n9868 ) ;
  assign n9870 = n583 & n7098 ;
  assign n9871 = x119 & n587 ;
  assign n9872 = x120 | n9871 ;
  assign n9873 = ( n589 & n9871 ) | ( n589 & n9872 ) | ( n9871 & n9872 ) ;
  assign n9874 = x118 & n676 ;
  assign n9875 = n9873 | n9874 ;
  assign n9876 = ( x14 & n9870 ) | ( x14 & ~n9875 ) | ( n9870 & ~n9875 ) ;
  assign n9877 = ( ~x14 & n9875 ) | ( ~x14 & n9876 ) | ( n9875 & n9876 ) ;
  assign n9878 = ( ~n9870 & n9876 ) | ( ~n9870 & n9877 ) | ( n9876 & n9877 ) ;
  assign n9879 = n810 & n6201 ;
  assign n9880 = x116 & n814 ;
  assign n9881 = x117 | n9880 ;
  assign n9882 = ( n816 & n9880 ) | ( n816 & n9881 ) | ( n9880 & n9881 ) ;
  assign n9883 = x115 & n885 ;
  assign n9884 = n9882 | n9883 ;
  assign n9885 = ( x17 & n9879 ) | ( x17 & ~n9884 ) | ( n9879 & ~n9884 ) ;
  assign n9886 = ( ~x17 & n9884 ) | ( ~x17 & n9885 ) | ( n9884 & n9885 ) ;
  assign n9887 = ( ~n9879 & n9885 ) | ( ~n9879 & n9886 ) | ( n9885 & n9886 ) ;
  assign n9888 = n1016 & n5750 ;
  assign n9889 = x113 & n1020 ;
  assign n9890 = x114 | n9889 ;
  assign n9891 = ( n1022 & n9889 ) | ( n1022 & n9890 ) | ( n9889 & n9890 ) ;
  assign n9892 = x112 & n1145 ;
  assign n9893 = n9891 | n9892 ;
  assign n9894 = ( x20 & n9888 ) | ( x20 & ~n9893 ) | ( n9888 & ~n9893 ) ;
  assign n9895 = ( ~x20 & n9893 ) | ( ~x20 & n9894 ) | ( n9893 & n9894 ) ;
  assign n9896 = ( ~n9888 & n9894 ) | ( ~n9888 & n9895 ) | ( n9894 & n9895 ) ;
  assign n9897 = n1297 & n5130 ;
  assign n9898 = x110 & n1301 ;
  assign n9899 = x111 | n9898 ;
  assign n9900 = ( n1303 & n9898 ) | ( n1303 & n9899 ) | ( n9898 & n9899 ) ;
  assign n9901 = x109 & n1426 ;
  assign n9902 = n9900 | n9901 ;
  assign n9903 = ( x23 & n9897 ) | ( x23 & ~n9902 ) | ( n9897 & ~n9902 ) ;
  assign n9904 = ( ~x23 & n9902 ) | ( ~x23 & n9903 ) | ( n9902 & n9903 ) ;
  assign n9905 = ( ~n9897 & n9903 ) | ( ~n9897 & n9904 ) | ( n9903 & n9904 ) ;
  assign n9906 = n1949 & n3998 ;
  assign n9907 = x104 & n1953 ;
  assign n9908 = x105 | n9907 ;
  assign n9909 = ( n1955 & n9907 ) | ( n1955 & n9908 ) | ( n9907 & n9908 ) ;
  assign n9910 = x103 & n2114 ;
  assign n9911 = n9909 | n9910 ;
  assign n9912 = ( x29 & n9906 ) | ( x29 & ~n9911 ) | ( n9906 & ~n9911 ) ;
  assign n9913 = ( ~x29 & n9911 ) | ( ~x29 & n9912 ) | ( n9911 & n9912 ) ;
  assign n9914 = ( ~n9906 & n9912 ) | ( ~n9906 & n9913 ) | ( n9912 & n9913 ) ;
  assign n9915 = n2320 & n3486 ;
  assign n9916 = x101 & n2324 ;
  assign n9917 = x102 | n9916 ;
  assign n9918 = ( n2326 & n9916 ) | ( n2326 & n9917 ) | ( n9916 & n9917 ) ;
  assign n9919 = x100 & n2497 ;
  assign n9920 = n9918 | n9919 ;
  assign n9921 = ( x32 & n9915 ) | ( x32 & ~n9920 ) | ( n9915 & ~n9920 ) ;
  assign n9922 = ( ~x32 & n9920 ) | ( ~x32 & n9921 ) | ( n9920 & n9921 ) ;
  assign n9923 = ( ~n9915 & n9921 ) | ( ~n9915 & n9922 ) | ( n9921 & n9922 ) ;
  assign n9924 = n346 & n8154 ;
  assign n9925 = x71 & n8158 ;
  assign n9926 = x72 | n9925 ;
  assign n9927 = ( n8160 & n9925 ) | ( n8160 & n9926 ) | ( n9925 & n9926 ) ;
  assign n9928 = x70 & n8439 ;
  assign n9929 = n9927 | n9928 ;
  assign n9930 = ( x62 & n9924 ) | ( x62 & ~n9929 ) | ( n9924 & ~n9929 ) ;
  assign n9931 = ( ~x62 & n9929 ) | ( ~x62 & n9930 ) | ( n9929 & n9930 ) ;
  assign n9932 = ( ~n9924 & n9930 ) | ( ~n9924 & n9931 ) | ( n9930 & n9931 ) ;
  assign n9933 = x68 & n8927 ;
  assign n9934 = ( ~x69 & n8693 ) | ( ~x69 & n8927 ) | ( n8693 & n8927 ) ;
  assign n9935 = ( n8693 & n9933 ) | ( n8693 & ~n9934 ) | ( n9933 & ~n9934 ) ;
  assign n9936 = ( x2 & n9932 ) | ( x2 & n9935 ) | ( n9932 & n9935 ) ;
  assign n9937 = ( ~x2 & n9932 ) | ( ~x2 & n9935 ) | ( n9932 & n9935 ) ;
  assign n9938 = ( x2 & ~n9936 ) | ( x2 & n9937 ) | ( ~n9936 & n9937 ) ;
  assign n9939 = n461 & n7423 ;
  assign n9940 = x74 & n7427 ;
  assign n9941 = x75 | n9940 ;
  assign n9942 = ( n7429 & n9940 ) | ( n7429 & n9941 ) | ( n9940 & n9941 ) ;
  assign n9943 = x73 & n7708 ;
  assign n9944 = n9942 | n9943 ;
  assign n9945 = ( x59 & n9939 ) | ( x59 & ~n9944 ) | ( n9939 & ~n9944 ) ;
  assign n9946 = ( ~x59 & n9944 ) | ( ~x59 & n9945 ) | ( n9944 & n9945 ) ;
  assign n9947 = ( ~n9939 & n9945 ) | ( ~n9939 & n9946 ) | ( n9945 & n9946 ) ;
  assign n9948 = ( n9674 & n9938 ) | ( n9674 & n9947 ) | ( n9938 & n9947 ) ;
  assign n9949 = ( ~n9674 & n9938 ) | ( ~n9674 & n9947 ) | ( n9938 & n9947 ) ;
  assign n9950 = ( n9674 & ~n9948 ) | ( n9674 & n9949 ) | ( ~n9948 & n9949 ) ;
  assign n9951 = n637 & n6713 ;
  assign n9952 = x77 & n6717 ;
  assign n9953 = x78 | n9952 ;
  assign n9954 = ( n6719 & n9952 ) | ( n6719 & n9953 ) | ( n9952 & n9953 ) ;
  assign n9955 = x76 & n6980 ;
  assign n9956 = n9954 | n9955 ;
  assign n9957 = ( x56 & n9951 ) | ( x56 & ~n9956 ) | ( n9951 & ~n9956 ) ;
  assign n9958 = ( ~x56 & n9956 ) | ( ~x56 & n9957 ) | ( n9956 & n9957 ) ;
  assign n9959 = ( ~n9951 & n9957 ) | ( ~n9951 & n9958 ) | ( n9957 & n9958 ) ;
  assign n9960 = ( n9686 & n9950 ) | ( n9686 & n9959 ) | ( n9950 & n9959 ) ;
  assign n9961 = ( n9686 & ~n9950 ) | ( n9686 & n9959 ) | ( ~n9950 & n9959 ) ;
  assign n9962 = ( n9950 & ~n9960 ) | ( n9950 & n9961 ) | ( ~n9960 & n9961 ) ;
  assign n9963 = n910 & n6027 ;
  assign n9964 = x80 & n6031 ;
  assign n9965 = x81 | n9964 ;
  assign n9966 = ( n6033 & n9964 ) | ( n6033 & n9965 ) | ( n9964 & n9965 ) ;
  assign n9967 = x79 & n6303 ;
  assign n9968 = n9966 | n9967 ;
  assign n9969 = ( x53 & n9963 ) | ( x53 & ~n9968 ) | ( n9963 & ~n9968 ) ;
  assign n9970 = ( ~x53 & n9968 ) | ( ~x53 & n9969 ) | ( n9968 & n9969 ) ;
  assign n9971 = ( ~n9963 & n9969 ) | ( ~n9963 & n9970 ) | ( n9969 & n9970 ) ;
  assign n9972 = ( n9698 & n9962 ) | ( n9698 & n9971 ) | ( n9962 & n9971 ) ;
  assign n9973 = ( ~n9698 & n9962 ) | ( ~n9698 & n9971 ) | ( n9962 & n9971 ) ;
  assign n9974 = ( n9698 & ~n9972 ) | ( n9698 & n9973 ) | ( ~n9972 & n9973 ) ;
  assign n9975 = n1097 & n5374 ;
  assign n9976 = x83 & n5378 ;
  assign n9977 = x84 | n9976 ;
  assign n9978 = ( n5380 & n9976 ) | ( n5380 & n9977 ) | ( n9976 & n9977 ) ;
  assign n9979 = x82 & n5638 ;
  assign n9980 = n9978 | n9979 ;
  assign n9981 = ( x50 & n9975 ) | ( x50 & ~n9980 ) | ( n9975 & ~n9980 ) ;
  assign n9982 = ( ~x50 & n9980 ) | ( ~x50 & n9981 ) | ( n9980 & n9981 ) ;
  assign n9983 = ( ~n9975 & n9981 ) | ( ~n9975 & n9982 ) | ( n9981 & n9982 ) ;
  assign n9984 = ( n9710 & n9974 ) | ( n9710 & n9983 ) | ( n9974 & n9983 ) ;
  assign n9985 = ( ~n9710 & n9974 ) | ( ~n9710 & n9983 ) | ( n9974 & n9983 ) ;
  assign n9986 = ( n9710 & ~n9984 ) | ( n9710 & n9985 ) | ( ~n9984 & n9985 ) ;
  assign n9987 = n1466 & n4787 ;
  assign n9988 = x86 & n4791 ;
  assign n9989 = x87 | n9988 ;
  assign n9990 = ( n4793 & n9988 ) | ( n4793 & n9989 ) | ( n9988 & n9989 ) ;
  assign n9991 = x85 & n5030 ;
  assign n9992 = n9990 | n9991 ;
  assign n9993 = ( x47 & n9987 ) | ( x47 & ~n9992 ) | ( n9987 & ~n9992 ) ;
  assign n9994 = ( ~x47 & n9992 ) | ( ~x47 & n9993 ) | ( n9992 & n9993 ) ;
  assign n9995 = ( ~n9987 & n9993 ) | ( ~n9987 & n9994 ) | ( n9993 & n9994 ) ;
  assign n9996 = ( n9722 & n9986 ) | ( n9722 & n9995 ) | ( n9986 & n9995 ) ;
  assign n9997 = ( n9722 & ~n9986 ) | ( n9722 & n9995 ) | ( ~n9986 & n9995 ) ;
  assign n9998 = ( n9986 & ~n9996 ) | ( n9986 & n9997 ) | ( ~n9996 & n9997 ) ;
  assign n9999 = n1701 & n4227 ;
  assign n10000 = x89 & n4231 ;
  assign n10001 = x90 | n10000 ;
  assign n10002 = ( n4233 & n10000 ) | ( n4233 & n10001 ) | ( n10000 & n10001 ) ;
  assign n10003 = x88 & n4470 ;
  assign n10004 = n10002 | n10003 ;
  assign n10005 = ( x44 & n9999 ) | ( x44 & ~n10004 ) | ( n9999 & ~n10004 ) ;
  assign n10006 = ( ~x44 & n10004 ) | ( ~x44 & n10005 ) | ( n10004 & n10005 ) ;
  assign n10007 = ( ~n9999 & n10005 ) | ( ~n9999 & n10006 ) | ( n10005 & n10006 ) ;
  assign n10008 = ( n9734 & n9998 ) | ( n9734 & n10007 ) | ( n9998 & n10007 ) ;
  assign n10009 = ( ~n9734 & n9998 ) | ( ~n9734 & n10007 ) | ( n9998 & n10007 ) ;
  assign n10010 = ( n9734 & ~n10008 ) | ( n9734 & n10009 ) | ( ~n10008 & n10009 ) ;
  assign n10011 = n2057 & n3715 ;
  assign n10012 = x92 & n3719 ;
  assign n10013 = x93 | n10012 ;
  assign n10014 = ( n3721 & n10012 ) | ( n3721 & n10013 ) | ( n10012 & n10013 ) ;
  assign n10015 = x91 & n3922 ;
  assign n10016 = n10014 | n10015 ;
  assign n10017 = ( x41 & n10011 ) | ( x41 & ~n10016 ) | ( n10011 & ~n10016 ) ;
  assign n10018 = ( ~x41 & n10016 ) | ( ~x41 & n10017 ) | ( n10016 & n10017 ) ;
  assign n10019 = ( ~n10011 & n10017 ) | ( ~n10011 & n10018 ) | ( n10017 & n10018 ) ;
  assign n10020 = ( n9746 & n10010 ) | ( n9746 & n10019 ) | ( n10010 & n10019 ) ;
  assign n10021 = ( ~n9746 & n10010 ) | ( ~n9746 & n10019 ) | ( n10010 & n10019 ) ;
  assign n10022 = ( n9746 & ~n10020 ) | ( n9746 & n10021 ) | ( ~n10020 & n10021 ) ;
  assign n10023 = n2449 & n3224 ;
  assign n10024 = x95 & n3228 ;
  assign n10025 = x96 | n10024 ;
  assign n10026 = ( n3230 & n10024 ) | ( n3230 & n10025 ) | ( n10024 & n10025 ) ;
  assign n10027 = x94 & n3413 ;
  assign n10028 = n10026 | n10027 ;
  assign n10029 = ( x38 & n10023 ) | ( x38 & ~n10028 ) | ( n10023 & ~n10028 ) ;
  assign n10030 = ( ~x38 & n10028 ) | ( ~x38 & n10029 ) | ( n10028 & n10029 ) ;
  assign n10031 = ( ~n10023 & n10029 ) | ( ~n10023 & n10030 ) | ( n10029 & n10030 ) ;
  assign n10032 = ( n9758 & n10022 ) | ( n9758 & n10031 ) | ( n10022 & n10031 ) ;
  assign n10033 = ( ~n9758 & n10022 ) | ( ~n9758 & n10031 ) | ( n10022 & n10031 ) ;
  assign n10034 = ( n9758 & ~n10032 ) | ( n9758 & n10033 ) | ( ~n10032 & n10033 ) ;
  assign n10035 = n2766 & n2877 ;
  assign n10036 = x98 & n2770 ;
  assign n10037 = x99 | n10036 ;
  assign n10038 = ( n2772 & n10036 ) | ( n2772 & n10037 ) | ( n10036 & n10037 ) ;
  assign n10039 = x97 & n2943 ;
  assign n10040 = n10038 | n10039 ;
  assign n10041 = ( x35 & n10035 ) | ( x35 & ~n10040 ) | ( n10035 & ~n10040 ) ;
  assign n10042 = ( ~x35 & n10040 ) | ( ~x35 & n10041 ) | ( n10040 & n10041 ) ;
  assign n10043 = ( ~n10035 & n10041 ) | ( ~n10035 & n10042 ) | ( n10041 & n10042 ) ;
  assign n10044 = ( n9770 & n10034 ) | ( n9770 & n10043 ) | ( n10034 & n10043 ) ;
  assign n10045 = ( n9770 & ~n10034 ) | ( n9770 & n10043 ) | ( ~n10034 & n10043 ) ;
  assign n10046 = ( n10034 & ~n10044 ) | ( n10034 & n10045 ) | ( ~n10044 & n10045 ) ;
  assign n10047 = ( n9773 & n9923 ) | ( n9773 & n10046 ) | ( n9923 & n10046 ) ;
  assign n10048 = ( ~n9773 & n9923 ) | ( ~n9773 & n10046 ) | ( n9923 & n10046 ) ;
  assign n10049 = ( n9773 & ~n10047 ) | ( n9773 & n10048 ) | ( ~n10047 & n10048 ) ;
  assign n10050 = ( n9776 & n9914 ) | ( n9776 & n10049 ) | ( n9914 & n10049 ) ;
  assign n10051 = ( n9776 & ~n9914 ) | ( n9776 & n10049 ) | ( ~n9914 & n10049 ) ;
  assign n10052 = ( n9914 & ~n10050 ) | ( n9914 & n10051 ) | ( ~n10050 & n10051 ) ;
  assign n10053 = n1617 & n4377 ;
  assign n10054 = x107 & n1621 ;
  assign n10055 = x108 | n10054 ;
  assign n10056 = ( n1623 & n10054 ) | ( n1623 & n10055 ) | ( n10054 & n10055 ) ;
  assign n10057 = x106 & n1749 ;
  assign n10058 = n10056 | n10057 ;
  assign n10059 = ( x26 & n10053 ) | ( x26 & ~n10058 ) | ( n10053 & ~n10058 ) ;
  assign n10060 = ( ~x26 & n10058 ) | ( ~x26 & n10059 ) | ( n10058 & n10059 ) ;
  assign n10061 = ( ~n10053 & n10059 ) | ( ~n10053 & n10060 ) | ( n10059 & n10060 ) ;
  assign n10062 = ( n9788 & n10052 ) | ( n9788 & n10061 ) | ( n10052 & n10061 ) ;
  assign n10063 = ( n9788 & ~n10052 ) | ( n9788 & n10061 ) | ( ~n10052 & n10061 ) ;
  assign n10064 = ( n10052 & ~n10062 ) | ( n10052 & n10063 ) | ( ~n10062 & n10063 ) ;
  assign n10065 = ( n9791 & n9905 ) | ( n9791 & n10064 ) | ( n9905 & n10064 ) ;
  assign n10066 = ( n9791 & ~n9905 ) | ( n9791 & n10064 ) | ( ~n9905 & n10064 ) ;
  assign n10067 = ( n9905 & ~n10065 ) | ( n9905 & n10066 ) | ( ~n10065 & n10066 ) ;
  assign n10068 = ( n9803 & n9896 ) | ( n9803 & n10067 ) | ( n9896 & n10067 ) ;
  assign n10069 = ( n9803 & ~n9896 ) | ( n9803 & n10067 ) | ( ~n9896 & n10067 ) ;
  assign n10070 = ( n9896 & ~n10068 ) | ( n9896 & n10069 ) | ( ~n10068 & n10069 ) ;
  assign n10071 = ( n9806 & n9887 ) | ( n9806 & n10070 ) | ( n9887 & n10070 ) ;
  assign n10072 = ( ~n9806 & n9887 ) | ( ~n9806 & n10070 ) | ( n9887 & n10070 ) ;
  assign n10073 = ( n9806 & ~n10071 ) | ( n9806 & n10072 ) | ( ~n10071 & n10072 ) ;
  assign n10074 = ( n9818 & n9878 ) | ( n9818 & n10073 ) | ( n9878 & n10073 ) ;
  assign n10075 = ( n9818 & ~n9878 ) | ( n9818 & n10073 ) | ( ~n9878 & n10073 ) ;
  assign n10076 = ( n9878 & ~n10074 ) | ( n9878 & n10075 ) | ( ~n10074 & n10075 ) ;
  assign n10077 = ( n9821 & n9869 ) | ( n9821 & n10076 ) | ( n9869 & n10076 ) ;
  assign n10078 = ( n9821 & ~n9869 ) | ( n9821 & n10076 ) | ( ~n9869 & n10076 ) ;
  assign n10079 = ( n9869 & ~n10077 ) | ( n9869 & n10078 ) | ( ~n10077 & n10078 ) ;
  assign n10080 = n291 & n8587 ;
  assign n10081 = x125 & n295 ;
  assign n10082 = x126 | n10081 ;
  assign n10083 = ( n297 & n10081 ) | ( n297 & n10082 ) | ( n10081 & n10082 ) ;
  assign n10084 = x124 & n330 ;
  assign n10085 = n10083 | n10084 ;
  assign n10086 = ( x8 & n10080 ) | ( x8 & ~n10085 ) | ( n10080 & ~n10085 ) ;
  assign n10087 = ( ~x8 & n10085 ) | ( ~x8 & n10086 ) | ( n10085 & n10086 ) ;
  assign n10088 = ( ~n10080 & n10086 ) | ( ~n10080 & n10087 ) | ( n10086 & n10087 ) ;
  assign n10089 = ( n9833 & n10079 ) | ( n9833 & n10088 ) | ( n10079 & n10088 ) ;
  assign n10090 = ( n9833 & ~n10079 ) | ( n9833 & n10088 ) | ( ~n10079 & n10088 ) ;
  assign n10091 = ( n10079 & ~n10089 ) | ( n10079 & n10090 ) | ( ~n10089 & n10090 ) ;
  assign n10092 = n186 & n8862 ;
  assign n10093 = ( x127 & n220 ) | ( x127 & n10092 ) | ( n220 & n10092 ) ;
  assign n10094 = x5 | n10093 ;
  assign n10095 = ~x5 & n10093 ;
  assign n10096 = ( ~n10093 & n10094 ) | ( ~n10093 & n10095 ) | ( n10094 & n10095 ) ;
  assign n10097 = ( n9845 & n10091 ) | ( n9845 & n10096 ) | ( n10091 & n10096 ) ;
  assign n10098 = ( n9845 & ~n10091 ) | ( n9845 & n10096 ) | ( ~n10091 & n10096 ) ;
  assign n10099 = ( n10091 & ~n10097 ) | ( n10091 & n10098 ) | ( ~n10097 & n10098 ) ;
  assign n10100 = ( n9855 & n9858 ) | ( n9855 & n10099 ) | ( n9858 & n10099 ) ;
  assign n10101 = ( n9855 & ~n9858 ) | ( n9855 & n10099 ) | ( ~n9858 & n10099 ) ;
  assign n10102 = ( n9858 & ~n10100 ) | ( n9858 & n10101 ) | ( ~n10100 & n10101 ) ;
  assign n10103 = n407 & n7841 ;
  assign n10104 = x123 & n411 ;
  assign n10105 = x124 | n10104 ;
  assign n10106 = ( n413 & n10104 ) | ( n413 & n10105 ) | ( n10104 & n10105 ) ;
  assign n10107 = x122 & n491 ;
  assign n10108 = n10106 | n10107 ;
  assign n10109 = ( x11 & n10103 ) | ( x11 & ~n10108 ) | ( n10103 & ~n10108 ) ;
  assign n10110 = ( ~x11 & n10108 ) | ( ~x11 & n10109 ) | ( n10108 & n10109 ) ;
  assign n10111 = ( ~n10103 & n10109 ) | ( ~n10103 & n10110 ) | ( n10109 & n10110 ) ;
  assign n10112 = n1016 & n5765 ;
  assign n10113 = x114 & n1020 ;
  assign n10114 = x115 | n10113 ;
  assign n10115 = ( n1022 & n10113 ) | ( n1022 & n10114 ) | ( n10113 & n10114 ) ;
  assign n10116 = x113 & n1145 ;
  assign n10117 = n10115 | n10116 ;
  assign n10118 = ( x20 & n10112 ) | ( x20 & ~n10117 ) | ( n10112 & ~n10117 ) ;
  assign n10119 = ( ~x20 & n10117 ) | ( ~x20 & n10118 ) | ( n10117 & n10118 ) ;
  assign n10120 = ( ~n10112 & n10118 ) | ( ~n10112 & n10119 ) | ( n10118 & n10119 ) ;
  assign n10121 = n1297 & n5145 ;
  assign n10122 = x111 & n1301 ;
  assign n10123 = x112 | n10122 ;
  assign n10124 = ( n1303 & n10122 ) | ( n1303 & n10123 ) | ( n10122 & n10123 ) ;
  assign n10125 = x110 & n1426 ;
  assign n10126 = n10124 | n10125 ;
  assign n10127 = ( x23 & n10121 ) | ( x23 & ~n10126 ) | ( n10121 & ~n10126 ) ;
  assign n10128 = ( ~x23 & n10126 ) | ( ~x23 & n10127 ) | ( n10126 & n10127 ) ;
  assign n10129 = ( ~n10121 & n10127 ) | ( ~n10121 & n10128 ) | ( n10127 & n10128 ) ;
  assign n10130 = n1949 & n4013 ;
  assign n10131 = x105 & n1953 ;
  assign n10132 = x106 | n10131 ;
  assign n10133 = ( n1955 & n10131 ) | ( n1955 & n10132 ) | ( n10131 & n10132 ) ;
  assign n10134 = x104 & n2114 ;
  assign n10135 = n10133 | n10134 ;
  assign n10136 = ( x29 & n10130 ) | ( x29 & ~n10135 ) | ( n10130 & ~n10135 ) ;
  assign n10137 = ( ~x29 & n10135 ) | ( ~x29 & n10136 ) | ( n10135 & n10136 ) ;
  assign n10138 = ( ~n10130 & n10136 ) | ( ~n10130 & n10137 ) | ( n10136 & n10137 ) ;
  assign n10139 = n2766 & n3162 ;
  assign n10140 = x99 & n2770 ;
  assign n10141 = x100 | n10140 ;
  assign n10142 = ( n2772 & n10140 ) | ( n2772 & n10141 ) | ( n10140 & n10141 ) ;
  assign n10143 = x98 & n2943 ;
  assign n10144 = n10142 | n10143 ;
  assign n10145 = ( x35 & n10139 ) | ( x35 & ~n10144 ) | ( n10139 & ~n10144 ) ;
  assign n10146 = ( ~x35 & n10144 ) | ( ~x35 & n10145 ) | ( n10144 & n10145 ) ;
  assign n10147 = ( ~n10139 & n10145 ) | ( ~n10139 & n10146 ) | ( n10145 & n10146 ) ;
  assign n10148 = n2585 & n3224 ;
  assign n10149 = x96 & n3228 ;
  assign n10150 = x97 | n10149 ;
  assign n10151 = ( n3230 & n10149 ) | ( n3230 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10152 = x95 & n3413 ;
  assign n10153 = n10151 | n10152 ;
  assign n10154 = ( x38 & n10148 ) | ( x38 & ~n10153 ) | ( n10148 & ~n10153 ) ;
  assign n10155 = ( ~x38 & n10153 ) | ( ~x38 & n10154 ) | ( n10153 & n10154 ) ;
  assign n10156 = ( ~n10148 & n10154 ) | ( ~n10148 & n10155 ) | ( n10154 & n10155 ) ;
  assign n10157 = n1481 & n4787 ;
  assign n10158 = x87 & n4791 ;
  assign n10159 = x88 | n10158 ;
  assign n10160 = ( n4793 & n10158 ) | ( n4793 & n10159 ) | ( n10158 & n10159 ) ;
  assign n10161 = x86 & n5030 ;
  assign n10162 = n10160 | n10161 ;
  assign n10163 = ( x47 & n10157 ) | ( x47 & ~n10162 ) | ( n10157 & ~n10162 ) ;
  assign n10164 = ( ~x47 & n10162 ) | ( ~x47 & n10163 ) | ( n10162 & n10163 ) ;
  assign n10165 = ( ~n10157 & n10163 ) | ( ~n10157 & n10164 ) | ( n10163 & n10164 ) ;
  assign n10166 = n554 & n7423 ;
  assign n10167 = x75 & n7427 ;
  assign n10168 = x76 | n10167 ;
  assign n10169 = ( n7429 & n10167 ) | ( n7429 & n10168 ) | ( n10167 & n10168 ) ;
  assign n10170 = x74 & n7708 ;
  assign n10171 = n10169 | n10170 ;
  assign n10172 = ( x59 & n10166 ) | ( x59 & ~n10171 ) | ( n10166 & ~n10171 ) ;
  assign n10173 = ( ~x59 & n10171 ) | ( ~x59 & n10172 ) | ( n10171 & n10172 ) ;
  assign n10174 = ( ~n10166 & n10172 ) | ( ~n10166 & n10173 ) | ( n10172 & n10173 ) ;
  assign n10175 = x69 & n8927 ;
  assign n10176 = ( ~x70 & n8693 ) | ( ~x70 & n8927 ) | ( n8693 & n8927 ) ;
  assign n10177 = ( n8693 & n10175 ) | ( n8693 & ~n10176 ) | ( n10175 & ~n10176 ) ;
  assign n10178 = ( x2 & x5 ) | ( x2 & ~n10177 ) | ( x5 & ~n10177 ) ;
  assign n10179 = ( x2 & ~x5 ) | ( x2 & n10177 ) | ( ~x5 & n10177 ) ;
  assign n10180 = ( ~x2 & n10178 ) | ( ~x2 & n10179 ) | ( n10178 & n10179 ) ;
  assign n10181 = n390 & n8154 ;
  assign n10182 = x72 & n8158 ;
  assign n10183 = x73 | n10182 ;
  assign n10184 = ( n8160 & n10182 ) | ( n8160 & n10183 ) | ( n10182 & n10183 ) ;
  assign n10185 = x71 & n8439 ;
  assign n10186 = n10184 | n10185 ;
  assign n10187 = ( x62 & n10181 ) | ( x62 & ~n10186 ) | ( n10181 & ~n10186 ) ;
  assign n10188 = ( ~x62 & n10186 ) | ( ~x62 & n10187 ) | ( n10186 & n10187 ) ;
  assign n10189 = ( ~n10181 & n10187 ) | ( ~n10181 & n10188 ) | ( n10187 & n10188 ) ;
  assign n10190 = ( n9936 & n10180 ) | ( n9936 & n10189 ) | ( n10180 & n10189 ) ;
  assign n10191 = ( ~n9936 & n10180 ) | ( ~n9936 & n10189 ) | ( n10180 & n10189 ) ;
  assign n10192 = ( n9936 & ~n10190 ) | ( n9936 & n10191 ) | ( ~n10190 & n10191 ) ;
  assign n10193 = ( n9948 & n10174 ) | ( n9948 & n10192 ) | ( n10174 & n10192 ) ;
  assign n10194 = ( ~n9948 & n10174 ) | ( ~n9948 & n10192 ) | ( n10174 & n10192 ) ;
  assign n10195 = ( n9948 & ~n10193 ) | ( n9948 & n10194 ) | ( ~n10193 & n10194 ) ;
  assign n10196 = n701 & n6713 ;
  assign n10197 = x78 & n6717 ;
  assign n10198 = x79 | n10197 ;
  assign n10199 = ( n6719 & n10197 ) | ( n6719 & n10198 ) | ( n10197 & n10198 ) ;
  assign n10200 = x77 & n6980 ;
  assign n10201 = n10199 | n10200 ;
  assign n10202 = ( x56 & n10196 ) | ( x56 & ~n10201 ) | ( n10196 & ~n10201 ) ;
  assign n10203 = ( ~x56 & n10201 ) | ( ~x56 & n10202 ) | ( n10201 & n10202 ) ;
  assign n10204 = ( ~n10196 & n10202 ) | ( ~n10196 & n10203 ) | ( n10202 & n10203 ) ;
  assign n10205 = ( n9960 & n10195 ) | ( n9960 & n10204 ) | ( n10195 & n10204 ) ;
  assign n10206 = ( ~n9960 & n10195 ) | ( ~n9960 & n10204 ) | ( n10195 & n10204 ) ;
  assign n10207 = ( n9960 & ~n10205 ) | ( n9960 & n10206 ) | ( ~n10205 & n10206 ) ;
  assign n10208 = n990 & n6027 ;
  assign n10209 = x81 & n6031 ;
  assign n10210 = x82 | n10209 ;
  assign n10211 = ( n6033 & n10209 ) | ( n6033 & n10210 ) | ( n10209 & n10210 ) ;
  assign n10212 = x80 & n6303 ;
  assign n10213 = n10211 | n10212 ;
  assign n10214 = ( x53 & n10208 ) | ( x53 & ~n10213 ) | ( n10208 & ~n10213 ) ;
  assign n10215 = ( ~x53 & n10213 ) | ( ~x53 & n10214 ) | ( n10213 & n10214 ) ;
  assign n10216 = ( ~n10208 & n10214 ) | ( ~n10208 & n10215 ) | ( n10214 & n10215 ) ;
  assign n10217 = ( n9972 & n10207 ) | ( n9972 & n10216 ) | ( n10207 & n10216 ) ;
  assign n10218 = ( ~n9972 & n10207 ) | ( ~n9972 & n10216 ) | ( n10207 & n10216 ) ;
  assign n10219 = ( n9972 & ~n10217 ) | ( n9972 & n10218 ) | ( ~n10217 & n10218 ) ;
  assign n10220 = n1262 & n5374 ;
  assign n10221 = x84 & n5378 ;
  assign n10222 = x85 | n10221 ;
  assign n10223 = ( n5380 & n10221 ) | ( n5380 & n10222 ) | ( n10221 & n10222 ) ;
  assign n10224 = x83 & n5638 ;
  assign n10225 = n10223 | n10224 ;
  assign n10226 = ( x50 & n10220 ) | ( x50 & ~n10225 ) | ( n10220 & ~n10225 ) ;
  assign n10227 = ( ~x50 & n10225 ) | ( ~x50 & n10226 ) | ( n10225 & n10226 ) ;
  assign n10228 = ( ~n10220 & n10226 ) | ( ~n10220 & n10227 ) | ( n10226 & n10227 ) ;
  assign n10229 = ( n9984 & n10219 ) | ( n9984 & n10228 ) | ( n10219 & n10228 ) ;
  assign n10230 = ( ~n9984 & n10219 ) | ( ~n9984 & n10228 ) | ( n10219 & n10228 ) ;
  assign n10231 = ( n9984 & ~n10229 ) | ( n9984 & n10230 ) | ( ~n10229 & n10230 ) ;
  assign n10232 = ( n9996 & n10165 ) | ( n9996 & n10231 ) | ( n10165 & n10231 ) ;
  assign n10233 = ( ~n9996 & n10165 ) | ( ~n9996 & n10231 ) | ( n10165 & n10231 ) ;
  assign n10234 = ( n9996 & ~n10232 ) | ( n9996 & n10233 ) | ( ~n10232 & n10233 ) ;
  assign n10235 = n1914 & n4227 ;
  assign n10236 = x90 & n4231 ;
  assign n10237 = x91 | n10236 ;
  assign n10238 = ( n4233 & n10236 ) | ( n4233 & n10237 ) | ( n10236 & n10237 ) ;
  assign n10239 = x89 & n4470 ;
  assign n10240 = n10238 | n10239 ;
  assign n10241 = ( x44 & n10235 ) | ( x44 & ~n10240 ) | ( n10235 & ~n10240 ) ;
  assign n10242 = ( ~x44 & n10240 ) | ( ~x44 & n10241 ) | ( n10240 & n10241 ) ;
  assign n10243 = ( ~n10235 & n10241 ) | ( ~n10235 & n10242 ) | ( n10241 & n10242 ) ;
  assign n10244 = ( n10008 & n10234 ) | ( n10008 & n10243 ) | ( n10234 & n10243 ) ;
  assign n10245 = ( ~n10008 & n10234 ) | ( ~n10008 & n10243 ) | ( n10234 & n10243 ) ;
  assign n10246 = ( n10008 & ~n10244 ) | ( n10008 & n10245 ) | ( ~n10244 & n10245 ) ;
  assign n10247 = n2294 & n3715 ;
  assign n10248 = x93 & n3719 ;
  assign n10249 = x94 | n10248 ;
  assign n10250 = ( n3721 & n10248 ) | ( n3721 & n10249 ) | ( n10248 & n10249 ) ;
  assign n10251 = x92 & n3922 ;
  assign n10252 = n10250 | n10251 ;
  assign n10253 = ( x41 & n10247 ) | ( x41 & ~n10252 ) | ( n10247 & ~n10252 ) ;
  assign n10254 = ( ~x41 & n10252 ) | ( ~x41 & n10253 ) | ( n10252 & n10253 ) ;
  assign n10255 = ( ~n10247 & n10253 ) | ( ~n10247 & n10254 ) | ( n10253 & n10254 ) ;
  assign n10256 = ( n10020 & n10246 ) | ( n10020 & n10255 ) | ( n10246 & n10255 ) ;
  assign n10257 = ( ~n10020 & n10246 ) | ( ~n10020 & n10255 ) | ( n10246 & n10255 ) ;
  assign n10258 = ( n10020 & ~n10256 ) | ( n10020 & n10257 ) | ( ~n10256 & n10257 ) ;
  assign n10259 = ( n10032 & n10156 ) | ( n10032 & n10258 ) | ( n10156 & n10258 ) ;
  assign n10260 = ( ~n10032 & n10156 ) | ( ~n10032 & n10258 ) | ( n10156 & n10258 ) ;
  assign n10261 = ( n10032 & ~n10259 ) | ( n10032 & n10260 ) | ( ~n10259 & n10260 ) ;
  assign n10262 = ( n10044 & n10147 ) | ( n10044 & n10261 ) | ( n10147 & n10261 ) ;
  assign n10263 = ( ~n10044 & n10147 ) | ( ~n10044 & n10261 ) | ( n10147 & n10261 ) ;
  assign n10264 = ( n10044 & ~n10262 ) | ( n10044 & n10263 ) | ( ~n10262 & n10263 ) ;
  assign n10265 = n2320 & n3650 ;
  assign n10266 = x102 & n2324 ;
  assign n10267 = x103 | n10266 ;
  assign n10268 = ( n2326 & n10266 ) | ( n2326 & n10267 ) | ( n10266 & n10267 ) ;
  assign n10269 = x101 & n2497 ;
  assign n10270 = n10268 | n10269 ;
  assign n10271 = ( x32 & n10265 ) | ( x32 & ~n10270 ) | ( n10265 & ~n10270 ) ;
  assign n10272 = ( ~x32 & n10270 ) | ( ~x32 & n10271 ) | ( n10270 & n10271 ) ;
  assign n10273 = ( ~n10265 & n10271 ) | ( ~n10265 & n10272 ) | ( n10271 & n10272 ) ;
  assign n10274 = ( n10047 & n10264 ) | ( n10047 & n10273 ) | ( n10264 & n10273 ) ;
  assign n10275 = ( n10047 & ~n10264 ) | ( n10047 & n10273 ) | ( ~n10264 & n10273 ) ;
  assign n10276 = ( n10264 & ~n10274 ) | ( n10264 & n10275 ) | ( ~n10274 & n10275 ) ;
  assign n10277 = ( n10050 & n10138 ) | ( n10050 & n10276 ) | ( n10138 & n10276 ) ;
  assign n10278 = ( n10050 & ~n10138 ) | ( n10050 & n10276 ) | ( ~n10138 & n10276 ) ;
  assign n10279 = ( n10138 & ~n10277 ) | ( n10138 & n10278 ) | ( ~n10277 & n10278 ) ;
  assign n10280 = n1617 & n4734 ;
  assign n10281 = x108 & n1621 ;
  assign n10282 = x109 | n10281 ;
  assign n10283 = ( n1623 & n10281 ) | ( n1623 & n10282 ) | ( n10281 & n10282 ) ;
  assign n10284 = x107 & n1749 ;
  assign n10285 = n10283 | n10284 ;
  assign n10286 = ( x26 & n10280 ) | ( x26 & ~n10285 ) | ( n10280 & ~n10285 ) ;
  assign n10287 = ( ~x26 & n10285 ) | ( ~x26 & n10286 ) | ( n10285 & n10286 ) ;
  assign n10288 = ( ~n10280 & n10286 ) | ( ~n10280 & n10287 ) | ( n10286 & n10287 ) ;
  assign n10289 = ( n10062 & n10279 ) | ( n10062 & n10288 ) | ( n10279 & n10288 ) ;
  assign n10290 = ( n10062 & ~n10279 ) | ( n10062 & n10288 ) | ( ~n10279 & n10288 ) ;
  assign n10291 = ( n10279 & ~n10289 ) | ( n10279 & n10290 ) | ( ~n10289 & n10290 ) ;
  assign n10292 = ( n10065 & n10129 ) | ( n10065 & n10291 ) | ( n10129 & n10291 ) ;
  assign n10293 = ( n10065 & ~n10129 ) | ( n10065 & n10291 ) | ( ~n10129 & n10291 ) ;
  assign n10294 = ( n10129 & ~n10292 ) | ( n10129 & n10293 ) | ( ~n10292 & n10293 ) ;
  assign n10295 = ( n10068 & n10120 ) | ( n10068 & n10294 ) | ( n10120 & n10294 ) ;
  assign n10296 = ( n10068 & ~n10120 ) | ( n10068 & n10294 ) | ( ~n10120 & n10294 ) ;
  assign n10297 = ( n10120 & ~n10295 ) | ( n10120 & n10296 ) | ( ~n10295 & n10296 ) ;
  assign n10298 = n810 & n6421 ;
  assign n10299 = x117 & n814 ;
  assign n10300 = x118 | n10299 ;
  assign n10301 = ( n816 & n10299 ) | ( n816 & n10300 ) | ( n10299 & n10300 ) ;
  assign n10302 = x116 & n885 ;
  assign n10303 = n10301 | n10302 ;
  assign n10304 = ( x17 & n10298 ) | ( x17 & ~n10303 ) | ( n10298 & ~n10303 ) ;
  assign n10305 = ( ~x17 & n10303 ) | ( ~x17 & n10304 ) | ( n10303 & n10304 ) ;
  assign n10306 = ( ~n10298 & n10304 ) | ( ~n10298 & n10305 ) | ( n10304 & n10305 ) ;
  assign n10307 = ( n10071 & n10297 ) | ( n10071 & n10306 ) | ( n10297 & n10306 ) ;
  assign n10308 = ( n10071 & ~n10297 ) | ( n10071 & n10306 ) | ( ~n10297 & n10306 ) ;
  assign n10309 = ( n10297 & ~n10307 ) | ( n10297 & n10308 ) | ( ~n10307 & n10308 ) ;
  assign n10310 = n583 & n7113 ;
  assign n10311 = x120 & n587 ;
  assign n10312 = x121 | n10311 ;
  assign n10313 = ( n589 & n10311 ) | ( n589 & n10312 ) | ( n10311 & n10312 ) ;
  assign n10314 = x119 & n676 ;
  assign n10315 = n10313 | n10314 ;
  assign n10316 = ( x14 & n10310 ) | ( x14 & ~n10315 ) | ( n10310 & ~n10315 ) ;
  assign n10317 = ( ~x14 & n10315 ) | ( ~x14 & n10316 ) | ( n10315 & n10316 ) ;
  assign n10318 = ( ~n10310 & n10316 ) | ( ~n10310 & n10317 ) | ( n10316 & n10317 ) ;
  assign n10319 = ( n10074 & n10309 ) | ( n10074 & n10318 ) | ( n10309 & n10318 ) ;
  assign n10320 = ( n10074 & ~n10309 ) | ( n10074 & n10318 ) | ( ~n10309 & n10318 ) ;
  assign n10321 = ( n10309 & ~n10319 ) | ( n10309 & n10320 ) | ( ~n10319 & n10320 ) ;
  assign n10322 = ( n10077 & n10111 ) | ( n10077 & n10321 ) | ( n10111 & n10321 ) ;
  assign n10323 = ( n10077 & ~n10111 ) | ( n10077 & n10321 ) | ( ~n10111 & n10321 ) ;
  assign n10324 = ( n10111 & ~n10322 ) | ( n10111 & n10323 ) | ( ~n10322 & n10323 ) ;
  assign n10325 = n291 & n8846 ;
  assign n10326 = x126 & n295 ;
  assign n10327 = x127 | n10326 ;
  assign n10328 = ( n297 & n10326 ) | ( n297 & n10327 ) | ( n10326 & n10327 ) ;
  assign n10329 = x125 & n330 ;
  assign n10330 = n10328 | n10329 ;
  assign n10331 = ( x8 & n10325 ) | ( x8 & ~n10330 ) | ( n10325 & ~n10330 ) ;
  assign n10332 = ( ~x8 & n10330 ) | ( ~x8 & n10331 ) | ( n10330 & n10331 ) ;
  assign n10333 = ( ~n10325 & n10331 ) | ( ~n10325 & n10332 ) | ( n10331 & n10332 ) ;
  assign n10334 = ( n10089 & n10324 ) | ( n10089 & n10333 ) | ( n10324 & n10333 ) ;
  assign n10335 = ( n10089 & ~n10324 ) | ( n10089 & n10333 ) | ( ~n10324 & n10333 ) ;
  assign n10336 = ( n10324 & ~n10334 ) | ( n10324 & n10335 ) | ( ~n10334 & n10335 ) ;
  assign n10337 = ( n10097 & n10100 ) | ( n10097 & n10336 ) | ( n10100 & n10336 ) ;
  assign n10338 = ( n10097 & ~n10100 ) | ( n10097 & n10336 ) | ( ~n10100 & n10336 ) ;
  assign n10339 = ( n10100 & ~n10337 ) | ( n10100 & n10338 ) | ( ~n10337 & n10338 ) ;
  assign n10340 = n291 & n8865 ;
  assign n10341 = x127 & n295 ;
  assign n10342 = x126 | n10341 ;
  assign n10343 = ( n330 & n10341 ) | ( n330 & n10342 ) | ( n10341 & n10342 ) ;
  assign n10344 = ( x8 & n10340 ) | ( x8 & ~n10343 ) | ( n10340 & ~n10343 ) ;
  assign n10345 = ( ~x8 & n10343 ) | ( ~x8 & n10344 ) | ( n10343 & n10344 ) ;
  assign n10346 = ( ~n10340 & n10344 ) | ( ~n10340 & n10345 ) | ( n10344 & n10345 ) ;
  assign n10347 = n407 & n8331 ;
  assign n10348 = x124 & n411 ;
  assign n10349 = x125 | n10348 ;
  assign n10350 = ( n413 & n10348 ) | ( n413 & n10349 ) | ( n10348 & n10349 ) ;
  assign n10351 = x123 & n491 ;
  assign n10352 = n10350 | n10351 ;
  assign n10353 = ( x11 & n10347 ) | ( x11 & ~n10352 ) | ( n10347 & ~n10352 ) ;
  assign n10354 = ( ~x11 & n10352 ) | ( ~x11 & n10353 ) | ( n10352 & n10353 ) ;
  assign n10355 = ( ~n10347 & n10353 ) | ( ~n10347 & n10354 ) | ( n10353 & n10354 ) ;
  assign n10356 = n583 & n7582 ;
  assign n10357 = x121 & n587 ;
  assign n10358 = x122 | n10357 ;
  assign n10359 = ( n589 & n10357 ) | ( n589 & n10358 ) | ( n10357 & n10358 ) ;
  assign n10360 = x120 & n676 ;
  assign n10361 = n10359 | n10360 ;
  assign n10362 = ( x14 & n10356 ) | ( x14 & ~n10361 ) | ( n10356 & ~n10361 ) ;
  assign n10363 = ( ~x14 & n10361 ) | ( ~x14 & n10362 ) | ( n10361 & n10362 ) ;
  assign n10364 = ( ~n10356 & n10362 ) | ( ~n10356 & n10363 ) | ( n10362 & n10363 ) ;
  assign n10365 = n810 & n6645 ;
  assign n10366 = x118 & n814 ;
  assign n10367 = x119 | n10366 ;
  assign n10368 = ( n816 & n10366 ) | ( n816 & n10367 ) | ( n10366 & n10367 ) ;
  assign n10369 = x117 & n885 ;
  assign n10370 = n10368 | n10369 ;
  assign n10371 = ( x17 & n10365 ) | ( x17 & ~n10370 ) | ( n10365 & ~n10370 ) ;
  assign n10372 = ( ~x17 & n10370 ) | ( ~x17 & n10371 ) | ( n10370 & n10371 ) ;
  assign n10373 = ( ~n10365 & n10371 ) | ( ~n10365 & n10372 ) | ( n10371 & n10372 ) ;
  assign n10374 = n1016 & n5977 ;
  assign n10375 = x115 & n1020 ;
  assign n10376 = x116 | n10375 ;
  assign n10377 = ( n1022 & n10375 ) | ( n1022 & n10376 ) | ( n10375 & n10376 ) ;
  assign n10378 = x114 & n1145 ;
  assign n10379 = n10377 | n10378 ;
  assign n10380 = ( x20 & n10374 ) | ( x20 & ~n10379 ) | ( n10374 & ~n10379 ) ;
  assign n10381 = ( ~x20 & n10379 ) | ( ~x20 & n10380 ) | ( n10379 & n10380 ) ;
  assign n10382 = ( ~n10374 & n10380 ) | ( ~n10374 & n10381 ) | ( n10380 & n10381 ) ;
  assign n10383 = n1297 & n5542 ;
  assign n10384 = x112 & n1301 ;
  assign n10385 = x113 | n10384 ;
  assign n10386 = ( n1303 & n10384 ) | ( n1303 & n10385 ) | ( n10384 & n10385 ) ;
  assign n10387 = x111 & n1426 ;
  assign n10388 = n10386 | n10387 ;
  assign n10389 = ( x23 & n10383 ) | ( x23 & ~n10388 ) | ( n10383 & ~n10388 ) ;
  assign n10390 = ( ~x23 & n10388 ) | ( ~x23 & n10389 ) | ( n10388 & n10389 ) ;
  assign n10391 = ( ~n10383 & n10389 ) | ( ~n10383 & n10390 ) | ( n10389 & n10390 ) ;
  assign n10392 = n1617 & n4934 ;
  assign n10393 = x109 & n1621 ;
  assign n10394 = x110 | n10393 ;
  assign n10395 = ( n1623 & n10393 ) | ( n1623 & n10394 ) | ( n10393 & n10394 ) ;
  assign n10396 = x108 & n1749 ;
  assign n10397 = n10395 | n10396 ;
  assign n10398 = ( x26 & n10392 ) | ( x26 & ~n10397 ) | ( n10392 & ~n10397 ) ;
  assign n10399 = ( ~x26 & n10397 ) | ( ~x26 & n10398 ) | ( n10397 & n10398 ) ;
  assign n10400 = ( ~n10392 & n10398 ) | ( ~n10392 & n10399 ) | ( n10398 & n10399 ) ;
  assign n10401 = n1949 & n4362 ;
  assign n10402 = x106 & n1953 ;
  assign n10403 = x107 | n10402 ;
  assign n10404 = ( n1955 & n10402 ) | ( n1955 & n10403 ) | ( n10402 & n10403 ) ;
  assign n10405 = x105 & n2114 ;
  assign n10406 = n10404 | n10405 ;
  assign n10407 = ( x29 & n10401 ) | ( x29 & ~n10406 ) | ( n10401 & ~n10406 ) ;
  assign n10408 = ( ~x29 & n10406 ) | ( ~x29 & n10407 ) | ( n10406 & n10407 ) ;
  assign n10409 = ( ~n10401 & n10407 ) | ( ~n10401 & n10408 ) | ( n10407 & n10408 ) ;
  assign n10410 = n2320 & n3665 ;
  assign n10411 = x103 & n2324 ;
  assign n10412 = x104 | n10411 ;
  assign n10413 = ( n2326 & n10411 ) | ( n2326 & n10412 ) | ( n10411 & n10412 ) ;
  assign n10414 = x102 & n2497 ;
  assign n10415 = n10413 | n10414 ;
  assign n10416 = ( x32 & n10410 ) | ( x32 & ~n10415 ) | ( n10410 & ~n10415 ) ;
  assign n10417 = ( ~x32 & n10415 ) | ( ~x32 & n10416 ) | ( n10415 & n10416 ) ;
  assign n10418 = ( ~n10410 & n10416 ) | ( ~n10410 & n10417 ) | ( n10416 & n10417 ) ;
  assign n10419 = n2766 & n3326 ;
  assign n10420 = x100 & n2770 ;
  assign n10421 = x101 | n10420 ;
  assign n10422 = ( n2772 & n10420 ) | ( n2772 & n10421 ) | ( n10420 & n10421 ) ;
  assign n10423 = x99 & n2943 ;
  assign n10424 = n10422 | n10423 ;
  assign n10425 = ( x35 & n10419 ) | ( x35 & ~n10424 ) | ( n10419 & ~n10424 ) ;
  assign n10426 = ( ~x35 & n10424 ) | ( ~x35 & n10425 ) | ( n10424 & n10425 ) ;
  assign n10427 = ( ~n10419 & n10425 ) | ( ~n10419 & n10426 ) | ( n10425 & n10426 ) ;
  assign n10428 = n2725 & n3224 ;
  assign n10429 = x97 & n3228 ;
  assign n10430 = x98 | n10429 ;
  assign n10431 = ( n3230 & n10429 ) | ( n3230 & n10430 ) | ( n10429 & n10430 ) ;
  assign n10432 = x96 & n3413 ;
  assign n10433 = n10431 | n10432 ;
  assign n10434 = ( x38 & n10428 ) | ( x38 & ~n10433 ) | ( n10428 & ~n10433 ) ;
  assign n10435 = ( ~x38 & n10433 ) | ( ~x38 & n10434 ) | ( n10433 & n10434 ) ;
  assign n10436 = ( ~n10428 & n10434 ) | ( ~n10428 & n10435 ) | ( n10434 & n10435 ) ;
  assign n10437 = n446 & n8154 ;
  assign n10438 = x73 & n8158 ;
  assign n10439 = x74 | n10438 ;
  assign n10440 = ( n8160 & n10438 ) | ( n8160 & n10439 ) | ( n10438 & n10439 ) ;
  assign n10441 = x72 & n8439 ;
  assign n10442 = n10440 | n10441 ;
  assign n10443 = ( x62 & n10437 ) | ( x62 & ~n10442 ) | ( n10437 & ~n10442 ) ;
  assign n10444 = ( ~x62 & n10442 ) | ( ~x62 & n10443 ) | ( n10442 & n10443 ) ;
  assign n10445 = ( ~n10437 & n10443 ) | ( ~n10437 & n10444 ) | ( n10443 & n10444 ) ;
  assign n10446 = x70 & n8927 ;
  assign n10447 = ( ~x71 & n8693 ) | ( ~x71 & n8927 ) | ( n8693 & n8927 ) ;
  assign n10448 = ( n8693 & n10446 ) | ( n8693 & ~n10447 ) | ( n10446 & ~n10447 ) ;
  assign n10449 = ( n10178 & n10445 ) | ( n10178 & n10448 ) | ( n10445 & n10448 ) ;
  assign n10450 = ( n10178 & ~n10445 ) | ( n10178 & n10448 ) | ( ~n10445 & n10448 ) ;
  assign n10451 = ( n10445 & ~n10449 ) | ( n10445 & n10450 ) | ( ~n10449 & n10450 ) ;
  assign n10452 = n569 & n7423 ;
  assign n10453 = x76 & n7427 ;
  assign n10454 = x77 | n10453 ;
  assign n10455 = ( n7429 & n10453 ) | ( n7429 & n10454 ) | ( n10453 & n10454 ) ;
  assign n10456 = x75 & n7708 ;
  assign n10457 = n10455 | n10456 ;
  assign n10458 = ( x59 & n10452 ) | ( x59 & ~n10457 ) | ( n10452 & ~n10457 ) ;
  assign n10459 = ( ~x59 & n10457 ) | ( ~x59 & n10458 ) | ( n10457 & n10458 ) ;
  assign n10460 = ( ~n10452 & n10458 ) | ( ~n10452 & n10459 ) | ( n10458 & n10459 ) ;
  assign n10461 = ( n10190 & n10451 ) | ( n10190 & n10460 ) | ( n10451 & n10460 ) ;
  assign n10462 = ( ~n10190 & n10451 ) | ( ~n10190 & n10460 ) | ( n10451 & n10460 ) ;
  assign n10463 = ( n10190 & ~n10461 ) | ( n10190 & n10462 ) | ( ~n10461 & n10462 ) ;
  assign n10464 = n769 & n6713 ;
  assign n10465 = x79 & n6717 ;
  assign n10466 = x80 | n10465 ;
  assign n10467 = ( n6719 & n10465 ) | ( n6719 & n10466 ) | ( n10465 & n10466 ) ;
  assign n10468 = x78 & n6980 ;
  assign n10469 = n10467 | n10468 ;
  assign n10470 = ( x56 & n10464 ) | ( x56 & ~n10469 ) | ( n10464 & ~n10469 ) ;
  assign n10471 = ( ~x56 & n10469 ) | ( ~x56 & n10470 ) | ( n10469 & n10470 ) ;
  assign n10472 = ( ~n10464 & n10470 ) | ( ~n10464 & n10471 ) | ( n10470 & n10471 ) ;
  assign n10473 = ( n10193 & n10463 ) | ( n10193 & n10472 ) | ( n10463 & n10472 ) ;
  assign n10474 = ( n10193 & ~n10463 ) | ( n10193 & n10472 ) | ( ~n10463 & n10472 ) ;
  assign n10475 = ( n10463 & ~n10473 ) | ( n10463 & n10474 ) | ( ~n10473 & n10474 ) ;
  assign n10476 = n1082 & n6027 ;
  assign n10477 = x82 & n6031 ;
  assign n10478 = x83 | n10477 ;
  assign n10479 = ( n6033 & n10477 ) | ( n6033 & n10478 ) | ( n10477 & n10478 ) ;
  assign n10480 = x81 & n6303 ;
  assign n10481 = n10479 | n10480 ;
  assign n10482 = ( x53 & n10476 ) | ( x53 & ~n10481 ) | ( n10476 & ~n10481 ) ;
  assign n10483 = ( ~x53 & n10481 ) | ( ~x53 & n10482 ) | ( n10481 & n10482 ) ;
  assign n10484 = ( ~n10476 & n10482 ) | ( ~n10476 & n10483 ) | ( n10482 & n10483 ) ;
  assign n10485 = ( n10205 & n10475 ) | ( n10205 & n10484 ) | ( n10475 & n10484 ) ;
  assign n10486 = ( ~n10205 & n10475 ) | ( ~n10205 & n10484 ) | ( n10475 & n10484 ) ;
  assign n10487 = ( n10205 & ~n10485 ) | ( n10205 & n10486 ) | ( ~n10485 & n10486 ) ;
  assign n10488 = n1366 & n5374 ;
  assign n10489 = x85 & n5378 ;
  assign n10490 = x86 | n10489 ;
  assign n10491 = ( n5380 & n10489 ) | ( n5380 & n10490 ) | ( n10489 & n10490 ) ;
  assign n10492 = x84 & n5638 ;
  assign n10493 = n10491 | n10492 ;
  assign n10494 = ( x50 & n10488 ) | ( x50 & ~n10493 ) | ( n10488 & ~n10493 ) ;
  assign n10495 = ( ~x50 & n10493 ) | ( ~x50 & n10494 ) | ( n10493 & n10494 ) ;
  assign n10496 = ( ~n10488 & n10494 ) | ( ~n10488 & n10495 ) | ( n10494 & n10495 ) ;
  assign n10497 = ( n10217 & n10487 ) | ( n10217 & n10496 ) | ( n10487 & n10496 ) ;
  assign n10498 = ( n10217 & ~n10487 ) | ( n10217 & n10496 ) | ( ~n10487 & n10496 ) ;
  assign n10499 = ( n10487 & ~n10497 ) | ( n10487 & n10498 ) | ( ~n10497 & n10498 ) ;
  assign n10500 = n1585 & n4787 ;
  assign n10501 = x88 & n4791 ;
  assign n10502 = x89 | n10501 ;
  assign n10503 = ( n4793 & n10501 ) | ( n4793 & n10502 ) | ( n10501 & n10502 ) ;
  assign n10504 = x87 & n5030 ;
  assign n10505 = n10503 | n10504 ;
  assign n10506 = ( x47 & n10500 ) | ( x47 & ~n10505 ) | ( n10500 & ~n10505 ) ;
  assign n10507 = ( ~x47 & n10505 ) | ( ~x47 & n10506 ) | ( n10505 & n10506 ) ;
  assign n10508 = ( ~n10500 & n10506 ) | ( ~n10500 & n10507 ) | ( n10506 & n10507 ) ;
  assign n10509 = ( n10229 & n10499 ) | ( n10229 & n10508 ) | ( n10499 & n10508 ) ;
  assign n10510 = ( ~n10229 & n10499 ) | ( ~n10229 & n10508 ) | ( n10499 & n10508 ) ;
  assign n10511 = ( n10229 & ~n10509 ) | ( n10229 & n10510 ) | ( ~n10509 & n10510 ) ;
  assign n10512 = n2042 & n4227 ;
  assign n10513 = x91 & n4231 ;
  assign n10514 = x92 | n10513 ;
  assign n10515 = ( n4233 & n10513 ) | ( n4233 & n10514 ) | ( n10513 & n10514 ) ;
  assign n10516 = x90 & n4470 ;
  assign n10517 = n10515 | n10516 ;
  assign n10518 = ( x44 & n10512 ) | ( x44 & ~n10517 ) | ( n10512 & ~n10517 ) ;
  assign n10519 = ( ~x44 & n10517 ) | ( ~x44 & n10518 ) | ( n10517 & n10518 ) ;
  assign n10520 = ( ~n10512 & n10518 ) | ( ~n10512 & n10519 ) | ( n10518 & n10519 ) ;
  assign n10521 = ( n10232 & n10511 ) | ( n10232 & n10520 ) | ( n10511 & n10520 ) ;
  assign n10522 = ( n10232 & ~n10511 ) | ( n10232 & n10520 ) | ( ~n10511 & n10520 ) ;
  assign n10523 = ( n10511 & ~n10521 ) | ( n10511 & n10522 ) | ( ~n10521 & n10522 ) ;
  assign n10524 = n2434 & n3715 ;
  assign n10525 = x94 & n3719 ;
  assign n10526 = x95 | n10525 ;
  assign n10527 = ( n3721 & n10525 ) | ( n3721 & n10526 ) | ( n10525 & n10526 ) ;
  assign n10528 = x93 & n3922 ;
  assign n10529 = n10527 | n10528 ;
  assign n10530 = ( x41 & n10524 ) | ( x41 & ~n10529 ) | ( n10524 & ~n10529 ) ;
  assign n10531 = ( ~x41 & n10529 ) | ( ~x41 & n10530 ) | ( n10529 & n10530 ) ;
  assign n10532 = ( ~n10524 & n10530 ) | ( ~n10524 & n10531 ) | ( n10530 & n10531 ) ;
  assign n10533 = ( n10244 & n10523 ) | ( n10244 & n10532 ) | ( n10523 & n10532 ) ;
  assign n10534 = ( ~n10244 & n10523 ) | ( ~n10244 & n10532 ) | ( n10523 & n10532 ) ;
  assign n10535 = ( n10244 & ~n10533 ) | ( n10244 & n10534 ) | ( ~n10533 & n10534 ) ;
  assign n10536 = ( n10256 & n10436 ) | ( n10256 & n10535 ) | ( n10436 & n10535 ) ;
  assign n10537 = ( n10256 & ~n10436 ) | ( n10256 & n10535 ) | ( ~n10436 & n10535 ) ;
  assign n10538 = ( n10436 & ~n10536 ) | ( n10436 & n10537 ) | ( ~n10536 & n10537 ) ;
  assign n10539 = ( n10259 & n10427 ) | ( n10259 & n10538 ) | ( n10427 & n10538 ) ;
  assign n10540 = ( n10259 & ~n10427 ) | ( n10259 & n10538 ) | ( ~n10427 & n10538 ) ;
  assign n10541 = ( n10427 & ~n10539 ) | ( n10427 & n10540 ) | ( ~n10539 & n10540 ) ;
  assign n10542 = ( n10262 & n10418 ) | ( n10262 & n10541 ) | ( n10418 & n10541 ) ;
  assign n10543 = ( n10262 & ~n10418 ) | ( n10262 & n10541 ) | ( ~n10418 & n10541 ) ;
  assign n10544 = ( n10418 & ~n10542 ) | ( n10418 & n10543 ) | ( ~n10542 & n10543 ) ;
  assign n10545 = ( n10274 & n10409 ) | ( n10274 & n10544 ) | ( n10409 & n10544 ) ;
  assign n10546 = ( n10274 & ~n10409 ) | ( n10274 & n10544 ) | ( ~n10409 & n10544 ) ;
  assign n10547 = ( n10409 & ~n10545 ) | ( n10409 & n10546 ) | ( ~n10545 & n10546 ) ;
  assign n10548 = ( n10277 & n10400 ) | ( n10277 & n10547 ) | ( n10400 & n10547 ) ;
  assign n10549 = ( ~n10277 & n10400 ) | ( ~n10277 & n10547 ) | ( n10400 & n10547 ) ;
  assign n10550 = ( n10277 & ~n10548 ) | ( n10277 & n10549 ) | ( ~n10548 & n10549 ) ;
  assign n10551 = ( n10289 & n10391 ) | ( n10289 & n10550 ) | ( n10391 & n10550 ) ;
  assign n10552 = ( n10289 & ~n10391 ) | ( n10289 & n10550 ) | ( ~n10391 & n10550 ) ;
  assign n10553 = ( n10391 & ~n10551 ) | ( n10391 & n10552 ) | ( ~n10551 & n10552 ) ;
  assign n10554 = ( n10292 & n10382 ) | ( n10292 & n10553 ) | ( n10382 & n10553 ) ;
  assign n10555 = ( n10292 & ~n10382 ) | ( n10292 & n10553 ) | ( ~n10382 & n10553 ) ;
  assign n10556 = ( n10382 & ~n10554 ) | ( n10382 & n10555 ) | ( ~n10554 & n10555 ) ;
  assign n10557 = ( n10295 & n10373 ) | ( n10295 & n10556 ) | ( n10373 & n10556 ) ;
  assign n10558 = ( n10295 & ~n10373 ) | ( n10295 & n10556 ) | ( ~n10373 & n10556 ) ;
  assign n10559 = ( n10373 & ~n10557 ) | ( n10373 & n10558 ) | ( ~n10557 & n10558 ) ;
  assign n10560 = ( n10307 & n10364 ) | ( n10307 & n10559 ) | ( n10364 & n10559 ) ;
  assign n10561 = ( ~n10307 & n10364 ) | ( ~n10307 & n10559 ) | ( n10364 & n10559 ) ;
  assign n10562 = ( n10307 & ~n10560 ) | ( n10307 & n10561 ) | ( ~n10560 & n10561 ) ;
  assign n10563 = ( n10319 & n10355 ) | ( n10319 & n10562 ) | ( n10355 & n10562 ) ;
  assign n10564 = ( n10319 & ~n10355 ) | ( n10319 & n10562 ) | ( ~n10355 & n10562 ) ;
  assign n10565 = ( n10355 & ~n10563 ) | ( n10355 & n10564 ) | ( ~n10563 & n10564 ) ;
  assign n10566 = ( n10322 & n10346 ) | ( n10322 & n10565 ) | ( n10346 & n10565 ) ;
  assign n10567 = ( ~n10322 & n10346 ) | ( ~n10322 & n10565 ) | ( n10346 & n10565 ) ;
  assign n10568 = ( n10322 & ~n10566 ) | ( n10322 & n10567 ) | ( ~n10566 & n10567 ) ;
  assign n10569 = ( n10334 & n10337 ) | ( n10334 & n10568 ) | ( n10337 & n10568 ) ;
  assign n10570 = ( n10334 & ~n10337 ) | ( n10334 & n10568 ) | ( ~n10337 & n10568 ) ;
  assign n10571 = ( n10337 & ~n10569 ) | ( n10337 & n10570 ) | ( ~n10569 & n10570 ) ;
  assign n10572 = n810 & n7098 ;
  assign n10573 = x119 & n814 ;
  assign n10574 = x120 | n10573 ;
  assign n10575 = ( n816 & n10573 ) | ( n816 & n10574 ) | ( n10573 & n10574 ) ;
  assign n10576 = x118 & n885 ;
  assign n10577 = n10575 | n10576 ;
  assign n10578 = ( x17 & n10572 ) | ( x17 & ~n10577 ) | ( n10572 & ~n10577 ) ;
  assign n10579 = ( ~x17 & n10577 ) | ( ~x17 & n10578 ) | ( n10577 & n10578 ) ;
  assign n10580 = ( ~n10572 & n10578 ) | ( ~n10572 & n10579 ) | ( n10578 & n10579 ) ;
  assign n10581 = n1297 & n5750 ;
  assign n10582 = x113 & n1301 ;
  assign n10583 = x114 | n10582 ;
  assign n10584 = ( n1303 & n10582 ) | ( n1303 & n10583 ) | ( n10582 & n10583 ) ;
  assign n10585 = x112 & n1426 ;
  assign n10586 = n10584 | n10585 ;
  assign n10587 = ( x23 & n10581 ) | ( x23 & ~n10586 ) | ( n10581 & ~n10586 ) ;
  assign n10588 = ( ~x23 & n10586 ) | ( ~x23 & n10587 ) | ( n10586 & n10587 ) ;
  assign n10589 = ( ~n10581 & n10587 ) | ( ~n10581 & n10588 ) | ( n10587 & n10588 ) ;
  assign n10590 = n2320 & n3998 ;
  assign n10591 = x104 & n2324 ;
  assign n10592 = x105 | n10591 ;
  assign n10593 = ( n2326 & n10591 ) | ( n2326 & n10592 ) | ( n10591 & n10592 ) ;
  assign n10594 = x103 & n2497 ;
  assign n10595 = n10593 | n10594 ;
  assign n10596 = ( x32 & n10590 ) | ( x32 & ~n10595 ) | ( n10590 & ~n10595 ) ;
  assign n10597 = ( ~x32 & n10595 ) | ( ~x32 & n10596 ) | ( n10595 & n10596 ) ;
  assign n10598 = ( ~n10590 & n10596 ) | ( ~n10590 & n10597 ) | ( n10596 & n10597 ) ;
  assign n10599 = n1466 & n5374 ;
  assign n10600 = x86 & n5378 ;
  assign n10601 = x87 | n10600 ;
  assign n10602 = ( n5380 & n10600 ) | ( n5380 & n10601 ) | ( n10600 & n10601 ) ;
  assign n10603 = x85 & n5638 ;
  assign n10604 = n10602 | n10603 ;
  assign n10605 = ( x50 & n10599 ) | ( x50 & ~n10604 ) | ( n10599 & ~n10604 ) ;
  assign n10606 = ( ~x50 & n10604 ) | ( ~x50 & n10605 ) | ( n10604 & n10605 ) ;
  assign n10607 = ( ~n10599 & n10605 ) | ( ~n10599 & n10606 ) | ( n10605 & n10606 ) ;
  assign n10608 = n637 & n7423 ;
  assign n10609 = x77 & n7427 ;
  assign n10610 = x78 | n10609 ;
  assign n10611 = ( n7429 & n10609 ) | ( n7429 & n10610 ) | ( n10609 & n10610 ) ;
  assign n10612 = x76 & n7708 ;
  assign n10613 = n10611 | n10612 ;
  assign n10614 = ( x59 & n10608 ) | ( x59 & ~n10613 ) | ( n10608 & ~n10613 ) ;
  assign n10615 = ( ~x59 & n10613 ) | ( ~x59 & n10614 ) | ( n10613 & n10614 ) ;
  assign n10616 = ( ~n10608 & n10614 ) | ( ~n10608 & n10615 ) | ( n10614 & n10615 ) ;
  assign n10617 = n461 & n8154 ;
  assign n10618 = x74 & n8158 ;
  assign n10619 = x75 | n10618 ;
  assign n10620 = ( n8160 & n10618 ) | ( n8160 & n10619 ) | ( n10618 & n10619 ) ;
  assign n10621 = x73 & n8439 ;
  assign n10622 = n10620 | n10621 ;
  assign n10623 = ( x62 & n10617 ) | ( x62 & ~n10622 ) | ( n10617 & ~n10622 ) ;
  assign n10624 = ( ~x62 & n10622 ) | ( ~x62 & n10623 ) | ( n10622 & n10623 ) ;
  assign n10625 = ( ~n10617 & n10623 ) | ( ~n10617 & n10624 ) | ( n10623 & n10624 ) ;
  assign n10626 = x71 & n8927 ;
  assign n10627 = ( ~x72 & n8693 ) | ( ~x72 & n8927 ) | ( n8693 & n8927 ) ;
  assign n10628 = ( n8693 & n10626 ) | ( n8693 & ~n10627 ) | ( n10626 & ~n10627 ) ;
  assign n10629 = ( ~n10448 & n10450 ) | ( ~n10448 & n10628 ) | ( n10450 & n10628 ) ;
  assign n10630 = ( n10448 & n10450 ) | ( n10448 & ~n10628 ) | ( n10450 & ~n10628 ) ;
  assign n10631 = ( ~n10450 & n10629 ) | ( ~n10450 & n10630 ) | ( n10629 & n10630 ) ;
  assign n10632 = ( n10616 & n10625 ) | ( n10616 & n10631 ) | ( n10625 & n10631 ) ;
  assign n10633 = ( ~n10616 & n10625 ) | ( ~n10616 & n10631 ) | ( n10625 & n10631 ) ;
  assign n10634 = ( n10616 & ~n10632 ) | ( n10616 & n10633 ) | ( ~n10632 & n10633 ) ;
  assign n10635 = n910 & n6713 ;
  assign n10636 = x80 & n6717 ;
  assign n10637 = x81 | n10636 ;
  assign n10638 = ( n6719 & n10636 ) | ( n6719 & n10637 ) | ( n10636 & n10637 ) ;
  assign n10639 = x79 & n6980 ;
  assign n10640 = n10638 | n10639 ;
  assign n10641 = ( x56 & n10635 ) | ( x56 & ~n10640 ) | ( n10635 & ~n10640 ) ;
  assign n10642 = ( ~x56 & n10640 ) | ( ~x56 & n10641 ) | ( n10640 & n10641 ) ;
  assign n10643 = ( ~n10635 & n10641 ) | ( ~n10635 & n10642 ) | ( n10641 & n10642 ) ;
  assign n10644 = ( n10461 & n10634 ) | ( n10461 & n10643 ) | ( n10634 & n10643 ) ;
  assign n10645 = ( n10461 & ~n10634 ) | ( n10461 & n10643 ) | ( ~n10634 & n10643 ) ;
  assign n10646 = ( n10634 & ~n10644 ) | ( n10634 & n10645 ) | ( ~n10644 & n10645 ) ;
  assign n10647 = n1097 & n6027 ;
  assign n10648 = x83 & n6031 ;
  assign n10649 = x84 | n10648 ;
  assign n10650 = ( n6033 & n10648 ) | ( n6033 & n10649 ) | ( n10648 & n10649 ) ;
  assign n10651 = x82 & n6303 ;
  assign n10652 = n10650 | n10651 ;
  assign n10653 = ( x53 & n10647 ) | ( x53 & ~n10652 ) | ( n10647 & ~n10652 ) ;
  assign n10654 = ( ~x53 & n10652 ) | ( ~x53 & n10653 ) | ( n10652 & n10653 ) ;
  assign n10655 = ( ~n10647 & n10653 ) | ( ~n10647 & n10654 ) | ( n10653 & n10654 ) ;
  assign n10656 = ( n10473 & n10646 ) | ( n10473 & n10655 ) | ( n10646 & n10655 ) ;
  assign n10657 = ( ~n10473 & n10646 ) | ( ~n10473 & n10655 ) | ( n10646 & n10655 ) ;
  assign n10658 = ( n10473 & ~n10656 ) | ( n10473 & n10657 ) | ( ~n10656 & n10657 ) ;
  assign n10659 = ( n10485 & n10607 ) | ( n10485 & n10658 ) | ( n10607 & n10658 ) ;
  assign n10660 = ( n10485 & ~n10607 ) | ( n10485 & n10658 ) | ( ~n10607 & n10658 ) ;
  assign n10661 = ( n10607 & ~n10659 ) | ( n10607 & n10660 ) | ( ~n10659 & n10660 ) ;
  assign n10662 = n1701 & n4787 ;
  assign n10663 = x89 & n4791 ;
  assign n10664 = x90 | n10663 ;
  assign n10665 = ( n4793 & n10663 ) | ( n4793 & n10664 ) | ( n10663 & n10664 ) ;
  assign n10666 = x88 & n5030 ;
  assign n10667 = n10665 | n10666 ;
  assign n10668 = ( x47 & n10662 ) | ( x47 & ~n10667 ) | ( n10662 & ~n10667 ) ;
  assign n10669 = ( ~x47 & n10667 ) | ( ~x47 & n10668 ) | ( n10667 & n10668 ) ;
  assign n10670 = ( ~n10662 & n10668 ) | ( ~n10662 & n10669 ) | ( n10668 & n10669 ) ;
  assign n10671 = ( n10497 & n10661 ) | ( n10497 & n10670 ) | ( n10661 & n10670 ) ;
  assign n10672 = ( ~n10497 & n10661 ) | ( ~n10497 & n10670 ) | ( n10661 & n10670 ) ;
  assign n10673 = ( n10497 & ~n10671 ) | ( n10497 & n10672 ) | ( ~n10671 & n10672 ) ;
  assign n10674 = n2057 & n4227 ;
  assign n10675 = x92 & n4231 ;
  assign n10676 = x93 | n10675 ;
  assign n10677 = ( n4233 & n10675 ) | ( n4233 & n10676 ) | ( n10675 & n10676 ) ;
  assign n10678 = x91 & n4470 ;
  assign n10679 = n10677 | n10678 ;
  assign n10680 = ( x44 & n10674 ) | ( x44 & ~n10679 ) | ( n10674 & ~n10679 ) ;
  assign n10681 = ( ~x44 & n10679 ) | ( ~x44 & n10680 ) | ( n10679 & n10680 ) ;
  assign n10682 = ( ~n10674 & n10680 ) | ( ~n10674 & n10681 ) | ( n10680 & n10681 ) ;
  assign n10683 = ( n10509 & n10673 ) | ( n10509 & n10682 ) | ( n10673 & n10682 ) ;
  assign n10684 = ( n10509 & ~n10673 ) | ( n10509 & n10682 ) | ( ~n10673 & n10682 ) ;
  assign n10685 = ( n10673 & ~n10683 ) | ( n10673 & n10684 ) | ( ~n10683 & n10684 ) ;
  assign n10686 = n2449 & n3715 ;
  assign n10687 = x95 & n3719 ;
  assign n10688 = x96 | n10687 ;
  assign n10689 = ( n3721 & n10687 ) | ( n3721 & n10688 ) | ( n10687 & n10688 ) ;
  assign n10690 = x94 & n3922 ;
  assign n10691 = n10689 | n10690 ;
  assign n10692 = ( x41 & n10686 ) | ( x41 & ~n10691 ) | ( n10686 & ~n10691 ) ;
  assign n10693 = ( ~x41 & n10691 ) | ( ~x41 & n10692 ) | ( n10691 & n10692 ) ;
  assign n10694 = ( ~n10686 & n10692 ) | ( ~n10686 & n10693 ) | ( n10692 & n10693 ) ;
  assign n10695 = ( n10521 & n10685 ) | ( n10521 & n10694 ) | ( n10685 & n10694 ) ;
  assign n10696 = ( ~n10521 & n10685 ) | ( ~n10521 & n10694 ) | ( n10685 & n10694 ) ;
  assign n10697 = ( n10521 & ~n10695 ) | ( n10521 & n10696 ) | ( ~n10695 & n10696 ) ;
  assign n10698 = n2877 & n3224 ;
  assign n10699 = x98 & n3228 ;
  assign n10700 = x99 | n10699 ;
  assign n10701 = ( n3230 & n10699 ) | ( n3230 & n10700 ) | ( n10699 & n10700 ) ;
  assign n10702 = x97 & n3413 ;
  assign n10703 = n10701 | n10702 ;
  assign n10704 = ( x38 & n10698 ) | ( x38 & ~n10703 ) | ( n10698 & ~n10703 ) ;
  assign n10705 = ( ~x38 & n10703 ) | ( ~x38 & n10704 ) | ( n10703 & n10704 ) ;
  assign n10706 = ( ~n10698 & n10704 ) | ( ~n10698 & n10705 ) | ( n10704 & n10705 ) ;
  assign n10707 = ( n10533 & n10697 ) | ( n10533 & n10706 ) | ( n10697 & n10706 ) ;
  assign n10708 = ( n10533 & ~n10697 ) | ( n10533 & n10706 ) | ( ~n10697 & n10706 ) ;
  assign n10709 = ( n10697 & ~n10707 ) | ( n10697 & n10708 ) | ( ~n10707 & n10708 ) ;
  assign n10710 = n2766 & n3486 ;
  assign n10711 = x101 & n2770 ;
  assign n10712 = x102 | n10711 ;
  assign n10713 = ( n2772 & n10711 ) | ( n2772 & n10712 ) | ( n10711 & n10712 ) ;
  assign n10714 = x100 & n2943 ;
  assign n10715 = n10713 | n10714 ;
  assign n10716 = ( x35 & n10710 ) | ( x35 & ~n10715 ) | ( n10710 & ~n10715 ) ;
  assign n10717 = ( ~x35 & n10715 ) | ( ~x35 & n10716 ) | ( n10715 & n10716 ) ;
  assign n10718 = ( ~n10710 & n10716 ) | ( ~n10710 & n10717 ) | ( n10716 & n10717 ) ;
  assign n10719 = ( n10536 & n10709 ) | ( n10536 & n10718 ) | ( n10709 & n10718 ) ;
  assign n10720 = ( ~n10536 & n10709 ) | ( ~n10536 & n10718 ) | ( n10709 & n10718 ) ;
  assign n10721 = ( n10536 & ~n10719 ) | ( n10536 & n10720 ) | ( ~n10719 & n10720 ) ;
  assign n10722 = ( n10539 & n10598 ) | ( n10539 & n10721 ) | ( n10598 & n10721 ) ;
  assign n10723 = ( n10539 & ~n10598 ) | ( n10539 & n10721 ) | ( ~n10598 & n10721 ) ;
  assign n10724 = ( n10598 & ~n10722 ) | ( n10598 & n10723 ) | ( ~n10722 & n10723 ) ;
  assign n10725 = n1949 & n4377 ;
  assign n10726 = x107 & n1953 ;
  assign n10727 = x108 | n10726 ;
  assign n10728 = ( n1955 & n10726 ) | ( n1955 & n10727 ) | ( n10726 & n10727 ) ;
  assign n10729 = x106 & n2114 ;
  assign n10730 = n10728 | n10729 ;
  assign n10731 = ( x29 & n10725 ) | ( x29 & ~n10730 ) | ( n10725 & ~n10730 ) ;
  assign n10732 = ( ~x29 & n10730 ) | ( ~x29 & n10731 ) | ( n10730 & n10731 ) ;
  assign n10733 = ( ~n10725 & n10731 ) | ( ~n10725 & n10732 ) | ( n10731 & n10732 ) ;
  assign n10734 = ( n10542 & n10724 ) | ( n10542 & n10733 ) | ( n10724 & n10733 ) ;
  assign n10735 = ( n10542 & ~n10724 ) | ( n10542 & n10733 ) | ( ~n10724 & n10733 ) ;
  assign n10736 = ( n10724 & ~n10734 ) | ( n10724 & n10735 ) | ( ~n10734 & n10735 ) ;
  assign n10737 = n1617 & n5130 ;
  assign n10738 = x110 & n1621 ;
  assign n10739 = x111 | n10738 ;
  assign n10740 = ( n1623 & n10738 ) | ( n1623 & n10739 ) | ( n10738 & n10739 ) ;
  assign n10741 = x109 & n1749 ;
  assign n10742 = n10740 | n10741 ;
  assign n10743 = ( x26 & n10737 ) | ( x26 & ~n10742 ) | ( n10737 & ~n10742 ) ;
  assign n10744 = ( ~x26 & n10742 ) | ( ~x26 & n10743 ) | ( n10742 & n10743 ) ;
  assign n10745 = ( ~n10737 & n10743 ) | ( ~n10737 & n10744 ) | ( n10743 & n10744 ) ;
  assign n10746 = ( n10545 & n10736 ) | ( n10545 & n10745 ) | ( n10736 & n10745 ) ;
  assign n10747 = ( n10545 & ~n10736 ) | ( n10545 & n10745 ) | ( ~n10736 & n10745 ) ;
  assign n10748 = ( n10736 & ~n10746 ) | ( n10736 & n10747 ) | ( ~n10746 & n10747 ) ;
  assign n10749 = ( n10548 & n10589 ) | ( n10548 & n10748 ) | ( n10589 & n10748 ) ;
  assign n10750 = ( n10548 & ~n10589 ) | ( n10548 & n10748 ) | ( ~n10589 & n10748 ) ;
  assign n10751 = ( n10589 & ~n10749 ) | ( n10589 & n10750 ) | ( ~n10749 & n10750 ) ;
  assign n10752 = n1016 & n6201 ;
  assign n10753 = x116 & n1020 ;
  assign n10754 = x117 | n10753 ;
  assign n10755 = ( n1022 & n10753 ) | ( n1022 & n10754 ) | ( n10753 & n10754 ) ;
  assign n10756 = x115 & n1145 ;
  assign n10757 = n10755 | n10756 ;
  assign n10758 = ( x20 & n10752 ) | ( x20 & ~n10757 ) | ( n10752 & ~n10757 ) ;
  assign n10759 = ( ~x20 & n10757 ) | ( ~x20 & n10758 ) | ( n10757 & n10758 ) ;
  assign n10760 = ( ~n10752 & n10758 ) | ( ~n10752 & n10759 ) | ( n10758 & n10759 ) ;
  assign n10761 = ( n10551 & n10751 ) | ( n10551 & n10760 ) | ( n10751 & n10760 ) ;
  assign n10762 = ( n10551 & ~n10751 ) | ( n10551 & n10760 ) | ( ~n10751 & n10760 ) ;
  assign n10763 = ( n10751 & ~n10761 ) | ( n10751 & n10762 ) | ( ~n10761 & n10762 ) ;
  assign n10764 = ( n10554 & n10580 ) | ( n10554 & n10763 ) | ( n10580 & n10763 ) ;
  assign n10765 = ( n10554 & ~n10580 ) | ( n10554 & n10763 ) | ( ~n10580 & n10763 ) ;
  assign n10766 = ( n10580 & ~n10764 ) | ( n10580 & n10765 ) | ( ~n10764 & n10765 ) ;
  assign n10767 = n583 & n7597 ;
  assign n10768 = x122 & n587 ;
  assign n10769 = x123 | n10768 ;
  assign n10770 = ( n589 & n10768 ) | ( n589 & n10769 ) | ( n10768 & n10769 ) ;
  assign n10771 = x121 & n676 ;
  assign n10772 = n10770 | n10771 ;
  assign n10773 = ( x14 & n10767 ) | ( x14 & ~n10772 ) | ( n10767 & ~n10772 ) ;
  assign n10774 = ( ~x14 & n10772 ) | ( ~x14 & n10773 ) | ( n10772 & n10773 ) ;
  assign n10775 = ( ~n10767 & n10773 ) | ( ~n10767 & n10774 ) | ( n10773 & n10774 ) ;
  assign n10776 = ( n10557 & n10766 ) | ( n10557 & n10775 ) | ( n10766 & n10775 ) ;
  assign n10777 = ( n10557 & ~n10766 ) | ( n10557 & n10775 ) | ( ~n10766 & n10775 ) ;
  assign n10778 = ( n10766 & ~n10776 ) | ( n10766 & n10777 ) | ( ~n10776 & n10777 ) ;
  assign n10779 = n407 & n8587 ;
  assign n10780 = x125 & n411 ;
  assign n10781 = x126 | n10780 ;
  assign n10782 = ( n413 & n10780 ) | ( n413 & n10781 ) | ( n10780 & n10781 ) ;
  assign n10783 = x124 & n491 ;
  assign n10784 = n10782 | n10783 ;
  assign n10785 = ( x11 & n10779 ) | ( x11 & ~n10784 ) | ( n10779 & ~n10784 ) ;
  assign n10786 = ( ~x11 & n10784 ) | ( ~x11 & n10785 ) | ( n10784 & n10785 ) ;
  assign n10787 = ( ~n10779 & n10785 ) | ( ~n10779 & n10786 ) | ( n10785 & n10786 ) ;
  assign n10788 = ( n10560 & n10778 ) | ( n10560 & n10787 ) | ( n10778 & n10787 ) ;
  assign n10789 = ( n10560 & ~n10778 ) | ( n10560 & n10787 ) | ( ~n10778 & n10787 ) ;
  assign n10790 = ( n10778 & ~n10788 ) | ( n10778 & n10789 ) | ( ~n10788 & n10789 ) ;
  assign n10791 = n291 & n8862 ;
  assign n10792 = ( x127 & n330 ) | ( x127 & n10791 ) | ( n330 & n10791 ) ;
  assign n10793 = x8 | n10792 ;
  assign n10794 = ~x8 & n10792 ;
  assign n10795 = ( ~n10792 & n10793 ) | ( ~n10792 & n10794 ) | ( n10793 & n10794 ) ;
  assign n10796 = ( n10563 & n10790 ) | ( n10563 & n10795 ) | ( n10790 & n10795 ) ;
  assign n10797 = ( n10563 & ~n10790 ) | ( n10563 & n10795 ) | ( ~n10790 & n10795 ) ;
  assign n10798 = ( n10790 & ~n10796 ) | ( n10790 & n10797 ) | ( ~n10796 & n10797 ) ;
  assign n10799 = ( n10566 & n10569 ) | ( n10566 & n10798 ) | ( n10569 & n10798 ) ;
  assign n10800 = ( n10566 & ~n10569 ) | ( n10566 & n10798 ) | ( ~n10569 & n10798 ) ;
  assign n10801 = ( n10569 & ~n10799 ) | ( n10569 & n10800 ) | ( ~n10799 & n10800 ) ;
  assign n10802 = n810 & n7113 ;
  assign n10803 = x120 & n814 ;
  assign n10804 = x121 | n10803 ;
  assign n10805 = ( n816 & n10803 ) | ( n816 & n10804 ) | ( n10803 & n10804 ) ;
  assign n10806 = x119 & n885 ;
  assign n10807 = n10805 | n10806 ;
  assign n10808 = ( x17 & n10802 ) | ( x17 & ~n10807 ) | ( n10802 & ~n10807 ) ;
  assign n10809 = ( ~x17 & n10807 ) | ( ~x17 & n10808 ) | ( n10807 & n10808 ) ;
  assign n10810 = ( ~n10802 & n10808 ) | ( ~n10802 & n10809 ) | ( n10808 & n10809 ) ;
  assign n10811 = n1297 & n5765 ;
  assign n10812 = x114 & n1301 ;
  assign n10813 = x115 | n10812 ;
  assign n10814 = ( n1303 & n10812 ) | ( n1303 & n10813 ) | ( n10812 & n10813 ) ;
  assign n10815 = x113 & n1426 ;
  assign n10816 = n10814 | n10815 ;
  assign n10817 = ( x23 & n10811 ) | ( x23 & ~n10816 ) | ( n10811 & ~n10816 ) ;
  assign n10818 = ( ~x23 & n10816 ) | ( ~x23 & n10817 ) | ( n10816 & n10817 ) ;
  assign n10819 = ( ~n10811 & n10817 ) | ( ~n10811 & n10818 ) | ( n10817 & n10818 ) ;
  assign n10820 = n1617 & n5145 ;
  assign n10821 = x111 & n1621 ;
  assign n10822 = x112 | n10821 ;
  assign n10823 = ( n1623 & n10821 ) | ( n1623 & n10822 ) | ( n10821 & n10822 ) ;
  assign n10824 = x110 & n1749 ;
  assign n10825 = n10823 | n10824 ;
  assign n10826 = ( x26 & n10820 ) | ( x26 & ~n10825 ) | ( n10820 & ~n10825 ) ;
  assign n10827 = ( ~x26 & n10825 ) | ( ~x26 & n10826 ) | ( n10825 & n10826 ) ;
  assign n10828 = ( ~n10820 & n10826 ) | ( ~n10820 & n10827 ) | ( n10826 & n10827 ) ;
  assign n10829 = n3162 & n3224 ;
  assign n10830 = x99 & n3228 ;
  assign n10831 = x100 | n10830 ;
  assign n10832 = ( n3230 & n10830 ) | ( n3230 & n10831 ) | ( n10830 & n10831 ) ;
  assign n10833 = x98 & n3413 ;
  assign n10834 = n10832 | n10833 ;
  assign n10835 = ( x38 & n10829 ) | ( x38 & ~n10834 ) | ( n10829 & ~n10834 ) ;
  assign n10836 = ( ~x38 & n10834 ) | ( ~x38 & n10835 ) | ( n10834 & n10835 ) ;
  assign n10837 = ( ~n10829 & n10835 ) | ( ~n10829 & n10836 ) | ( n10835 & n10836 ) ;
  assign n10838 = n2585 & n3715 ;
  assign n10839 = x96 & n3719 ;
  assign n10840 = x97 | n10839 ;
  assign n10841 = ( n3721 & n10839 ) | ( n3721 & n10840 ) | ( n10839 & n10840 ) ;
  assign n10842 = x95 & n3922 ;
  assign n10843 = n10841 | n10842 ;
  assign n10844 = ( x41 & n10838 ) | ( x41 & ~n10843 ) | ( n10838 & ~n10843 ) ;
  assign n10845 = ( ~x41 & n10843 ) | ( ~x41 & n10844 ) | ( n10843 & n10844 ) ;
  assign n10846 = ( ~n10838 & n10844 ) | ( ~n10838 & n10845 ) | ( n10844 & n10845 ) ;
  assign n10847 = n1481 & n5374 ;
  assign n10848 = x87 & n5378 ;
  assign n10849 = x88 | n10848 ;
  assign n10850 = ( n5380 & n10848 ) | ( n5380 & n10849 ) | ( n10848 & n10849 ) ;
  assign n10851 = x86 & n5638 ;
  assign n10852 = n10850 | n10851 ;
  assign n10853 = ( x50 & n10847 ) | ( x50 & ~n10852 ) | ( n10847 & ~n10852 ) ;
  assign n10854 = ( ~x50 & n10852 ) | ( ~x50 & n10853 ) | ( n10852 & n10853 ) ;
  assign n10855 = ( ~n10847 & n10853 ) | ( ~n10847 & n10854 ) | ( n10853 & n10854 ) ;
  assign n10856 = n554 & n8154 ;
  assign n10857 = x75 & n8158 ;
  assign n10858 = x76 | n10857 ;
  assign n10859 = ( n8160 & n10857 ) | ( n8160 & n10858 ) | ( n10857 & n10858 ) ;
  assign n10860 = x74 & n8439 ;
  assign n10861 = n10859 | n10860 ;
  assign n10862 = ( x62 & n10856 ) | ( x62 & ~n10861 ) | ( n10856 & ~n10861 ) ;
  assign n10863 = ( ~x62 & n10861 ) | ( ~x62 & n10862 ) | ( n10861 & n10862 ) ;
  assign n10864 = ( ~n10856 & n10862 ) | ( ~n10856 & n10863 ) | ( n10862 & n10863 ) ;
  assign n10865 = x72 & n8927 ;
  assign n10866 = ( ~x73 & n8693 ) | ( ~x73 & n8927 ) | ( n8693 & n8927 ) ;
  assign n10867 = ( n8693 & n10865 ) | ( n8693 & ~n10866 ) | ( n10865 & ~n10866 ) ;
  assign n10868 = ( ~x8 & n10628 ) | ( ~x8 & n10867 ) | ( n10628 & n10867 ) ;
  assign n10869 = ( n10628 & n10867 ) | ( n10628 & ~n10868 ) | ( n10867 & ~n10868 ) ;
  assign n10870 = ( x8 & n10868 ) | ( x8 & ~n10869 ) | ( n10868 & ~n10869 ) ;
  assign n10871 = ( n10629 & ~n10864 ) | ( n10629 & n10870 ) | ( ~n10864 & n10870 ) ;
  assign n10872 = ( n10629 & n10864 ) | ( n10629 & n10870 ) | ( n10864 & n10870 ) ;
  assign n10873 = ( n10864 & n10871 ) | ( n10864 & ~n10872 ) | ( n10871 & ~n10872 ) ;
  assign n10874 = n701 & n7423 ;
  assign n10875 = x78 & n7427 ;
  assign n10876 = x79 | n10875 ;
  assign n10877 = ( n7429 & n10875 ) | ( n7429 & n10876 ) | ( n10875 & n10876 ) ;
  assign n10878 = x77 & n7708 ;
  assign n10879 = n10877 | n10878 ;
  assign n10880 = ( x59 & n10874 ) | ( x59 & ~n10879 ) | ( n10874 & ~n10879 ) ;
  assign n10881 = ( ~x59 & n10879 ) | ( ~x59 & n10880 ) | ( n10879 & n10880 ) ;
  assign n10882 = ( ~n10874 & n10880 ) | ( ~n10874 & n10881 ) | ( n10880 & n10881 ) ;
  assign n10883 = ( n10632 & n10873 ) | ( n10632 & n10882 ) | ( n10873 & n10882 ) ;
  assign n10884 = ( ~n10632 & n10873 ) | ( ~n10632 & n10882 ) | ( n10873 & n10882 ) ;
  assign n10885 = ( n10632 & ~n10883 ) | ( n10632 & n10884 ) | ( ~n10883 & n10884 ) ;
  assign n10886 = n990 & n6713 ;
  assign n10887 = x81 & n6717 ;
  assign n10888 = x82 | n10887 ;
  assign n10889 = ( n6719 & n10887 ) | ( n6719 & n10888 ) | ( n10887 & n10888 ) ;
  assign n10890 = x80 & n6980 ;
  assign n10891 = n10889 | n10890 ;
  assign n10892 = ( x56 & n10886 ) | ( x56 & ~n10891 ) | ( n10886 & ~n10891 ) ;
  assign n10893 = ( ~x56 & n10891 ) | ( ~x56 & n10892 ) | ( n10891 & n10892 ) ;
  assign n10894 = ( ~n10886 & n10892 ) | ( ~n10886 & n10893 ) | ( n10892 & n10893 ) ;
  assign n10895 = ( n10644 & n10885 ) | ( n10644 & n10894 ) | ( n10885 & n10894 ) ;
  assign n10896 = ( ~n10644 & n10885 ) | ( ~n10644 & n10894 ) | ( n10885 & n10894 ) ;
  assign n10897 = ( n10644 & ~n10895 ) | ( n10644 & n10896 ) | ( ~n10895 & n10896 ) ;
  assign n10898 = n1262 & n6027 ;
  assign n10899 = x84 & n6031 ;
  assign n10900 = x85 | n10899 ;
  assign n10901 = ( n6033 & n10899 ) | ( n6033 & n10900 ) | ( n10899 & n10900 ) ;
  assign n10902 = x83 & n6303 ;
  assign n10903 = n10901 | n10902 ;
  assign n10904 = ( x53 & n10898 ) | ( x53 & ~n10903 ) | ( n10898 & ~n10903 ) ;
  assign n10905 = ( ~x53 & n10903 ) | ( ~x53 & n10904 ) | ( n10903 & n10904 ) ;
  assign n10906 = ( ~n10898 & n10904 ) | ( ~n10898 & n10905 ) | ( n10904 & n10905 ) ;
  assign n10907 = ( n10656 & n10897 ) | ( n10656 & n10906 ) | ( n10897 & n10906 ) ;
  assign n10908 = ( ~n10656 & n10897 ) | ( ~n10656 & n10906 ) | ( n10897 & n10906 ) ;
  assign n10909 = ( n10656 & ~n10907 ) | ( n10656 & n10908 ) | ( ~n10907 & n10908 ) ;
  assign n10910 = ( n10659 & n10855 ) | ( n10659 & n10909 ) | ( n10855 & n10909 ) ;
  assign n10911 = ( ~n10659 & n10855 ) | ( ~n10659 & n10909 ) | ( n10855 & n10909 ) ;
  assign n10912 = ( n10659 & ~n10910 ) | ( n10659 & n10911 ) | ( ~n10910 & n10911 ) ;
  assign n10913 = n1914 & n4787 ;
  assign n10914 = x90 & n4791 ;
  assign n10915 = x91 | n10914 ;
  assign n10916 = ( n4793 & n10914 ) | ( n4793 & n10915 ) | ( n10914 & n10915 ) ;
  assign n10917 = x89 & n5030 ;
  assign n10918 = n10916 | n10917 ;
  assign n10919 = ( x47 & n10913 ) | ( x47 & ~n10918 ) | ( n10913 & ~n10918 ) ;
  assign n10920 = ( ~x47 & n10918 ) | ( ~x47 & n10919 ) | ( n10918 & n10919 ) ;
  assign n10921 = ( ~n10913 & n10919 ) | ( ~n10913 & n10920 ) | ( n10919 & n10920 ) ;
  assign n10922 = ( n10671 & n10912 ) | ( n10671 & n10921 ) | ( n10912 & n10921 ) ;
  assign n10923 = ( ~n10671 & n10912 ) | ( ~n10671 & n10921 ) | ( n10912 & n10921 ) ;
  assign n10924 = ( n10671 & ~n10922 ) | ( n10671 & n10923 ) | ( ~n10922 & n10923 ) ;
  assign n10925 = n2294 & n4227 ;
  assign n10926 = x93 & n4231 ;
  assign n10927 = x94 | n10926 ;
  assign n10928 = ( n4233 & n10926 ) | ( n4233 & n10927 ) | ( n10926 & n10927 ) ;
  assign n10929 = x92 & n4470 ;
  assign n10930 = n10928 | n10929 ;
  assign n10931 = ( x44 & n10925 ) | ( x44 & ~n10930 ) | ( n10925 & ~n10930 ) ;
  assign n10932 = ( ~x44 & n10930 ) | ( ~x44 & n10931 ) | ( n10930 & n10931 ) ;
  assign n10933 = ( ~n10925 & n10931 ) | ( ~n10925 & n10932 ) | ( n10931 & n10932 ) ;
  assign n10934 = ( n10683 & n10924 ) | ( n10683 & n10933 ) | ( n10924 & n10933 ) ;
  assign n10935 = ( ~n10683 & n10924 ) | ( ~n10683 & n10933 ) | ( n10924 & n10933 ) ;
  assign n10936 = ( n10683 & ~n10934 ) | ( n10683 & n10935 ) | ( ~n10934 & n10935 ) ;
  assign n10937 = ( n10695 & n10846 ) | ( n10695 & n10936 ) | ( n10846 & n10936 ) ;
  assign n10938 = ( ~n10695 & n10846 ) | ( ~n10695 & n10936 ) | ( n10846 & n10936 ) ;
  assign n10939 = ( n10695 & ~n10937 ) | ( n10695 & n10938 ) | ( ~n10937 & n10938 ) ;
  assign n10940 = ( n10707 & n10837 ) | ( n10707 & n10939 ) | ( n10837 & n10939 ) ;
  assign n10941 = ( ~n10707 & n10837 ) | ( ~n10707 & n10939 ) | ( n10837 & n10939 ) ;
  assign n10942 = ( n10707 & ~n10940 ) | ( n10707 & n10941 ) | ( ~n10940 & n10941 ) ;
  assign n10943 = n2766 & n3650 ;
  assign n10944 = x102 & n2770 ;
  assign n10945 = x103 | n10944 ;
  assign n10946 = ( n2772 & n10944 ) | ( n2772 & n10945 ) | ( n10944 & n10945 ) ;
  assign n10947 = x101 & n2943 ;
  assign n10948 = n10946 | n10947 ;
  assign n10949 = ( x35 & n10943 ) | ( x35 & ~n10948 ) | ( n10943 & ~n10948 ) ;
  assign n10950 = ( ~x35 & n10948 ) | ( ~x35 & n10949 ) | ( n10948 & n10949 ) ;
  assign n10951 = ( ~n10943 & n10949 ) | ( ~n10943 & n10950 ) | ( n10949 & n10950 ) ;
  assign n10952 = ( n10719 & n10942 ) | ( n10719 & n10951 ) | ( n10942 & n10951 ) ;
  assign n10953 = ( ~n10719 & n10942 ) | ( ~n10719 & n10951 ) | ( n10942 & n10951 ) ;
  assign n10954 = ( n10719 & ~n10952 ) | ( n10719 & n10953 ) | ( ~n10952 & n10953 ) ;
  assign n10955 = n2320 & n4013 ;
  assign n10956 = x105 & n2324 ;
  assign n10957 = x106 | n10956 ;
  assign n10958 = ( n2326 & n10956 ) | ( n2326 & n10957 ) | ( n10956 & n10957 ) ;
  assign n10959 = x104 & n2497 ;
  assign n10960 = n10958 | n10959 ;
  assign n10961 = ( x32 & n10955 ) | ( x32 & ~n10960 ) | ( n10955 & ~n10960 ) ;
  assign n10962 = ( ~x32 & n10960 ) | ( ~x32 & n10961 ) | ( n10960 & n10961 ) ;
  assign n10963 = ( ~n10955 & n10961 ) | ( ~n10955 & n10962 ) | ( n10961 & n10962 ) ;
  assign n10964 = ( n10722 & n10954 ) | ( n10722 & n10963 ) | ( n10954 & n10963 ) ;
  assign n10965 = ( n10722 & ~n10954 ) | ( n10722 & n10963 ) | ( ~n10954 & n10963 ) ;
  assign n10966 = ( n10954 & ~n10964 ) | ( n10954 & n10965 ) | ( ~n10964 & n10965 ) ;
  assign n10967 = n1949 & n4734 ;
  assign n10968 = x108 & n1953 ;
  assign n10969 = x109 | n10968 ;
  assign n10970 = ( n1955 & n10968 ) | ( n1955 & n10969 ) | ( n10968 & n10969 ) ;
  assign n10971 = x107 & n2114 ;
  assign n10972 = n10970 | n10971 ;
  assign n10973 = ( x29 & n10967 ) | ( x29 & ~n10972 ) | ( n10967 & ~n10972 ) ;
  assign n10974 = ( ~x29 & n10972 ) | ( ~x29 & n10973 ) | ( n10972 & n10973 ) ;
  assign n10975 = ( ~n10967 & n10973 ) | ( ~n10967 & n10974 ) | ( n10973 & n10974 ) ;
  assign n10976 = ( n10734 & n10966 ) | ( n10734 & n10975 ) | ( n10966 & n10975 ) ;
  assign n10977 = ( n10734 & ~n10966 ) | ( n10734 & n10975 ) | ( ~n10966 & n10975 ) ;
  assign n10978 = ( n10966 & ~n10976 ) | ( n10966 & n10977 ) | ( ~n10976 & n10977 ) ;
  assign n10979 = ( n10746 & n10828 ) | ( n10746 & n10978 ) | ( n10828 & n10978 ) ;
  assign n10980 = ( n10746 & ~n10828 ) | ( n10746 & n10978 ) | ( ~n10828 & n10978 ) ;
  assign n10981 = ( n10828 & ~n10979 ) | ( n10828 & n10980 ) | ( ~n10979 & n10980 ) ;
  assign n10982 = ( n10749 & n10819 ) | ( n10749 & n10981 ) | ( n10819 & n10981 ) ;
  assign n10983 = ( n10749 & ~n10819 ) | ( n10749 & n10981 ) | ( ~n10819 & n10981 ) ;
  assign n10984 = ( n10819 & ~n10982 ) | ( n10819 & n10983 ) | ( ~n10982 & n10983 ) ;
  assign n10985 = n1016 & n6421 ;
  assign n10986 = x117 & n1020 ;
  assign n10987 = x118 | n10986 ;
  assign n10988 = ( n1022 & n10986 ) | ( n1022 & n10987 ) | ( n10986 & n10987 ) ;
  assign n10989 = x116 & n1145 ;
  assign n10990 = n10988 | n10989 ;
  assign n10991 = ( x20 & n10985 ) | ( x20 & ~n10990 ) | ( n10985 & ~n10990 ) ;
  assign n10992 = ( ~x20 & n10990 ) | ( ~x20 & n10991 ) | ( n10990 & n10991 ) ;
  assign n10993 = ( ~n10985 & n10991 ) | ( ~n10985 & n10992 ) | ( n10991 & n10992 ) ;
  assign n10994 = ( n10761 & n10984 ) | ( n10761 & n10993 ) | ( n10984 & n10993 ) ;
  assign n10995 = ( n10761 & ~n10984 ) | ( n10761 & n10993 ) | ( ~n10984 & n10993 ) ;
  assign n10996 = ( n10984 & ~n10994 ) | ( n10984 & n10995 ) | ( ~n10994 & n10995 ) ;
  assign n10997 = ( n10764 & n10810 ) | ( n10764 & n10996 ) | ( n10810 & n10996 ) ;
  assign n10998 = ( n10764 & ~n10810 ) | ( n10764 & n10996 ) | ( ~n10810 & n10996 ) ;
  assign n10999 = ( n10810 & ~n10997 ) | ( n10810 & n10998 ) | ( ~n10997 & n10998 ) ;
  assign n11000 = n583 & n7841 ;
  assign n11001 = x123 & n587 ;
  assign n11002 = x124 | n11001 ;
  assign n11003 = ( n589 & n11001 ) | ( n589 & n11002 ) | ( n11001 & n11002 ) ;
  assign n11004 = x122 & n676 ;
  assign n11005 = n11003 | n11004 ;
  assign n11006 = ( x14 & n11000 ) | ( x14 & ~n11005 ) | ( n11000 & ~n11005 ) ;
  assign n11007 = ( ~x14 & n11005 ) | ( ~x14 & n11006 ) | ( n11005 & n11006 ) ;
  assign n11008 = ( ~n11000 & n11006 ) | ( ~n11000 & n11007 ) | ( n11006 & n11007 ) ;
  assign n11009 = ( n10776 & n10999 ) | ( n10776 & n11008 ) | ( n10999 & n11008 ) ;
  assign n11010 = ( n10776 & ~n10999 ) | ( n10776 & n11008 ) | ( ~n10999 & n11008 ) ;
  assign n11011 = ( n10999 & ~n11009 ) | ( n10999 & n11010 ) | ( ~n11009 & n11010 ) ;
  assign n11012 = n407 & n8846 ;
  assign n11013 = x126 & n411 ;
  assign n11014 = x127 | n11013 ;
  assign n11015 = ( n413 & n11013 ) | ( n413 & n11014 ) | ( n11013 & n11014 ) ;
  assign n11016 = x125 & n491 ;
  assign n11017 = n11015 | n11016 ;
  assign n11018 = ( x11 & n11012 ) | ( x11 & ~n11017 ) | ( n11012 & ~n11017 ) ;
  assign n11019 = ( ~x11 & n11017 ) | ( ~x11 & n11018 ) | ( n11017 & n11018 ) ;
  assign n11020 = ( ~n11012 & n11018 ) | ( ~n11012 & n11019 ) | ( n11018 & n11019 ) ;
  assign n11021 = ( n10788 & n11011 ) | ( n10788 & n11020 ) | ( n11011 & n11020 ) ;
  assign n11022 = ( n10788 & ~n11011 ) | ( n10788 & n11020 ) | ( ~n11011 & n11020 ) ;
  assign n11023 = ( n11011 & ~n11021 ) | ( n11011 & n11022 ) | ( ~n11021 & n11022 ) ;
  assign n11024 = ( n10796 & n10799 ) | ( n10796 & n11023 ) | ( n10799 & n11023 ) ;
  assign n11025 = ( n10796 & ~n10799 ) | ( n10796 & n11023 ) | ( ~n10799 & n11023 ) ;
  assign n11026 = ( n10799 & ~n11024 ) | ( n10799 & n11025 ) | ( ~n11024 & n11025 ) ;
  assign n11027 = n407 & n8865 ;
  assign n11028 = x127 & n411 ;
  assign n11029 = x126 | n11028 ;
  assign n11030 = ( n491 & n11028 ) | ( n491 & n11029 ) | ( n11028 & n11029 ) ;
  assign n11031 = ( x11 & n11027 ) | ( x11 & ~n11030 ) | ( n11027 & ~n11030 ) ;
  assign n11032 = ( ~x11 & n11030 ) | ( ~x11 & n11031 ) | ( n11030 & n11031 ) ;
  assign n11033 = ( ~n11027 & n11031 ) | ( ~n11027 & n11032 ) | ( n11031 & n11032 ) ;
  assign n11034 = n583 & n8331 ;
  assign n11035 = x124 & n587 ;
  assign n11036 = x125 | n11035 ;
  assign n11037 = ( n589 & n11035 ) | ( n589 & n11036 ) | ( n11035 & n11036 ) ;
  assign n11038 = x123 & n676 ;
  assign n11039 = n11037 | n11038 ;
  assign n11040 = ( x14 & n11034 ) | ( x14 & ~n11039 ) | ( n11034 & ~n11039 ) ;
  assign n11041 = ( ~x14 & n11039 ) | ( ~x14 & n11040 ) | ( n11039 & n11040 ) ;
  assign n11042 = ( ~n11034 & n11040 ) | ( ~n11034 & n11041 ) | ( n11040 & n11041 ) ;
  assign n11043 = n1016 & n6645 ;
  assign n11044 = x118 & n1020 ;
  assign n11045 = x119 | n11044 ;
  assign n11046 = ( n1022 & n11044 ) | ( n1022 & n11045 ) | ( n11044 & n11045 ) ;
  assign n11047 = x117 & n1145 ;
  assign n11048 = n11046 | n11047 ;
  assign n11049 = ( x20 & n11043 ) | ( x20 & ~n11048 ) | ( n11043 & ~n11048 ) ;
  assign n11050 = ( ~x20 & n11048 ) | ( ~x20 & n11049 ) | ( n11048 & n11049 ) ;
  assign n11051 = ( ~n11043 & n11049 ) | ( ~n11043 & n11050 ) | ( n11049 & n11050 ) ;
  assign n11052 = n1297 & n5977 ;
  assign n11053 = x115 & n1301 ;
  assign n11054 = x116 | n11053 ;
  assign n11055 = ( n1303 & n11053 ) | ( n1303 & n11054 ) | ( n11053 & n11054 ) ;
  assign n11056 = x114 & n1426 ;
  assign n11057 = n11055 | n11056 ;
  assign n11058 = ( x23 & n11052 ) | ( x23 & ~n11057 ) | ( n11052 & ~n11057 ) ;
  assign n11059 = ( ~x23 & n11057 ) | ( ~x23 & n11058 ) | ( n11057 & n11058 ) ;
  assign n11060 = ( ~n11052 & n11058 ) | ( ~n11052 & n11059 ) | ( n11058 & n11059 ) ;
  assign n11061 = n1617 & n5542 ;
  assign n11062 = x112 & n1621 ;
  assign n11063 = x113 | n11062 ;
  assign n11064 = ( n1623 & n11062 ) | ( n1623 & n11063 ) | ( n11062 & n11063 ) ;
  assign n11065 = x111 & n1749 ;
  assign n11066 = n11064 | n11065 ;
  assign n11067 = ( x26 & n11061 ) | ( x26 & ~n11066 ) | ( n11061 & ~n11066 ) ;
  assign n11068 = ( ~x26 & n11066 ) | ( ~x26 & n11067 ) | ( n11066 & n11067 ) ;
  assign n11069 = ( ~n11061 & n11067 ) | ( ~n11061 & n11068 ) | ( n11067 & n11068 ) ;
  assign n11070 = n2320 & n4362 ;
  assign n11071 = x106 & n2324 ;
  assign n11072 = x107 | n11071 ;
  assign n11073 = ( n2326 & n11071 ) | ( n2326 & n11072 ) | ( n11071 & n11072 ) ;
  assign n11074 = x105 & n2497 ;
  assign n11075 = n11073 | n11074 ;
  assign n11076 = ( x32 & n11070 ) | ( x32 & ~n11075 ) | ( n11070 & ~n11075 ) ;
  assign n11077 = ( ~x32 & n11075 ) | ( ~x32 & n11076 ) | ( n11075 & n11076 ) ;
  assign n11078 = ( ~n11070 & n11076 ) | ( ~n11070 & n11077 ) | ( n11076 & n11077 ) ;
  assign n11079 = n2766 & n3665 ;
  assign n11080 = x103 & n2770 ;
  assign n11081 = x104 | n11080 ;
  assign n11082 = ( n2772 & n11080 ) | ( n2772 & n11081 ) | ( n11080 & n11081 ) ;
  assign n11083 = x102 & n2943 ;
  assign n11084 = n11082 | n11083 ;
  assign n11085 = ( x35 & n11079 ) | ( x35 & ~n11084 ) | ( n11079 & ~n11084 ) ;
  assign n11086 = ( ~x35 & n11084 ) | ( ~x35 & n11085 ) | ( n11084 & n11085 ) ;
  assign n11087 = ( ~n11079 & n11085 ) | ( ~n11079 & n11086 ) | ( n11085 & n11086 ) ;
  assign n11088 = n3224 & n3326 ;
  assign n11089 = x100 & n3228 ;
  assign n11090 = x101 | n11089 ;
  assign n11091 = ( n3230 & n11089 ) | ( n3230 & n11090 ) | ( n11089 & n11090 ) ;
  assign n11092 = x99 & n3413 ;
  assign n11093 = n11091 | n11092 ;
  assign n11094 = ( x38 & n11088 ) | ( x38 & ~n11093 ) | ( n11088 & ~n11093 ) ;
  assign n11095 = ( ~x38 & n11093 ) | ( ~x38 & n11094 ) | ( n11093 & n11094 ) ;
  assign n11096 = ( ~n11088 & n11094 ) | ( ~n11088 & n11095 ) | ( n11094 & n11095 ) ;
  assign n11097 = n2725 & n3715 ;
  assign n11098 = x97 & n3719 ;
  assign n11099 = x98 | n11098 ;
  assign n11100 = ( n3721 & n11098 ) | ( n3721 & n11099 ) | ( n11098 & n11099 ) ;
  assign n11101 = x96 & n3922 ;
  assign n11102 = n11100 | n11101 ;
  assign n11103 = ( x41 & n11097 ) | ( x41 & ~n11102 ) | ( n11097 & ~n11102 ) ;
  assign n11104 = ( ~x41 & n11102 ) | ( ~x41 & n11103 ) | ( n11102 & n11103 ) ;
  assign n11105 = ( ~n11097 & n11103 ) | ( ~n11097 & n11104 ) | ( n11103 & n11104 ) ;
  assign n11106 = n769 & n7423 ;
  assign n11107 = x79 & n7427 ;
  assign n11108 = x80 | n11107 ;
  assign n11109 = ( n7429 & n11107 ) | ( n7429 & n11108 ) | ( n11107 & n11108 ) ;
  assign n11110 = x78 & n7708 ;
  assign n11111 = n11109 | n11110 ;
  assign n11112 = ( x59 & n11106 ) | ( x59 & ~n11111 ) | ( n11106 & ~n11111 ) ;
  assign n11113 = ( ~x59 & n11111 ) | ( ~x59 & n11112 ) | ( n11111 & n11112 ) ;
  assign n11114 = ( ~n11106 & n11112 ) | ( ~n11106 & n11113 ) | ( n11112 & n11113 ) ;
  assign n11115 = n569 & n8154 ;
  assign n11116 = x76 & n8158 ;
  assign n11117 = x77 | n11116 ;
  assign n11118 = ( n8160 & n11116 ) | ( n8160 & n11117 ) | ( n11116 & n11117 ) ;
  assign n11119 = x75 & n8439 ;
  assign n11120 = n11118 | n11119 ;
  assign n11121 = ( x62 & n11115 ) | ( x62 & ~n11120 ) | ( n11115 & ~n11120 ) ;
  assign n11122 = ( ~x62 & n11120 ) | ( ~x62 & n11121 ) | ( n11120 & n11121 ) ;
  assign n11123 = ( ~n11115 & n11121 ) | ( ~n11115 & n11122 ) | ( n11121 & n11122 ) ;
  assign n11124 = x73 & n8927 ;
  assign n11125 = ( ~x74 & n8693 ) | ( ~x74 & n8927 ) | ( n8693 & n8927 ) ;
  assign n11126 = ( n8693 & n11124 ) | ( n8693 & ~n11125 ) | ( n11124 & ~n11125 ) ;
  assign n11127 = ( n10868 & n11123 ) | ( n10868 & ~n11126 ) | ( n11123 & ~n11126 ) ;
  assign n11128 = ( ~n10868 & n11123 ) | ( ~n10868 & n11126 ) | ( n11123 & n11126 ) ;
  assign n11129 = ( ~n11123 & n11127 ) | ( ~n11123 & n11128 ) | ( n11127 & n11128 ) ;
  assign n11130 = ( n10871 & ~n11114 ) | ( n10871 & n11129 ) | ( ~n11114 & n11129 ) ;
  assign n11131 = ( n10871 & n11114 ) | ( n10871 & n11129 ) | ( n11114 & n11129 ) ;
  assign n11132 = ( n11114 & n11130 ) | ( n11114 & ~n11131 ) | ( n11130 & ~n11131 ) ;
  assign n11133 = n1082 & n6713 ;
  assign n11134 = x82 & n6717 ;
  assign n11135 = x83 | n11134 ;
  assign n11136 = ( n6719 & n11134 ) | ( n6719 & n11135 ) | ( n11134 & n11135 ) ;
  assign n11137 = x81 & n6980 ;
  assign n11138 = n11136 | n11137 ;
  assign n11139 = ( x56 & n11133 ) | ( x56 & ~n11138 ) | ( n11133 & ~n11138 ) ;
  assign n11140 = ( ~x56 & n11138 ) | ( ~x56 & n11139 ) | ( n11138 & n11139 ) ;
  assign n11141 = ( ~n11133 & n11139 ) | ( ~n11133 & n11140 ) | ( n11139 & n11140 ) ;
  assign n11142 = ( n10883 & n11132 ) | ( n10883 & n11141 ) | ( n11132 & n11141 ) ;
  assign n11143 = ( ~n10883 & n11132 ) | ( ~n10883 & n11141 ) | ( n11132 & n11141 ) ;
  assign n11144 = ( n10883 & ~n11142 ) | ( n10883 & n11143 ) | ( ~n11142 & n11143 ) ;
  assign n11145 = n1366 & n6027 ;
  assign n11146 = x85 & n6031 ;
  assign n11147 = x86 | n11146 ;
  assign n11148 = ( n6033 & n11146 ) | ( n6033 & n11147 ) | ( n11146 & n11147 ) ;
  assign n11149 = x84 & n6303 ;
  assign n11150 = n11148 | n11149 ;
  assign n11151 = ( x53 & n11145 ) | ( x53 & ~n11150 ) | ( n11145 & ~n11150 ) ;
  assign n11152 = ( ~x53 & n11150 ) | ( ~x53 & n11151 ) | ( n11150 & n11151 ) ;
  assign n11153 = ( ~n11145 & n11151 ) | ( ~n11145 & n11152 ) | ( n11151 & n11152 ) ;
  assign n11154 = ( n10895 & n11144 ) | ( n10895 & n11153 ) | ( n11144 & n11153 ) ;
  assign n11155 = ( ~n10895 & n11144 ) | ( ~n10895 & n11153 ) | ( n11144 & n11153 ) ;
  assign n11156 = ( n10895 & ~n11154 ) | ( n10895 & n11155 ) | ( ~n11154 & n11155 ) ;
  assign n11157 = n1585 & n5374 ;
  assign n11158 = x88 & n5378 ;
  assign n11159 = x89 | n11158 ;
  assign n11160 = ( n5380 & n11158 ) | ( n5380 & n11159 ) | ( n11158 & n11159 ) ;
  assign n11161 = x87 & n5638 ;
  assign n11162 = n11160 | n11161 ;
  assign n11163 = ( x50 & n11157 ) | ( x50 & ~n11162 ) | ( n11157 & ~n11162 ) ;
  assign n11164 = ( ~x50 & n11162 ) | ( ~x50 & n11163 ) | ( n11162 & n11163 ) ;
  assign n11165 = ( ~n11157 & n11163 ) | ( ~n11157 & n11164 ) | ( n11163 & n11164 ) ;
  assign n11166 = ( n10907 & n11156 ) | ( n10907 & n11165 ) | ( n11156 & n11165 ) ;
  assign n11167 = ( ~n10907 & n11156 ) | ( ~n10907 & n11165 ) | ( n11156 & n11165 ) ;
  assign n11168 = ( n10907 & ~n11166 ) | ( n10907 & n11167 ) | ( ~n11166 & n11167 ) ;
  assign n11169 = n2042 & n4787 ;
  assign n11170 = x91 & n4791 ;
  assign n11171 = x92 | n11170 ;
  assign n11172 = ( n4793 & n11170 ) | ( n4793 & n11171 ) | ( n11170 & n11171 ) ;
  assign n11173 = x90 & n5030 ;
  assign n11174 = n11172 | n11173 ;
  assign n11175 = ( x47 & n11169 ) | ( x47 & ~n11174 ) | ( n11169 & ~n11174 ) ;
  assign n11176 = ( ~x47 & n11174 ) | ( ~x47 & n11175 ) | ( n11174 & n11175 ) ;
  assign n11177 = ( ~n11169 & n11175 ) | ( ~n11169 & n11176 ) | ( n11175 & n11176 ) ;
  assign n11178 = ( n10910 & n11168 ) | ( n10910 & n11177 ) | ( n11168 & n11177 ) ;
  assign n11179 = ( ~n10910 & n11168 ) | ( ~n10910 & n11177 ) | ( n11168 & n11177 ) ;
  assign n11180 = ( n10910 & ~n11178 ) | ( n10910 & n11179 ) | ( ~n11178 & n11179 ) ;
  assign n11181 = n2434 & n4227 ;
  assign n11182 = x94 & n4231 ;
  assign n11183 = x95 | n11182 ;
  assign n11184 = ( n4233 & n11182 ) | ( n4233 & n11183 ) | ( n11182 & n11183 ) ;
  assign n11185 = x93 & n4470 ;
  assign n11186 = n11184 | n11185 ;
  assign n11187 = ( x44 & n11181 ) | ( x44 & ~n11186 ) | ( n11181 & ~n11186 ) ;
  assign n11188 = ( ~x44 & n11186 ) | ( ~x44 & n11187 ) | ( n11186 & n11187 ) ;
  assign n11189 = ( ~n11181 & n11187 ) | ( ~n11181 & n11188 ) | ( n11187 & n11188 ) ;
  assign n11190 = ( n10922 & n11180 ) | ( n10922 & n11189 ) | ( n11180 & n11189 ) ;
  assign n11191 = ( ~n10922 & n11180 ) | ( ~n10922 & n11189 ) | ( n11180 & n11189 ) ;
  assign n11192 = ( n10922 & ~n11190 ) | ( n10922 & n11191 ) | ( ~n11190 & n11191 ) ;
  assign n11193 = ( n10934 & n11105 ) | ( n10934 & n11192 ) | ( n11105 & n11192 ) ;
  assign n11194 = ( n10934 & ~n11105 ) | ( n10934 & n11192 ) | ( ~n11105 & n11192 ) ;
  assign n11195 = ( n11105 & ~n11193 ) | ( n11105 & n11194 ) | ( ~n11193 & n11194 ) ;
  assign n11196 = ( n10937 & n11096 ) | ( n10937 & n11195 ) | ( n11096 & n11195 ) ;
  assign n11197 = ( n10937 & ~n11096 ) | ( n10937 & n11195 ) | ( ~n11096 & n11195 ) ;
  assign n11198 = ( n11096 & ~n11196 ) | ( n11096 & n11197 ) | ( ~n11196 & n11197 ) ;
  assign n11199 = ( n10940 & n11087 ) | ( n10940 & n11198 ) | ( n11087 & n11198 ) ;
  assign n11200 = ( n10940 & ~n11087 ) | ( n10940 & n11198 ) | ( ~n11087 & n11198 ) ;
  assign n11201 = ( n11087 & ~n11199 ) | ( n11087 & n11200 ) | ( ~n11199 & n11200 ) ;
  assign n11202 = ( n10952 & n11078 ) | ( n10952 & n11201 ) | ( n11078 & n11201 ) ;
  assign n11203 = ( n10952 & ~n11078 ) | ( n10952 & n11201 ) | ( ~n11078 & n11201 ) ;
  assign n11204 = ( n11078 & ~n11202 ) | ( n11078 & n11203 ) | ( ~n11202 & n11203 ) ;
  assign n11205 = n1949 & n4934 ;
  assign n11206 = x109 & n1953 ;
  assign n11207 = x110 | n11206 ;
  assign n11208 = ( n1955 & n11206 ) | ( n1955 & n11207 ) | ( n11206 & n11207 ) ;
  assign n11209 = x108 & n2114 ;
  assign n11210 = n11208 | n11209 ;
  assign n11211 = ( x29 & n11205 ) | ( x29 & ~n11210 ) | ( n11205 & ~n11210 ) ;
  assign n11212 = ( ~x29 & n11210 ) | ( ~x29 & n11211 ) | ( n11210 & n11211 ) ;
  assign n11213 = ( ~n11205 & n11211 ) | ( ~n11205 & n11212 ) | ( n11211 & n11212 ) ;
  assign n11214 = ( n10964 & n11204 ) | ( n10964 & n11213 ) | ( n11204 & n11213 ) ;
  assign n11215 = ( n10964 & ~n11204 ) | ( n10964 & n11213 ) | ( ~n11204 & n11213 ) ;
  assign n11216 = ( n11204 & ~n11214 ) | ( n11204 & n11215 ) | ( ~n11214 & n11215 ) ;
  assign n11217 = ( n10976 & n11069 ) | ( n10976 & n11216 ) | ( n11069 & n11216 ) ;
  assign n11218 = ( n10976 & ~n11069 ) | ( n10976 & n11216 ) | ( ~n11069 & n11216 ) ;
  assign n11219 = ( n11069 & ~n11217 ) | ( n11069 & n11218 ) | ( ~n11217 & n11218 ) ;
  assign n11220 = ( n10979 & n11060 ) | ( n10979 & n11219 ) | ( n11060 & n11219 ) ;
  assign n11221 = ( n10979 & ~n11060 ) | ( n10979 & n11219 ) | ( ~n11060 & n11219 ) ;
  assign n11222 = ( n11060 & ~n11220 ) | ( n11060 & n11221 ) | ( ~n11220 & n11221 ) ;
  assign n11223 = ( n10982 & n11051 ) | ( n10982 & n11222 ) | ( n11051 & n11222 ) ;
  assign n11224 = ( n10982 & ~n11051 ) | ( n10982 & n11222 ) | ( ~n11051 & n11222 ) ;
  assign n11225 = ( n11051 & ~n11223 ) | ( n11051 & n11224 ) | ( ~n11223 & n11224 ) ;
  assign n11226 = n810 & n7582 ;
  assign n11227 = x121 & n814 ;
  assign n11228 = x122 | n11227 ;
  assign n11229 = ( n816 & n11227 ) | ( n816 & n11228 ) | ( n11227 & n11228 ) ;
  assign n11230 = x120 & n885 ;
  assign n11231 = n11229 | n11230 ;
  assign n11232 = ( x17 & n11226 ) | ( x17 & ~n11231 ) | ( n11226 & ~n11231 ) ;
  assign n11233 = ( ~x17 & n11231 ) | ( ~x17 & n11232 ) | ( n11231 & n11232 ) ;
  assign n11234 = ( ~n11226 & n11232 ) | ( ~n11226 & n11233 ) | ( n11232 & n11233 ) ;
  assign n11235 = ( n10994 & n11225 ) | ( n10994 & n11234 ) | ( n11225 & n11234 ) ;
  assign n11236 = ( n10994 & ~n11225 ) | ( n10994 & n11234 ) | ( ~n11225 & n11234 ) ;
  assign n11237 = ( n11225 & ~n11235 ) | ( n11225 & n11236 ) | ( ~n11235 & n11236 ) ;
  assign n11238 = ( n10997 & n11042 ) | ( n10997 & n11237 ) | ( n11042 & n11237 ) ;
  assign n11239 = ( n10997 & ~n11042 ) | ( n10997 & n11237 ) | ( ~n11042 & n11237 ) ;
  assign n11240 = ( n11042 & ~n11238 ) | ( n11042 & n11239 ) | ( ~n11238 & n11239 ) ;
  assign n11241 = ( n11009 & n11033 ) | ( n11009 & n11240 ) | ( n11033 & n11240 ) ;
  assign n11242 = ( ~n11009 & n11033 ) | ( ~n11009 & n11240 ) | ( n11033 & n11240 ) ;
  assign n11243 = ( n11009 & ~n11241 ) | ( n11009 & n11242 ) | ( ~n11241 & n11242 ) ;
  assign n11244 = ( n11021 & n11024 ) | ( n11021 & n11243 ) | ( n11024 & n11243 ) ;
  assign n11245 = ( n11021 & ~n11024 ) | ( n11021 & n11243 ) | ( ~n11024 & n11243 ) ;
  assign n11246 = ( n11024 & ~n11244 ) | ( n11024 & n11245 ) | ( ~n11244 & n11245 ) ;
  assign n11247 = n583 & n8587 ;
  assign n11248 = x125 & n587 ;
  assign n11249 = x126 | n11248 ;
  assign n11250 = ( n589 & n11248 ) | ( n589 & n11249 ) | ( n11248 & n11249 ) ;
  assign n11251 = x124 & n676 ;
  assign n11252 = n11250 | n11251 ;
  assign n11253 = ( x14 & n11247 ) | ( x14 & ~n11252 ) | ( n11247 & ~n11252 ) ;
  assign n11254 = ( ~x14 & n11252 ) | ( ~x14 & n11253 ) | ( n11252 & n11253 ) ;
  assign n11255 = ( ~n11247 & n11253 ) | ( ~n11247 & n11254 ) | ( n11253 & n11254 ) ;
  assign n11256 = n810 & n7597 ;
  assign n11257 = x122 & n814 ;
  assign n11258 = x123 | n11257 ;
  assign n11259 = ( n816 & n11257 ) | ( n816 & n11258 ) | ( n11257 & n11258 ) ;
  assign n11260 = x121 & n885 ;
  assign n11261 = n11259 | n11260 ;
  assign n11262 = ( x17 & n11256 ) | ( x17 & ~n11261 ) | ( n11256 & ~n11261 ) ;
  assign n11263 = ( ~x17 & n11261 ) | ( ~x17 & n11262 ) | ( n11261 & n11262 ) ;
  assign n11264 = ( ~n11256 & n11262 ) | ( ~n11256 & n11263 ) | ( n11262 & n11263 ) ;
  assign n11265 = n1016 & n7098 ;
  assign n11266 = x119 & n1020 ;
  assign n11267 = x120 | n11266 ;
  assign n11268 = ( n1022 & n11266 ) | ( n1022 & n11267 ) | ( n11266 & n11267 ) ;
  assign n11269 = x118 & n1145 ;
  assign n11270 = n11268 | n11269 ;
  assign n11271 = ( x20 & n11265 ) | ( x20 & ~n11270 ) | ( n11265 & ~n11270 ) ;
  assign n11272 = ( ~x20 & n11270 ) | ( ~x20 & n11271 ) | ( n11270 & n11271 ) ;
  assign n11273 = ( ~n11265 & n11271 ) | ( ~n11265 & n11272 ) | ( n11271 & n11272 ) ;
  assign n11274 = n1617 & n5750 ;
  assign n11275 = x113 & n1621 ;
  assign n11276 = x114 | n11275 ;
  assign n11277 = ( n1623 & n11275 ) | ( n1623 & n11276 ) | ( n11275 & n11276 ) ;
  assign n11278 = x112 & n1749 ;
  assign n11279 = n11277 | n11278 ;
  assign n11280 = ( x26 & n11274 ) | ( x26 & ~n11279 ) | ( n11274 & ~n11279 ) ;
  assign n11281 = ( ~x26 & n11279 ) | ( ~x26 & n11280 ) | ( n11279 & n11280 ) ;
  assign n11282 = ( ~n11274 & n11280 ) | ( ~n11274 & n11281 ) | ( n11280 & n11281 ) ;
  assign n11283 = n1949 & n5130 ;
  assign n11284 = x110 & n1953 ;
  assign n11285 = x111 | n11284 ;
  assign n11286 = ( n1955 & n11284 ) | ( n1955 & n11285 ) | ( n11284 & n11285 ) ;
  assign n11287 = x109 & n2114 ;
  assign n11288 = n11286 | n11287 ;
  assign n11289 = ( x29 & n11283 ) | ( x29 & ~n11288 ) | ( n11283 & ~n11288 ) ;
  assign n11290 = ( ~x29 & n11288 ) | ( ~x29 & n11289 ) | ( n11288 & n11289 ) ;
  assign n11291 = ( ~n11283 & n11289 ) | ( ~n11283 & n11290 ) | ( n11289 & n11290 ) ;
  assign n11292 = n2320 & n4377 ;
  assign n11293 = x107 & n2324 ;
  assign n11294 = x108 | n11293 ;
  assign n11295 = ( n2326 & n11293 ) | ( n2326 & n11294 ) | ( n11293 & n11294 ) ;
  assign n11296 = x106 & n2497 ;
  assign n11297 = n11295 | n11296 ;
  assign n11298 = ( x32 & n11292 ) | ( x32 & ~n11297 ) | ( n11292 & ~n11297 ) ;
  assign n11299 = ( ~x32 & n11297 ) | ( ~x32 & n11298 ) | ( n11297 & n11298 ) ;
  assign n11300 = ( ~n11292 & n11298 ) | ( ~n11292 & n11299 ) | ( n11298 & n11299 ) ;
  assign n11301 = n2766 & n3998 ;
  assign n11302 = x104 & n2770 ;
  assign n11303 = x105 | n11302 ;
  assign n11304 = ( n2772 & n11302 ) | ( n2772 & n11303 ) | ( n11302 & n11303 ) ;
  assign n11305 = x103 & n2943 ;
  assign n11306 = n11304 | n11305 ;
  assign n11307 = ( x35 & n11301 ) | ( x35 & ~n11306 ) | ( n11301 & ~n11306 ) ;
  assign n11308 = ( ~x35 & n11306 ) | ( ~x35 & n11307 ) | ( n11306 & n11307 ) ;
  assign n11309 = ( ~n11301 & n11307 ) | ( ~n11301 & n11308 ) | ( n11307 & n11308 ) ;
  assign n11310 = n1701 & n5374 ;
  assign n11311 = x89 & n5378 ;
  assign n11312 = x90 | n11311 ;
  assign n11313 = ( n5380 & n11311 ) | ( n5380 & n11312 ) | ( n11311 & n11312 ) ;
  assign n11314 = x88 & n5638 ;
  assign n11315 = n11313 | n11314 ;
  assign n11316 = ( x50 & n11310 ) | ( x50 & ~n11315 ) | ( n11310 & ~n11315 ) ;
  assign n11317 = ( ~x50 & n11315 ) | ( ~x50 & n11316 ) | ( n11315 & n11316 ) ;
  assign n11318 = ( ~n11310 & n11316 ) | ( ~n11310 & n11317 ) | ( n11316 & n11317 ) ;
  assign n11319 = n1466 & n6027 ;
  assign n11320 = x86 & n6031 ;
  assign n11321 = x87 | n11320 ;
  assign n11322 = ( n6033 & n11320 ) | ( n6033 & n11321 ) | ( n11320 & n11321 ) ;
  assign n11323 = x85 & n6303 ;
  assign n11324 = n11322 | n11323 ;
  assign n11325 = ( x53 & n11319 ) | ( x53 & ~n11324 ) | ( n11319 & ~n11324 ) ;
  assign n11326 = ( ~x53 & n11324 ) | ( ~x53 & n11325 ) | ( n11324 & n11325 ) ;
  assign n11327 = ( ~n11319 & n11325 ) | ( ~n11319 & n11326 ) | ( n11325 & n11326 ) ;
  assign n11328 = x74 & n8927 ;
  assign n11329 = ( ~x75 & n8693 ) | ( ~x75 & n8927 ) | ( n8693 & n8927 ) ;
  assign n11330 = ( n8693 & n11328 ) | ( n8693 & ~n11329 ) | ( n11328 & ~n11329 ) ;
  assign n11331 = ( ~n11126 & n11127 ) | ( ~n11126 & n11330 ) | ( n11127 & n11330 ) ;
  assign n11332 = ( n11126 & n11127 ) | ( n11126 & n11330 ) | ( n11127 & n11330 ) ;
  assign n11333 = ( n11126 & n11331 ) | ( n11126 & ~n11332 ) | ( n11331 & ~n11332 ) ;
  assign n11334 = n910 & n7423 ;
  assign n11335 = x80 & n7427 ;
  assign n11336 = x81 | n11335 ;
  assign n11337 = ( n7429 & n11335 ) | ( n7429 & n11336 ) | ( n11335 & n11336 ) ;
  assign n11338 = x79 & n7708 ;
  assign n11339 = n11337 | n11338 ;
  assign n11340 = ( x59 & n11334 ) | ( x59 & ~n11339 ) | ( n11334 & ~n11339 ) ;
  assign n11341 = ( ~x59 & n11339 ) | ( ~x59 & n11340 ) | ( n11339 & n11340 ) ;
  assign n11342 = ( ~n11334 & n11340 ) | ( ~n11334 & n11341 ) | ( n11340 & n11341 ) ;
  assign n11343 = n637 & n8154 ;
  assign n11344 = x77 & n8158 ;
  assign n11345 = x78 | n11344 ;
  assign n11346 = ( n8160 & n11344 ) | ( n8160 & n11345 ) | ( n11344 & n11345 ) ;
  assign n11347 = x76 & n8439 ;
  assign n11348 = n11346 | n11347 ;
  assign n11349 = ( x62 & n11343 ) | ( x62 & ~n11348 ) | ( n11343 & ~n11348 ) ;
  assign n11350 = ( ~x62 & n11348 ) | ( ~x62 & n11349 ) | ( n11348 & n11349 ) ;
  assign n11351 = ( ~n11343 & n11349 ) | ( ~n11343 & n11350 ) | ( n11349 & n11350 ) ;
  assign n11352 = ( ~n11333 & n11342 ) | ( ~n11333 & n11351 ) | ( n11342 & n11351 ) ;
  assign n11353 = ( n11342 & n11351 ) | ( n11342 & ~n11352 ) | ( n11351 & ~n11352 ) ;
  assign n11354 = ( n11333 & n11352 ) | ( n11333 & ~n11353 ) | ( n11352 & ~n11353 ) ;
  assign n11355 = n1097 & n6713 ;
  assign n11356 = x83 & n6717 ;
  assign n11357 = x84 | n11356 ;
  assign n11358 = ( n6719 & n11356 ) | ( n6719 & n11357 ) | ( n11356 & n11357 ) ;
  assign n11359 = x82 & n6980 ;
  assign n11360 = n11358 | n11359 ;
  assign n11361 = ( x56 & n11355 ) | ( x56 & ~n11360 ) | ( n11355 & ~n11360 ) ;
  assign n11362 = ( ~x56 & n11360 ) | ( ~x56 & n11361 ) | ( n11360 & n11361 ) ;
  assign n11363 = ( ~n11355 & n11361 ) | ( ~n11355 & n11362 ) | ( n11361 & n11362 ) ;
  assign n11364 = ( n11130 & n11354 ) | ( n11130 & ~n11363 ) | ( n11354 & ~n11363 ) ;
  assign n11365 = ( ~n11130 & n11354 ) | ( ~n11130 & n11363 ) | ( n11354 & n11363 ) ;
  assign n11366 = ( ~n11354 & n11364 ) | ( ~n11354 & n11365 ) | ( n11364 & n11365 ) ;
  assign n11367 = ( n11142 & n11327 ) | ( n11142 & n11366 ) | ( n11327 & n11366 ) ;
  assign n11368 = ( n11142 & ~n11327 ) | ( n11142 & n11366 ) | ( ~n11327 & n11366 ) ;
  assign n11369 = ( n11327 & ~n11367 ) | ( n11327 & n11368 ) | ( ~n11367 & n11368 ) ;
  assign n11370 = ( n11154 & n11318 ) | ( n11154 & n11369 ) | ( n11318 & n11369 ) ;
  assign n11371 = ( n11154 & ~n11318 ) | ( n11154 & n11369 ) | ( ~n11318 & n11369 ) ;
  assign n11372 = ( n11318 & ~n11370 ) | ( n11318 & n11371 ) | ( ~n11370 & n11371 ) ;
  assign n11373 = n2057 & n4787 ;
  assign n11374 = x92 & n4791 ;
  assign n11375 = x93 | n11374 ;
  assign n11376 = ( n4793 & n11374 ) | ( n4793 & n11375 ) | ( n11374 & n11375 ) ;
  assign n11377 = x91 & n5030 ;
  assign n11378 = n11376 | n11377 ;
  assign n11379 = ( x47 & n11373 ) | ( x47 & ~n11378 ) | ( n11373 & ~n11378 ) ;
  assign n11380 = ( ~x47 & n11378 ) | ( ~x47 & n11379 ) | ( n11378 & n11379 ) ;
  assign n11381 = ( ~n11373 & n11379 ) | ( ~n11373 & n11380 ) | ( n11379 & n11380 ) ;
  assign n11382 = ( n11166 & n11372 ) | ( n11166 & n11381 ) | ( n11372 & n11381 ) ;
  assign n11383 = ( ~n11166 & n11372 ) | ( ~n11166 & n11381 ) | ( n11372 & n11381 ) ;
  assign n11384 = ( n11166 & ~n11382 ) | ( n11166 & n11383 ) | ( ~n11382 & n11383 ) ;
  assign n11385 = n2449 & n4227 ;
  assign n11386 = x95 & n4231 ;
  assign n11387 = x96 | n11386 ;
  assign n11388 = ( n4233 & n11386 ) | ( n4233 & n11387 ) | ( n11386 & n11387 ) ;
  assign n11389 = x94 & n4470 ;
  assign n11390 = n11388 | n11389 ;
  assign n11391 = ( x44 & n11385 ) | ( x44 & ~n11390 ) | ( n11385 & ~n11390 ) ;
  assign n11392 = ( ~x44 & n11390 ) | ( ~x44 & n11391 ) | ( n11390 & n11391 ) ;
  assign n11393 = ( ~n11385 & n11391 ) | ( ~n11385 & n11392 ) | ( n11391 & n11392 ) ;
  assign n11394 = ( n11178 & n11384 ) | ( n11178 & n11393 ) | ( n11384 & n11393 ) ;
  assign n11395 = ( ~n11178 & n11384 ) | ( ~n11178 & n11393 ) | ( n11384 & n11393 ) ;
  assign n11396 = ( n11178 & ~n11394 ) | ( n11178 & n11395 ) | ( ~n11394 & n11395 ) ;
  assign n11397 = n2877 & n3715 ;
  assign n11398 = x98 & n3719 ;
  assign n11399 = x99 | n11398 ;
  assign n11400 = ( n3721 & n11398 ) | ( n3721 & n11399 ) | ( n11398 & n11399 ) ;
  assign n11401 = x97 & n3922 ;
  assign n11402 = n11400 | n11401 ;
  assign n11403 = ( x41 & n11397 ) | ( x41 & ~n11402 ) | ( n11397 & ~n11402 ) ;
  assign n11404 = ( ~x41 & n11402 ) | ( ~x41 & n11403 ) | ( n11402 & n11403 ) ;
  assign n11405 = ( ~n11397 & n11403 ) | ( ~n11397 & n11404 ) | ( n11403 & n11404 ) ;
  assign n11406 = ( n11190 & n11396 ) | ( n11190 & n11405 ) | ( n11396 & n11405 ) ;
  assign n11407 = ( n11190 & ~n11396 ) | ( n11190 & n11405 ) | ( ~n11396 & n11405 ) ;
  assign n11408 = ( n11396 & ~n11406 ) | ( n11396 & n11407 ) | ( ~n11406 & n11407 ) ;
  assign n11409 = n3224 & n3486 ;
  assign n11410 = x101 & n3228 ;
  assign n11411 = x102 | n11410 ;
  assign n11412 = ( n3230 & n11410 ) | ( n3230 & n11411 ) | ( n11410 & n11411 ) ;
  assign n11413 = x100 & n3413 ;
  assign n11414 = n11412 | n11413 ;
  assign n11415 = ( x38 & n11409 ) | ( x38 & ~n11414 ) | ( n11409 & ~n11414 ) ;
  assign n11416 = ( ~x38 & n11414 ) | ( ~x38 & n11415 ) | ( n11414 & n11415 ) ;
  assign n11417 = ( ~n11409 & n11415 ) | ( ~n11409 & n11416 ) | ( n11415 & n11416 ) ;
  assign n11418 = ( n11193 & n11408 ) | ( n11193 & n11417 ) | ( n11408 & n11417 ) ;
  assign n11419 = ( ~n11193 & n11408 ) | ( ~n11193 & n11417 ) | ( n11408 & n11417 ) ;
  assign n11420 = ( n11193 & ~n11418 ) | ( n11193 & n11419 ) | ( ~n11418 & n11419 ) ;
  assign n11421 = ( n11196 & n11309 ) | ( n11196 & n11420 ) | ( n11309 & n11420 ) ;
  assign n11422 = ( n11196 & ~n11309 ) | ( n11196 & n11420 ) | ( ~n11309 & n11420 ) ;
  assign n11423 = ( n11309 & ~n11421 ) | ( n11309 & n11422 ) | ( ~n11421 & n11422 ) ;
  assign n11424 = ( n11199 & n11300 ) | ( n11199 & n11423 ) | ( n11300 & n11423 ) ;
  assign n11425 = ( n11199 & ~n11300 ) | ( n11199 & n11423 ) | ( ~n11300 & n11423 ) ;
  assign n11426 = ( n11300 & ~n11424 ) | ( n11300 & n11425 ) | ( ~n11424 & n11425 ) ;
  assign n11427 = ( n11202 & n11291 ) | ( n11202 & n11426 ) | ( n11291 & n11426 ) ;
  assign n11428 = ( n11202 & ~n11291 ) | ( n11202 & n11426 ) | ( ~n11291 & n11426 ) ;
  assign n11429 = ( n11291 & ~n11427 ) | ( n11291 & n11428 ) | ( ~n11427 & n11428 ) ;
  assign n11430 = ( n11214 & n11282 ) | ( n11214 & n11429 ) | ( n11282 & n11429 ) ;
  assign n11431 = ( ~n11214 & n11282 ) | ( ~n11214 & n11429 ) | ( n11282 & n11429 ) ;
  assign n11432 = ( n11214 & ~n11430 ) | ( n11214 & n11431 ) | ( ~n11430 & n11431 ) ;
  assign n11433 = n1297 & n6201 ;
  assign n11434 = x116 & n1301 ;
  assign n11435 = x117 | n11434 ;
  assign n11436 = ( n1303 & n11434 ) | ( n1303 & n11435 ) | ( n11434 & n11435 ) ;
  assign n11437 = x115 & n1426 ;
  assign n11438 = n11436 | n11437 ;
  assign n11439 = ( x23 & n11433 ) | ( x23 & ~n11438 ) | ( n11433 & ~n11438 ) ;
  assign n11440 = ( ~x23 & n11438 ) | ( ~x23 & n11439 ) | ( n11438 & n11439 ) ;
  assign n11441 = ( ~n11433 & n11439 ) | ( ~n11433 & n11440 ) | ( n11439 & n11440 ) ;
  assign n11442 = ( n11217 & n11432 ) | ( n11217 & n11441 ) | ( n11432 & n11441 ) ;
  assign n11443 = ( n11217 & ~n11432 ) | ( n11217 & n11441 ) | ( ~n11432 & n11441 ) ;
  assign n11444 = ( n11432 & ~n11442 ) | ( n11432 & n11443 ) | ( ~n11442 & n11443 ) ;
  assign n11445 = ( n11220 & n11273 ) | ( n11220 & n11444 ) | ( n11273 & n11444 ) ;
  assign n11446 = ( n11220 & ~n11273 ) | ( n11220 & n11444 ) | ( ~n11273 & n11444 ) ;
  assign n11447 = ( n11273 & ~n11445 ) | ( n11273 & n11446 ) | ( ~n11445 & n11446 ) ;
  assign n11448 = ( n11223 & n11264 ) | ( n11223 & n11447 ) | ( n11264 & n11447 ) ;
  assign n11449 = ( n11223 & ~n11264 ) | ( n11223 & n11447 ) | ( ~n11264 & n11447 ) ;
  assign n11450 = ( n11264 & ~n11448 ) | ( n11264 & n11449 ) | ( ~n11448 & n11449 ) ;
  assign n11451 = ( n11235 & n11255 ) | ( n11235 & n11450 ) | ( n11255 & n11450 ) ;
  assign n11452 = ( ~n11235 & n11255 ) | ( ~n11235 & n11450 ) | ( n11255 & n11450 ) ;
  assign n11453 = ( n11235 & ~n11451 ) | ( n11235 & n11452 ) | ( ~n11451 & n11452 ) ;
  assign n11454 = n407 & n8862 ;
  assign n11455 = ( x127 & n491 ) | ( x127 & n11454 ) | ( n491 & n11454 ) ;
  assign n11456 = x11 | n11455 ;
  assign n11457 = ~x11 & n11455 ;
  assign n11458 = ( ~n11455 & n11456 ) | ( ~n11455 & n11457 ) | ( n11456 & n11457 ) ;
  assign n11459 = ( n11238 & n11453 ) | ( n11238 & n11458 ) | ( n11453 & n11458 ) ;
  assign n11460 = ( n11238 & ~n11453 ) | ( n11238 & n11458 ) | ( ~n11453 & n11458 ) ;
  assign n11461 = ( n11453 & ~n11459 ) | ( n11453 & n11460 ) | ( ~n11459 & n11460 ) ;
  assign n11462 = ( n11241 & n11244 ) | ( n11241 & n11461 ) | ( n11244 & n11461 ) ;
  assign n11463 = ( n11241 & ~n11244 ) | ( n11241 & n11461 ) | ( ~n11244 & n11461 ) ;
  assign n11464 = ( n11244 & ~n11462 ) | ( n11244 & n11463 ) | ( ~n11462 & n11463 ) ;
  assign n11465 = n1016 & n7113 ;
  assign n11466 = x120 & n1020 ;
  assign n11467 = x121 | n11466 ;
  assign n11468 = ( n1022 & n11466 ) | ( n1022 & n11467 ) | ( n11466 & n11467 ) ;
  assign n11469 = x119 & n1145 ;
  assign n11470 = n11468 | n11469 ;
  assign n11471 = ( x20 & n11465 ) | ( x20 & ~n11470 ) | ( n11465 & ~n11470 ) ;
  assign n11472 = ( ~x20 & n11470 ) | ( ~x20 & n11471 ) | ( n11470 & n11471 ) ;
  assign n11473 = ( ~n11465 & n11471 ) | ( ~n11465 & n11472 ) | ( n11471 & n11472 ) ;
  assign n11474 = n1617 & n5765 ;
  assign n11475 = x114 & n1621 ;
  assign n11476 = x115 | n11475 ;
  assign n11477 = ( n1623 & n11475 ) | ( n1623 & n11476 ) | ( n11475 & n11476 ) ;
  assign n11478 = x113 & n1749 ;
  assign n11479 = n11477 | n11478 ;
  assign n11480 = ( x26 & n11474 ) | ( x26 & ~n11479 ) | ( n11474 & ~n11479 ) ;
  assign n11481 = ( ~x26 & n11479 ) | ( ~x26 & n11480 ) | ( n11479 & n11480 ) ;
  assign n11482 = ( ~n11474 & n11480 ) | ( ~n11474 & n11481 ) | ( n11480 & n11481 ) ;
  assign n11483 = n2766 & n4013 ;
  assign n11484 = x105 & n2770 ;
  assign n11485 = x106 | n11484 ;
  assign n11486 = ( n2772 & n11484 ) | ( n2772 & n11485 ) | ( n11484 & n11485 ) ;
  assign n11487 = x104 & n2943 ;
  assign n11488 = n11486 | n11487 ;
  assign n11489 = ( x35 & n11483 ) | ( x35 & ~n11488 ) | ( n11483 & ~n11488 ) ;
  assign n11490 = ( ~x35 & n11488 ) | ( ~x35 & n11489 ) | ( n11488 & n11489 ) ;
  assign n11491 = ( ~n11483 & n11489 ) | ( ~n11483 & n11490 ) | ( n11489 & n11490 ) ;
  assign n11492 = n3162 & n3715 ;
  assign n11493 = x99 & n3719 ;
  assign n11494 = x100 | n11493 ;
  assign n11495 = ( n3721 & n11493 ) | ( n3721 & n11494 ) | ( n11493 & n11494 ) ;
  assign n11496 = x98 & n3922 ;
  assign n11497 = n11495 | n11496 ;
  assign n11498 = ( x41 & n11492 ) | ( x41 & ~n11497 ) | ( n11492 & ~n11497 ) ;
  assign n11499 = ( ~x41 & n11497 ) | ( ~x41 & n11498 ) | ( n11497 & n11498 ) ;
  assign n11500 = ( ~n11492 & n11498 ) | ( ~n11492 & n11499 ) | ( n11498 & n11499 ) ;
  assign n11501 = n2585 & n4227 ;
  assign n11502 = x96 & n4231 ;
  assign n11503 = x97 | n11502 ;
  assign n11504 = ( n4233 & n11502 ) | ( n4233 & n11503 ) | ( n11502 & n11503 ) ;
  assign n11505 = x95 & n4470 ;
  assign n11506 = n11504 | n11505 ;
  assign n11507 = ( x44 & n11501 ) | ( x44 & ~n11506 ) | ( n11501 & ~n11506 ) ;
  assign n11508 = ( ~x44 & n11506 ) | ( ~x44 & n11507 ) | ( n11506 & n11507 ) ;
  assign n11509 = ( ~n11501 & n11507 ) | ( ~n11501 & n11508 ) | ( n11507 & n11508 ) ;
  assign n11510 = n1481 & n6027 ;
  assign n11511 = x87 & n6031 ;
  assign n11512 = x88 | n11511 ;
  assign n11513 = ( n6033 & n11511 ) | ( n6033 & n11512 ) | ( n11511 & n11512 ) ;
  assign n11514 = x86 & n6303 ;
  assign n11515 = n11513 | n11514 ;
  assign n11516 = ( x53 & n11510 ) | ( x53 & ~n11515 ) | ( n11510 & ~n11515 ) ;
  assign n11517 = ( ~x53 & n11515 ) | ( ~x53 & n11516 ) | ( n11515 & n11516 ) ;
  assign n11518 = ( ~n11510 & n11516 ) | ( ~n11510 & n11517 ) | ( n11516 & n11517 ) ;
  assign n11519 = n990 & n7423 ;
  assign n11520 = x81 & n7427 ;
  assign n11521 = x82 | n11520 ;
  assign n11522 = ( n7429 & n11520 ) | ( n7429 & n11521 ) | ( n11520 & n11521 ) ;
  assign n11523 = x80 & n7708 ;
  assign n11524 = n11522 | n11523 ;
  assign n11525 = ( x59 & n11519 ) | ( x59 & ~n11524 ) | ( n11519 & ~n11524 ) ;
  assign n11526 = ( ~x59 & n11524 ) | ( ~x59 & n11525 ) | ( n11524 & n11525 ) ;
  assign n11527 = ( ~n11519 & n11525 ) | ( ~n11519 & n11526 ) | ( n11525 & n11526 ) ;
  assign n11528 = n701 & n8154 ;
  assign n11529 = x78 & n8158 ;
  assign n11530 = x79 | n11529 ;
  assign n11531 = ( n8160 & n11529 ) | ( n8160 & n11530 ) | ( n11529 & n11530 ) ;
  assign n11532 = x77 & n8439 ;
  assign n11533 = n11531 | n11532 ;
  assign n11534 = ( x62 & n11528 ) | ( x62 & ~n11533 ) | ( n11528 & ~n11533 ) ;
  assign n11535 = ( ~x62 & n11533 ) | ( ~x62 & n11534 ) | ( n11533 & n11534 ) ;
  assign n11536 = ( ~n11528 & n11534 ) | ( ~n11528 & n11535 ) | ( n11534 & n11535 ) ;
  assign n11537 = x75 & n8927 ;
  assign n11538 = ( ~x76 & n8693 ) | ( ~x76 & n8927 ) | ( n8693 & n8927 ) ;
  assign n11539 = ( n8693 & n11537 ) | ( n8693 & ~n11538 ) | ( n11537 & ~n11538 ) ;
  assign n11540 = ( ~x11 & n11126 ) | ( ~x11 & n11539 ) | ( n11126 & n11539 ) ;
  assign n11541 = ( n11126 & n11539 ) | ( n11126 & ~n11540 ) | ( n11539 & ~n11540 ) ;
  assign n11542 = ( x11 & n11540 ) | ( x11 & ~n11541 ) | ( n11540 & ~n11541 ) ;
  assign n11543 = ( n11331 & n11536 ) | ( n11331 & ~n11542 ) | ( n11536 & ~n11542 ) ;
  assign n11544 = ( ~n11331 & n11536 ) | ( ~n11331 & n11542 ) | ( n11536 & n11542 ) ;
  assign n11545 = ( ~n11536 & n11543 ) | ( ~n11536 & n11544 ) | ( n11543 & n11544 ) ;
  assign n11546 = ( n11352 & n11527 ) | ( n11352 & ~n11545 ) | ( n11527 & ~n11545 ) ;
  assign n11547 = ( ~n11352 & n11527 ) | ( ~n11352 & n11545 ) | ( n11527 & n11545 ) ;
  assign n11548 = ( ~n11527 & n11546 ) | ( ~n11527 & n11547 ) | ( n11546 & n11547 ) ;
  assign n11549 = n1262 & n6713 ;
  assign n11550 = x84 & n6717 ;
  assign n11551 = x85 | n11550 ;
  assign n11552 = ( n6719 & n11550 ) | ( n6719 & n11551 ) | ( n11550 & n11551 ) ;
  assign n11553 = x83 & n6980 ;
  assign n11554 = n11552 | n11553 ;
  assign n11555 = ( x56 & n11549 ) | ( x56 & ~n11554 ) | ( n11549 & ~n11554 ) ;
  assign n11556 = ( ~x56 & n11554 ) | ( ~x56 & n11555 ) | ( n11554 & n11555 ) ;
  assign n11557 = ( ~n11549 & n11555 ) | ( ~n11549 & n11556 ) | ( n11555 & n11556 ) ;
  assign n11558 = ( n11364 & n11548 ) | ( n11364 & ~n11557 ) | ( n11548 & ~n11557 ) ;
  assign n11559 = ( ~n11364 & n11548 ) | ( ~n11364 & n11557 ) | ( n11548 & n11557 ) ;
  assign n11560 = ( ~n11548 & n11558 ) | ( ~n11548 & n11559 ) | ( n11558 & n11559 ) ;
  assign n11561 = ( n11367 & n11518 ) | ( n11367 & n11560 ) | ( n11518 & n11560 ) ;
  assign n11562 = ( ~n11367 & n11518 ) | ( ~n11367 & n11560 ) | ( n11518 & n11560 ) ;
  assign n11563 = ( n11367 & ~n11561 ) | ( n11367 & n11562 ) | ( ~n11561 & n11562 ) ;
  assign n11564 = n1914 & n5374 ;
  assign n11565 = x90 & n5378 ;
  assign n11566 = x91 | n11565 ;
  assign n11567 = ( n5380 & n11565 ) | ( n5380 & n11566 ) | ( n11565 & n11566 ) ;
  assign n11568 = x89 & n5638 ;
  assign n11569 = n11567 | n11568 ;
  assign n11570 = ( x50 & n11564 ) | ( x50 & ~n11569 ) | ( n11564 & ~n11569 ) ;
  assign n11571 = ( ~x50 & n11569 ) | ( ~x50 & n11570 ) | ( n11569 & n11570 ) ;
  assign n11572 = ( ~n11564 & n11570 ) | ( ~n11564 & n11571 ) | ( n11570 & n11571 ) ;
  assign n11573 = ( n11370 & n11563 ) | ( n11370 & n11572 ) | ( n11563 & n11572 ) ;
  assign n11574 = ( ~n11370 & n11563 ) | ( ~n11370 & n11572 ) | ( n11563 & n11572 ) ;
  assign n11575 = ( n11370 & ~n11573 ) | ( n11370 & n11574 ) | ( ~n11573 & n11574 ) ;
  assign n11576 = n2294 & n4787 ;
  assign n11577 = x93 & n4791 ;
  assign n11578 = x94 | n11577 ;
  assign n11579 = ( n4793 & n11577 ) | ( n4793 & n11578 ) | ( n11577 & n11578 ) ;
  assign n11580 = x92 & n5030 ;
  assign n11581 = n11579 | n11580 ;
  assign n11582 = ( x47 & n11576 ) | ( x47 & ~n11581 ) | ( n11576 & ~n11581 ) ;
  assign n11583 = ( ~x47 & n11581 ) | ( ~x47 & n11582 ) | ( n11581 & n11582 ) ;
  assign n11584 = ( ~n11576 & n11582 ) | ( ~n11576 & n11583 ) | ( n11582 & n11583 ) ;
  assign n11585 = ( n11382 & n11575 ) | ( n11382 & n11584 ) | ( n11575 & n11584 ) ;
  assign n11586 = ( ~n11382 & n11575 ) | ( ~n11382 & n11584 ) | ( n11575 & n11584 ) ;
  assign n11587 = ( n11382 & ~n11585 ) | ( n11382 & n11586 ) | ( ~n11585 & n11586 ) ;
  assign n11588 = ( n11394 & n11509 ) | ( n11394 & n11587 ) | ( n11509 & n11587 ) ;
  assign n11589 = ( ~n11394 & n11509 ) | ( ~n11394 & n11587 ) | ( n11509 & n11587 ) ;
  assign n11590 = ( n11394 & ~n11588 ) | ( n11394 & n11589 ) | ( ~n11588 & n11589 ) ;
  assign n11591 = ( n11406 & n11500 ) | ( n11406 & n11590 ) | ( n11500 & n11590 ) ;
  assign n11592 = ( ~n11406 & n11500 ) | ( ~n11406 & n11590 ) | ( n11500 & n11590 ) ;
  assign n11593 = ( n11406 & ~n11591 ) | ( n11406 & n11592 ) | ( ~n11591 & n11592 ) ;
  assign n11594 = n3224 & n3650 ;
  assign n11595 = x102 & n3228 ;
  assign n11596 = x103 | n11595 ;
  assign n11597 = ( n3230 & n11595 ) | ( n3230 & n11596 ) | ( n11595 & n11596 ) ;
  assign n11598 = x101 & n3413 ;
  assign n11599 = n11597 | n11598 ;
  assign n11600 = ( x38 & n11594 ) | ( x38 & ~n11599 ) | ( n11594 & ~n11599 ) ;
  assign n11601 = ( ~x38 & n11599 ) | ( ~x38 & n11600 ) | ( n11599 & n11600 ) ;
  assign n11602 = ( ~n11594 & n11600 ) | ( ~n11594 & n11601 ) | ( n11600 & n11601 ) ;
  assign n11603 = ( n11418 & n11593 ) | ( n11418 & n11602 ) | ( n11593 & n11602 ) ;
  assign n11604 = ( ~n11418 & n11593 ) | ( ~n11418 & n11602 ) | ( n11593 & n11602 ) ;
  assign n11605 = ( n11418 & ~n11603 ) | ( n11418 & n11604 ) | ( ~n11603 & n11604 ) ;
  assign n11606 = ( n11421 & n11491 ) | ( n11421 & n11605 ) | ( n11491 & n11605 ) ;
  assign n11607 = ( ~n11421 & n11491 ) | ( ~n11421 & n11605 ) | ( n11491 & n11605 ) ;
  assign n11608 = ( n11421 & ~n11606 ) | ( n11421 & n11607 ) | ( ~n11606 & n11607 ) ;
  assign n11609 = n2320 & n4734 ;
  assign n11610 = x108 & n2324 ;
  assign n11611 = x109 | n11610 ;
  assign n11612 = ( n2326 & n11610 ) | ( n2326 & n11611 ) | ( n11610 & n11611 ) ;
  assign n11613 = x107 & n2497 ;
  assign n11614 = n11612 | n11613 ;
  assign n11615 = ( x32 & n11609 ) | ( x32 & ~n11614 ) | ( n11609 & ~n11614 ) ;
  assign n11616 = ( ~x32 & n11614 ) | ( ~x32 & n11615 ) | ( n11614 & n11615 ) ;
  assign n11617 = ( ~n11609 & n11615 ) | ( ~n11609 & n11616 ) | ( n11615 & n11616 ) ;
  assign n11618 = ( n11424 & n11608 ) | ( n11424 & n11617 ) | ( n11608 & n11617 ) ;
  assign n11619 = ( n11424 & ~n11608 ) | ( n11424 & n11617 ) | ( ~n11608 & n11617 ) ;
  assign n11620 = ( n11608 & ~n11618 ) | ( n11608 & n11619 ) | ( ~n11618 & n11619 ) ;
  assign n11621 = n1949 & n5145 ;
  assign n11622 = x111 & n1953 ;
  assign n11623 = x112 | n11622 ;
  assign n11624 = ( n1955 & n11622 ) | ( n1955 & n11623 ) | ( n11622 & n11623 ) ;
  assign n11625 = x110 & n2114 ;
  assign n11626 = n11624 | n11625 ;
  assign n11627 = ( x29 & n11621 ) | ( x29 & ~n11626 ) | ( n11621 & ~n11626 ) ;
  assign n11628 = ( ~x29 & n11626 ) | ( ~x29 & n11627 ) | ( n11626 & n11627 ) ;
  assign n11629 = ( ~n11621 & n11627 ) | ( ~n11621 & n11628 ) | ( n11627 & n11628 ) ;
  assign n11630 = ( n11427 & n11620 ) | ( n11427 & n11629 ) | ( n11620 & n11629 ) ;
  assign n11631 = ( n11427 & ~n11620 ) | ( n11427 & n11629 ) | ( ~n11620 & n11629 ) ;
  assign n11632 = ( n11620 & ~n11630 ) | ( n11620 & n11631 ) | ( ~n11630 & n11631 ) ;
  assign n11633 = ( n11430 & n11482 ) | ( n11430 & n11632 ) | ( n11482 & n11632 ) ;
  assign n11634 = ( n11430 & ~n11482 ) | ( n11430 & n11632 ) | ( ~n11482 & n11632 ) ;
  assign n11635 = ( n11482 & ~n11633 ) | ( n11482 & n11634 ) | ( ~n11633 & n11634 ) ;
  assign n11636 = n1297 & n6421 ;
  assign n11637 = x117 & n1301 ;
  assign n11638 = x118 | n11637 ;
  assign n11639 = ( n1303 & n11637 ) | ( n1303 & n11638 ) | ( n11637 & n11638 ) ;
  assign n11640 = x116 & n1426 ;
  assign n11641 = n11639 | n11640 ;
  assign n11642 = ( x23 & n11636 ) | ( x23 & ~n11641 ) | ( n11636 & ~n11641 ) ;
  assign n11643 = ( ~x23 & n11641 ) | ( ~x23 & n11642 ) | ( n11641 & n11642 ) ;
  assign n11644 = ( ~n11636 & n11642 ) | ( ~n11636 & n11643 ) | ( n11642 & n11643 ) ;
  assign n11645 = ( n11442 & n11635 ) | ( n11442 & n11644 ) | ( n11635 & n11644 ) ;
  assign n11646 = ( n11442 & ~n11635 ) | ( n11442 & n11644 ) | ( ~n11635 & n11644 ) ;
  assign n11647 = ( n11635 & ~n11645 ) | ( n11635 & n11646 ) | ( ~n11645 & n11646 ) ;
  assign n11648 = ( n11445 & n11473 ) | ( n11445 & n11647 ) | ( n11473 & n11647 ) ;
  assign n11649 = ( n11445 & ~n11473 ) | ( n11445 & n11647 ) | ( ~n11473 & n11647 ) ;
  assign n11650 = ( n11473 & ~n11648 ) | ( n11473 & n11649 ) | ( ~n11648 & n11649 ) ;
  assign n11651 = n810 & n7841 ;
  assign n11652 = x123 & n814 ;
  assign n11653 = x124 | n11652 ;
  assign n11654 = ( n816 & n11652 ) | ( n816 & n11653 ) | ( n11652 & n11653 ) ;
  assign n11655 = x122 & n885 ;
  assign n11656 = n11654 | n11655 ;
  assign n11657 = ( x17 & n11651 ) | ( x17 & ~n11656 ) | ( n11651 & ~n11656 ) ;
  assign n11658 = ( ~x17 & n11656 ) | ( ~x17 & n11657 ) | ( n11656 & n11657 ) ;
  assign n11659 = ( ~n11651 & n11657 ) | ( ~n11651 & n11658 ) | ( n11657 & n11658 ) ;
  assign n11660 = ( n11448 & n11650 ) | ( n11448 & n11659 ) | ( n11650 & n11659 ) ;
  assign n11661 = ( n11448 & ~n11650 ) | ( n11448 & n11659 ) | ( ~n11650 & n11659 ) ;
  assign n11662 = ( n11650 & ~n11660 ) | ( n11650 & n11661 ) | ( ~n11660 & n11661 ) ;
  assign n11663 = n583 & n8846 ;
  assign n11664 = x126 & n587 ;
  assign n11665 = x127 | n11664 ;
  assign n11666 = ( n589 & n11664 ) | ( n589 & n11665 ) | ( n11664 & n11665 ) ;
  assign n11667 = x125 & n676 ;
  assign n11668 = n11666 | n11667 ;
  assign n11669 = ( x14 & n11663 ) | ( x14 & ~n11668 ) | ( n11663 & ~n11668 ) ;
  assign n11670 = ( ~x14 & n11668 ) | ( ~x14 & n11669 ) | ( n11668 & n11669 ) ;
  assign n11671 = ( ~n11663 & n11669 ) | ( ~n11663 & n11670 ) | ( n11669 & n11670 ) ;
  assign n11672 = ( n11451 & n11662 ) | ( n11451 & n11671 ) | ( n11662 & n11671 ) ;
  assign n11673 = ( n11451 & ~n11662 ) | ( n11451 & n11671 ) | ( ~n11662 & n11671 ) ;
  assign n11674 = ( n11662 & ~n11672 ) | ( n11662 & n11673 ) | ( ~n11672 & n11673 ) ;
  assign n11675 = ( n11459 & n11462 ) | ( n11459 & n11674 ) | ( n11462 & n11674 ) ;
  assign n11676 = ( n11459 & ~n11462 ) | ( n11459 & n11674 ) | ( ~n11462 & n11674 ) ;
  assign n11677 = ( n11462 & ~n11675 ) | ( n11462 & n11676 ) | ( ~n11675 & n11676 ) ;
  assign n11678 = n583 & n8865 ;
  assign n11679 = x127 & n587 ;
  assign n11680 = x126 | n11679 ;
  assign n11681 = ( n676 & n11679 ) | ( n676 & n11680 ) | ( n11679 & n11680 ) ;
  assign n11682 = ( x14 & n11678 ) | ( x14 & ~n11681 ) | ( n11678 & ~n11681 ) ;
  assign n11683 = ( ~x14 & n11681 ) | ( ~x14 & n11682 ) | ( n11681 & n11682 ) ;
  assign n11684 = ( ~n11678 & n11682 ) | ( ~n11678 & n11683 ) | ( n11682 & n11683 ) ;
  assign n11685 = n810 & n8331 ;
  assign n11686 = x124 & n814 ;
  assign n11687 = x125 | n11686 ;
  assign n11688 = ( n816 & n11686 ) | ( n816 & n11687 ) | ( n11686 & n11687 ) ;
  assign n11689 = x123 & n885 ;
  assign n11690 = n11688 | n11689 ;
  assign n11691 = ( x17 & n11685 ) | ( x17 & ~n11690 ) | ( n11685 & ~n11690 ) ;
  assign n11692 = ( ~x17 & n11690 ) | ( ~x17 & n11691 ) | ( n11690 & n11691 ) ;
  assign n11693 = ( ~n11685 & n11691 ) | ( ~n11685 & n11692 ) | ( n11691 & n11692 ) ;
  assign n11694 = n1297 & n6645 ;
  assign n11695 = x118 & n1301 ;
  assign n11696 = x119 | n11695 ;
  assign n11697 = ( n1303 & n11695 ) | ( n1303 & n11696 ) | ( n11695 & n11696 ) ;
  assign n11698 = x117 & n1426 ;
  assign n11699 = n11697 | n11698 ;
  assign n11700 = ( x23 & n11694 ) | ( x23 & ~n11699 ) | ( n11694 & ~n11699 ) ;
  assign n11701 = ( ~x23 & n11699 ) | ( ~x23 & n11700 ) | ( n11699 & n11700 ) ;
  assign n11702 = ( ~n11694 & n11700 ) | ( ~n11694 & n11701 ) | ( n11700 & n11701 ) ;
  assign n11703 = n1617 & n5977 ;
  assign n11704 = x115 & n1621 ;
  assign n11705 = x116 | n11704 ;
  assign n11706 = ( n1623 & n11704 ) | ( n1623 & n11705 ) | ( n11704 & n11705 ) ;
  assign n11707 = x114 & n1749 ;
  assign n11708 = n11706 | n11707 ;
  assign n11709 = ( x26 & n11703 ) | ( x26 & ~n11708 ) | ( n11703 & ~n11708 ) ;
  assign n11710 = ( ~x26 & n11708 ) | ( ~x26 & n11709 ) | ( n11708 & n11709 ) ;
  assign n11711 = ( ~n11703 & n11709 ) | ( ~n11703 & n11710 ) | ( n11709 & n11710 ) ;
  assign n11712 = n1949 & n5542 ;
  assign n11713 = x112 & n1953 ;
  assign n11714 = x113 | n11713 ;
  assign n11715 = ( n1955 & n11713 ) | ( n1955 & n11714 ) | ( n11713 & n11714 ) ;
  assign n11716 = x111 & n2114 ;
  assign n11717 = n11715 | n11716 ;
  assign n11718 = ( x29 & n11712 ) | ( x29 & ~n11717 ) | ( n11712 & ~n11717 ) ;
  assign n11719 = ( ~x29 & n11717 ) | ( ~x29 & n11718 ) | ( n11717 & n11718 ) ;
  assign n11720 = ( ~n11712 & n11718 ) | ( ~n11712 & n11719 ) | ( n11718 & n11719 ) ;
  assign n11721 = n3224 & n3665 ;
  assign n11722 = x103 & n3228 ;
  assign n11723 = x104 | n11722 ;
  assign n11724 = ( n3230 & n11722 ) | ( n3230 & n11723 ) | ( n11722 & n11723 ) ;
  assign n11725 = x102 & n3413 ;
  assign n11726 = n11724 | n11725 ;
  assign n11727 = ( x38 & n11721 ) | ( x38 & ~n11726 ) | ( n11721 & ~n11726 ) ;
  assign n11728 = ( ~x38 & n11726 ) | ( ~x38 & n11727 ) | ( n11726 & n11727 ) ;
  assign n11729 = ( ~n11721 & n11727 ) | ( ~n11721 & n11728 ) | ( n11727 & n11728 ) ;
  assign n11730 = n3326 & n3715 ;
  assign n11731 = x100 & n3719 ;
  assign n11732 = x101 | n11731 ;
  assign n11733 = ( n3721 & n11731 ) | ( n3721 & n11732 ) | ( n11731 & n11732 ) ;
  assign n11734 = x99 & n3922 ;
  assign n11735 = n11733 | n11734 ;
  assign n11736 = ( x41 & n11730 ) | ( x41 & ~n11735 ) | ( n11730 & ~n11735 ) ;
  assign n11737 = ( ~x41 & n11735 ) | ( ~x41 & n11736 ) | ( n11735 & n11736 ) ;
  assign n11738 = ( ~n11730 & n11736 ) | ( ~n11730 & n11737 ) | ( n11736 & n11737 ) ;
  assign n11739 = n2725 & n4227 ;
  assign n11740 = x97 & n4231 ;
  assign n11741 = x98 | n11740 ;
  assign n11742 = ( n4233 & n11740 ) | ( n4233 & n11741 ) | ( n11740 & n11741 ) ;
  assign n11743 = x96 & n4470 ;
  assign n11744 = n11742 | n11743 ;
  assign n11745 = ( x44 & n11739 ) | ( x44 & ~n11744 ) | ( n11739 & ~n11744 ) ;
  assign n11746 = ( ~x44 & n11744 ) | ( ~x44 & n11745 ) | ( n11744 & n11745 ) ;
  assign n11747 = ( ~n11739 & n11745 ) | ( ~n11739 & n11746 ) | ( n11745 & n11746 ) ;
  assign n11748 = n2434 & n4787 ;
  assign n11749 = x94 & n4791 ;
  assign n11750 = x95 | n11749 ;
  assign n11751 = ( n4793 & n11749 ) | ( n4793 & n11750 ) | ( n11749 & n11750 ) ;
  assign n11752 = x93 & n5030 ;
  assign n11753 = n11751 | n11752 ;
  assign n11754 = ( x47 & n11748 ) | ( x47 & ~n11753 ) | ( n11748 & ~n11753 ) ;
  assign n11755 = ( ~x47 & n11753 ) | ( ~x47 & n11754 ) | ( n11753 & n11754 ) ;
  assign n11756 = ( ~n11748 & n11754 ) | ( ~n11748 & n11755 ) | ( n11754 & n11755 ) ;
  assign n11757 = n1082 & n7423 ;
  assign n11758 = x82 & n7427 ;
  assign n11759 = x83 | n11758 ;
  assign n11760 = ( n7429 & n11758 ) | ( n7429 & n11759 ) | ( n11758 & n11759 ) ;
  assign n11761 = x81 & n7708 ;
  assign n11762 = n11760 | n11761 ;
  assign n11763 = ( x59 & n11757 ) | ( x59 & ~n11762 ) | ( n11757 & ~n11762 ) ;
  assign n11764 = ( ~x59 & n11762 ) | ( ~x59 & n11763 ) | ( n11762 & n11763 ) ;
  assign n11765 = ( ~n11757 & n11763 ) | ( ~n11757 & n11764 ) | ( n11763 & n11764 ) ;
  assign n11766 = n769 & n8154 ;
  assign n11767 = x79 & n8158 ;
  assign n11768 = x80 | n11767 ;
  assign n11769 = ( n8160 & n11767 ) | ( n8160 & n11768 ) | ( n11767 & n11768 ) ;
  assign n11770 = x78 & n8439 ;
  assign n11771 = n11769 | n11770 ;
  assign n11772 = ( x62 & n11766 ) | ( x62 & ~n11771 ) | ( n11766 & ~n11771 ) ;
  assign n11773 = ( ~x62 & n11771 ) | ( ~x62 & n11772 ) | ( n11771 & n11772 ) ;
  assign n11774 = ( ~n11766 & n11772 ) | ( ~n11766 & n11773 ) | ( n11772 & n11773 ) ;
  assign n11775 = x76 & n8927 ;
  assign n11776 = ( ~x77 & n8693 ) | ( ~x77 & n8927 ) | ( n8693 & n8927 ) ;
  assign n11777 = ( n8693 & n11775 ) | ( n8693 & ~n11776 ) | ( n11775 & ~n11776 ) ;
  assign n11778 = ( n11540 & n11774 ) | ( n11540 & ~n11777 ) | ( n11774 & ~n11777 ) ;
  assign n11779 = ( ~n11540 & n11774 ) | ( ~n11540 & n11777 ) | ( n11774 & n11777 ) ;
  assign n11780 = ( ~n11774 & n11778 ) | ( ~n11774 & n11779 ) | ( n11778 & n11779 ) ;
  assign n11781 = ( n11543 & n11765 ) | ( n11543 & ~n11780 ) | ( n11765 & ~n11780 ) ;
  assign n11782 = ( ~n11543 & n11765 ) | ( ~n11543 & n11780 ) | ( n11765 & n11780 ) ;
  assign n11783 = ( ~n11765 & n11781 ) | ( ~n11765 & n11782 ) | ( n11781 & n11782 ) ;
  assign n11784 = n1366 & n6713 ;
  assign n11785 = x85 & n6717 ;
  assign n11786 = x86 | n11785 ;
  assign n11787 = ( n6719 & n11785 ) | ( n6719 & n11786 ) | ( n11785 & n11786 ) ;
  assign n11788 = x84 & n6980 ;
  assign n11789 = n11787 | n11788 ;
  assign n11790 = ( x56 & n11784 ) | ( x56 & ~n11789 ) | ( n11784 & ~n11789 ) ;
  assign n11791 = ( ~x56 & n11789 ) | ( ~x56 & n11790 ) | ( n11789 & n11790 ) ;
  assign n11792 = ( ~n11784 & n11790 ) | ( ~n11784 & n11791 ) | ( n11790 & n11791 ) ;
  assign n11793 = ( n11546 & ~n11783 ) | ( n11546 & n11792 ) | ( ~n11783 & n11792 ) ;
  assign n11794 = ( n11546 & n11783 ) | ( n11546 & n11792 ) | ( n11783 & n11792 ) ;
  assign n11795 = ( n11783 & n11793 ) | ( n11783 & ~n11794 ) | ( n11793 & ~n11794 ) ;
  assign n11796 = n1585 & n6027 ;
  assign n11797 = x88 & n6031 ;
  assign n11798 = x89 | n11797 ;
  assign n11799 = ( n6033 & n11797 ) | ( n6033 & n11798 ) | ( n11797 & n11798 ) ;
  assign n11800 = x87 & n6303 ;
  assign n11801 = n11799 | n11800 ;
  assign n11802 = ( x53 & n11796 ) | ( x53 & ~n11801 ) | ( n11796 & ~n11801 ) ;
  assign n11803 = ( ~x53 & n11801 ) | ( ~x53 & n11802 ) | ( n11801 & n11802 ) ;
  assign n11804 = ( ~n11796 & n11802 ) | ( ~n11796 & n11803 ) | ( n11802 & n11803 ) ;
  assign n11805 = ( n11558 & n11795 ) | ( n11558 & ~n11804 ) | ( n11795 & ~n11804 ) ;
  assign n11806 = ( ~n11558 & n11795 ) | ( ~n11558 & n11804 ) | ( n11795 & n11804 ) ;
  assign n11807 = ( ~n11795 & n11805 ) | ( ~n11795 & n11806 ) | ( n11805 & n11806 ) ;
  assign n11808 = n2042 & n5374 ;
  assign n11809 = x91 & n5378 ;
  assign n11810 = x92 | n11809 ;
  assign n11811 = ( n5380 & n11809 ) | ( n5380 & n11810 ) | ( n11809 & n11810 ) ;
  assign n11812 = x90 & n5638 ;
  assign n11813 = n11811 | n11812 ;
  assign n11814 = ( x50 & n11808 ) | ( x50 & ~n11813 ) | ( n11808 & ~n11813 ) ;
  assign n11815 = ( ~x50 & n11813 ) | ( ~x50 & n11814 ) | ( n11813 & n11814 ) ;
  assign n11816 = ( ~n11808 & n11814 ) | ( ~n11808 & n11815 ) | ( n11814 & n11815 ) ;
  assign n11817 = ( n11561 & n11807 ) | ( n11561 & n11816 ) | ( n11807 & n11816 ) ;
  assign n11818 = ( n11561 & ~n11807 ) | ( n11561 & n11816 ) | ( ~n11807 & n11816 ) ;
  assign n11819 = ( n11807 & ~n11817 ) | ( n11807 & n11818 ) | ( ~n11817 & n11818 ) ;
  assign n11820 = ( n11573 & n11756 ) | ( n11573 & n11819 ) | ( n11756 & n11819 ) ;
  assign n11821 = ( n11573 & ~n11756 ) | ( n11573 & n11819 ) | ( ~n11756 & n11819 ) ;
  assign n11822 = ( n11756 & ~n11820 ) | ( n11756 & n11821 ) | ( ~n11820 & n11821 ) ;
  assign n11823 = ( n11585 & n11747 ) | ( n11585 & n11822 ) | ( n11747 & n11822 ) ;
  assign n11824 = ( n11585 & ~n11747 ) | ( n11585 & n11822 ) | ( ~n11747 & n11822 ) ;
  assign n11825 = ( n11747 & ~n11823 ) | ( n11747 & n11824 ) | ( ~n11823 & n11824 ) ;
  assign n11826 = ( n11588 & n11738 ) | ( n11588 & n11825 ) | ( n11738 & n11825 ) ;
  assign n11827 = ( n11588 & ~n11738 ) | ( n11588 & n11825 ) | ( ~n11738 & n11825 ) ;
  assign n11828 = ( n11738 & ~n11826 ) | ( n11738 & n11827 ) | ( ~n11826 & n11827 ) ;
  assign n11829 = ( n11591 & n11729 ) | ( n11591 & n11828 ) | ( n11729 & n11828 ) ;
  assign n11830 = ( n11591 & ~n11729 ) | ( n11591 & n11828 ) | ( ~n11729 & n11828 ) ;
  assign n11831 = ( n11729 & ~n11829 ) | ( n11729 & n11830 ) | ( ~n11829 & n11830 ) ;
  assign n11832 = n2766 & n4362 ;
  assign n11833 = x106 & n2770 ;
  assign n11834 = x107 | n11833 ;
  assign n11835 = ( n2772 & n11833 ) | ( n2772 & n11834 ) | ( n11833 & n11834 ) ;
  assign n11836 = x105 & n2943 ;
  assign n11837 = n11835 | n11836 ;
  assign n11838 = ( x35 & n11832 ) | ( x35 & ~n11837 ) | ( n11832 & ~n11837 ) ;
  assign n11839 = ( ~x35 & n11837 ) | ( ~x35 & n11838 ) | ( n11837 & n11838 ) ;
  assign n11840 = ( ~n11832 & n11838 ) | ( ~n11832 & n11839 ) | ( n11838 & n11839 ) ;
  assign n11841 = ( n11603 & n11831 ) | ( n11603 & n11840 ) | ( n11831 & n11840 ) ;
  assign n11842 = ( ~n11603 & n11831 ) | ( ~n11603 & n11840 ) | ( n11831 & n11840 ) ;
  assign n11843 = ( n11603 & ~n11841 ) | ( n11603 & n11842 ) | ( ~n11841 & n11842 ) ;
  assign n11844 = n2320 & n4934 ;
  assign n11845 = x109 & n2324 ;
  assign n11846 = x110 | n11845 ;
  assign n11847 = ( n2326 & n11845 ) | ( n2326 & n11846 ) | ( n11845 & n11846 ) ;
  assign n11848 = x108 & n2497 ;
  assign n11849 = n11847 | n11848 ;
  assign n11850 = ( x32 & n11844 ) | ( x32 & ~n11849 ) | ( n11844 & ~n11849 ) ;
  assign n11851 = ( ~x32 & n11849 ) | ( ~x32 & n11850 ) | ( n11849 & n11850 ) ;
  assign n11852 = ( ~n11844 & n11850 ) | ( ~n11844 & n11851 ) | ( n11850 & n11851 ) ;
  assign n11853 = ( n11606 & n11843 ) | ( n11606 & n11852 ) | ( n11843 & n11852 ) ;
  assign n11854 = ( n11606 & ~n11843 ) | ( n11606 & n11852 ) | ( ~n11843 & n11852 ) ;
  assign n11855 = ( n11843 & ~n11853 ) | ( n11843 & n11854 ) | ( ~n11853 & n11854 ) ;
  assign n11856 = ( n11618 & n11720 ) | ( n11618 & n11855 ) | ( n11720 & n11855 ) ;
  assign n11857 = ( n11618 & ~n11720 ) | ( n11618 & n11855 ) | ( ~n11720 & n11855 ) ;
  assign n11858 = ( n11720 & ~n11856 ) | ( n11720 & n11857 ) | ( ~n11856 & n11857 ) ;
  assign n11859 = ( n11630 & n11711 ) | ( n11630 & n11858 ) | ( n11711 & n11858 ) ;
  assign n11860 = ( ~n11630 & n11711 ) | ( ~n11630 & n11858 ) | ( n11711 & n11858 ) ;
  assign n11861 = ( n11630 & ~n11859 ) | ( n11630 & n11860 ) | ( ~n11859 & n11860 ) ;
  assign n11862 = ( n11633 & n11702 ) | ( n11633 & n11861 ) | ( n11702 & n11861 ) ;
  assign n11863 = ( n11633 & ~n11702 ) | ( n11633 & n11861 ) | ( ~n11702 & n11861 ) ;
  assign n11864 = ( n11702 & ~n11862 ) | ( n11702 & n11863 ) | ( ~n11862 & n11863 ) ;
  assign n11865 = n1016 & n7582 ;
  assign n11866 = x121 & n1020 ;
  assign n11867 = x122 | n11866 ;
  assign n11868 = ( n1022 & n11866 ) | ( n1022 & n11867 ) | ( n11866 & n11867 ) ;
  assign n11869 = x120 & n1145 ;
  assign n11870 = n11868 | n11869 ;
  assign n11871 = ( x20 & n11865 ) | ( x20 & ~n11870 ) | ( n11865 & ~n11870 ) ;
  assign n11872 = ( ~x20 & n11870 ) | ( ~x20 & n11871 ) | ( n11870 & n11871 ) ;
  assign n11873 = ( ~n11865 & n11871 ) | ( ~n11865 & n11872 ) | ( n11871 & n11872 ) ;
  assign n11874 = ( n11645 & n11864 ) | ( n11645 & n11873 ) | ( n11864 & n11873 ) ;
  assign n11875 = ( n11645 & ~n11864 ) | ( n11645 & n11873 ) | ( ~n11864 & n11873 ) ;
  assign n11876 = ( n11864 & ~n11874 ) | ( n11864 & n11875 ) | ( ~n11874 & n11875 ) ;
  assign n11877 = ( n11648 & n11693 ) | ( n11648 & n11876 ) | ( n11693 & n11876 ) ;
  assign n11878 = ( n11648 & ~n11693 ) | ( n11648 & n11876 ) | ( ~n11693 & n11876 ) ;
  assign n11879 = ( n11693 & ~n11877 ) | ( n11693 & n11878 ) | ( ~n11877 & n11878 ) ;
  assign n11880 = ( n11660 & n11684 ) | ( n11660 & n11879 ) | ( n11684 & n11879 ) ;
  assign n11881 = ( ~n11660 & n11684 ) | ( ~n11660 & n11879 ) | ( n11684 & n11879 ) ;
  assign n11882 = ( n11660 & ~n11880 ) | ( n11660 & n11881 ) | ( ~n11880 & n11881 ) ;
  assign n11883 = ( n11672 & n11675 ) | ( n11672 & n11882 ) | ( n11675 & n11882 ) ;
  assign n11884 = ( n11672 & ~n11675 ) | ( n11672 & n11882 ) | ( ~n11675 & n11882 ) ;
  assign n11885 = ( n11675 & ~n11883 ) | ( n11675 & n11884 ) | ( ~n11883 & n11884 ) ;
  assign n11886 = n1016 & n7597 ;
  assign n11887 = x122 & n1020 ;
  assign n11888 = x123 | n11887 ;
  assign n11889 = ( n1022 & n11887 ) | ( n1022 & n11888 ) | ( n11887 & n11888 ) ;
  assign n11890 = x121 & n1145 ;
  assign n11891 = n11889 | n11890 ;
  assign n11892 = ( x20 & n11886 ) | ( x20 & ~n11891 ) | ( n11886 & ~n11891 ) ;
  assign n11893 = ( ~x20 & n11891 ) | ( ~x20 & n11892 ) | ( n11891 & n11892 ) ;
  assign n11894 = ( ~n11886 & n11892 ) | ( ~n11886 & n11893 ) | ( n11892 & n11893 ) ;
  assign n11895 = n1297 & n7098 ;
  assign n11896 = x119 & n1301 ;
  assign n11897 = x120 | n11896 ;
  assign n11898 = ( n1303 & n11896 ) | ( n1303 & n11897 ) | ( n11896 & n11897 ) ;
  assign n11899 = x118 & n1426 ;
  assign n11900 = n11898 | n11899 ;
  assign n11901 = ( x23 & n11895 ) | ( x23 & ~n11900 ) | ( n11895 & ~n11900 ) ;
  assign n11902 = ( ~x23 & n11900 ) | ( ~x23 & n11901 ) | ( n11900 & n11901 ) ;
  assign n11903 = ( ~n11895 & n11901 ) | ( ~n11895 & n11902 ) | ( n11901 & n11902 ) ;
  assign n11904 = n1617 & n6201 ;
  assign n11905 = x116 & n1621 ;
  assign n11906 = x117 | n11905 ;
  assign n11907 = ( n1623 & n11905 ) | ( n1623 & n11906 ) | ( n11905 & n11906 ) ;
  assign n11908 = x115 & n1749 ;
  assign n11909 = n11907 | n11908 ;
  assign n11910 = ( x26 & n11904 ) | ( x26 & ~n11909 ) | ( n11904 & ~n11909 ) ;
  assign n11911 = ( ~x26 & n11909 ) | ( ~x26 & n11910 ) | ( n11909 & n11910 ) ;
  assign n11912 = ( ~n11904 & n11910 ) | ( ~n11904 & n11911 ) | ( n11910 & n11911 ) ;
  assign n11913 = n1949 & n5750 ;
  assign n11914 = x113 & n1953 ;
  assign n11915 = x114 | n11914 ;
  assign n11916 = ( n1955 & n11914 ) | ( n1955 & n11915 ) | ( n11914 & n11915 ) ;
  assign n11917 = x112 & n2114 ;
  assign n11918 = n11916 | n11917 ;
  assign n11919 = ( x29 & n11913 ) | ( x29 & ~n11918 ) | ( n11913 & ~n11918 ) ;
  assign n11920 = ( ~x29 & n11918 ) | ( ~x29 & n11919 ) | ( n11918 & n11919 ) ;
  assign n11921 = ( ~n11913 & n11919 ) | ( ~n11913 & n11920 ) | ( n11919 & n11920 ) ;
  assign n11922 = n2320 & n5130 ;
  assign n11923 = x110 & n2324 ;
  assign n11924 = x111 | n11923 ;
  assign n11925 = ( n2326 & n11923 ) | ( n2326 & n11924 ) | ( n11923 & n11924 ) ;
  assign n11926 = x109 & n2497 ;
  assign n11927 = n11925 | n11926 ;
  assign n11928 = ( x32 & n11922 ) | ( x32 & ~n11927 ) | ( n11922 & ~n11927 ) ;
  assign n11929 = ( ~x32 & n11927 ) | ( ~x32 & n11928 ) | ( n11927 & n11928 ) ;
  assign n11930 = ( ~n11922 & n11928 ) | ( ~n11922 & n11929 ) | ( n11928 & n11929 ) ;
  assign n11931 = n2766 & n4377 ;
  assign n11932 = x107 & n2770 ;
  assign n11933 = x108 | n11932 ;
  assign n11934 = ( n2772 & n11932 ) | ( n2772 & n11933 ) | ( n11932 & n11933 ) ;
  assign n11935 = x106 & n2943 ;
  assign n11936 = n11934 | n11935 ;
  assign n11937 = ( x35 & n11931 ) | ( x35 & ~n11936 ) | ( n11931 & ~n11936 ) ;
  assign n11938 = ( ~x35 & n11936 ) | ( ~x35 & n11937 ) | ( n11936 & n11937 ) ;
  assign n11939 = ( ~n11931 & n11937 ) | ( ~n11931 & n11938 ) | ( n11937 & n11938 ) ;
  assign n11940 = n3224 & n3998 ;
  assign n11941 = x104 & n3228 ;
  assign n11942 = x105 | n11941 ;
  assign n11943 = ( n3230 & n11941 ) | ( n3230 & n11942 ) | ( n11941 & n11942 ) ;
  assign n11944 = x103 & n3413 ;
  assign n11945 = n11943 | n11944 ;
  assign n11946 = ( x38 & n11940 ) | ( x38 & ~n11945 ) | ( n11940 & ~n11945 ) ;
  assign n11947 = ( ~x38 & n11945 ) | ( ~x38 & n11946 ) | ( n11945 & n11946 ) ;
  assign n11948 = ( ~n11940 & n11946 ) | ( ~n11940 & n11947 ) | ( n11946 & n11947 ) ;
  assign n11949 = n2449 & n4787 ;
  assign n11950 = x95 & n4791 ;
  assign n11951 = x96 | n11950 ;
  assign n11952 = ( n4793 & n11950 ) | ( n4793 & n11951 ) | ( n11950 & n11951 ) ;
  assign n11953 = x94 & n5030 ;
  assign n11954 = n11952 | n11953 ;
  assign n11955 = ( x47 & n11949 ) | ( x47 & ~n11954 ) | ( n11949 & ~n11954 ) ;
  assign n11956 = ( ~x47 & n11954 ) | ( ~x47 & n11955 ) | ( n11954 & n11955 ) ;
  assign n11957 = ( ~n11949 & n11955 ) | ( ~n11949 & n11956 ) | ( n11955 & n11956 ) ;
  assign n11958 = n1701 & n6027 ;
  assign n11959 = x89 & n6031 ;
  assign n11960 = x90 | n11959 ;
  assign n11961 = ( n6033 & n11959 ) | ( n6033 & n11960 ) | ( n11959 & n11960 ) ;
  assign n11962 = x88 & n6303 ;
  assign n11963 = n11961 | n11962 ;
  assign n11964 = ( x53 & n11958 ) | ( x53 & ~n11963 ) | ( n11958 & ~n11963 ) ;
  assign n11965 = ( ~x53 & n11963 ) | ( ~x53 & n11964 ) | ( n11963 & n11964 ) ;
  assign n11966 = ( ~n11958 & n11964 ) | ( ~n11958 & n11965 ) | ( n11964 & n11965 ) ;
  assign n11967 = n1097 & n7423 ;
  assign n11968 = x83 & n7427 ;
  assign n11969 = x84 | n11968 ;
  assign n11970 = ( n7429 & n11968 ) | ( n7429 & n11969 ) | ( n11968 & n11969 ) ;
  assign n11971 = x82 & n7708 ;
  assign n11972 = n11970 | n11971 ;
  assign n11973 = ( x59 & n11967 ) | ( x59 & ~n11972 ) | ( n11967 & ~n11972 ) ;
  assign n11974 = ( ~x59 & n11972 ) | ( ~x59 & n11973 ) | ( n11972 & n11973 ) ;
  assign n11975 = ( ~n11967 & n11973 ) | ( ~n11967 & n11974 ) | ( n11973 & n11974 ) ;
  assign n11976 = x77 & n8927 ;
  assign n11977 = ( ~x78 & n8693 ) | ( ~x78 & n8927 ) | ( n8693 & n8927 ) ;
  assign n11978 = ( n8693 & n11976 ) | ( n8693 & ~n11977 ) | ( n11976 & ~n11977 ) ;
  assign n11979 = n910 & n8154 ;
  assign n11980 = x80 & n8158 ;
  assign n11981 = x81 | n11980 ;
  assign n11982 = ( n8160 & n11980 ) | ( n8160 & n11981 ) | ( n11980 & n11981 ) ;
  assign n11983 = x79 & n8439 ;
  assign n11984 = n11982 | n11983 ;
  assign n11985 = ( x62 & n11979 ) | ( x62 & ~n11984 ) | ( n11979 & ~n11984 ) ;
  assign n11986 = ( ~x62 & n11984 ) | ( ~x62 & n11985 ) | ( n11984 & n11985 ) ;
  assign n11987 = ( ~n11979 & n11985 ) | ( ~n11979 & n11986 ) | ( n11985 & n11986 ) ;
  assign n11988 = ( ~n11777 & n11978 ) | ( ~n11777 & n11987 ) | ( n11978 & n11987 ) ;
  assign n11989 = ( n11978 & n11987 ) | ( n11978 & ~n11988 ) | ( n11987 & ~n11988 ) ;
  assign n11990 = ( n11777 & n11988 ) | ( n11777 & ~n11989 ) | ( n11988 & ~n11989 ) ;
  assign n11991 = ( n11778 & n11975 ) | ( n11778 & ~n11990 ) | ( n11975 & ~n11990 ) ;
  assign n11992 = ( ~n11778 & n11975 ) | ( ~n11778 & n11990 ) | ( n11975 & n11990 ) ;
  assign n11993 = ( ~n11975 & n11991 ) | ( ~n11975 & n11992 ) | ( n11991 & n11992 ) ;
  assign n11994 = n1466 & n6713 ;
  assign n11995 = x86 & n6717 ;
  assign n11996 = x87 | n11995 ;
  assign n11997 = ( n6719 & n11995 ) | ( n6719 & n11996 ) | ( n11995 & n11996 ) ;
  assign n11998 = x85 & n6980 ;
  assign n11999 = n11997 | n11998 ;
  assign n12000 = ( x56 & n11994 ) | ( x56 & ~n11999 ) | ( n11994 & ~n11999 ) ;
  assign n12001 = ( ~x56 & n11999 ) | ( ~x56 & n12000 ) | ( n11999 & n12000 ) ;
  assign n12002 = ( ~n11994 & n12000 ) | ( ~n11994 & n12001 ) | ( n12000 & n12001 ) ;
  assign n12003 = ( n11781 & ~n11993 ) | ( n11781 & n12002 ) | ( ~n11993 & n12002 ) ;
  assign n12004 = ( n11781 & n11993 ) | ( n11781 & n12002 ) | ( n11993 & n12002 ) ;
  assign n12005 = ( n11993 & n12003 ) | ( n11993 & ~n12004 ) | ( n12003 & ~n12004 ) ;
  assign n12006 = ( n11793 & n11966 ) | ( n11793 & ~n12005 ) | ( n11966 & ~n12005 ) ;
  assign n12007 = ( ~n11793 & n11966 ) | ( ~n11793 & n12005 ) | ( n11966 & n12005 ) ;
  assign n12008 = ( ~n11966 & n12006 ) | ( ~n11966 & n12007 ) | ( n12006 & n12007 ) ;
  assign n12009 = n2057 & n5374 ;
  assign n12010 = x92 & n5378 ;
  assign n12011 = x93 | n12010 ;
  assign n12012 = ( n5380 & n12010 ) | ( n5380 & n12011 ) | ( n12010 & n12011 ) ;
  assign n12013 = x91 & n5638 ;
  assign n12014 = n12012 | n12013 ;
  assign n12015 = ( x50 & n12009 ) | ( x50 & ~n12014 ) | ( n12009 & ~n12014 ) ;
  assign n12016 = ( ~x50 & n12014 ) | ( ~x50 & n12015 ) | ( n12014 & n12015 ) ;
  assign n12017 = ( ~n12009 & n12015 ) | ( ~n12009 & n12016 ) | ( n12015 & n12016 ) ;
  assign n12018 = ( n11805 & n12008 ) | ( n11805 & ~n12017 ) | ( n12008 & ~n12017 ) ;
  assign n12019 = ( ~n11805 & n12008 ) | ( ~n11805 & n12017 ) | ( n12008 & n12017 ) ;
  assign n12020 = ( ~n12008 & n12018 ) | ( ~n12008 & n12019 ) | ( n12018 & n12019 ) ;
  assign n12021 = ( n11817 & n11957 ) | ( n11817 & n12020 ) | ( n11957 & n12020 ) ;
  assign n12022 = ( n11817 & ~n11957 ) | ( n11817 & n12020 ) | ( ~n11957 & n12020 ) ;
  assign n12023 = ( n11957 & ~n12021 ) | ( n11957 & n12022 ) | ( ~n12021 & n12022 ) ;
  assign n12024 = n2877 & n4227 ;
  assign n12025 = x98 & n4231 ;
  assign n12026 = x99 | n12025 ;
  assign n12027 = ( n4233 & n12025 ) | ( n4233 & n12026 ) | ( n12025 & n12026 ) ;
  assign n12028 = x97 & n4470 ;
  assign n12029 = n12027 | n12028 ;
  assign n12030 = ( x44 & n12024 ) | ( x44 & ~n12029 ) | ( n12024 & ~n12029 ) ;
  assign n12031 = ( ~x44 & n12029 ) | ( ~x44 & n12030 ) | ( n12029 & n12030 ) ;
  assign n12032 = ( ~n12024 & n12030 ) | ( ~n12024 & n12031 ) | ( n12030 & n12031 ) ;
  assign n12033 = ( n11820 & n12023 ) | ( n11820 & n12032 ) | ( n12023 & n12032 ) ;
  assign n12034 = ( ~n11820 & n12023 ) | ( ~n11820 & n12032 ) | ( n12023 & n12032 ) ;
  assign n12035 = ( n11820 & ~n12033 ) | ( n11820 & n12034 ) | ( ~n12033 & n12034 ) ;
  assign n12036 = n3486 & n3715 ;
  assign n12037 = x101 & n3719 ;
  assign n12038 = x102 | n12037 ;
  assign n12039 = ( n3721 & n12037 ) | ( n3721 & n12038 ) | ( n12037 & n12038 ) ;
  assign n12040 = x100 & n3922 ;
  assign n12041 = n12039 | n12040 ;
  assign n12042 = ( x41 & n12036 ) | ( x41 & ~n12041 ) | ( n12036 & ~n12041 ) ;
  assign n12043 = ( ~x41 & n12041 ) | ( ~x41 & n12042 ) | ( n12041 & n12042 ) ;
  assign n12044 = ( ~n12036 & n12042 ) | ( ~n12036 & n12043 ) | ( n12042 & n12043 ) ;
  assign n12045 = ( n11823 & n12035 ) | ( n11823 & n12044 ) | ( n12035 & n12044 ) ;
  assign n12046 = ( ~n11823 & n12035 ) | ( ~n11823 & n12044 ) | ( n12035 & n12044 ) ;
  assign n12047 = ( n11823 & ~n12045 ) | ( n11823 & n12046 ) | ( ~n12045 & n12046 ) ;
  assign n12048 = ( n11826 & n11948 ) | ( n11826 & n12047 ) | ( n11948 & n12047 ) ;
  assign n12049 = ( n11826 & ~n11948 ) | ( n11826 & n12047 ) | ( ~n11948 & n12047 ) ;
  assign n12050 = ( n11948 & ~n12048 ) | ( n11948 & n12049 ) | ( ~n12048 & n12049 ) ;
  assign n12051 = ( n11829 & n11939 ) | ( n11829 & n12050 ) | ( n11939 & n12050 ) ;
  assign n12052 = ( n11829 & ~n11939 ) | ( n11829 & n12050 ) | ( ~n11939 & n12050 ) ;
  assign n12053 = ( n11939 & ~n12051 ) | ( n11939 & n12052 ) | ( ~n12051 & n12052 ) ;
  assign n12054 = ( n11841 & n11930 ) | ( n11841 & n12053 ) | ( n11930 & n12053 ) ;
  assign n12055 = ( ~n11841 & n11930 ) | ( ~n11841 & n12053 ) | ( n11930 & n12053 ) ;
  assign n12056 = ( n11841 & ~n12054 ) | ( n11841 & n12055 ) | ( ~n12054 & n12055 ) ;
  assign n12057 = ( n11853 & n11921 ) | ( n11853 & n12056 ) | ( n11921 & n12056 ) ;
  assign n12058 = ( ~n11853 & n11921 ) | ( ~n11853 & n12056 ) | ( n11921 & n12056 ) ;
  assign n12059 = ( n11853 & ~n12057 ) | ( n11853 & n12058 ) | ( ~n12057 & n12058 ) ;
  assign n12060 = ( n11856 & n11912 ) | ( n11856 & n12059 ) | ( n11912 & n12059 ) ;
  assign n12061 = ( n11856 & ~n11912 ) | ( n11856 & n12059 ) | ( ~n11912 & n12059 ) ;
  assign n12062 = ( n11912 & ~n12060 ) | ( n11912 & n12061 ) | ( ~n12060 & n12061 ) ;
  assign n12063 = ( n11859 & n11903 ) | ( n11859 & n12062 ) | ( n11903 & n12062 ) ;
  assign n12064 = ( n11859 & ~n11903 ) | ( n11859 & n12062 ) | ( ~n11903 & n12062 ) ;
  assign n12065 = ( n11903 & ~n12063 ) | ( n11903 & n12064 ) | ( ~n12063 & n12064 ) ;
  assign n12066 = ( n11862 & n11894 ) | ( n11862 & n12065 ) | ( n11894 & n12065 ) ;
  assign n12067 = ( n11862 & ~n11894 ) | ( n11862 & n12065 ) | ( ~n11894 & n12065 ) ;
  assign n12068 = ( n11894 & ~n12066 ) | ( n11894 & n12067 ) | ( ~n12066 & n12067 ) ;
  assign n12069 = n810 & n8587 ;
  assign n12070 = x125 & n814 ;
  assign n12071 = x126 | n12070 ;
  assign n12072 = ( n816 & n12070 ) | ( n816 & n12071 ) | ( n12070 & n12071 ) ;
  assign n12073 = x124 & n885 ;
  assign n12074 = n12072 | n12073 ;
  assign n12075 = ( x17 & n12069 ) | ( x17 & ~n12074 ) | ( n12069 & ~n12074 ) ;
  assign n12076 = ( ~x17 & n12074 ) | ( ~x17 & n12075 ) | ( n12074 & n12075 ) ;
  assign n12077 = ( ~n12069 & n12075 ) | ( ~n12069 & n12076 ) | ( n12075 & n12076 ) ;
  assign n12078 = ( n11874 & n12068 ) | ( n11874 & n12077 ) | ( n12068 & n12077 ) ;
  assign n12079 = ( n11874 & ~n12068 ) | ( n11874 & n12077 ) | ( ~n12068 & n12077 ) ;
  assign n12080 = ( n12068 & ~n12078 ) | ( n12068 & n12079 ) | ( ~n12078 & n12079 ) ;
  assign n12081 = n583 & n8862 ;
  assign n12082 = ( x127 & n676 ) | ( x127 & n12081 ) | ( n676 & n12081 ) ;
  assign n12083 = x14 | n12082 ;
  assign n12084 = ~x14 & n12082 ;
  assign n12085 = ( ~n12082 & n12083 ) | ( ~n12082 & n12084 ) | ( n12083 & n12084 ) ;
  assign n12086 = ( n11877 & n12080 ) | ( n11877 & n12085 ) | ( n12080 & n12085 ) ;
  assign n12087 = ( n11877 & ~n12080 ) | ( n11877 & n12085 ) | ( ~n12080 & n12085 ) ;
  assign n12088 = ( n12080 & ~n12086 ) | ( n12080 & n12087 ) | ( ~n12086 & n12087 ) ;
  assign n12089 = ( n11880 & n11883 ) | ( n11880 & n12088 ) | ( n11883 & n12088 ) ;
  assign n12090 = ( n11880 & ~n11883 ) | ( n11880 & n12088 ) | ( ~n11883 & n12088 ) ;
  assign n12091 = ( n11883 & ~n12089 ) | ( n11883 & n12090 ) | ( ~n12089 & n12090 ) ;
  assign n12092 = n1016 & n7841 ;
  assign n12093 = x123 & n1020 ;
  assign n12094 = x124 | n12093 ;
  assign n12095 = ( n1022 & n12093 ) | ( n1022 & n12094 ) | ( n12093 & n12094 ) ;
  assign n12096 = x122 & n1145 ;
  assign n12097 = n12095 | n12096 ;
  assign n12098 = ( x20 & n12092 ) | ( x20 & ~n12097 ) | ( n12092 & ~n12097 ) ;
  assign n12099 = ( ~x20 & n12097 ) | ( ~x20 & n12098 ) | ( n12097 & n12098 ) ;
  assign n12100 = ( ~n12092 & n12098 ) | ( ~n12092 & n12099 ) | ( n12098 & n12099 ) ;
  assign n12101 = n1617 & n6421 ;
  assign n12102 = x117 & n1621 ;
  assign n12103 = x118 | n12102 ;
  assign n12104 = ( n1623 & n12102 ) | ( n1623 & n12103 ) | ( n12102 & n12103 ) ;
  assign n12105 = x116 & n1749 ;
  assign n12106 = n12104 | n12105 ;
  assign n12107 = ( x26 & n12101 ) | ( x26 & ~n12106 ) | ( n12101 & ~n12106 ) ;
  assign n12108 = ( ~x26 & n12106 ) | ( ~x26 & n12107 ) | ( n12106 & n12107 ) ;
  assign n12109 = ( ~n12101 & n12107 ) | ( ~n12101 & n12108 ) | ( n12107 & n12108 ) ;
  assign n12110 = n1949 & n5765 ;
  assign n12111 = x114 & n1953 ;
  assign n12112 = x115 | n12111 ;
  assign n12113 = ( n1955 & n12111 ) | ( n1955 & n12112 ) | ( n12111 & n12112 ) ;
  assign n12114 = x113 & n2114 ;
  assign n12115 = n12113 | n12114 ;
  assign n12116 = ( x29 & n12110 ) | ( x29 & ~n12115 ) | ( n12110 & ~n12115 ) ;
  assign n12117 = ( ~x29 & n12115 ) | ( ~x29 & n12116 ) | ( n12115 & n12116 ) ;
  assign n12118 = ( ~n12110 & n12116 ) | ( ~n12110 & n12117 ) | ( n12116 & n12117 ) ;
  assign n12119 = n3224 & n4013 ;
  assign n12120 = x105 & n3228 ;
  assign n12121 = x106 | n12120 ;
  assign n12122 = ( n3230 & n12120 ) | ( n3230 & n12121 ) | ( n12120 & n12121 ) ;
  assign n12123 = x104 & n3413 ;
  assign n12124 = n12122 | n12123 ;
  assign n12125 = ( x38 & n12119 ) | ( x38 & ~n12124 ) | ( n12119 & ~n12124 ) ;
  assign n12126 = ( ~x38 & n12124 ) | ( ~x38 & n12125 ) | ( n12124 & n12125 ) ;
  assign n12127 = ( ~n12119 & n12125 ) | ( ~n12119 & n12126 ) | ( n12125 & n12126 ) ;
  assign n12128 = n1914 & n6027 ;
  assign n12129 = x90 & n6031 ;
  assign n12130 = x91 | n12129 ;
  assign n12131 = ( n6033 & n12129 ) | ( n6033 & n12130 ) | ( n12129 & n12130 ) ;
  assign n12132 = x89 & n6303 ;
  assign n12133 = n12131 | n12132 ;
  assign n12134 = ( x53 & n12128 ) | ( x53 & ~n12133 ) | ( n12128 & ~n12133 ) ;
  assign n12135 = ( ~x53 & n12133 ) | ( ~x53 & n12134 ) | ( n12133 & n12134 ) ;
  assign n12136 = ( ~n12128 & n12134 ) | ( ~n12128 & n12135 ) | ( n12134 & n12135 ) ;
  assign n12137 = n1481 & n6713 ;
  assign n12138 = x87 & n6717 ;
  assign n12139 = x88 | n12138 ;
  assign n12140 = ( n6719 & n12138 ) | ( n6719 & n12139 ) | ( n12138 & n12139 ) ;
  assign n12141 = x86 & n6980 ;
  assign n12142 = n12140 | n12141 ;
  assign n12143 = ( x56 & n12137 ) | ( x56 & ~n12142 ) | ( n12137 & ~n12142 ) ;
  assign n12144 = ( ~x56 & n12142 ) | ( ~x56 & n12143 ) | ( n12142 & n12143 ) ;
  assign n12145 = ( ~n12137 & n12143 ) | ( ~n12137 & n12144 ) | ( n12143 & n12144 ) ;
  assign n12146 = n1262 & n7423 ;
  assign n12147 = x84 & n7427 ;
  assign n12148 = x85 | n12147 ;
  assign n12149 = ( n7429 & n12147 ) | ( n7429 & n12148 ) | ( n12147 & n12148 ) ;
  assign n12150 = x83 & n7708 ;
  assign n12151 = n12149 | n12150 ;
  assign n12152 = ( x59 & n12146 ) | ( x59 & ~n12151 ) | ( n12146 & ~n12151 ) ;
  assign n12153 = ( ~x59 & n12151 ) | ( ~x59 & n12152 ) | ( n12151 & n12152 ) ;
  assign n12154 = ( ~n12146 & n12152 ) | ( ~n12146 & n12153 ) | ( n12152 & n12153 ) ;
  assign n12155 = n990 & n8154 ;
  assign n12156 = x81 & n8158 ;
  assign n12157 = x82 | n12156 ;
  assign n12158 = ( n8160 & n12156 ) | ( n8160 & n12157 ) | ( n12156 & n12157 ) ;
  assign n12159 = x80 & n8439 ;
  assign n12160 = n12158 | n12159 ;
  assign n12161 = ( x62 & n12155 ) | ( x62 & ~n12160 ) | ( n12155 & ~n12160 ) ;
  assign n12162 = ( ~x62 & n12160 ) | ( ~x62 & n12161 ) | ( n12160 & n12161 ) ;
  assign n12163 = ( ~n12155 & n12161 ) | ( ~n12155 & n12162 ) | ( n12161 & n12162 ) ;
  assign n12164 = x78 & n8927 ;
  assign n12165 = ( ~x79 & n8693 ) | ( ~x79 & n8927 ) | ( n8693 & n8927 ) ;
  assign n12166 = ( n8693 & n12164 ) | ( n8693 & ~n12165 ) | ( n12164 & ~n12165 ) ;
  assign n12167 = ( ~x14 & n11777 ) | ( ~x14 & n12166 ) | ( n11777 & n12166 ) ;
  assign n12168 = ( n11777 & n12166 ) | ( n11777 & ~n12167 ) | ( n12166 & ~n12167 ) ;
  assign n12169 = ( x14 & n12167 ) | ( x14 & ~n12168 ) | ( n12167 & ~n12168 ) ;
  assign n12170 = ( n11988 & n12163 ) | ( n11988 & ~n12169 ) | ( n12163 & ~n12169 ) ;
  assign n12171 = ( ~n11988 & n12163 ) | ( ~n11988 & n12169 ) | ( n12163 & n12169 ) ;
  assign n12172 = ( ~n12163 & n12170 ) | ( ~n12163 & n12171 ) | ( n12170 & n12171 ) ;
  assign n12173 = ( n11991 & n12154 ) | ( n11991 & ~n12172 ) | ( n12154 & ~n12172 ) ;
  assign n12174 = ( ~n11991 & n12154 ) | ( ~n11991 & n12172 ) | ( n12154 & n12172 ) ;
  assign n12175 = ( ~n12154 & n12173 ) | ( ~n12154 & n12174 ) | ( n12173 & n12174 ) ;
  assign n12176 = ( n12003 & n12145 ) | ( n12003 & ~n12175 ) | ( n12145 & ~n12175 ) ;
  assign n12177 = ( ~n12003 & n12145 ) | ( ~n12003 & n12175 ) | ( n12145 & n12175 ) ;
  assign n12178 = ( ~n12145 & n12176 ) | ( ~n12145 & n12177 ) | ( n12176 & n12177 ) ;
  assign n12179 = ( n12006 & n12136 ) | ( n12006 & ~n12178 ) | ( n12136 & ~n12178 ) ;
  assign n12180 = ( ~n12006 & n12136 ) | ( ~n12006 & n12178 ) | ( n12136 & n12178 ) ;
  assign n12181 = ( ~n12136 & n12179 ) | ( ~n12136 & n12180 ) | ( n12179 & n12180 ) ;
  assign n12182 = n2294 & n5374 ;
  assign n12183 = x93 & n5378 ;
  assign n12184 = x94 | n12183 ;
  assign n12185 = ( n5380 & n12183 ) | ( n5380 & n12184 ) | ( n12183 & n12184 ) ;
  assign n12186 = x92 & n5638 ;
  assign n12187 = n12185 | n12186 ;
  assign n12188 = ( x50 & n12182 ) | ( x50 & ~n12187 ) | ( n12182 & ~n12187 ) ;
  assign n12189 = ( ~x50 & n12187 ) | ( ~x50 & n12188 ) | ( n12187 & n12188 ) ;
  assign n12190 = ( ~n12182 & n12188 ) | ( ~n12182 & n12189 ) | ( n12188 & n12189 ) ;
  assign n12191 = ( n12018 & n12181 ) | ( n12018 & ~n12190 ) | ( n12181 & ~n12190 ) ;
  assign n12192 = ( ~n12018 & n12181 ) | ( ~n12018 & n12190 ) | ( n12181 & n12190 ) ;
  assign n12193 = ( ~n12181 & n12191 ) | ( ~n12181 & n12192 ) | ( n12191 & n12192 ) ;
  assign n12194 = n2585 & n4787 ;
  assign n12195 = x96 & n4791 ;
  assign n12196 = x97 | n12195 ;
  assign n12197 = ( n4793 & n12195 ) | ( n4793 & n12196 ) | ( n12195 & n12196 ) ;
  assign n12198 = x95 & n5030 ;
  assign n12199 = n12197 | n12198 ;
  assign n12200 = ( x47 & n12194 ) | ( x47 & ~n12199 ) | ( n12194 & ~n12199 ) ;
  assign n12201 = ( ~x47 & n12199 ) | ( ~x47 & n12200 ) | ( n12199 & n12200 ) ;
  assign n12202 = ( ~n12194 & n12200 ) | ( ~n12194 & n12201 ) | ( n12200 & n12201 ) ;
  assign n12203 = ( n12021 & n12193 ) | ( n12021 & n12202 ) | ( n12193 & n12202 ) ;
  assign n12204 = ( ~n12021 & n12193 ) | ( ~n12021 & n12202 ) | ( n12193 & n12202 ) ;
  assign n12205 = ( n12021 & ~n12203 ) | ( n12021 & n12204 ) | ( ~n12203 & n12204 ) ;
  assign n12206 = n3162 & n4227 ;
  assign n12207 = x99 & n4231 ;
  assign n12208 = x100 | n12207 ;
  assign n12209 = ( n4233 & n12207 ) | ( n4233 & n12208 ) | ( n12207 & n12208 ) ;
  assign n12210 = x98 & n4470 ;
  assign n12211 = n12209 | n12210 ;
  assign n12212 = ( x44 & n12206 ) | ( x44 & ~n12211 ) | ( n12206 & ~n12211 ) ;
  assign n12213 = ( ~x44 & n12211 ) | ( ~x44 & n12212 ) | ( n12211 & n12212 ) ;
  assign n12214 = ( ~n12206 & n12212 ) | ( ~n12206 & n12213 ) | ( n12212 & n12213 ) ;
  assign n12215 = ( n12033 & n12205 ) | ( n12033 & n12214 ) | ( n12205 & n12214 ) ;
  assign n12216 = ( ~n12033 & n12205 ) | ( ~n12033 & n12214 ) | ( n12205 & n12214 ) ;
  assign n12217 = ( n12033 & ~n12215 ) | ( n12033 & n12216 ) | ( ~n12215 & n12216 ) ;
  assign n12218 = n3650 & n3715 ;
  assign n12219 = x102 & n3719 ;
  assign n12220 = x103 | n12219 ;
  assign n12221 = ( n3721 & n12219 ) | ( n3721 & n12220 ) | ( n12219 & n12220 ) ;
  assign n12222 = x101 & n3922 ;
  assign n12223 = n12221 | n12222 ;
  assign n12224 = ( x41 & n12218 ) | ( x41 & ~n12223 ) | ( n12218 & ~n12223 ) ;
  assign n12225 = ( ~x41 & n12223 ) | ( ~x41 & n12224 ) | ( n12223 & n12224 ) ;
  assign n12226 = ( ~n12218 & n12224 ) | ( ~n12218 & n12225 ) | ( n12224 & n12225 ) ;
  assign n12227 = ( n12045 & n12217 ) | ( n12045 & n12226 ) | ( n12217 & n12226 ) ;
  assign n12228 = ( ~n12045 & n12217 ) | ( ~n12045 & n12226 ) | ( n12217 & n12226 ) ;
  assign n12229 = ( n12045 & ~n12227 ) | ( n12045 & n12228 ) | ( ~n12227 & n12228 ) ;
  assign n12230 = ( n12048 & n12127 ) | ( n12048 & n12229 ) | ( n12127 & n12229 ) ;
  assign n12231 = ( ~n12048 & n12127 ) | ( ~n12048 & n12229 ) | ( n12127 & n12229 ) ;
  assign n12232 = ( n12048 & ~n12230 ) | ( n12048 & n12231 ) | ( ~n12230 & n12231 ) ;
  assign n12233 = n2766 & n4734 ;
  assign n12234 = x108 & n2770 ;
  assign n12235 = x109 | n12234 ;
  assign n12236 = ( n2772 & n12234 ) | ( n2772 & n12235 ) | ( n12234 & n12235 ) ;
  assign n12237 = x107 & n2943 ;
  assign n12238 = n12236 | n12237 ;
  assign n12239 = ( x35 & n12233 ) | ( x35 & ~n12238 ) | ( n12233 & ~n12238 ) ;
  assign n12240 = ( ~x35 & n12238 ) | ( ~x35 & n12239 ) | ( n12238 & n12239 ) ;
  assign n12241 = ( ~n12233 & n12239 ) | ( ~n12233 & n12240 ) | ( n12239 & n12240 ) ;
  assign n12242 = ( n12051 & n12232 ) | ( n12051 & n12241 ) | ( n12232 & n12241 ) ;
  assign n12243 = ( ~n12051 & n12232 ) | ( ~n12051 & n12241 ) | ( n12232 & n12241 ) ;
  assign n12244 = ( n12051 & ~n12242 ) | ( n12051 & n12243 ) | ( ~n12242 & n12243 ) ;
  assign n12245 = n2320 & n5145 ;
  assign n12246 = x111 & n2324 ;
  assign n12247 = x112 | n12246 ;
  assign n12248 = ( n2326 & n12246 ) | ( n2326 & n12247 ) | ( n12246 & n12247 ) ;
  assign n12249 = x110 & n2497 ;
  assign n12250 = n12248 | n12249 ;
  assign n12251 = ( x32 & n12245 ) | ( x32 & ~n12250 ) | ( n12245 & ~n12250 ) ;
  assign n12252 = ( ~x32 & n12250 ) | ( ~x32 & n12251 ) | ( n12250 & n12251 ) ;
  assign n12253 = ( ~n12245 & n12251 ) | ( ~n12245 & n12252 ) | ( n12251 & n12252 ) ;
  assign n12254 = ( n12054 & n12244 ) | ( n12054 & n12253 ) | ( n12244 & n12253 ) ;
  assign n12255 = ( n12054 & ~n12244 ) | ( n12054 & n12253 ) | ( ~n12244 & n12253 ) ;
  assign n12256 = ( n12244 & ~n12254 ) | ( n12244 & n12255 ) | ( ~n12254 & n12255 ) ;
  assign n12257 = ( n12057 & n12118 ) | ( n12057 & n12256 ) | ( n12118 & n12256 ) ;
  assign n12258 = ( n12057 & ~n12118 ) | ( n12057 & n12256 ) | ( ~n12118 & n12256 ) ;
  assign n12259 = ( n12118 & ~n12257 ) | ( n12118 & n12258 ) | ( ~n12257 & n12258 ) ;
  assign n12260 = ( n12060 & n12109 ) | ( n12060 & n12259 ) | ( n12109 & n12259 ) ;
  assign n12261 = ( n12060 & ~n12109 ) | ( n12060 & n12259 ) | ( ~n12109 & n12259 ) ;
  assign n12262 = ( n12109 & ~n12260 ) | ( n12109 & n12261 ) | ( ~n12260 & n12261 ) ;
  assign n12263 = n1297 & n7113 ;
  assign n12264 = x120 & n1301 ;
  assign n12265 = x121 | n12264 ;
  assign n12266 = ( n1303 & n12264 ) | ( n1303 & n12265 ) | ( n12264 & n12265 ) ;
  assign n12267 = x119 & n1426 ;
  assign n12268 = n12266 | n12267 ;
  assign n12269 = ( x23 & n12263 ) | ( x23 & ~n12268 ) | ( n12263 & ~n12268 ) ;
  assign n12270 = ( ~x23 & n12268 ) | ( ~x23 & n12269 ) | ( n12268 & n12269 ) ;
  assign n12271 = ( ~n12263 & n12269 ) | ( ~n12263 & n12270 ) | ( n12269 & n12270 ) ;
  assign n12272 = ( n12063 & n12262 ) | ( n12063 & n12271 ) | ( n12262 & n12271 ) ;
  assign n12273 = ( n12063 & ~n12262 ) | ( n12063 & n12271 ) | ( ~n12262 & n12271 ) ;
  assign n12274 = ( n12262 & ~n12272 ) | ( n12262 & n12273 ) | ( ~n12272 & n12273 ) ;
  assign n12275 = ( n12066 & n12100 ) | ( n12066 & n12274 ) | ( n12100 & n12274 ) ;
  assign n12276 = ( n12066 & ~n12100 ) | ( n12066 & n12274 ) | ( ~n12100 & n12274 ) ;
  assign n12277 = ( n12100 & ~n12275 ) | ( n12100 & n12276 ) | ( ~n12275 & n12276 ) ;
  assign n12278 = n810 & n8846 ;
  assign n12279 = x126 & n814 ;
  assign n12280 = x127 | n12279 ;
  assign n12281 = ( n816 & n12279 ) | ( n816 & n12280 ) | ( n12279 & n12280 ) ;
  assign n12282 = x125 & n885 ;
  assign n12283 = n12281 | n12282 ;
  assign n12284 = ( x17 & n12278 ) | ( x17 & ~n12283 ) | ( n12278 & ~n12283 ) ;
  assign n12285 = ( ~x17 & n12283 ) | ( ~x17 & n12284 ) | ( n12283 & n12284 ) ;
  assign n12286 = ( ~n12278 & n12284 ) | ( ~n12278 & n12285 ) | ( n12284 & n12285 ) ;
  assign n12287 = ( n12078 & n12277 ) | ( n12078 & n12286 ) | ( n12277 & n12286 ) ;
  assign n12288 = ( n12078 & ~n12277 ) | ( n12078 & n12286 ) | ( ~n12277 & n12286 ) ;
  assign n12289 = ( n12277 & ~n12287 ) | ( n12277 & n12288 ) | ( ~n12287 & n12288 ) ;
  assign n12290 = ( n12086 & n12089 ) | ( n12086 & n12289 ) | ( n12089 & n12289 ) ;
  assign n12291 = ( ~n12086 & n12089 ) | ( ~n12086 & n12289 ) | ( n12089 & n12289 ) ;
  assign n12292 = ( n12086 & ~n12290 ) | ( n12086 & n12291 ) | ( ~n12290 & n12291 ) ;
  assign n12293 = n810 & n8865 ;
  assign n12294 = x127 & n814 ;
  assign n12295 = x126 | n12294 ;
  assign n12296 = ( n885 & n12294 ) | ( n885 & n12295 ) | ( n12294 & n12295 ) ;
  assign n12297 = ( x17 & n12293 ) | ( x17 & ~n12296 ) | ( n12293 & ~n12296 ) ;
  assign n12298 = ( ~x17 & n12296 ) | ( ~x17 & n12297 ) | ( n12296 & n12297 ) ;
  assign n12299 = ( ~n12293 & n12297 ) | ( ~n12293 & n12298 ) | ( n12297 & n12298 ) ;
  assign n12300 = n1016 & n8331 ;
  assign n12301 = x124 & n1020 ;
  assign n12302 = x125 | n12301 ;
  assign n12303 = ( n1022 & n12301 ) | ( n1022 & n12302 ) | ( n12301 & n12302 ) ;
  assign n12304 = x123 & n1145 ;
  assign n12305 = n12303 | n12304 ;
  assign n12306 = ( x20 & n12300 ) | ( x20 & ~n12305 ) | ( n12300 & ~n12305 ) ;
  assign n12307 = ( ~x20 & n12305 ) | ( ~x20 & n12306 ) | ( n12305 & n12306 ) ;
  assign n12308 = ( ~n12300 & n12306 ) | ( ~n12300 & n12307 ) | ( n12306 & n12307 ) ;
  assign n12309 = n1297 & n7582 ;
  assign n12310 = x121 & n1301 ;
  assign n12311 = x122 | n12310 ;
  assign n12312 = ( n1303 & n12310 ) | ( n1303 & n12311 ) | ( n12310 & n12311 ) ;
  assign n12313 = x120 & n1426 ;
  assign n12314 = n12312 | n12313 ;
  assign n12315 = ( x23 & n12309 ) | ( x23 & ~n12314 ) | ( n12309 & ~n12314 ) ;
  assign n12316 = ( ~x23 & n12314 ) | ( ~x23 & n12315 ) | ( n12314 & n12315 ) ;
  assign n12317 = ( ~n12309 & n12315 ) | ( ~n12309 & n12316 ) | ( n12315 & n12316 ) ;
  assign n12318 = n1617 & n6645 ;
  assign n12319 = x118 & n1621 ;
  assign n12320 = x119 | n12319 ;
  assign n12321 = ( n1623 & n12319 ) | ( n1623 & n12320 ) | ( n12319 & n12320 ) ;
  assign n12322 = x117 & n1749 ;
  assign n12323 = n12321 | n12322 ;
  assign n12324 = ( x26 & n12318 ) | ( x26 & ~n12323 ) | ( n12318 & ~n12323 ) ;
  assign n12325 = ( ~x26 & n12323 ) | ( ~x26 & n12324 ) | ( n12323 & n12324 ) ;
  assign n12326 = ( ~n12318 & n12324 ) | ( ~n12318 & n12325 ) | ( n12324 & n12325 ) ;
  assign n12327 = n1949 & n5977 ;
  assign n12328 = x115 & n1953 ;
  assign n12329 = x116 | n12328 ;
  assign n12330 = ( n1955 & n12328 ) | ( n1955 & n12329 ) | ( n12328 & n12329 ) ;
  assign n12331 = x114 & n2114 ;
  assign n12332 = n12330 | n12331 ;
  assign n12333 = ( x29 & n12327 ) | ( x29 & ~n12332 ) | ( n12327 & ~n12332 ) ;
  assign n12334 = ( ~x29 & n12332 ) | ( ~x29 & n12333 ) | ( n12332 & n12333 ) ;
  assign n12335 = ( ~n12327 & n12333 ) | ( ~n12327 & n12334 ) | ( n12333 & n12334 ) ;
  assign n12336 = n2320 & n5542 ;
  assign n12337 = x112 & n2324 ;
  assign n12338 = x113 | n12337 ;
  assign n12339 = ( n2326 & n12337 ) | ( n2326 & n12338 ) | ( n12337 & n12338 ) ;
  assign n12340 = x111 & n2497 ;
  assign n12341 = n12339 | n12340 ;
  assign n12342 = ( x32 & n12336 ) | ( x32 & ~n12341 ) | ( n12336 & ~n12341 ) ;
  assign n12343 = ( ~x32 & n12341 ) | ( ~x32 & n12342 ) | ( n12341 & n12342 ) ;
  assign n12344 = ( ~n12336 & n12342 ) | ( ~n12336 & n12343 ) | ( n12342 & n12343 ) ;
  assign n12345 = n3665 & n3715 ;
  assign n12346 = x103 & n3719 ;
  assign n12347 = x104 | n12346 ;
  assign n12348 = ( n3721 & n12346 ) | ( n3721 & n12347 ) | ( n12346 & n12347 ) ;
  assign n12349 = x102 & n3922 ;
  assign n12350 = n12348 | n12349 ;
  assign n12351 = ( x41 & n12345 ) | ( x41 & ~n12350 ) | ( n12345 & ~n12350 ) ;
  assign n12352 = ( ~x41 & n12350 ) | ( ~x41 & n12351 ) | ( n12350 & n12351 ) ;
  assign n12353 = ( ~n12345 & n12351 ) | ( ~n12345 & n12352 ) | ( n12351 & n12352 ) ;
  assign n12354 = n3326 & n4227 ;
  assign n12355 = x100 & n4231 ;
  assign n12356 = x101 | n12355 ;
  assign n12357 = ( n4233 & n12355 ) | ( n4233 & n12356 ) | ( n12355 & n12356 ) ;
  assign n12358 = x99 & n4470 ;
  assign n12359 = n12357 | n12358 ;
  assign n12360 = ( x44 & n12354 ) | ( x44 & ~n12359 ) | ( n12354 & ~n12359 ) ;
  assign n12361 = ( ~x44 & n12359 ) | ( ~x44 & n12360 ) | ( n12359 & n12360 ) ;
  assign n12362 = ( ~n12354 & n12360 ) | ( ~n12354 & n12361 ) | ( n12360 & n12361 ) ;
  assign n12363 = n2042 & n6027 ;
  assign n12364 = x91 & n6031 ;
  assign n12365 = x92 | n12364 ;
  assign n12366 = ( n6033 & n12364 ) | ( n6033 & n12365 ) | ( n12364 & n12365 ) ;
  assign n12367 = x90 & n6303 ;
  assign n12368 = n12366 | n12367 ;
  assign n12369 = ( x53 & n12363 ) | ( x53 & ~n12368 ) | ( n12363 & ~n12368 ) ;
  assign n12370 = ( ~x53 & n12368 ) | ( ~x53 & n12369 ) | ( n12368 & n12369 ) ;
  assign n12371 = ( ~n12363 & n12369 ) | ( ~n12363 & n12370 ) | ( n12369 & n12370 ) ;
  assign n12372 = n1585 & n6713 ;
  assign n12373 = x88 & n6717 ;
  assign n12374 = x89 | n12373 ;
  assign n12375 = ( n6719 & n12373 ) | ( n6719 & n12374 ) | ( n12373 & n12374 ) ;
  assign n12376 = x87 & n6980 ;
  assign n12377 = n12375 | n12376 ;
  assign n12378 = ( x56 & n12372 ) | ( x56 & ~n12377 ) | ( n12372 & ~n12377 ) ;
  assign n12379 = ( ~x56 & n12377 ) | ( ~x56 & n12378 ) | ( n12377 & n12378 ) ;
  assign n12380 = ( ~n12372 & n12378 ) | ( ~n12372 & n12379 ) | ( n12378 & n12379 ) ;
  assign n12381 = n1366 & n7423 ;
  assign n12382 = x85 & n7427 ;
  assign n12383 = x86 | n12382 ;
  assign n12384 = ( n7429 & n12382 ) | ( n7429 & n12383 ) | ( n12382 & n12383 ) ;
  assign n12385 = x84 & n7708 ;
  assign n12386 = n12384 | n12385 ;
  assign n12387 = ( x59 & n12381 ) | ( x59 & ~n12386 ) | ( n12381 & ~n12386 ) ;
  assign n12388 = ( ~x59 & n12386 ) | ( ~x59 & n12387 ) | ( n12386 & n12387 ) ;
  assign n12389 = ( ~n12381 & n12387 ) | ( ~n12381 & n12388 ) | ( n12387 & n12388 ) ;
  assign n12390 = x79 & n8927 ;
  assign n12391 = ( ~x80 & n8693 ) | ( ~x80 & n8927 ) | ( n8693 & n8927 ) ;
  assign n12392 = ( n8693 & n12390 ) | ( n8693 & ~n12391 ) | ( n12390 & ~n12391 ) ;
  assign n12393 = n1082 & n8154 ;
  assign n12394 = x82 & n8158 ;
  assign n12395 = x83 | n12394 ;
  assign n12396 = ( n8160 & n12394 ) | ( n8160 & n12395 ) | ( n12394 & n12395 ) ;
  assign n12397 = x81 & n8439 ;
  assign n12398 = n12396 | n12397 ;
  assign n12399 = ( x62 & n12393 ) | ( x62 & ~n12398 ) | ( n12393 & ~n12398 ) ;
  assign n12400 = ( ~x62 & n12398 ) | ( ~x62 & n12399 ) | ( n12398 & n12399 ) ;
  assign n12401 = ( ~n12393 & n12399 ) | ( ~n12393 & n12400 ) | ( n12399 & n12400 ) ;
  assign n12402 = ( n12167 & ~n12392 ) | ( n12167 & n12401 ) | ( ~n12392 & n12401 ) ;
  assign n12403 = ( n12167 & n12392 ) | ( n12167 & n12401 ) | ( n12392 & n12401 ) ;
  assign n12404 = ( n12392 & n12402 ) | ( n12392 & ~n12403 ) | ( n12402 & ~n12403 ) ;
  assign n12405 = ( n12170 & n12389 ) | ( n12170 & ~n12404 ) | ( n12389 & ~n12404 ) ;
  assign n12406 = ( ~n12170 & n12389 ) | ( ~n12170 & n12404 ) | ( n12389 & n12404 ) ;
  assign n12407 = ( ~n12389 & n12405 ) | ( ~n12389 & n12406 ) | ( n12405 & n12406 ) ;
  assign n12408 = ( n12173 & n12380 ) | ( n12173 & ~n12407 ) | ( n12380 & ~n12407 ) ;
  assign n12409 = ( ~n12173 & n12380 ) | ( ~n12173 & n12407 ) | ( n12380 & n12407 ) ;
  assign n12410 = ( ~n12380 & n12408 ) | ( ~n12380 & n12409 ) | ( n12408 & n12409 ) ;
  assign n12411 = ( n12176 & n12371 ) | ( n12176 & ~n12410 ) | ( n12371 & ~n12410 ) ;
  assign n12412 = ( ~n12176 & n12371 ) | ( ~n12176 & n12410 ) | ( n12371 & n12410 ) ;
  assign n12413 = ( ~n12371 & n12411 ) | ( ~n12371 & n12412 ) | ( n12411 & n12412 ) ;
  assign n12414 = n2434 & n5374 ;
  assign n12415 = x94 & n5378 ;
  assign n12416 = x95 | n12415 ;
  assign n12417 = ( n5380 & n12415 ) | ( n5380 & n12416 ) | ( n12415 & n12416 ) ;
  assign n12418 = x93 & n5638 ;
  assign n12419 = n12417 | n12418 ;
  assign n12420 = ( x50 & n12414 ) | ( x50 & ~n12419 ) | ( n12414 & ~n12419 ) ;
  assign n12421 = ( ~x50 & n12419 ) | ( ~x50 & n12420 ) | ( n12419 & n12420 ) ;
  assign n12422 = ( ~n12414 & n12420 ) | ( ~n12414 & n12421 ) | ( n12420 & n12421 ) ;
  assign n12423 = ( n12179 & ~n12413 ) | ( n12179 & n12422 ) | ( ~n12413 & n12422 ) ;
  assign n12424 = ( n12179 & n12413 ) | ( n12179 & n12422 ) | ( n12413 & n12422 ) ;
  assign n12425 = ( n12413 & n12423 ) | ( n12413 & ~n12424 ) | ( n12423 & ~n12424 ) ;
  assign n12426 = n2725 & n4787 ;
  assign n12427 = x97 & n4791 ;
  assign n12428 = x98 | n12427 ;
  assign n12429 = ( n4793 & n12427 ) | ( n4793 & n12428 ) | ( n12427 & n12428 ) ;
  assign n12430 = x96 & n5030 ;
  assign n12431 = n12429 | n12430 ;
  assign n12432 = ( x47 & n12426 ) | ( x47 & ~n12431 ) | ( n12426 & ~n12431 ) ;
  assign n12433 = ( ~x47 & n12431 ) | ( ~x47 & n12432 ) | ( n12431 & n12432 ) ;
  assign n12434 = ( ~n12426 & n12432 ) | ( ~n12426 & n12433 ) | ( n12432 & n12433 ) ;
  assign n12435 = ( n12191 & n12425 ) | ( n12191 & ~n12434 ) | ( n12425 & ~n12434 ) ;
  assign n12436 = ( ~n12191 & n12425 ) | ( ~n12191 & n12434 ) | ( n12425 & n12434 ) ;
  assign n12437 = ( ~n12425 & n12435 ) | ( ~n12425 & n12436 ) | ( n12435 & n12436 ) ;
  assign n12438 = ( n12203 & n12362 ) | ( n12203 & n12437 ) | ( n12362 & n12437 ) ;
  assign n12439 = ( n12203 & ~n12362 ) | ( n12203 & n12437 ) | ( ~n12362 & n12437 ) ;
  assign n12440 = ( n12362 & ~n12438 ) | ( n12362 & n12439 ) | ( ~n12438 & n12439 ) ;
  assign n12441 = ( n12215 & n12353 ) | ( n12215 & n12440 ) | ( n12353 & n12440 ) ;
  assign n12442 = ( n12215 & ~n12353 ) | ( n12215 & n12440 ) | ( ~n12353 & n12440 ) ;
  assign n12443 = ( n12353 & ~n12441 ) | ( n12353 & n12442 ) | ( ~n12441 & n12442 ) ;
  assign n12444 = n3224 & n4362 ;
  assign n12445 = x106 & n3228 ;
  assign n12446 = x107 | n12445 ;
  assign n12447 = ( n3230 & n12445 ) | ( n3230 & n12446 ) | ( n12445 & n12446 ) ;
  assign n12448 = x105 & n3413 ;
  assign n12449 = n12447 | n12448 ;
  assign n12450 = ( x38 & n12444 ) | ( x38 & ~n12449 ) | ( n12444 & ~n12449 ) ;
  assign n12451 = ( ~x38 & n12449 ) | ( ~x38 & n12450 ) | ( n12449 & n12450 ) ;
  assign n12452 = ( ~n12444 & n12450 ) | ( ~n12444 & n12451 ) | ( n12450 & n12451 ) ;
  assign n12453 = ( n12227 & n12443 ) | ( n12227 & n12452 ) | ( n12443 & n12452 ) ;
  assign n12454 = ( ~n12227 & n12443 ) | ( ~n12227 & n12452 ) | ( n12443 & n12452 ) ;
  assign n12455 = ( n12227 & ~n12453 ) | ( n12227 & n12454 ) | ( ~n12453 & n12454 ) ;
  assign n12456 = n2766 & n4934 ;
  assign n12457 = x109 & n2770 ;
  assign n12458 = x110 | n12457 ;
  assign n12459 = ( n2772 & n12457 ) | ( n2772 & n12458 ) | ( n12457 & n12458 ) ;
  assign n12460 = x108 & n2943 ;
  assign n12461 = n12459 | n12460 ;
  assign n12462 = ( x35 & n12456 ) | ( x35 & ~n12461 ) | ( n12456 & ~n12461 ) ;
  assign n12463 = ( ~x35 & n12461 ) | ( ~x35 & n12462 ) | ( n12461 & n12462 ) ;
  assign n12464 = ( ~n12456 & n12462 ) | ( ~n12456 & n12463 ) | ( n12462 & n12463 ) ;
  assign n12465 = ( n12230 & n12455 ) | ( n12230 & n12464 ) | ( n12455 & n12464 ) ;
  assign n12466 = ( ~n12230 & n12455 ) | ( ~n12230 & n12464 ) | ( n12455 & n12464 ) ;
  assign n12467 = ( n12230 & ~n12465 ) | ( n12230 & n12466 ) | ( ~n12465 & n12466 ) ;
  assign n12468 = ( n12242 & n12344 ) | ( n12242 & n12467 ) | ( n12344 & n12467 ) ;
  assign n12469 = ( n12242 & ~n12344 ) | ( n12242 & n12467 ) | ( ~n12344 & n12467 ) ;
  assign n12470 = ( n12344 & ~n12468 ) | ( n12344 & n12469 ) | ( ~n12468 & n12469 ) ;
  assign n12471 = ( n12254 & n12335 ) | ( n12254 & n12470 ) | ( n12335 & n12470 ) ;
  assign n12472 = ( n12254 & ~n12335 ) | ( n12254 & n12470 ) | ( ~n12335 & n12470 ) ;
  assign n12473 = ( n12335 & ~n12471 ) | ( n12335 & n12472 ) | ( ~n12471 & n12472 ) ;
  assign n12474 = ( n12257 & n12326 ) | ( n12257 & n12473 ) | ( n12326 & n12473 ) ;
  assign n12475 = ( n12257 & ~n12326 ) | ( n12257 & n12473 ) | ( ~n12326 & n12473 ) ;
  assign n12476 = ( n12326 & ~n12474 ) | ( n12326 & n12475 ) | ( ~n12474 & n12475 ) ;
  assign n12477 = ( n12260 & n12317 ) | ( n12260 & n12476 ) | ( n12317 & n12476 ) ;
  assign n12478 = ( ~n12260 & n12317 ) | ( ~n12260 & n12476 ) | ( n12317 & n12476 ) ;
  assign n12479 = ( n12260 & ~n12477 ) | ( n12260 & n12478 ) | ( ~n12477 & n12478 ) ;
  assign n12480 = ( n12272 & n12308 ) | ( n12272 & n12479 ) | ( n12308 & n12479 ) ;
  assign n12481 = ( n12272 & ~n12308 ) | ( n12272 & n12479 ) | ( ~n12308 & n12479 ) ;
  assign n12482 = ( n12308 & ~n12480 ) | ( n12308 & n12481 ) | ( ~n12480 & n12481 ) ;
  assign n12483 = ( n12275 & n12299 ) | ( n12275 & n12482 ) | ( n12299 & n12482 ) ;
  assign n12484 = ( ~n12275 & n12299 ) | ( ~n12275 & n12482 ) | ( n12299 & n12482 ) ;
  assign n12485 = ( n12275 & ~n12483 ) | ( n12275 & n12484 ) | ( ~n12483 & n12484 ) ;
  assign n12486 = ( n12287 & n12290 ) | ( n12287 & n12485 ) | ( n12290 & n12485 ) ;
  assign n12487 = ( ~n12287 & n12290 ) | ( ~n12287 & n12485 ) | ( n12290 & n12485 ) ;
  assign n12488 = ( n12287 & ~n12486 ) | ( n12287 & n12487 ) | ( ~n12486 & n12487 ) ;
  assign n12489 = n1016 & n8587 ;
  assign n12490 = x125 & n1020 ;
  assign n12491 = x126 | n12490 ;
  assign n12492 = ( n1022 & n12490 ) | ( n1022 & n12491 ) | ( n12490 & n12491 ) ;
  assign n12493 = x124 & n1145 ;
  assign n12494 = n12492 | n12493 ;
  assign n12495 = ( x20 & n12489 ) | ( x20 & ~n12494 ) | ( n12489 & ~n12494 ) ;
  assign n12496 = ( ~x20 & n12494 ) | ( ~x20 & n12495 ) | ( n12494 & n12495 ) ;
  assign n12497 = ( ~n12489 & n12495 ) | ( ~n12489 & n12496 ) | ( n12495 & n12496 ) ;
  assign n12498 = n1617 & n7098 ;
  assign n12499 = x119 & n1621 ;
  assign n12500 = x120 | n12499 ;
  assign n12501 = ( n1623 & n12499 ) | ( n1623 & n12500 ) | ( n12499 & n12500 ) ;
  assign n12502 = x118 & n1749 ;
  assign n12503 = n12501 | n12502 ;
  assign n12504 = ( x26 & n12498 ) | ( x26 & ~n12503 ) | ( n12498 & ~n12503 ) ;
  assign n12505 = ( ~x26 & n12503 ) | ( ~x26 & n12504 ) | ( n12503 & n12504 ) ;
  assign n12506 = ( ~n12498 & n12504 ) | ( ~n12498 & n12505 ) | ( n12504 & n12505 ) ;
  assign n12507 = n2320 & n5750 ;
  assign n12508 = x113 & n2324 ;
  assign n12509 = x114 | n12508 ;
  assign n12510 = ( n2326 & n12508 ) | ( n2326 & n12509 ) | ( n12508 & n12509 ) ;
  assign n12511 = x112 & n2497 ;
  assign n12512 = n12510 | n12511 ;
  assign n12513 = ( x32 & n12507 ) | ( x32 & ~n12512 ) | ( n12507 & ~n12512 ) ;
  assign n12514 = ( ~x32 & n12512 ) | ( ~x32 & n12513 ) | ( n12512 & n12513 ) ;
  assign n12515 = ( ~n12507 & n12513 ) | ( ~n12507 & n12514 ) | ( n12513 & n12514 ) ;
  assign n12516 = n3224 & n4377 ;
  assign n12517 = x107 & n3228 ;
  assign n12518 = x108 | n12517 ;
  assign n12519 = ( n3230 & n12517 ) | ( n3230 & n12518 ) | ( n12517 & n12518 ) ;
  assign n12520 = x106 & n3413 ;
  assign n12521 = n12519 | n12520 ;
  assign n12522 = ( x38 & n12516 ) | ( x38 & ~n12521 ) | ( n12516 & ~n12521 ) ;
  assign n12523 = ( ~x38 & n12521 ) | ( ~x38 & n12522 ) | ( n12521 & n12522 ) ;
  assign n12524 = ( ~n12516 & n12522 ) | ( ~n12516 & n12523 ) | ( n12522 & n12523 ) ;
  assign n12525 = n3715 & n3998 ;
  assign n12526 = x104 & n3719 ;
  assign n12527 = x105 | n12526 ;
  assign n12528 = ( n3721 & n12526 ) | ( n3721 & n12527 ) | ( n12526 & n12527 ) ;
  assign n12529 = x103 & n3922 ;
  assign n12530 = n12528 | n12529 ;
  assign n12531 = ( x41 & n12525 ) | ( x41 & ~n12530 ) | ( n12525 & ~n12530 ) ;
  assign n12532 = ( ~x41 & n12530 ) | ( ~x41 & n12531 ) | ( n12530 & n12531 ) ;
  assign n12533 = ( ~n12525 & n12531 ) | ( ~n12525 & n12532 ) | ( n12531 & n12532 ) ;
  assign n12534 = n3486 & n4227 ;
  assign n12535 = x101 & n4231 ;
  assign n12536 = x102 | n12535 ;
  assign n12537 = ( n4233 & n12535 ) | ( n4233 & n12536 ) | ( n12535 & n12536 ) ;
  assign n12538 = x100 & n4470 ;
  assign n12539 = n12537 | n12538 ;
  assign n12540 = ( x44 & n12534 ) | ( x44 & ~n12539 ) | ( n12534 & ~n12539 ) ;
  assign n12541 = ( ~x44 & n12539 ) | ( ~x44 & n12540 ) | ( n12539 & n12540 ) ;
  assign n12542 = ( ~n12534 & n12540 ) | ( ~n12534 & n12541 ) | ( n12540 & n12541 ) ;
  assign n12543 = n2449 & n5374 ;
  assign n12544 = x95 & n5378 ;
  assign n12545 = x96 | n12544 ;
  assign n12546 = ( n5380 & n12544 ) | ( n5380 & n12545 ) | ( n12544 & n12545 ) ;
  assign n12547 = x94 & n5638 ;
  assign n12548 = n12546 | n12547 ;
  assign n12549 = ( x50 & n12543 ) | ( x50 & ~n12548 ) | ( n12543 & ~n12548 ) ;
  assign n12550 = ( ~x50 & n12548 ) | ( ~x50 & n12549 ) | ( n12548 & n12549 ) ;
  assign n12551 = ( ~n12543 & n12549 ) | ( ~n12543 & n12550 ) | ( n12549 & n12550 ) ;
  assign n12552 = n2057 & n6027 ;
  assign n12553 = x92 & n6031 ;
  assign n12554 = x93 | n12553 ;
  assign n12555 = ( n6033 & n12553 ) | ( n6033 & n12554 ) | ( n12553 & n12554 ) ;
  assign n12556 = x91 & n6303 ;
  assign n12557 = n12555 | n12556 ;
  assign n12558 = ( x53 & n12552 ) | ( x53 & ~n12557 ) | ( n12552 & ~n12557 ) ;
  assign n12559 = ( ~x53 & n12557 ) | ( ~x53 & n12558 ) | ( n12557 & n12558 ) ;
  assign n12560 = ( ~n12552 & n12558 ) | ( ~n12552 & n12559 ) | ( n12558 & n12559 ) ;
  assign n12561 = n1701 & n6713 ;
  assign n12562 = x89 & n6717 ;
  assign n12563 = x90 | n12562 ;
  assign n12564 = ( n6719 & n12562 ) | ( n6719 & n12563 ) | ( n12562 & n12563 ) ;
  assign n12565 = x88 & n6980 ;
  assign n12566 = n12564 | n12565 ;
  assign n12567 = ( x56 & n12561 ) | ( x56 & ~n12566 ) | ( n12561 & ~n12566 ) ;
  assign n12568 = ( ~x56 & n12566 ) | ( ~x56 & n12567 ) | ( n12566 & n12567 ) ;
  assign n12569 = ( ~n12561 & n12567 ) | ( ~n12561 & n12568 ) | ( n12567 & n12568 ) ;
  assign n12570 = n1466 & n7423 ;
  assign n12571 = x86 & n7427 ;
  assign n12572 = x87 | n12571 ;
  assign n12573 = ( n7429 & n12571 ) | ( n7429 & n12572 ) | ( n12571 & n12572 ) ;
  assign n12574 = x85 & n7708 ;
  assign n12575 = n12573 | n12574 ;
  assign n12576 = ( x59 & n12570 ) | ( x59 & ~n12575 ) | ( n12570 & ~n12575 ) ;
  assign n12577 = ( ~x59 & n12575 ) | ( ~x59 & n12576 ) | ( n12575 & n12576 ) ;
  assign n12578 = ( ~n12570 & n12576 ) | ( ~n12570 & n12577 ) | ( n12576 & n12577 ) ;
  assign n12579 = n1097 & n8154 ;
  assign n12580 = x83 & n8158 ;
  assign n12581 = x84 | n12580 ;
  assign n12582 = ( n8160 & n12580 ) | ( n8160 & n12581 ) | ( n12580 & n12581 ) ;
  assign n12583 = x82 & n8439 ;
  assign n12584 = n12582 | n12583 ;
  assign n12585 = ( x62 & n12579 ) | ( x62 & ~n12584 ) | ( n12579 & ~n12584 ) ;
  assign n12586 = ( ~x62 & n12584 ) | ( ~x62 & n12585 ) | ( n12584 & n12585 ) ;
  assign n12587 = ( ~n12579 & n12585 ) | ( ~n12579 & n12586 ) | ( n12585 & n12586 ) ;
  assign n12588 = x80 & n8927 ;
  assign n12589 = ( ~x81 & n8693 ) | ( ~x81 & n8927 ) | ( n8693 & n8927 ) ;
  assign n12590 = ( n8693 & n12588 ) | ( n8693 & ~n12589 ) | ( n12588 & ~n12589 ) ;
  assign n12591 = ( n12392 & n12587 ) | ( n12392 & ~n12590 ) | ( n12587 & ~n12590 ) ;
  assign n12592 = ( ~n12392 & n12587 ) | ( ~n12392 & n12590 ) | ( n12587 & n12590 ) ;
  assign n12593 = ( ~n12587 & n12591 ) | ( ~n12587 & n12592 ) | ( n12591 & n12592 ) ;
  assign n12594 = ( n12402 & n12578 ) | ( n12402 & ~n12593 ) | ( n12578 & ~n12593 ) ;
  assign n12595 = ( ~n12402 & n12578 ) | ( ~n12402 & n12593 ) | ( n12578 & n12593 ) ;
  assign n12596 = ( ~n12578 & n12594 ) | ( ~n12578 & n12595 ) | ( n12594 & n12595 ) ;
  assign n12597 = ( n12405 & n12569 ) | ( n12405 & ~n12596 ) | ( n12569 & ~n12596 ) ;
  assign n12598 = ( ~n12405 & n12569 ) | ( ~n12405 & n12596 ) | ( n12569 & n12596 ) ;
  assign n12599 = ( ~n12569 & n12597 ) | ( ~n12569 & n12598 ) | ( n12597 & n12598 ) ;
  assign n12600 = ( n12408 & n12560 ) | ( n12408 & ~n12599 ) | ( n12560 & ~n12599 ) ;
  assign n12601 = ( ~n12408 & n12560 ) | ( ~n12408 & n12599 ) | ( n12560 & n12599 ) ;
  assign n12602 = ( ~n12560 & n12600 ) | ( ~n12560 & n12601 ) | ( n12600 & n12601 ) ;
  assign n12603 = ( n12411 & n12551 ) | ( n12411 & ~n12602 ) | ( n12551 & ~n12602 ) ;
  assign n12604 = ( ~n12411 & n12551 ) | ( ~n12411 & n12602 ) | ( n12551 & n12602 ) ;
  assign n12605 = ( ~n12551 & n12603 ) | ( ~n12551 & n12604 ) | ( n12603 & n12604 ) ;
  assign n12606 = n2877 & n4787 ;
  assign n12607 = x98 & n4791 ;
  assign n12608 = x99 | n12607 ;
  assign n12609 = ( n4793 & n12607 ) | ( n4793 & n12608 ) | ( n12607 & n12608 ) ;
  assign n12610 = x97 & n5030 ;
  assign n12611 = n12609 | n12610 ;
  assign n12612 = ( x47 & n12606 ) | ( x47 & ~n12611 ) | ( n12606 & ~n12611 ) ;
  assign n12613 = ( ~x47 & n12611 ) | ( ~x47 & n12612 ) | ( n12611 & n12612 ) ;
  assign n12614 = ( ~n12606 & n12612 ) | ( ~n12606 & n12613 ) | ( n12612 & n12613 ) ;
  assign n12615 = ( n12423 & ~n12605 ) | ( n12423 & n12614 ) | ( ~n12605 & n12614 ) ;
  assign n12616 = ( n12423 & n12605 ) | ( n12423 & n12614 ) | ( n12605 & n12614 ) ;
  assign n12617 = ( n12605 & n12615 ) | ( n12605 & ~n12616 ) | ( n12615 & ~n12616 ) ;
  assign n12618 = ( n12435 & ~n12542 ) | ( n12435 & n12617 ) | ( ~n12542 & n12617 ) ;
  assign n12619 = ( n12435 & n12542 ) | ( n12435 & n12617 ) | ( n12542 & n12617 ) ;
  assign n12620 = ( n12542 & n12618 ) | ( n12542 & ~n12619 ) | ( n12618 & ~n12619 ) ;
  assign n12621 = ( n12438 & n12533 ) | ( n12438 & n12620 ) | ( n12533 & n12620 ) ;
  assign n12622 = ( n12438 & ~n12533 ) | ( n12438 & n12620 ) | ( ~n12533 & n12620 ) ;
  assign n12623 = ( n12533 & ~n12621 ) | ( n12533 & n12622 ) | ( ~n12621 & n12622 ) ;
  assign n12624 = ( n12441 & n12524 ) | ( n12441 & n12623 ) | ( n12524 & n12623 ) ;
  assign n12625 = ( n12441 & ~n12524 ) | ( n12441 & n12623 ) | ( ~n12524 & n12623 ) ;
  assign n12626 = ( n12524 & ~n12624 ) | ( n12524 & n12625 ) | ( ~n12624 & n12625 ) ;
  assign n12627 = n2766 & n5130 ;
  assign n12628 = x110 & n2770 ;
  assign n12629 = x111 | n12628 ;
  assign n12630 = ( n2772 & n12628 ) | ( n2772 & n12629 ) | ( n12628 & n12629 ) ;
  assign n12631 = x109 & n2943 ;
  assign n12632 = n12630 | n12631 ;
  assign n12633 = ( x35 & n12627 ) | ( x35 & ~n12632 ) | ( n12627 & ~n12632 ) ;
  assign n12634 = ( ~x35 & n12632 ) | ( ~x35 & n12633 ) | ( n12632 & n12633 ) ;
  assign n12635 = ( ~n12627 & n12633 ) | ( ~n12627 & n12634 ) | ( n12633 & n12634 ) ;
  assign n12636 = ( n12453 & n12626 ) | ( n12453 & n12635 ) | ( n12626 & n12635 ) ;
  assign n12637 = ( ~n12453 & n12626 ) | ( ~n12453 & n12635 ) | ( n12626 & n12635 ) ;
  assign n12638 = ( n12453 & ~n12636 ) | ( n12453 & n12637 ) | ( ~n12636 & n12637 ) ;
  assign n12639 = ( n12465 & n12515 ) | ( n12465 & n12638 ) | ( n12515 & n12638 ) ;
  assign n12640 = ( n12465 & ~n12515 ) | ( n12465 & n12638 ) | ( ~n12515 & n12638 ) ;
  assign n12641 = ( n12515 & ~n12639 ) | ( n12515 & n12640 ) | ( ~n12639 & n12640 ) ;
  assign n12642 = n1949 & n6201 ;
  assign n12643 = x116 & n1953 ;
  assign n12644 = x117 | n12643 ;
  assign n12645 = ( n1955 & n12643 ) | ( n1955 & n12644 ) | ( n12643 & n12644 ) ;
  assign n12646 = x115 & n2114 ;
  assign n12647 = n12645 | n12646 ;
  assign n12648 = ( x29 & n12642 ) | ( x29 & ~n12647 ) | ( n12642 & ~n12647 ) ;
  assign n12649 = ( ~x29 & n12647 ) | ( ~x29 & n12648 ) | ( n12647 & n12648 ) ;
  assign n12650 = ( ~n12642 & n12648 ) | ( ~n12642 & n12649 ) | ( n12648 & n12649 ) ;
  assign n12651 = ( n12468 & n12641 ) | ( n12468 & n12650 ) | ( n12641 & n12650 ) ;
  assign n12652 = ( n12468 & ~n12641 ) | ( n12468 & n12650 ) | ( ~n12641 & n12650 ) ;
  assign n12653 = ( n12641 & ~n12651 ) | ( n12641 & n12652 ) | ( ~n12651 & n12652 ) ;
  assign n12654 = ( n12471 & n12506 ) | ( n12471 & n12653 ) | ( n12506 & n12653 ) ;
  assign n12655 = ( n12471 & ~n12506 ) | ( n12471 & n12653 ) | ( ~n12506 & n12653 ) ;
  assign n12656 = ( n12506 & ~n12654 ) | ( n12506 & n12655 ) | ( ~n12654 & n12655 ) ;
  assign n12657 = n1297 & n7597 ;
  assign n12658 = x122 & n1301 ;
  assign n12659 = x123 | n12658 ;
  assign n12660 = ( n1303 & n12658 ) | ( n1303 & n12659 ) | ( n12658 & n12659 ) ;
  assign n12661 = x121 & n1426 ;
  assign n12662 = n12660 | n12661 ;
  assign n12663 = ( x23 & n12657 ) | ( x23 & ~n12662 ) | ( n12657 & ~n12662 ) ;
  assign n12664 = ( ~x23 & n12662 ) | ( ~x23 & n12663 ) | ( n12662 & n12663 ) ;
  assign n12665 = ( ~n12657 & n12663 ) | ( ~n12657 & n12664 ) | ( n12663 & n12664 ) ;
  assign n12666 = ( n12474 & n12656 ) | ( n12474 & n12665 ) | ( n12656 & n12665 ) ;
  assign n12667 = ( n12474 & ~n12656 ) | ( n12474 & n12665 ) | ( ~n12656 & n12665 ) ;
  assign n12668 = ( n12656 & ~n12666 ) | ( n12656 & n12667 ) | ( ~n12666 & n12667 ) ;
  assign n12669 = ( n12477 & n12497 ) | ( n12477 & n12668 ) | ( n12497 & n12668 ) ;
  assign n12670 = ( n12477 & ~n12497 ) | ( n12477 & n12668 ) | ( ~n12497 & n12668 ) ;
  assign n12671 = ( n12497 & ~n12669 ) | ( n12497 & n12670 ) | ( ~n12669 & n12670 ) ;
  assign n12672 = n810 & n8862 ;
  assign n12673 = ( x127 & n885 ) | ( x127 & n12672 ) | ( n885 & n12672 ) ;
  assign n12674 = x17 | n12673 ;
  assign n12675 = ~x17 & n12673 ;
  assign n12676 = ( ~n12673 & n12674 ) | ( ~n12673 & n12675 ) | ( n12674 & n12675 ) ;
  assign n12677 = ( n12480 & n12671 ) | ( n12480 & n12676 ) | ( n12671 & n12676 ) ;
  assign n12678 = ( n12480 & ~n12671 ) | ( n12480 & n12676 ) | ( ~n12671 & n12676 ) ;
  assign n12679 = ( n12671 & ~n12677 ) | ( n12671 & n12678 ) | ( ~n12677 & n12678 ) ;
  assign n12680 = ( n12483 & n12486 ) | ( n12483 & n12679 ) | ( n12486 & n12679 ) ;
  assign n12681 = ( n12483 & ~n12486 ) | ( n12483 & n12679 ) | ( ~n12486 & n12679 ) ;
  assign n12682 = ( n12486 & ~n12680 ) | ( n12486 & n12681 ) | ( ~n12680 & n12681 ) ;
  assign n12683 = n1297 & n7841 ;
  assign n12684 = x123 & n1301 ;
  assign n12685 = x124 | n12684 ;
  assign n12686 = ( n1303 & n12684 ) | ( n1303 & n12685 ) | ( n12684 & n12685 ) ;
  assign n12687 = x122 & n1426 ;
  assign n12688 = n12686 | n12687 ;
  assign n12689 = ( x23 & n12683 ) | ( x23 & ~n12688 ) | ( n12683 & ~n12688 ) ;
  assign n12690 = ( ~x23 & n12688 ) | ( ~x23 & n12689 ) | ( n12688 & n12689 ) ;
  assign n12691 = ( ~n12683 & n12689 ) | ( ~n12683 & n12690 ) | ( n12689 & n12690 ) ;
  assign n12692 = n1617 & n7113 ;
  assign n12693 = x120 & n1621 ;
  assign n12694 = x121 | n12693 ;
  assign n12695 = ( n1623 & n12693 ) | ( n1623 & n12694 ) | ( n12693 & n12694 ) ;
  assign n12696 = x119 & n1749 ;
  assign n12697 = n12695 | n12696 ;
  assign n12698 = ( x26 & n12692 ) | ( x26 & ~n12697 ) | ( n12692 & ~n12697 ) ;
  assign n12699 = ( ~x26 & n12697 ) | ( ~x26 & n12698 ) | ( n12697 & n12698 ) ;
  assign n12700 = ( ~n12692 & n12698 ) | ( ~n12692 & n12699 ) | ( n12698 & n12699 ) ;
  assign n12701 = n1949 & n6421 ;
  assign n12702 = x117 & n1953 ;
  assign n12703 = x118 | n12702 ;
  assign n12704 = ( n1955 & n12702 ) | ( n1955 & n12703 ) | ( n12702 & n12703 ) ;
  assign n12705 = x116 & n2114 ;
  assign n12706 = n12704 | n12705 ;
  assign n12707 = ( x29 & n12701 ) | ( x29 & ~n12706 ) | ( n12701 & ~n12706 ) ;
  assign n12708 = ( ~x29 & n12706 ) | ( ~x29 & n12707 ) | ( n12706 & n12707 ) ;
  assign n12709 = ( ~n12701 & n12707 ) | ( ~n12701 & n12708 ) | ( n12707 & n12708 ) ;
  assign n12710 = n3715 & n4013 ;
  assign n12711 = x105 & n3719 ;
  assign n12712 = x106 | n12711 ;
  assign n12713 = ( n3721 & n12711 ) | ( n3721 & n12712 ) | ( n12711 & n12712 ) ;
  assign n12714 = x104 & n3922 ;
  assign n12715 = n12713 | n12714 ;
  assign n12716 = ( x41 & n12710 ) | ( x41 & ~n12715 ) | ( n12710 & ~n12715 ) ;
  assign n12717 = ( ~x41 & n12715 ) | ( ~x41 & n12716 ) | ( n12715 & n12716 ) ;
  assign n12718 = ( ~n12710 & n12716 ) | ( ~n12710 & n12717 ) | ( n12716 & n12717 ) ;
  assign n12719 = n3162 & n4787 ;
  assign n12720 = x99 & n4791 ;
  assign n12721 = x100 | n12720 ;
  assign n12722 = ( n4793 & n12720 ) | ( n4793 & n12721 ) | ( n12720 & n12721 ) ;
  assign n12723 = x98 & n5030 ;
  assign n12724 = n12722 | n12723 ;
  assign n12725 = ( x47 & n12719 ) | ( x47 & ~n12724 ) | ( n12719 & ~n12724 ) ;
  assign n12726 = ( ~x47 & n12724 ) | ( ~x47 & n12725 ) | ( n12724 & n12725 ) ;
  assign n12727 = ( ~n12719 & n12725 ) | ( ~n12719 & n12726 ) | ( n12725 & n12726 ) ;
  assign n12728 = n2294 & n6027 ;
  assign n12729 = x93 & n6031 ;
  assign n12730 = x94 | n12729 ;
  assign n12731 = ( n6033 & n12729 ) | ( n6033 & n12730 ) | ( n12729 & n12730 ) ;
  assign n12732 = x92 & n6303 ;
  assign n12733 = n12731 | n12732 ;
  assign n12734 = ( x53 & n12728 ) | ( x53 & ~n12733 ) | ( n12728 & ~n12733 ) ;
  assign n12735 = ( ~x53 & n12733 ) | ( ~x53 & n12734 ) | ( n12733 & n12734 ) ;
  assign n12736 = ( ~n12728 & n12734 ) | ( ~n12728 & n12735 ) | ( n12734 & n12735 ) ;
  assign n12737 = n1914 & n6713 ;
  assign n12738 = x90 & n6717 ;
  assign n12739 = x91 | n12738 ;
  assign n12740 = ( n6719 & n12738 ) | ( n6719 & n12739 ) | ( n12738 & n12739 ) ;
  assign n12741 = x89 & n6980 ;
  assign n12742 = n12740 | n12741 ;
  assign n12743 = ( x56 & n12737 ) | ( x56 & ~n12742 ) | ( n12737 & ~n12742 ) ;
  assign n12744 = ( ~x56 & n12742 ) | ( ~x56 & n12743 ) | ( n12742 & n12743 ) ;
  assign n12745 = ( ~n12737 & n12743 ) | ( ~n12737 & n12744 ) | ( n12743 & n12744 ) ;
  assign n12746 = n1481 & n7423 ;
  assign n12747 = x87 & n7427 ;
  assign n12748 = x88 | n12747 ;
  assign n12749 = ( n7429 & n12747 ) | ( n7429 & n12748 ) | ( n12747 & n12748 ) ;
  assign n12750 = x86 & n7708 ;
  assign n12751 = n12749 | n12750 ;
  assign n12752 = ( x59 & n12746 ) | ( x59 & ~n12751 ) | ( n12746 & ~n12751 ) ;
  assign n12753 = ( ~x59 & n12751 ) | ( ~x59 & n12752 ) | ( n12751 & n12752 ) ;
  assign n12754 = ( ~n12746 & n12752 ) | ( ~n12746 & n12753 ) | ( n12752 & n12753 ) ;
  assign n12755 = n1262 & n8154 ;
  assign n12756 = x84 & n8158 ;
  assign n12757 = x85 | n12756 ;
  assign n12758 = ( n8160 & n12756 ) | ( n8160 & n12757 ) | ( n12756 & n12757 ) ;
  assign n12759 = x83 & n8439 ;
  assign n12760 = n12758 | n12759 ;
  assign n12761 = ( x62 & n12755 ) | ( x62 & ~n12760 ) | ( n12755 & ~n12760 ) ;
  assign n12762 = ( ~x62 & n12760 ) | ( ~x62 & n12761 ) | ( n12760 & n12761 ) ;
  assign n12763 = ( ~n12755 & n12761 ) | ( ~n12755 & n12762 ) | ( n12761 & n12762 ) ;
  assign n12764 = x81 & n8927 ;
  assign n12765 = ( ~x82 & n8693 ) | ( ~x82 & n8927 ) | ( n8693 & n8927 ) ;
  assign n12766 = ( n8693 & n12764 ) | ( n8693 & ~n12765 ) | ( n12764 & ~n12765 ) ;
  assign n12767 = ( ~x17 & n12590 ) | ( ~x17 & n12766 ) | ( n12590 & n12766 ) ;
  assign n12768 = ( n12590 & n12766 ) | ( n12590 & ~n12767 ) | ( n12766 & ~n12767 ) ;
  assign n12769 = ( x17 & n12767 ) | ( x17 & ~n12768 ) | ( n12767 & ~n12768 ) ;
  assign n12770 = ( n12591 & n12763 ) | ( n12591 & ~n12769 ) | ( n12763 & ~n12769 ) ;
  assign n12771 = ( ~n12591 & n12763 ) | ( ~n12591 & n12769 ) | ( n12763 & n12769 ) ;
  assign n12772 = ( ~n12763 & n12770 ) | ( ~n12763 & n12771 ) | ( n12770 & n12771 ) ;
  assign n12773 = ( n12594 & n12754 ) | ( n12594 & ~n12772 ) | ( n12754 & ~n12772 ) ;
  assign n12774 = ( ~n12594 & n12754 ) | ( ~n12594 & n12772 ) | ( n12754 & n12772 ) ;
  assign n12775 = ( ~n12754 & n12773 ) | ( ~n12754 & n12774 ) | ( n12773 & n12774 ) ;
  assign n12776 = ( n12597 & n12745 ) | ( n12597 & ~n12775 ) | ( n12745 & ~n12775 ) ;
  assign n12777 = ( ~n12597 & n12745 ) | ( ~n12597 & n12775 ) | ( n12745 & n12775 ) ;
  assign n12778 = ( ~n12745 & n12776 ) | ( ~n12745 & n12777 ) | ( n12776 & n12777 ) ;
  assign n12779 = ( n12600 & n12736 ) | ( n12600 & ~n12778 ) | ( n12736 & ~n12778 ) ;
  assign n12780 = ( ~n12600 & n12736 ) | ( ~n12600 & n12778 ) | ( n12736 & n12778 ) ;
  assign n12781 = ( ~n12736 & n12779 ) | ( ~n12736 & n12780 ) | ( n12779 & n12780 ) ;
  assign n12782 = n2585 & n5374 ;
  assign n12783 = x96 & n5378 ;
  assign n12784 = x97 | n12783 ;
  assign n12785 = ( n5380 & n12783 ) | ( n5380 & n12784 ) | ( n12783 & n12784 ) ;
  assign n12786 = x95 & n5638 ;
  assign n12787 = n12785 | n12786 ;
  assign n12788 = ( x50 & n12782 ) | ( x50 & ~n12787 ) | ( n12782 & ~n12787 ) ;
  assign n12789 = ( ~x50 & n12787 ) | ( ~x50 & n12788 ) | ( n12787 & n12788 ) ;
  assign n12790 = ( ~n12782 & n12788 ) | ( ~n12782 & n12789 ) | ( n12788 & n12789 ) ;
  assign n12791 = ( n12603 & ~n12781 ) | ( n12603 & n12790 ) | ( ~n12781 & n12790 ) ;
  assign n12792 = ( n12603 & n12781 ) | ( n12603 & n12790 ) | ( n12781 & n12790 ) ;
  assign n12793 = ( n12781 & n12791 ) | ( n12781 & ~n12792 ) | ( n12791 & ~n12792 ) ;
  assign n12794 = ( n12615 & n12727 ) | ( n12615 & ~n12793 ) | ( n12727 & ~n12793 ) ;
  assign n12795 = ( ~n12615 & n12727 ) | ( ~n12615 & n12793 ) | ( n12727 & n12793 ) ;
  assign n12796 = ( ~n12727 & n12794 ) | ( ~n12727 & n12795 ) | ( n12794 & n12795 ) ;
  assign n12797 = n3650 & n4227 ;
  assign n12798 = x102 & n4231 ;
  assign n12799 = x103 | n12798 ;
  assign n12800 = ( n4233 & n12798 ) | ( n4233 & n12799 ) | ( n12798 & n12799 ) ;
  assign n12801 = x101 & n4470 ;
  assign n12802 = n12800 | n12801 ;
  assign n12803 = ( x44 & n12797 ) | ( x44 & ~n12802 ) | ( n12797 & ~n12802 ) ;
  assign n12804 = ( ~x44 & n12802 ) | ( ~x44 & n12803 ) | ( n12802 & n12803 ) ;
  assign n12805 = ( ~n12797 & n12803 ) | ( ~n12797 & n12804 ) | ( n12803 & n12804 ) ;
  assign n12806 = ( n12618 & n12796 ) | ( n12618 & ~n12805 ) | ( n12796 & ~n12805 ) ;
  assign n12807 = ( ~n12618 & n12796 ) | ( ~n12618 & n12805 ) | ( n12796 & n12805 ) ;
  assign n12808 = ( ~n12796 & n12806 ) | ( ~n12796 & n12807 ) | ( n12806 & n12807 ) ;
  assign n12809 = ( n12621 & n12718 ) | ( n12621 & n12808 ) | ( n12718 & n12808 ) ;
  assign n12810 = ( ~n12621 & n12718 ) | ( ~n12621 & n12808 ) | ( n12718 & n12808 ) ;
  assign n12811 = ( n12621 & ~n12809 ) | ( n12621 & n12810 ) | ( ~n12809 & n12810 ) ;
  assign n12812 = n3224 & n4734 ;
  assign n12813 = x108 & n3228 ;
  assign n12814 = x109 | n12813 ;
  assign n12815 = ( n3230 & n12813 ) | ( n3230 & n12814 ) | ( n12813 & n12814 ) ;
  assign n12816 = x107 & n3413 ;
  assign n12817 = n12815 | n12816 ;
  assign n12818 = ( x38 & n12812 ) | ( x38 & ~n12817 ) | ( n12812 & ~n12817 ) ;
  assign n12819 = ( ~x38 & n12817 ) | ( ~x38 & n12818 ) | ( n12817 & n12818 ) ;
  assign n12820 = ( ~n12812 & n12818 ) | ( ~n12812 & n12819 ) | ( n12818 & n12819 ) ;
  assign n12821 = ( n12624 & n12811 ) | ( n12624 & n12820 ) | ( n12811 & n12820 ) ;
  assign n12822 = ( ~n12624 & n12811 ) | ( ~n12624 & n12820 ) | ( n12811 & n12820 ) ;
  assign n12823 = ( n12624 & ~n12821 ) | ( n12624 & n12822 ) | ( ~n12821 & n12822 ) ;
  assign n12824 = n2766 & n5145 ;
  assign n12825 = x111 & n2770 ;
  assign n12826 = x112 | n12825 ;
  assign n12827 = ( n2772 & n12825 ) | ( n2772 & n12826 ) | ( n12825 & n12826 ) ;
  assign n12828 = x110 & n2943 ;
  assign n12829 = n12827 | n12828 ;
  assign n12830 = ( x35 & n12824 ) | ( x35 & ~n12829 ) | ( n12824 & ~n12829 ) ;
  assign n12831 = ( ~x35 & n12829 ) | ( ~x35 & n12830 ) | ( n12829 & n12830 ) ;
  assign n12832 = ( ~n12824 & n12830 ) | ( ~n12824 & n12831 ) | ( n12830 & n12831 ) ;
  assign n12833 = ( n12636 & n12823 ) | ( n12636 & n12832 ) | ( n12823 & n12832 ) ;
  assign n12834 = ( ~n12636 & n12823 ) | ( ~n12636 & n12832 ) | ( n12823 & n12832 ) ;
  assign n12835 = ( n12636 & ~n12833 ) | ( n12636 & n12834 ) | ( ~n12833 & n12834 ) ;
  assign n12836 = n2320 & n5765 ;
  assign n12837 = x114 & n2324 ;
  assign n12838 = x115 | n12837 ;
  assign n12839 = ( n2326 & n12837 ) | ( n2326 & n12838 ) | ( n12837 & n12838 ) ;
  assign n12840 = x113 & n2497 ;
  assign n12841 = n12839 | n12840 ;
  assign n12842 = ( x32 & n12836 ) | ( x32 & ~n12841 ) | ( n12836 & ~n12841 ) ;
  assign n12843 = ( ~x32 & n12841 ) | ( ~x32 & n12842 ) | ( n12841 & n12842 ) ;
  assign n12844 = ( ~n12836 & n12842 ) | ( ~n12836 & n12843 ) | ( n12842 & n12843 ) ;
  assign n12845 = ( n12639 & n12835 ) | ( n12639 & n12844 ) | ( n12835 & n12844 ) ;
  assign n12846 = ( n12639 & ~n12835 ) | ( n12639 & n12844 ) | ( ~n12835 & n12844 ) ;
  assign n12847 = ( n12835 & ~n12845 ) | ( n12835 & n12846 ) | ( ~n12845 & n12846 ) ;
  assign n12848 = ( n12651 & n12709 ) | ( n12651 & n12847 ) | ( n12709 & n12847 ) ;
  assign n12849 = ( n12651 & ~n12709 ) | ( n12651 & n12847 ) | ( ~n12709 & n12847 ) ;
  assign n12850 = ( n12709 & ~n12848 ) | ( n12709 & n12849 ) | ( ~n12848 & n12849 ) ;
  assign n12851 = ( n12654 & n12700 ) | ( n12654 & n12850 ) | ( n12700 & n12850 ) ;
  assign n12852 = ( n12654 & ~n12700 ) | ( n12654 & n12850 ) | ( ~n12700 & n12850 ) ;
  assign n12853 = ( n12700 & ~n12851 ) | ( n12700 & n12852 ) | ( ~n12851 & n12852 ) ;
  assign n12854 = ( n12666 & n12691 ) | ( n12666 & n12853 ) | ( n12691 & n12853 ) ;
  assign n12855 = ( n12666 & ~n12691 ) | ( n12666 & n12853 ) | ( ~n12691 & n12853 ) ;
  assign n12856 = ( n12691 & ~n12854 ) | ( n12691 & n12855 ) | ( ~n12854 & n12855 ) ;
  assign n12857 = n1016 & n8846 ;
  assign n12858 = x126 & n1020 ;
  assign n12859 = x127 | n12858 ;
  assign n12860 = ( n1022 & n12858 ) | ( n1022 & n12859 ) | ( n12858 & n12859 ) ;
  assign n12861 = x125 & n1145 ;
  assign n12862 = n12860 | n12861 ;
  assign n12863 = ( x20 & n12857 ) | ( x20 & ~n12862 ) | ( n12857 & ~n12862 ) ;
  assign n12864 = ( ~x20 & n12862 ) | ( ~x20 & n12863 ) | ( n12862 & n12863 ) ;
  assign n12865 = ( ~n12857 & n12863 ) | ( ~n12857 & n12864 ) | ( n12863 & n12864 ) ;
  assign n12866 = ( n12669 & n12856 ) | ( n12669 & n12865 ) | ( n12856 & n12865 ) ;
  assign n12867 = ( n12669 & ~n12856 ) | ( n12669 & n12865 ) | ( ~n12856 & n12865 ) ;
  assign n12868 = ( n12856 & ~n12866 ) | ( n12856 & n12867 ) | ( ~n12866 & n12867 ) ;
  assign n12869 = ( n12677 & n12680 ) | ( n12677 & n12868 ) | ( n12680 & n12868 ) ;
  assign n12870 = ( n12677 & ~n12680 ) | ( n12677 & n12868 ) | ( ~n12680 & n12868 ) ;
  assign n12871 = ( n12680 & ~n12869 ) | ( n12680 & n12870 ) | ( ~n12869 & n12870 ) ;
  assign n12872 = n1016 & n8865 ;
  assign n12873 = x127 & n1020 ;
  assign n12874 = x126 | n12873 ;
  assign n12875 = ( n1145 & n12873 ) | ( n1145 & n12874 ) | ( n12873 & n12874 ) ;
  assign n12876 = ( x20 & n12872 ) | ( x20 & ~n12875 ) | ( n12872 & ~n12875 ) ;
  assign n12877 = ( ~x20 & n12875 ) | ( ~x20 & n12876 ) | ( n12875 & n12876 ) ;
  assign n12878 = ( ~n12872 & n12876 ) | ( ~n12872 & n12877 ) | ( n12876 & n12877 ) ;
  assign n12879 = n1297 & n8331 ;
  assign n12880 = x124 & n1301 ;
  assign n12881 = x125 | n12880 ;
  assign n12882 = ( n1303 & n12880 ) | ( n1303 & n12881 ) | ( n12880 & n12881 ) ;
  assign n12883 = x123 & n1426 ;
  assign n12884 = n12882 | n12883 ;
  assign n12885 = ( x23 & n12879 ) | ( x23 & ~n12884 ) | ( n12879 & ~n12884 ) ;
  assign n12886 = ( ~x23 & n12884 ) | ( ~x23 & n12885 ) | ( n12884 & n12885 ) ;
  assign n12887 = ( ~n12879 & n12885 ) | ( ~n12879 & n12886 ) | ( n12885 & n12886 ) ;
  assign n12888 = n1617 & n7582 ;
  assign n12889 = x121 & n1621 ;
  assign n12890 = x122 | n12889 ;
  assign n12891 = ( n1623 & n12889 ) | ( n1623 & n12890 ) | ( n12889 & n12890 ) ;
  assign n12892 = x120 & n1749 ;
  assign n12893 = n12891 | n12892 ;
  assign n12894 = ( x26 & n12888 ) | ( x26 & ~n12893 ) | ( n12888 & ~n12893 ) ;
  assign n12895 = ( ~x26 & n12893 ) | ( ~x26 & n12894 ) | ( n12893 & n12894 ) ;
  assign n12896 = ( ~n12888 & n12894 ) | ( ~n12888 & n12895 ) | ( n12894 & n12895 ) ;
  assign n12897 = n1949 & n6645 ;
  assign n12898 = x118 & n1953 ;
  assign n12899 = x119 | n12898 ;
  assign n12900 = ( n1955 & n12898 ) | ( n1955 & n12899 ) | ( n12898 & n12899 ) ;
  assign n12901 = x117 & n2114 ;
  assign n12902 = n12900 | n12901 ;
  assign n12903 = ( x29 & n12897 ) | ( x29 & ~n12902 ) | ( n12897 & ~n12902 ) ;
  assign n12904 = ( ~x29 & n12902 ) | ( ~x29 & n12903 ) | ( n12902 & n12903 ) ;
  assign n12905 = ( ~n12897 & n12903 ) | ( ~n12897 & n12904 ) | ( n12903 & n12904 ) ;
  assign n12906 = n2320 & n5977 ;
  assign n12907 = x115 & n2324 ;
  assign n12908 = x116 | n12907 ;
  assign n12909 = ( n2326 & n12907 ) | ( n2326 & n12908 ) | ( n12907 & n12908 ) ;
  assign n12910 = x114 & n2497 ;
  assign n12911 = n12909 | n12910 ;
  assign n12912 = ( x32 & n12906 ) | ( x32 & ~n12911 ) | ( n12906 & ~n12911 ) ;
  assign n12913 = ( ~x32 & n12911 ) | ( ~x32 & n12912 ) | ( n12911 & n12912 ) ;
  assign n12914 = ( ~n12906 & n12912 ) | ( ~n12906 & n12913 ) | ( n12912 & n12913 ) ;
  assign n12915 = n3665 & n4227 ;
  assign n12916 = x103 & n4231 ;
  assign n12917 = x104 | n12916 ;
  assign n12918 = ( n4233 & n12916 ) | ( n4233 & n12917 ) | ( n12916 & n12917 ) ;
  assign n12919 = x102 & n4470 ;
  assign n12920 = n12918 | n12919 ;
  assign n12921 = ( x44 & n12915 ) | ( x44 & ~n12920 ) | ( n12915 & ~n12920 ) ;
  assign n12922 = ( ~x44 & n12920 ) | ( ~x44 & n12921 ) | ( n12920 & n12921 ) ;
  assign n12923 = ( ~n12915 & n12921 ) | ( ~n12915 & n12922 ) | ( n12921 & n12922 ) ;
  assign n12924 = n3326 & n4787 ;
  assign n12925 = x100 & n4791 ;
  assign n12926 = x101 | n12925 ;
  assign n12927 = ( n4793 & n12925 ) | ( n4793 & n12926 ) | ( n12925 & n12926 ) ;
  assign n12928 = x99 & n5030 ;
  assign n12929 = n12927 | n12928 ;
  assign n12930 = ( x47 & n12924 ) | ( x47 & ~n12929 ) | ( n12924 & ~n12929 ) ;
  assign n12931 = ( ~x47 & n12929 ) | ( ~x47 & n12930 ) | ( n12929 & n12930 ) ;
  assign n12932 = ( ~n12924 & n12930 ) | ( ~n12924 & n12931 ) | ( n12930 & n12931 ) ;
  assign n12933 = n2725 & n5374 ;
  assign n12934 = x97 & n5378 ;
  assign n12935 = x98 | n12934 ;
  assign n12936 = ( n5380 & n12934 ) | ( n5380 & n12935 ) | ( n12934 & n12935 ) ;
  assign n12937 = x96 & n5638 ;
  assign n12938 = n12936 | n12937 ;
  assign n12939 = ( x50 & n12933 ) | ( x50 & ~n12938 ) | ( n12933 & ~n12938 ) ;
  assign n12940 = ( ~x50 & n12938 ) | ( ~x50 & n12939 ) | ( n12938 & n12939 ) ;
  assign n12941 = ( ~n12933 & n12939 ) | ( ~n12933 & n12940 ) | ( n12939 & n12940 ) ;
  assign n12942 = n2042 & n6713 ;
  assign n12943 = x91 & n6717 ;
  assign n12944 = x92 | n12943 ;
  assign n12945 = ( n6719 & n12943 ) | ( n6719 & n12944 ) | ( n12943 & n12944 ) ;
  assign n12946 = x90 & n6980 ;
  assign n12947 = n12945 | n12946 ;
  assign n12948 = ( x56 & n12942 ) | ( x56 & ~n12947 ) | ( n12942 & ~n12947 ) ;
  assign n12949 = ( ~x56 & n12947 ) | ( ~x56 & n12948 ) | ( n12947 & n12948 ) ;
  assign n12950 = ( ~n12942 & n12948 ) | ( ~n12942 & n12949 ) | ( n12948 & n12949 ) ;
  assign n12951 = x82 & n8927 ;
  assign n12952 = ( ~x83 & n8693 ) | ( ~x83 & n8927 ) | ( n8693 & n8927 ) ;
  assign n12953 = ( n8693 & n12951 ) | ( n8693 & ~n12952 ) | ( n12951 & ~n12952 ) ;
  assign n12954 = n1366 & n8154 ;
  assign n12955 = x85 & n8158 ;
  assign n12956 = x86 | n12955 ;
  assign n12957 = ( n8160 & n12955 ) | ( n8160 & n12956 ) | ( n12955 & n12956 ) ;
  assign n12958 = x84 & n8439 ;
  assign n12959 = n12957 | n12958 ;
  assign n12960 = ( x62 & n12954 ) | ( x62 & ~n12959 ) | ( n12954 & ~n12959 ) ;
  assign n12961 = ( ~x62 & n12959 ) | ( ~x62 & n12960 ) | ( n12959 & n12960 ) ;
  assign n12962 = ( ~n12954 & n12960 ) | ( ~n12954 & n12961 ) | ( n12960 & n12961 ) ;
  assign n12963 = ( n12767 & ~n12953 ) | ( n12767 & n12962 ) | ( ~n12953 & n12962 ) ;
  assign n12964 = ( n12767 & n12953 ) | ( n12767 & n12962 ) | ( n12953 & n12962 ) ;
  assign n12965 = ( n12953 & n12963 ) | ( n12953 & ~n12964 ) | ( n12963 & ~n12964 ) ;
  assign n12966 = n1585 & n7423 ;
  assign n12967 = x88 & n7427 ;
  assign n12968 = x89 | n12967 ;
  assign n12969 = ( n7429 & n12967 ) | ( n7429 & n12968 ) | ( n12967 & n12968 ) ;
  assign n12970 = x87 & n7708 ;
  assign n12971 = n12969 | n12970 ;
  assign n12972 = ( x59 & n12966 ) | ( x59 & ~n12971 ) | ( n12966 & ~n12971 ) ;
  assign n12973 = ( ~x59 & n12971 ) | ( ~x59 & n12972 ) | ( n12971 & n12972 ) ;
  assign n12974 = ( ~n12966 & n12972 ) | ( ~n12966 & n12973 ) | ( n12972 & n12973 ) ;
  assign n12975 = ( n12770 & ~n12965 ) | ( n12770 & n12974 ) | ( ~n12965 & n12974 ) ;
  assign n12976 = ( n12770 & n12965 ) | ( n12770 & n12974 ) | ( n12965 & n12974 ) ;
  assign n12977 = ( n12965 & n12975 ) | ( n12965 & ~n12976 ) | ( n12975 & ~n12976 ) ;
  assign n12978 = ( n12773 & n12950 ) | ( n12773 & ~n12977 ) | ( n12950 & ~n12977 ) ;
  assign n12979 = ( ~n12773 & n12950 ) | ( ~n12773 & n12977 ) | ( n12950 & n12977 ) ;
  assign n12980 = ( ~n12950 & n12978 ) | ( ~n12950 & n12979 ) | ( n12978 & n12979 ) ;
  assign n12981 = n2434 & n6027 ;
  assign n12982 = x94 & n6031 ;
  assign n12983 = x95 | n12982 ;
  assign n12984 = ( n6033 & n12982 ) | ( n6033 & n12983 ) | ( n12982 & n12983 ) ;
  assign n12985 = x93 & n6303 ;
  assign n12986 = n12984 | n12985 ;
  assign n12987 = ( x53 & n12981 ) | ( x53 & ~n12986 ) | ( n12981 & ~n12986 ) ;
  assign n12988 = ( ~x53 & n12986 ) | ( ~x53 & n12987 ) | ( n12986 & n12987 ) ;
  assign n12989 = ( ~n12981 & n12987 ) | ( ~n12981 & n12988 ) | ( n12987 & n12988 ) ;
  assign n12990 = ( n12776 & ~n12980 ) | ( n12776 & n12989 ) | ( ~n12980 & n12989 ) ;
  assign n12991 = ( n12776 & n12980 ) | ( n12776 & n12989 ) | ( n12980 & n12989 ) ;
  assign n12992 = ( n12980 & n12990 ) | ( n12980 & ~n12991 ) | ( n12990 & ~n12991 ) ;
  assign n12993 = ( n12779 & n12941 ) | ( n12779 & ~n12992 ) | ( n12941 & ~n12992 ) ;
  assign n12994 = ( ~n12779 & n12941 ) | ( ~n12779 & n12992 ) | ( n12941 & n12992 ) ;
  assign n12995 = ( ~n12941 & n12993 ) | ( ~n12941 & n12994 ) | ( n12993 & n12994 ) ;
  assign n12996 = ( n12791 & n12932 ) | ( n12791 & ~n12995 ) | ( n12932 & ~n12995 ) ;
  assign n12997 = ( ~n12791 & n12932 ) | ( ~n12791 & n12995 ) | ( n12932 & n12995 ) ;
  assign n12998 = ( ~n12932 & n12996 ) | ( ~n12932 & n12997 ) | ( n12996 & n12997 ) ;
  assign n12999 = ( n12794 & n12923 ) | ( n12794 & ~n12998 ) | ( n12923 & ~n12998 ) ;
  assign n13000 = ( ~n12794 & n12923 ) | ( ~n12794 & n12998 ) | ( n12923 & n12998 ) ;
  assign n13001 = ( ~n12923 & n12999 ) | ( ~n12923 & n13000 ) | ( n12999 & n13000 ) ;
  assign n13002 = n3715 & n4362 ;
  assign n13003 = x106 & n3719 ;
  assign n13004 = x107 | n13003 ;
  assign n13005 = ( n3721 & n13003 ) | ( n3721 & n13004 ) | ( n13003 & n13004 ) ;
  assign n13006 = x105 & n3922 ;
  assign n13007 = n13005 | n13006 ;
  assign n13008 = ( x41 & n13002 ) | ( x41 & ~n13007 ) | ( n13002 & ~n13007 ) ;
  assign n13009 = ( ~x41 & n13007 ) | ( ~x41 & n13008 ) | ( n13007 & n13008 ) ;
  assign n13010 = ( ~n13002 & n13008 ) | ( ~n13002 & n13009 ) | ( n13008 & n13009 ) ;
  assign n13011 = ( n12806 & n13001 ) | ( n12806 & ~n13010 ) | ( n13001 & ~n13010 ) ;
  assign n13012 = ( ~n12806 & n13001 ) | ( ~n12806 & n13010 ) | ( n13001 & n13010 ) ;
  assign n13013 = ( ~n13001 & n13011 ) | ( ~n13001 & n13012 ) | ( n13011 & n13012 ) ;
  assign n13014 = n3224 & n4934 ;
  assign n13015 = x109 & n3228 ;
  assign n13016 = x110 | n13015 ;
  assign n13017 = ( n3230 & n13015 ) | ( n3230 & n13016 ) | ( n13015 & n13016 ) ;
  assign n13018 = x108 & n3413 ;
  assign n13019 = n13017 | n13018 ;
  assign n13020 = ( x38 & n13014 ) | ( x38 & ~n13019 ) | ( n13014 & ~n13019 ) ;
  assign n13021 = ( ~x38 & n13019 ) | ( ~x38 & n13020 ) | ( n13019 & n13020 ) ;
  assign n13022 = ( ~n13014 & n13020 ) | ( ~n13014 & n13021 ) | ( n13020 & n13021 ) ;
  assign n13023 = ( n12809 & n13013 ) | ( n12809 & n13022 ) | ( n13013 & n13022 ) ;
  assign n13024 = ( ~n12809 & n13013 ) | ( ~n12809 & n13022 ) | ( n13013 & n13022 ) ;
  assign n13025 = ( n12809 & ~n13023 ) | ( n12809 & n13024 ) | ( ~n13023 & n13024 ) ;
  assign n13026 = n2766 & n5542 ;
  assign n13027 = x112 & n2770 ;
  assign n13028 = x113 | n13027 ;
  assign n13029 = ( n2772 & n13027 ) | ( n2772 & n13028 ) | ( n13027 & n13028 ) ;
  assign n13030 = x111 & n2943 ;
  assign n13031 = n13029 | n13030 ;
  assign n13032 = ( x35 & n13026 ) | ( x35 & ~n13031 ) | ( n13026 & ~n13031 ) ;
  assign n13033 = ( ~x35 & n13031 ) | ( ~x35 & n13032 ) | ( n13031 & n13032 ) ;
  assign n13034 = ( ~n13026 & n13032 ) | ( ~n13026 & n13033 ) | ( n13032 & n13033 ) ;
  assign n13035 = ( n12821 & n13025 ) | ( n12821 & n13034 ) | ( n13025 & n13034 ) ;
  assign n13036 = ( ~n12821 & n13025 ) | ( ~n12821 & n13034 ) | ( n13025 & n13034 ) ;
  assign n13037 = ( n12821 & ~n13035 ) | ( n12821 & n13036 ) | ( ~n13035 & n13036 ) ;
  assign n13038 = ( n12833 & n12914 ) | ( n12833 & n13037 ) | ( n12914 & n13037 ) ;
  assign n13039 = ( n12833 & ~n12914 ) | ( n12833 & n13037 ) | ( ~n12914 & n13037 ) ;
  assign n13040 = ( n12914 & ~n13038 ) | ( n12914 & n13039 ) | ( ~n13038 & n13039 ) ;
  assign n13041 = ( n12845 & n12905 ) | ( n12845 & n13040 ) | ( n12905 & n13040 ) ;
  assign n13042 = ( n12845 & ~n12905 ) | ( n12845 & n13040 ) | ( ~n12905 & n13040 ) ;
  assign n13043 = ( n12905 & ~n13041 ) | ( n12905 & n13042 ) | ( ~n13041 & n13042 ) ;
  assign n13044 = ( n12848 & n12896 ) | ( n12848 & n13043 ) | ( n12896 & n13043 ) ;
  assign n13045 = ( n12848 & ~n12896 ) | ( n12848 & n13043 ) | ( ~n12896 & n13043 ) ;
  assign n13046 = ( n12896 & ~n13044 ) | ( n12896 & n13045 ) | ( ~n13044 & n13045 ) ;
  assign n13047 = ( n12851 & n12887 ) | ( n12851 & n13046 ) | ( n12887 & n13046 ) ;
  assign n13048 = ( n12851 & ~n12887 ) | ( n12851 & n13046 ) | ( ~n12887 & n13046 ) ;
  assign n13049 = ( n12887 & ~n13047 ) | ( n12887 & n13048 ) | ( ~n13047 & n13048 ) ;
  assign n13050 = ( n12854 & n12878 ) | ( n12854 & n13049 ) | ( n12878 & n13049 ) ;
  assign n13051 = ( ~n12854 & n12878 ) | ( ~n12854 & n13049 ) | ( n12878 & n13049 ) ;
  assign n13052 = ( n12854 & ~n13050 ) | ( n12854 & n13051 ) | ( ~n13050 & n13051 ) ;
  assign n13053 = ( n12866 & n12869 ) | ( n12866 & n13052 ) | ( n12869 & n13052 ) ;
  assign n13054 = ( n12866 & ~n12869 ) | ( n12866 & n13052 ) | ( ~n12869 & n13052 ) ;
  assign n13055 = ( n12869 & ~n13053 ) | ( n12869 & n13054 ) | ( ~n13053 & n13054 ) ;
  assign n13056 = n1016 & n8862 ;
  assign n13057 = ( x127 & n1145 ) | ( x127 & n13056 ) | ( n1145 & n13056 ) ;
  assign n13058 = x20 | n13057 ;
  assign n13059 = ~x20 & n13057 ;
  assign n13060 = ( ~n13057 & n13058 ) | ( ~n13057 & n13059 ) | ( n13058 & n13059 ) ;
  assign n13061 = n1297 & n8587 ;
  assign n13062 = x125 & n1301 ;
  assign n13063 = x126 | n13062 ;
  assign n13064 = ( n1303 & n13062 ) | ( n1303 & n13063 ) | ( n13062 & n13063 ) ;
  assign n13065 = x124 & n1426 ;
  assign n13066 = n13064 | n13065 ;
  assign n13067 = ( x23 & n13061 ) | ( x23 & ~n13066 ) | ( n13061 & ~n13066 ) ;
  assign n13068 = ( ~x23 & n13066 ) | ( ~x23 & n13067 ) | ( n13066 & n13067 ) ;
  assign n13069 = ( ~n13061 & n13067 ) | ( ~n13061 & n13068 ) | ( n13067 & n13068 ) ;
  assign n13070 = n1617 & n7597 ;
  assign n13071 = x122 & n1621 ;
  assign n13072 = x123 | n13071 ;
  assign n13073 = ( n1623 & n13071 ) | ( n1623 & n13072 ) | ( n13071 & n13072 ) ;
  assign n13074 = x121 & n1749 ;
  assign n13075 = n13073 | n13074 ;
  assign n13076 = ( x26 & n13070 ) | ( x26 & ~n13075 ) | ( n13070 & ~n13075 ) ;
  assign n13077 = ( ~x26 & n13075 ) | ( ~x26 & n13076 ) | ( n13075 & n13076 ) ;
  assign n13078 = ( ~n13070 & n13076 ) | ( ~n13070 & n13077 ) | ( n13076 & n13077 ) ;
  assign n13079 = n2320 & n6201 ;
  assign n13080 = x116 & n2324 ;
  assign n13081 = x117 | n13080 ;
  assign n13082 = ( n2326 & n13080 ) | ( n2326 & n13081 ) | ( n13080 & n13081 ) ;
  assign n13083 = x115 & n2497 ;
  assign n13084 = n13082 | n13083 ;
  assign n13085 = ( x32 & n13079 ) | ( x32 & ~n13084 ) | ( n13079 & ~n13084 ) ;
  assign n13086 = ( ~x32 & n13084 ) | ( ~x32 & n13085 ) | ( n13084 & n13085 ) ;
  assign n13087 = ( ~n13079 & n13085 ) | ( ~n13079 & n13086 ) | ( n13085 & n13086 ) ;
  assign n13088 = n3715 & n4377 ;
  assign n13089 = x107 & n3719 ;
  assign n13090 = x108 | n13089 ;
  assign n13091 = ( n3721 & n13089 ) | ( n3721 & n13090 ) | ( n13089 & n13090 ) ;
  assign n13092 = x106 & n3922 ;
  assign n13093 = n13091 | n13092 ;
  assign n13094 = ( x41 & n13088 ) | ( x41 & ~n13093 ) | ( n13088 & ~n13093 ) ;
  assign n13095 = ( ~x41 & n13093 ) | ( ~x41 & n13094 ) | ( n13093 & n13094 ) ;
  assign n13096 = ( ~n13088 & n13094 ) | ( ~n13088 & n13095 ) | ( n13094 & n13095 ) ;
  assign n13097 = n3998 & n4227 ;
  assign n13098 = x104 & n4231 ;
  assign n13099 = x105 | n13098 ;
  assign n13100 = ( n4233 & n13098 ) | ( n4233 & n13099 ) | ( n13098 & n13099 ) ;
  assign n13101 = x103 & n4470 ;
  assign n13102 = n13100 | n13101 ;
  assign n13103 = ( x44 & n13097 ) | ( x44 & ~n13102 ) | ( n13097 & ~n13102 ) ;
  assign n13104 = ( ~x44 & n13102 ) | ( ~x44 & n13103 ) | ( n13102 & n13103 ) ;
  assign n13105 = ( ~n13097 & n13103 ) | ( ~n13097 & n13104 ) | ( n13103 & n13104 ) ;
  assign n13106 = n3486 & n4787 ;
  assign n13107 = x101 & n4791 ;
  assign n13108 = x102 | n13107 ;
  assign n13109 = ( n4793 & n13107 ) | ( n4793 & n13108 ) | ( n13107 & n13108 ) ;
  assign n13110 = x100 & n5030 ;
  assign n13111 = n13109 | n13110 ;
  assign n13112 = ( x47 & n13106 ) | ( x47 & ~n13111 ) | ( n13106 & ~n13111 ) ;
  assign n13113 = ( ~x47 & n13111 ) | ( ~x47 & n13112 ) | ( n13111 & n13112 ) ;
  assign n13114 = ( ~n13106 & n13112 ) | ( ~n13106 & n13113 ) | ( n13112 & n13113 ) ;
  assign n13115 = n2877 & n5374 ;
  assign n13116 = x98 & n5378 ;
  assign n13117 = x99 | n13116 ;
  assign n13118 = ( n5380 & n13116 ) | ( n5380 & n13117 ) | ( n13116 & n13117 ) ;
  assign n13119 = x97 & n5638 ;
  assign n13120 = n13118 | n13119 ;
  assign n13121 = ( x50 & n13115 ) | ( x50 & ~n13120 ) | ( n13115 & ~n13120 ) ;
  assign n13122 = ( ~x50 & n13120 ) | ( ~x50 & n13121 ) | ( n13120 & n13121 ) ;
  assign n13123 = ( ~n13115 & n13121 ) | ( ~n13115 & n13122 ) | ( n13121 & n13122 ) ;
  assign n13124 = n2449 & n6027 ;
  assign n13125 = x95 & n6031 ;
  assign n13126 = x96 | n13125 ;
  assign n13127 = ( n6033 & n13125 ) | ( n6033 & n13126 ) | ( n13125 & n13126 ) ;
  assign n13128 = x94 & n6303 ;
  assign n13129 = n13127 | n13128 ;
  assign n13130 = ( x53 & n13124 ) | ( x53 & ~n13129 ) | ( n13124 & ~n13129 ) ;
  assign n13131 = ( ~x53 & n13129 ) | ( ~x53 & n13130 ) | ( n13129 & n13130 ) ;
  assign n13132 = ( ~n13124 & n13130 ) | ( ~n13124 & n13131 ) | ( n13130 & n13131 ) ;
  assign n13133 = n2057 & n6713 ;
  assign n13134 = x92 & n6717 ;
  assign n13135 = x93 | n13134 ;
  assign n13136 = ( n6719 & n13134 ) | ( n6719 & n13135 ) | ( n13134 & n13135 ) ;
  assign n13137 = x91 & n6980 ;
  assign n13138 = n13136 | n13137 ;
  assign n13139 = ( x56 & n13133 ) | ( x56 & ~n13138 ) | ( n13133 & ~n13138 ) ;
  assign n13140 = ( ~x56 & n13138 ) | ( ~x56 & n13139 ) | ( n13138 & n13139 ) ;
  assign n13141 = ( ~n13133 & n13139 ) | ( ~n13133 & n13140 ) | ( n13139 & n13140 ) ;
  assign n13142 = n1701 & n7423 ;
  assign n13143 = x89 & n7427 ;
  assign n13144 = x90 | n13143 ;
  assign n13145 = ( n7429 & n13143 ) | ( n7429 & n13144 ) | ( n13143 & n13144 ) ;
  assign n13146 = x88 & n7708 ;
  assign n13147 = n13145 | n13146 ;
  assign n13148 = ( x59 & n13142 ) | ( x59 & ~n13147 ) | ( n13142 & ~n13147 ) ;
  assign n13149 = ( ~x59 & n13147 ) | ( ~x59 & n13148 ) | ( n13147 & n13148 ) ;
  assign n13150 = ( ~n13142 & n13148 ) | ( ~n13142 & n13149 ) | ( n13148 & n13149 ) ;
  assign n13151 = n1466 & n8154 ;
  assign n13152 = x86 & n8158 ;
  assign n13153 = x87 | n13152 ;
  assign n13154 = ( n8160 & n13152 ) | ( n8160 & n13153 ) | ( n13152 & n13153 ) ;
  assign n13155 = x85 & n8439 ;
  assign n13156 = n13154 | n13155 ;
  assign n13157 = ( x62 & n13151 ) | ( x62 & ~n13156 ) | ( n13151 & ~n13156 ) ;
  assign n13158 = ( ~x62 & n13156 ) | ( ~x62 & n13157 ) | ( n13156 & n13157 ) ;
  assign n13159 = ( ~n13151 & n13157 ) | ( ~n13151 & n13158 ) | ( n13157 & n13158 ) ;
  assign n13160 = x83 & n8927 ;
  assign n13161 = ( ~x84 & n8693 ) | ( ~x84 & n8927 ) | ( n8693 & n8927 ) ;
  assign n13162 = ( n8693 & n13160 ) | ( n8693 & ~n13161 ) | ( n13160 & ~n13161 ) ;
  assign n13163 = ( n12953 & n13159 ) | ( n12953 & ~n13162 ) | ( n13159 & ~n13162 ) ;
  assign n13164 = ( ~n12953 & n13159 ) | ( ~n12953 & n13162 ) | ( n13159 & n13162 ) ;
  assign n13165 = ( ~n13159 & n13163 ) | ( ~n13159 & n13164 ) | ( n13163 & n13164 ) ;
  assign n13166 = ( n12963 & n13150 ) | ( n12963 & ~n13165 ) | ( n13150 & ~n13165 ) ;
  assign n13167 = ( ~n12963 & n13150 ) | ( ~n12963 & n13165 ) | ( n13150 & n13165 ) ;
  assign n13168 = ( ~n13150 & n13166 ) | ( ~n13150 & n13167 ) | ( n13166 & n13167 ) ;
  assign n13169 = ( n12975 & n13141 ) | ( n12975 & ~n13168 ) | ( n13141 & ~n13168 ) ;
  assign n13170 = ( ~n12975 & n13141 ) | ( ~n12975 & n13168 ) | ( n13141 & n13168 ) ;
  assign n13171 = ( ~n13141 & n13169 ) | ( ~n13141 & n13170 ) | ( n13169 & n13170 ) ;
  assign n13172 = ( n12978 & n13132 ) | ( n12978 & ~n13171 ) | ( n13132 & ~n13171 ) ;
  assign n13173 = ( ~n12978 & n13132 ) | ( ~n12978 & n13171 ) | ( n13132 & n13171 ) ;
  assign n13174 = ( ~n13132 & n13172 ) | ( ~n13132 & n13173 ) | ( n13172 & n13173 ) ;
  assign n13175 = ( n12990 & n13123 ) | ( n12990 & ~n13174 ) | ( n13123 & ~n13174 ) ;
  assign n13176 = ( ~n12990 & n13123 ) | ( ~n12990 & n13174 ) | ( n13123 & n13174 ) ;
  assign n13177 = ( ~n13123 & n13175 ) | ( ~n13123 & n13176 ) | ( n13175 & n13176 ) ;
  assign n13178 = ( n12993 & n13114 ) | ( n12993 & ~n13177 ) | ( n13114 & ~n13177 ) ;
  assign n13179 = ( ~n12993 & n13114 ) | ( ~n12993 & n13177 ) | ( n13114 & n13177 ) ;
  assign n13180 = ( ~n13114 & n13178 ) | ( ~n13114 & n13179 ) | ( n13178 & n13179 ) ;
  assign n13181 = ( n12996 & n13105 ) | ( n12996 & ~n13180 ) | ( n13105 & ~n13180 ) ;
  assign n13182 = ( ~n12996 & n13105 ) | ( ~n12996 & n13180 ) | ( n13105 & n13180 ) ;
  assign n13183 = ( ~n13105 & n13181 ) | ( ~n13105 & n13182 ) | ( n13181 & n13182 ) ;
  assign n13184 = ( n12999 & n13096 ) | ( n12999 & ~n13183 ) | ( n13096 & ~n13183 ) ;
  assign n13185 = ( ~n12999 & n13096 ) | ( ~n12999 & n13183 ) | ( n13096 & n13183 ) ;
  assign n13186 = ( ~n13096 & n13184 ) | ( ~n13096 & n13185 ) | ( n13184 & n13185 ) ;
  assign n13187 = n3224 & n5130 ;
  assign n13188 = x110 & n3228 ;
  assign n13189 = x111 | n13188 ;
  assign n13190 = ( n3230 & n13188 ) | ( n3230 & n13189 ) | ( n13188 & n13189 ) ;
  assign n13191 = x109 & n3413 ;
  assign n13192 = n13190 | n13191 ;
  assign n13193 = ( x38 & n13187 ) | ( x38 & ~n13192 ) | ( n13187 & ~n13192 ) ;
  assign n13194 = ( ~x38 & n13192 ) | ( ~x38 & n13193 ) | ( n13192 & n13193 ) ;
  assign n13195 = ( ~n13187 & n13193 ) | ( ~n13187 & n13194 ) | ( n13193 & n13194 ) ;
  assign n13196 = ( n13011 & n13186 ) | ( n13011 & ~n13195 ) | ( n13186 & ~n13195 ) ;
  assign n13197 = ( ~n13011 & n13186 ) | ( ~n13011 & n13195 ) | ( n13186 & n13195 ) ;
  assign n13198 = ( ~n13186 & n13196 ) | ( ~n13186 & n13197 ) | ( n13196 & n13197 ) ;
  assign n13199 = n2766 & n5750 ;
  assign n13200 = x113 & n2770 ;
  assign n13201 = x114 | n13200 ;
  assign n13202 = ( n2772 & n13200 ) | ( n2772 & n13201 ) | ( n13200 & n13201 ) ;
  assign n13203 = x112 & n2943 ;
  assign n13204 = n13202 | n13203 ;
  assign n13205 = ( x35 & n13199 ) | ( x35 & ~n13204 ) | ( n13199 & ~n13204 ) ;
  assign n13206 = ( ~x35 & n13204 ) | ( ~x35 & n13205 ) | ( n13204 & n13205 ) ;
  assign n13207 = ( ~n13199 & n13205 ) | ( ~n13199 & n13206 ) | ( n13205 & n13206 ) ;
  assign n13208 = ( n13023 & n13198 ) | ( n13023 & n13207 ) | ( n13198 & n13207 ) ;
  assign n13209 = ( ~n13023 & n13198 ) | ( ~n13023 & n13207 ) | ( n13198 & n13207 ) ;
  assign n13210 = ( n13023 & ~n13208 ) | ( n13023 & n13209 ) | ( ~n13208 & n13209 ) ;
  assign n13211 = ( n13035 & n13087 ) | ( n13035 & n13210 ) | ( n13087 & n13210 ) ;
  assign n13212 = ( n13035 & ~n13087 ) | ( n13035 & n13210 ) | ( ~n13087 & n13210 ) ;
  assign n13213 = ( n13087 & ~n13211 ) | ( n13087 & n13212 ) | ( ~n13211 & n13212 ) ;
  assign n13214 = n1949 & n7098 ;
  assign n13215 = x119 & n1953 ;
  assign n13216 = x120 | n13215 ;
  assign n13217 = ( n1955 & n13215 ) | ( n1955 & n13216 ) | ( n13215 & n13216 ) ;
  assign n13218 = x118 & n2114 ;
  assign n13219 = n13217 | n13218 ;
  assign n13220 = ( x29 & n13214 ) | ( x29 & ~n13219 ) | ( n13214 & ~n13219 ) ;
  assign n13221 = ( ~x29 & n13219 ) | ( ~x29 & n13220 ) | ( n13219 & n13220 ) ;
  assign n13222 = ( ~n13214 & n13220 ) | ( ~n13214 & n13221 ) | ( n13220 & n13221 ) ;
  assign n13223 = ( n13038 & n13213 ) | ( n13038 & n13222 ) | ( n13213 & n13222 ) ;
  assign n13224 = ( n13038 & ~n13213 ) | ( n13038 & n13222 ) | ( ~n13213 & n13222 ) ;
  assign n13225 = ( n13213 & ~n13223 ) | ( n13213 & n13224 ) | ( ~n13223 & n13224 ) ;
  assign n13226 = ( n13041 & n13078 ) | ( n13041 & n13225 ) | ( n13078 & n13225 ) ;
  assign n13227 = ( n13041 & ~n13078 ) | ( n13041 & n13225 ) | ( ~n13078 & n13225 ) ;
  assign n13228 = ( n13078 & ~n13226 ) | ( n13078 & n13227 ) | ( ~n13226 & n13227 ) ;
  assign n13229 = ( n13044 & n13069 ) | ( n13044 & n13228 ) | ( n13069 & n13228 ) ;
  assign n13230 = ( n13044 & ~n13069 ) | ( n13044 & n13228 ) | ( ~n13069 & n13228 ) ;
  assign n13231 = ( n13069 & ~n13229 ) | ( n13069 & n13230 ) | ( ~n13229 & n13230 ) ;
  assign n13232 = ( n13047 & n13060 ) | ( n13047 & n13231 ) | ( n13060 & n13231 ) ;
  assign n13233 = ( ~n13047 & n13060 ) | ( ~n13047 & n13231 ) | ( n13060 & n13231 ) ;
  assign n13234 = ( n13047 & ~n13232 ) | ( n13047 & n13233 ) | ( ~n13232 & n13233 ) ;
  assign n13235 = ( n13050 & n13053 ) | ( n13050 & n13234 ) | ( n13053 & n13234 ) ;
  assign n13236 = ( n13050 & ~n13053 ) | ( n13050 & n13234 ) | ( ~n13053 & n13234 ) ;
  assign n13237 = ( n13053 & ~n13235 ) | ( n13053 & n13236 ) | ( ~n13235 & n13236 ) ;
  assign n13238 = n1617 & n7841 ;
  assign n13239 = x123 & n1621 ;
  assign n13240 = x124 | n13239 ;
  assign n13241 = ( n1623 & n13239 ) | ( n1623 & n13240 ) | ( n13239 & n13240 ) ;
  assign n13242 = x122 & n1749 ;
  assign n13243 = n13241 | n13242 ;
  assign n13244 = ( x26 & n13238 ) | ( x26 & ~n13243 ) | ( n13238 & ~n13243 ) ;
  assign n13245 = ( ~x26 & n13243 ) | ( ~x26 & n13244 ) | ( n13243 & n13244 ) ;
  assign n13246 = ( ~n13238 & n13244 ) | ( ~n13238 & n13245 ) | ( n13244 & n13245 ) ;
  assign n13247 = n2320 & n6421 ;
  assign n13248 = x117 & n2324 ;
  assign n13249 = x118 | n13248 ;
  assign n13250 = ( n2326 & n13248 ) | ( n2326 & n13249 ) | ( n13248 & n13249 ) ;
  assign n13251 = x116 & n2497 ;
  assign n13252 = n13250 | n13251 ;
  assign n13253 = ( x32 & n13247 ) | ( x32 & ~n13252 ) | ( n13247 & ~n13252 ) ;
  assign n13254 = ( ~x32 & n13252 ) | ( ~x32 & n13253 ) | ( n13252 & n13253 ) ;
  assign n13255 = ( ~n13247 & n13253 ) | ( ~n13247 & n13254 ) | ( n13253 & n13254 ) ;
  assign n13256 = n3715 & n4734 ;
  assign n13257 = x108 & n3719 ;
  assign n13258 = x109 | n13257 ;
  assign n13259 = ( n3721 & n13257 ) | ( n3721 & n13258 ) | ( n13257 & n13258 ) ;
  assign n13260 = x107 & n3922 ;
  assign n13261 = n13259 | n13260 ;
  assign n13262 = ( x41 & n13256 ) | ( x41 & ~n13261 ) | ( n13256 & ~n13261 ) ;
  assign n13263 = ( ~x41 & n13261 ) | ( ~x41 & n13262 ) | ( n13261 & n13262 ) ;
  assign n13264 = ( ~n13256 & n13262 ) | ( ~n13256 & n13263 ) | ( n13262 & n13263 ) ;
  assign n13265 = n4013 & n4227 ;
  assign n13266 = x105 & n4231 ;
  assign n13267 = x106 | n13266 ;
  assign n13268 = ( n4233 & n13266 ) | ( n4233 & n13267 ) | ( n13266 & n13267 ) ;
  assign n13269 = x104 & n4470 ;
  assign n13270 = n13268 | n13269 ;
  assign n13271 = ( x44 & n13265 ) | ( x44 & ~n13270 ) | ( n13265 & ~n13270 ) ;
  assign n13272 = ( ~x44 & n13270 ) | ( ~x44 & n13271 ) | ( n13270 & n13271 ) ;
  assign n13273 = ( ~n13265 & n13271 ) | ( ~n13265 & n13272 ) | ( n13271 & n13272 ) ;
  assign n13274 = n3650 & n4787 ;
  assign n13275 = x102 & n4791 ;
  assign n13276 = x103 | n13275 ;
  assign n13277 = ( n4793 & n13275 ) | ( n4793 & n13276 ) | ( n13275 & n13276 ) ;
  assign n13278 = x101 & n5030 ;
  assign n13279 = n13277 | n13278 ;
  assign n13280 = ( x47 & n13274 ) | ( x47 & ~n13279 ) | ( n13274 & ~n13279 ) ;
  assign n13281 = ( ~x47 & n13279 ) | ( ~x47 & n13280 ) | ( n13279 & n13280 ) ;
  assign n13282 = ( ~n13274 & n13280 ) | ( ~n13274 & n13281 ) | ( n13280 & n13281 ) ;
  assign n13283 = n3162 & n5374 ;
  assign n13284 = x99 & n5378 ;
  assign n13285 = x100 | n13284 ;
  assign n13286 = ( n5380 & n13284 ) | ( n5380 & n13285 ) | ( n13284 & n13285 ) ;
  assign n13287 = x98 & n5638 ;
  assign n13288 = n13286 | n13287 ;
  assign n13289 = ( x50 & n13283 ) | ( x50 & ~n13288 ) | ( n13283 & ~n13288 ) ;
  assign n13290 = ( ~x50 & n13288 ) | ( ~x50 & n13289 ) | ( n13288 & n13289 ) ;
  assign n13291 = ( ~n13283 & n13289 ) | ( ~n13283 & n13290 ) | ( n13289 & n13290 ) ;
  assign n13292 = n2294 & n6713 ;
  assign n13293 = x93 & n6717 ;
  assign n13294 = x94 | n13293 ;
  assign n13295 = ( n6719 & n13293 ) | ( n6719 & n13294 ) | ( n13293 & n13294 ) ;
  assign n13296 = x92 & n6980 ;
  assign n13297 = n13295 | n13296 ;
  assign n13298 = ( x56 & n13292 ) | ( x56 & ~n13297 ) | ( n13292 & ~n13297 ) ;
  assign n13299 = ( ~x56 & n13297 ) | ( ~x56 & n13298 ) | ( n13297 & n13298 ) ;
  assign n13300 = ( ~n13292 & n13298 ) | ( ~n13292 & n13299 ) | ( n13298 & n13299 ) ;
  assign n13301 = n1914 & n7423 ;
  assign n13302 = x90 & n7427 ;
  assign n13303 = x91 | n13302 ;
  assign n13304 = ( n7429 & n13302 ) | ( n7429 & n13303 ) | ( n13302 & n13303 ) ;
  assign n13305 = x89 & n7708 ;
  assign n13306 = n13304 | n13305 ;
  assign n13307 = ( x59 & n13301 ) | ( x59 & ~n13306 ) | ( n13301 & ~n13306 ) ;
  assign n13308 = ( ~x59 & n13306 ) | ( ~x59 & n13307 ) | ( n13306 & n13307 ) ;
  assign n13309 = ( ~n13301 & n13307 ) | ( ~n13301 & n13308 ) | ( n13307 & n13308 ) ;
  assign n13310 = x84 & n8927 ;
  assign n13311 = ( ~x85 & n8693 ) | ( ~x85 & n8927 ) | ( n8693 & n8927 ) ;
  assign n13312 = ( n8693 & n13310 ) | ( n8693 & ~n13311 ) | ( n13310 & ~n13311 ) ;
  assign n13313 = ( ~x20 & n13162 ) | ( ~x20 & n13312 ) | ( n13162 & n13312 ) ;
  assign n13314 = ( n13162 & n13312 ) | ( n13162 & ~n13313 ) | ( n13312 & ~n13313 ) ;
  assign n13315 = ( x20 & n13313 ) | ( x20 & ~n13314 ) | ( n13313 & ~n13314 ) ;
  assign n13316 = n1481 & n8154 ;
  assign n13317 = x87 & n8158 ;
  assign n13318 = x88 | n13317 ;
  assign n13319 = ( n8160 & n13317 ) | ( n8160 & n13318 ) | ( n13317 & n13318 ) ;
  assign n13320 = x86 & n8439 ;
  assign n13321 = n13319 | n13320 ;
  assign n13322 = ( x62 & n13316 ) | ( x62 & ~n13321 ) | ( n13316 & ~n13321 ) ;
  assign n13323 = ( ~x62 & n13321 ) | ( ~x62 & n13322 ) | ( n13321 & n13322 ) ;
  assign n13324 = ( ~n13316 & n13322 ) | ( ~n13316 & n13323 ) | ( n13322 & n13323 ) ;
  assign n13325 = ( n13163 & ~n13315 ) | ( n13163 & n13324 ) | ( ~n13315 & n13324 ) ;
  assign n13326 = ( n13163 & n13315 ) | ( n13163 & n13324 ) | ( n13315 & n13324 ) ;
  assign n13327 = ( n13315 & n13325 ) | ( n13315 & ~n13326 ) | ( n13325 & ~n13326 ) ;
  assign n13328 = ( n13166 & n13309 ) | ( n13166 & ~n13327 ) | ( n13309 & ~n13327 ) ;
  assign n13329 = ( ~n13166 & n13309 ) | ( ~n13166 & n13327 ) | ( n13309 & n13327 ) ;
  assign n13330 = ( ~n13309 & n13328 ) | ( ~n13309 & n13329 ) | ( n13328 & n13329 ) ;
  assign n13331 = ( n13169 & n13300 ) | ( n13169 & ~n13330 ) | ( n13300 & ~n13330 ) ;
  assign n13332 = ( ~n13169 & n13300 ) | ( ~n13169 & n13330 ) | ( n13300 & n13330 ) ;
  assign n13333 = ( ~n13300 & n13331 ) | ( ~n13300 & n13332 ) | ( n13331 & n13332 ) ;
  assign n13334 = n2585 & n6027 ;
  assign n13335 = x96 & n6031 ;
  assign n13336 = x97 | n13335 ;
  assign n13337 = ( n6033 & n13335 ) | ( n6033 & n13336 ) | ( n13335 & n13336 ) ;
  assign n13338 = x95 & n6303 ;
  assign n13339 = n13337 | n13338 ;
  assign n13340 = ( x53 & n13334 ) | ( x53 & ~n13339 ) | ( n13334 & ~n13339 ) ;
  assign n13341 = ( ~x53 & n13339 ) | ( ~x53 & n13340 ) | ( n13339 & n13340 ) ;
  assign n13342 = ( ~n13334 & n13340 ) | ( ~n13334 & n13341 ) | ( n13340 & n13341 ) ;
  assign n13343 = ( n13172 & ~n13333 ) | ( n13172 & n13342 ) | ( ~n13333 & n13342 ) ;
  assign n13344 = ( n13172 & n13333 ) | ( n13172 & n13342 ) | ( n13333 & n13342 ) ;
  assign n13345 = ( n13333 & n13343 ) | ( n13333 & ~n13344 ) | ( n13343 & ~n13344 ) ;
  assign n13346 = ( n13175 & n13291 ) | ( n13175 & ~n13345 ) | ( n13291 & ~n13345 ) ;
  assign n13347 = ( ~n13175 & n13291 ) | ( ~n13175 & n13345 ) | ( n13291 & n13345 ) ;
  assign n13348 = ( ~n13291 & n13346 ) | ( ~n13291 & n13347 ) | ( n13346 & n13347 ) ;
  assign n13349 = ( n13178 & n13282 ) | ( n13178 & ~n13348 ) | ( n13282 & ~n13348 ) ;
  assign n13350 = ( ~n13178 & n13282 ) | ( ~n13178 & n13348 ) | ( n13282 & n13348 ) ;
  assign n13351 = ( ~n13282 & n13349 ) | ( ~n13282 & n13350 ) | ( n13349 & n13350 ) ;
  assign n13352 = ( n13181 & n13273 ) | ( n13181 & ~n13351 ) | ( n13273 & ~n13351 ) ;
  assign n13353 = ( ~n13181 & n13273 ) | ( ~n13181 & n13351 ) | ( n13273 & n13351 ) ;
  assign n13354 = ( ~n13273 & n13352 ) | ( ~n13273 & n13353 ) | ( n13352 & n13353 ) ;
  assign n13355 = ( n13184 & n13264 ) | ( n13184 & ~n13354 ) | ( n13264 & ~n13354 ) ;
  assign n13356 = ( ~n13184 & n13264 ) | ( ~n13184 & n13354 ) | ( n13264 & n13354 ) ;
  assign n13357 = ( ~n13264 & n13355 ) | ( ~n13264 & n13356 ) | ( n13355 & n13356 ) ;
  assign n13358 = n3224 & n5145 ;
  assign n13359 = x111 & n3228 ;
  assign n13360 = x112 | n13359 ;
  assign n13361 = ( n3230 & n13359 ) | ( n3230 & n13360 ) | ( n13359 & n13360 ) ;
  assign n13362 = x110 & n3413 ;
  assign n13363 = n13361 | n13362 ;
  assign n13364 = ( x38 & n13358 ) | ( x38 & ~n13363 ) | ( n13358 & ~n13363 ) ;
  assign n13365 = ( ~x38 & n13363 ) | ( ~x38 & n13364 ) | ( n13363 & n13364 ) ;
  assign n13366 = ( ~n13358 & n13364 ) | ( ~n13358 & n13365 ) | ( n13364 & n13365 ) ;
  assign n13367 = ( n13196 & n13357 ) | ( n13196 & ~n13366 ) | ( n13357 & ~n13366 ) ;
  assign n13368 = ( ~n13196 & n13357 ) | ( ~n13196 & n13366 ) | ( n13357 & n13366 ) ;
  assign n13369 = ( ~n13357 & n13367 ) | ( ~n13357 & n13368 ) | ( n13367 & n13368 ) ;
  assign n13370 = n2766 & n5765 ;
  assign n13371 = x114 & n2770 ;
  assign n13372 = x115 | n13371 ;
  assign n13373 = ( n2772 & n13371 ) | ( n2772 & n13372 ) | ( n13371 & n13372 ) ;
  assign n13374 = x113 & n2943 ;
  assign n13375 = n13373 | n13374 ;
  assign n13376 = ( x35 & n13370 ) | ( x35 & ~n13375 ) | ( n13370 & ~n13375 ) ;
  assign n13377 = ( ~x35 & n13375 ) | ( ~x35 & n13376 ) | ( n13375 & n13376 ) ;
  assign n13378 = ( ~n13370 & n13376 ) | ( ~n13370 & n13377 ) | ( n13376 & n13377 ) ;
  assign n13379 = ( n13208 & n13369 ) | ( n13208 & n13378 ) | ( n13369 & n13378 ) ;
  assign n13380 = ( ~n13208 & n13369 ) | ( ~n13208 & n13378 ) | ( n13369 & n13378 ) ;
  assign n13381 = ( n13208 & ~n13379 ) | ( n13208 & n13380 ) | ( ~n13379 & n13380 ) ;
  assign n13382 = ( n13211 & n13255 ) | ( n13211 & n13381 ) | ( n13255 & n13381 ) ;
  assign n13383 = ( n13211 & ~n13255 ) | ( n13211 & n13381 ) | ( ~n13255 & n13381 ) ;
  assign n13384 = ( n13255 & ~n13382 ) | ( n13255 & n13383 ) | ( ~n13382 & n13383 ) ;
  assign n13385 = n1949 & n7113 ;
  assign n13386 = x120 & n1953 ;
  assign n13387 = x121 | n13386 ;
  assign n13388 = ( n1955 & n13386 ) | ( n1955 & n13387 ) | ( n13386 & n13387 ) ;
  assign n13389 = x119 & n2114 ;
  assign n13390 = n13388 | n13389 ;
  assign n13391 = ( x29 & n13385 ) | ( x29 & ~n13390 ) | ( n13385 & ~n13390 ) ;
  assign n13392 = ( ~x29 & n13390 ) | ( ~x29 & n13391 ) | ( n13390 & n13391 ) ;
  assign n13393 = ( ~n13385 & n13391 ) | ( ~n13385 & n13392 ) | ( n13391 & n13392 ) ;
  assign n13394 = ( n13223 & n13384 ) | ( n13223 & n13393 ) | ( n13384 & n13393 ) ;
  assign n13395 = ( n13223 & ~n13384 ) | ( n13223 & n13393 ) | ( ~n13384 & n13393 ) ;
  assign n13396 = ( n13384 & ~n13394 ) | ( n13384 & n13395 ) | ( ~n13394 & n13395 ) ;
  assign n13397 = ( n13226 & n13246 ) | ( n13226 & n13396 ) | ( n13246 & n13396 ) ;
  assign n13398 = ( n13226 & ~n13246 ) | ( n13226 & n13396 ) | ( ~n13246 & n13396 ) ;
  assign n13399 = ( n13246 & ~n13397 ) | ( n13246 & n13398 ) | ( ~n13397 & n13398 ) ;
  assign n13400 = n1297 & n8846 ;
  assign n13401 = x126 & n1301 ;
  assign n13402 = x127 | n13401 ;
  assign n13403 = ( n1303 & n13401 ) | ( n1303 & n13402 ) | ( n13401 & n13402 ) ;
  assign n13404 = x125 & n1426 ;
  assign n13405 = n13403 | n13404 ;
  assign n13406 = ( x23 & n13400 ) | ( x23 & ~n13405 ) | ( n13400 & ~n13405 ) ;
  assign n13407 = ( ~x23 & n13405 ) | ( ~x23 & n13406 ) | ( n13405 & n13406 ) ;
  assign n13408 = ( ~n13400 & n13406 ) | ( ~n13400 & n13407 ) | ( n13406 & n13407 ) ;
  assign n13409 = ( n13229 & n13399 ) | ( n13229 & n13408 ) | ( n13399 & n13408 ) ;
  assign n13410 = ( n13229 & ~n13399 ) | ( n13229 & n13408 ) | ( ~n13399 & n13408 ) ;
  assign n13411 = ( n13399 & ~n13409 ) | ( n13399 & n13410 ) | ( ~n13409 & n13410 ) ;
  assign n13412 = ( n13232 & n13235 ) | ( n13232 & n13411 ) | ( n13235 & n13411 ) ;
  assign n13413 = ( ~n13232 & n13235 ) | ( ~n13232 & n13411 ) | ( n13235 & n13411 ) ;
  assign n13414 = ( n13232 & ~n13412 ) | ( n13232 & n13413 ) | ( ~n13412 & n13413 ) ;
  assign n13415 = n1297 & n8865 ;
  assign n13416 = x127 & n1301 ;
  assign n13417 = x126 | n13416 ;
  assign n13418 = ( n1426 & n13416 ) | ( n1426 & n13417 ) | ( n13416 & n13417 ) ;
  assign n13419 = ( x23 & n13415 ) | ( x23 & ~n13418 ) | ( n13415 & ~n13418 ) ;
  assign n13420 = ( ~x23 & n13418 ) | ( ~x23 & n13419 ) | ( n13418 & n13419 ) ;
  assign n13421 = ( ~n13415 & n13419 ) | ( ~n13415 & n13420 ) | ( n13419 & n13420 ) ;
  assign n13422 = n1617 & n8331 ;
  assign n13423 = x124 & n1621 ;
  assign n13424 = x125 | n13423 ;
  assign n13425 = ( n1623 & n13423 ) | ( n1623 & n13424 ) | ( n13423 & n13424 ) ;
  assign n13426 = x123 & n1749 ;
  assign n13427 = n13425 | n13426 ;
  assign n13428 = ( x26 & n13422 ) | ( x26 & ~n13427 ) | ( n13422 & ~n13427 ) ;
  assign n13429 = ( ~x26 & n13427 ) | ( ~x26 & n13428 ) | ( n13427 & n13428 ) ;
  assign n13430 = ( ~n13422 & n13428 ) | ( ~n13422 & n13429 ) | ( n13428 & n13429 ) ;
  assign n13431 = n1949 & n7582 ;
  assign n13432 = x121 & n1953 ;
  assign n13433 = x122 | n13432 ;
  assign n13434 = ( n1955 & n13432 ) | ( n1955 & n13433 ) | ( n13432 & n13433 ) ;
  assign n13435 = x120 & n2114 ;
  assign n13436 = n13434 | n13435 ;
  assign n13437 = ( x29 & n13431 ) | ( x29 & ~n13436 ) | ( n13431 & ~n13436 ) ;
  assign n13438 = ( ~x29 & n13436 ) | ( ~x29 & n13437 ) | ( n13436 & n13437 ) ;
  assign n13439 = ( ~n13431 & n13437 ) | ( ~n13431 & n13438 ) | ( n13437 & n13438 ) ;
  assign n13440 = n2320 & n6645 ;
  assign n13441 = x118 & n2324 ;
  assign n13442 = x119 | n13441 ;
  assign n13443 = ( n2326 & n13441 ) | ( n2326 & n13442 ) | ( n13441 & n13442 ) ;
  assign n13444 = x117 & n2497 ;
  assign n13445 = n13443 | n13444 ;
  assign n13446 = ( x32 & n13440 ) | ( x32 & ~n13445 ) | ( n13440 & ~n13445 ) ;
  assign n13447 = ( ~x32 & n13445 ) | ( ~x32 & n13446 ) | ( n13445 & n13446 ) ;
  assign n13448 = ( ~n13440 & n13446 ) | ( ~n13440 & n13447 ) | ( n13446 & n13447 ) ;
  assign n13449 = n3224 & n5542 ;
  assign n13450 = x112 & n3228 ;
  assign n13451 = x113 | n13450 ;
  assign n13452 = ( n3230 & n13450 ) | ( n3230 & n13451 ) | ( n13450 & n13451 ) ;
  assign n13453 = x111 & n3413 ;
  assign n13454 = n13452 | n13453 ;
  assign n13455 = ( x38 & n13449 ) | ( x38 & ~n13454 ) | ( n13449 & ~n13454 ) ;
  assign n13456 = ( ~x38 & n13454 ) | ( ~x38 & n13455 ) | ( n13454 & n13455 ) ;
  assign n13457 = ( ~n13449 & n13455 ) | ( ~n13449 & n13456 ) | ( n13455 & n13456 ) ;
  assign n13458 = n3715 & n4934 ;
  assign n13459 = x109 & n3719 ;
  assign n13460 = x110 | n13459 ;
  assign n13461 = ( n3721 & n13459 ) | ( n3721 & n13460 ) | ( n13459 & n13460 ) ;
  assign n13462 = x108 & n3922 ;
  assign n13463 = n13461 | n13462 ;
  assign n13464 = ( x41 & n13458 ) | ( x41 & ~n13463 ) | ( n13458 & ~n13463 ) ;
  assign n13465 = ( ~x41 & n13463 ) | ( ~x41 & n13464 ) | ( n13463 & n13464 ) ;
  assign n13466 = ( ~n13458 & n13464 ) | ( ~n13458 & n13465 ) | ( n13464 & n13465 ) ;
  assign n13467 = n4227 & n4362 ;
  assign n13468 = x106 & n4231 ;
  assign n13469 = x107 | n13468 ;
  assign n13470 = ( n4233 & n13468 ) | ( n4233 & n13469 ) | ( n13468 & n13469 ) ;
  assign n13471 = x105 & n4470 ;
  assign n13472 = n13470 | n13471 ;
  assign n13473 = ( x44 & n13467 ) | ( x44 & ~n13472 ) | ( n13467 & ~n13472 ) ;
  assign n13474 = ( ~x44 & n13472 ) | ( ~x44 & n13473 ) | ( n13472 & n13473 ) ;
  assign n13475 = ( ~n13467 & n13473 ) | ( ~n13467 & n13474 ) | ( n13473 & n13474 ) ;
  assign n13476 = n3665 & n4787 ;
  assign n13477 = x103 & n4791 ;
  assign n13478 = x104 | n13477 ;
  assign n13479 = ( n4793 & n13477 ) | ( n4793 & n13478 ) | ( n13477 & n13478 ) ;
  assign n13480 = x102 & n5030 ;
  assign n13481 = n13479 | n13480 ;
  assign n13482 = ( x47 & n13476 ) | ( x47 & ~n13481 ) | ( n13476 & ~n13481 ) ;
  assign n13483 = ( ~x47 & n13481 ) | ( ~x47 & n13482 ) | ( n13481 & n13482 ) ;
  assign n13484 = ( ~n13476 & n13482 ) | ( ~n13476 & n13483 ) | ( n13482 & n13483 ) ;
  assign n13485 = n3326 & n5374 ;
  assign n13486 = x100 & n5378 ;
  assign n13487 = x101 | n13486 ;
  assign n13488 = ( n5380 & n13486 ) | ( n5380 & n13487 ) | ( n13486 & n13487 ) ;
  assign n13489 = x99 & n5638 ;
  assign n13490 = n13488 | n13489 ;
  assign n13491 = ( x50 & n13485 ) | ( x50 & ~n13490 ) | ( n13485 & ~n13490 ) ;
  assign n13492 = ( ~x50 & n13490 ) | ( ~x50 & n13491 ) | ( n13490 & n13491 ) ;
  assign n13493 = ( ~n13485 & n13491 ) | ( ~n13485 & n13492 ) | ( n13491 & n13492 ) ;
  assign n13494 = n2725 & n6027 ;
  assign n13495 = x97 & n6031 ;
  assign n13496 = x98 | n13495 ;
  assign n13497 = ( n6033 & n13495 ) | ( n6033 & n13496 ) | ( n13495 & n13496 ) ;
  assign n13498 = x96 & n6303 ;
  assign n13499 = n13497 | n13498 ;
  assign n13500 = ( x53 & n13494 ) | ( x53 & ~n13499 ) | ( n13494 & ~n13499 ) ;
  assign n13501 = ( ~x53 & n13499 ) | ( ~x53 & n13500 ) | ( n13499 & n13500 ) ;
  assign n13502 = ( ~n13494 & n13500 ) | ( ~n13494 & n13501 ) | ( n13500 & n13501 ) ;
  assign n13503 = n2434 & n6713 ;
  assign n13504 = x94 & n6717 ;
  assign n13505 = x95 | n13504 ;
  assign n13506 = ( n6719 & n13504 ) | ( n6719 & n13505 ) | ( n13504 & n13505 ) ;
  assign n13507 = x93 & n6980 ;
  assign n13508 = n13506 | n13507 ;
  assign n13509 = ( x56 & n13503 ) | ( x56 & ~n13508 ) | ( n13503 & ~n13508 ) ;
  assign n13510 = ( ~x56 & n13508 ) | ( ~x56 & n13509 ) | ( n13508 & n13509 ) ;
  assign n13511 = ( ~n13503 & n13509 ) | ( ~n13503 & n13510 ) | ( n13509 & n13510 ) ;
  assign n13512 = n2042 & n7423 ;
  assign n13513 = x91 & n7427 ;
  assign n13514 = x92 | n13513 ;
  assign n13515 = ( n7429 & n13513 ) | ( n7429 & n13514 ) | ( n13513 & n13514 ) ;
  assign n13516 = x90 & n7708 ;
  assign n13517 = n13515 | n13516 ;
  assign n13518 = ( x59 & n13512 ) | ( x59 & ~n13517 ) | ( n13512 & ~n13517 ) ;
  assign n13519 = ( ~x59 & n13517 ) | ( ~x59 & n13518 ) | ( n13517 & n13518 ) ;
  assign n13520 = ( ~n13512 & n13518 ) | ( ~n13512 & n13519 ) | ( n13518 & n13519 ) ;
  assign n13521 = x85 & n8927 ;
  assign n13522 = ( ~x86 & n8693 ) | ( ~x86 & n8927 ) | ( n8693 & n8927 ) ;
  assign n13523 = ( n8693 & n13521 ) | ( n8693 & ~n13522 ) | ( n13521 & ~n13522 ) ;
  assign n13524 = n1585 & n8154 ;
  assign n13525 = x88 & n8158 ;
  assign n13526 = x89 | n13525 ;
  assign n13527 = ( n8160 & n13525 ) | ( n8160 & n13526 ) | ( n13525 & n13526 ) ;
  assign n13528 = x87 & n8439 ;
  assign n13529 = n13527 | n13528 ;
  assign n13530 = ( x62 & n13524 ) | ( x62 & ~n13529 ) | ( n13524 & ~n13529 ) ;
  assign n13531 = ( ~x62 & n13529 ) | ( ~x62 & n13530 ) | ( n13529 & n13530 ) ;
  assign n13532 = ( ~n13524 & n13530 ) | ( ~n13524 & n13531 ) | ( n13530 & n13531 ) ;
  assign n13533 = ( n13313 & ~n13523 ) | ( n13313 & n13532 ) | ( ~n13523 & n13532 ) ;
  assign n13534 = ( n13313 & n13523 ) | ( n13313 & n13532 ) | ( n13523 & n13532 ) ;
  assign n13535 = ( n13523 & n13533 ) | ( n13523 & ~n13534 ) | ( n13533 & ~n13534 ) ;
  assign n13536 = ( n13325 & n13520 ) | ( n13325 & ~n13535 ) | ( n13520 & ~n13535 ) ;
  assign n13537 = ( ~n13325 & n13520 ) | ( ~n13325 & n13535 ) | ( n13520 & n13535 ) ;
  assign n13538 = ( ~n13520 & n13536 ) | ( ~n13520 & n13537 ) | ( n13536 & n13537 ) ;
  assign n13539 = ( n13328 & n13511 ) | ( n13328 & ~n13538 ) | ( n13511 & ~n13538 ) ;
  assign n13540 = ( ~n13328 & n13511 ) | ( ~n13328 & n13538 ) | ( n13511 & n13538 ) ;
  assign n13541 = ( ~n13511 & n13539 ) | ( ~n13511 & n13540 ) | ( n13539 & n13540 ) ;
  assign n13542 = ( n13331 & n13502 ) | ( n13331 & ~n13541 ) | ( n13502 & ~n13541 ) ;
  assign n13543 = ( ~n13331 & n13502 ) | ( ~n13331 & n13541 ) | ( n13502 & n13541 ) ;
  assign n13544 = ( ~n13502 & n13542 ) | ( ~n13502 & n13543 ) | ( n13542 & n13543 ) ;
  assign n13545 = ( n13343 & n13493 ) | ( n13343 & ~n13544 ) | ( n13493 & ~n13544 ) ;
  assign n13546 = ( ~n13343 & n13493 ) | ( ~n13343 & n13544 ) | ( n13493 & n13544 ) ;
  assign n13547 = ( ~n13493 & n13545 ) | ( ~n13493 & n13546 ) | ( n13545 & n13546 ) ;
  assign n13548 = ( n13346 & n13484 ) | ( n13346 & ~n13547 ) | ( n13484 & ~n13547 ) ;
  assign n13549 = ( ~n13346 & n13484 ) | ( ~n13346 & n13547 ) | ( n13484 & n13547 ) ;
  assign n13550 = ( ~n13484 & n13548 ) | ( ~n13484 & n13549 ) | ( n13548 & n13549 ) ;
  assign n13551 = ( n13349 & n13475 ) | ( n13349 & ~n13550 ) | ( n13475 & ~n13550 ) ;
  assign n13552 = ( ~n13349 & n13475 ) | ( ~n13349 & n13550 ) | ( n13475 & n13550 ) ;
  assign n13553 = ( ~n13475 & n13551 ) | ( ~n13475 & n13552 ) | ( n13551 & n13552 ) ;
  assign n13554 = ( n13352 & n13466 ) | ( n13352 & ~n13553 ) | ( n13466 & ~n13553 ) ;
  assign n13555 = ( ~n13352 & n13466 ) | ( ~n13352 & n13553 ) | ( n13466 & n13553 ) ;
  assign n13556 = ( ~n13466 & n13554 ) | ( ~n13466 & n13555 ) | ( n13554 & n13555 ) ;
  assign n13557 = ( n13355 & n13457 ) | ( n13355 & ~n13556 ) | ( n13457 & ~n13556 ) ;
  assign n13558 = ( ~n13355 & n13457 ) | ( ~n13355 & n13556 ) | ( n13457 & n13556 ) ;
  assign n13559 = ( ~n13457 & n13557 ) | ( ~n13457 & n13558 ) | ( n13557 & n13558 ) ;
  assign n13560 = n2766 & n5977 ;
  assign n13561 = x115 & n2770 ;
  assign n13562 = x116 | n13561 ;
  assign n13563 = ( n2772 & n13561 ) | ( n2772 & n13562 ) | ( n13561 & n13562 ) ;
  assign n13564 = x114 & n2943 ;
  assign n13565 = n13563 | n13564 ;
  assign n13566 = ( x35 & n13560 ) | ( x35 & ~n13565 ) | ( n13560 & ~n13565 ) ;
  assign n13567 = ( ~x35 & n13565 ) | ( ~x35 & n13566 ) | ( n13565 & n13566 ) ;
  assign n13568 = ( ~n13560 & n13566 ) | ( ~n13560 & n13567 ) | ( n13566 & n13567 ) ;
  assign n13569 = ( n13367 & n13559 ) | ( n13367 & ~n13568 ) | ( n13559 & ~n13568 ) ;
  assign n13570 = ( ~n13367 & n13559 ) | ( ~n13367 & n13568 ) | ( n13559 & n13568 ) ;
  assign n13571 = ( ~n13559 & n13569 ) | ( ~n13559 & n13570 ) | ( n13569 & n13570 ) ;
  assign n13572 = ( n13379 & n13448 ) | ( n13379 & n13571 ) | ( n13448 & n13571 ) ;
  assign n13573 = ( n13379 & ~n13448 ) | ( n13379 & n13571 ) | ( ~n13448 & n13571 ) ;
  assign n13574 = ( n13448 & ~n13572 ) | ( n13448 & n13573 ) | ( ~n13572 & n13573 ) ;
  assign n13575 = ( n13382 & n13439 ) | ( n13382 & n13574 ) | ( n13439 & n13574 ) ;
  assign n13576 = ( ~n13382 & n13439 ) | ( ~n13382 & n13574 ) | ( n13439 & n13574 ) ;
  assign n13577 = ( n13382 & ~n13575 ) | ( n13382 & n13576 ) | ( ~n13575 & n13576 ) ;
  assign n13578 = ( n13394 & n13430 ) | ( n13394 & n13577 ) | ( n13430 & n13577 ) ;
  assign n13579 = ( n13394 & ~n13430 ) | ( n13394 & n13577 ) | ( ~n13430 & n13577 ) ;
  assign n13580 = ( n13430 & ~n13578 ) | ( n13430 & n13579 ) | ( ~n13578 & n13579 ) ;
  assign n13581 = ( n13397 & n13421 ) | ( n13397 & n13580 ) | ( n13421 & n13580 ) ;
  assign n13582 = ( ~n13397 & n13421 ) | ( ~n13397 & n13580 ) | ( n13421 & n13580 ) ;
  assign n13583 = ( n13397 & ~n13581 ) | ( n13397 & n13582 ) | ( ~n13581 & n13582 ) ;
  assign n13584 = ( n13409 & n13412 ) | ( n13409 & n13583 ) | ( n13412 & n13583 ) ;
  assign n13585 = ( ~n13409 & n13412 ) | ( ~n13409 & n13583 ) | ( n13412 & n13583 ) ;
  assign n13586 = ( n13409 & ~n13584 ) | ( n13409 & n13585 ) | ( ~n13584 & n13585 ) ;
  assign n13587 = n1297 & n8862 ;
  assign n13588 = ( x127 & n1426 ) | ( x127 & n13587 ) | ( n1426 & n13587 ) ;
  assign n13589 = x23 | n13588 ;
  assign n13590 = ~x23 & n13588 ;
  assign n13591 = ( ~n13588 & n13589 ) | ( ~n13588 & n13590 ) | ( n13589 & n13590 ) ;
  assign n13592 = n1617 & n8587 ;
  assign n13593 = x125 & n1621 ;
  assign n13594 = x126 | n13593 ;
  assign n13595 = ( n1623 & n13593 ) | ( n1623 & n13594 ) | ( n13593 & n13594 ) ;
  assign n13596 = x124 & n1749 ;
  assign n13597 = n13595 | n13596 ;
  assign n13598 = ( x26 & n13592 ) | ( x26 & ~n13597 ) | ( n13592 & ~n13597 ) ;
  assign n13599 = ( ~x26 & n13597 ) | ( ~x26 & n13598 ) | ( n13597 & n13598 ) ;
  assign n13600 = ( ~n13592 & n13598 ) | ( ~n13592 & n13599 ) | ( n13598 & n13599 ) ;
  assign n13601 = n1949 & n7597 ;
  assign n13602 = x122 & n1953 ;
  assign n13603 = x123 | n13602 ;
  assign n13604 = ( n1955 & n13602 ) | ( n1955 & n13603 ) | ( n13602 & n13603 ) ;
  assign n13605 = x121 & n2114 ;
  assign n13606 = n13604 | n13605 ;
  assign n13607 = ( x29 & n13601 ) | ( x29 & ~n13606 ) | ( n13601 & ~n13606 ) ;
  assign n13608 = ( ~x29 & n13606 ) | ( ~x29 & n13607 ) | ( n13606 & n13607 ) ;
  assign n13609 = ( ~n13601 & n13607 ) | ( ~n13601 & n13608 ) | ( n13607 & n13608 ) ;
  assign n13610 = n2320 & n7098 ;
  assign n13611 = x119 & n2324 ;
  assign n13612 = x120 | n13611 ;
  assign n13613 = ( n2326 & n13611 ) | ( n2326 & n13612 ) | ( n13611 & n13612 ) ;
  assign n13614 = x118 & n2497 ;
  assign n13615 = n13613 | n13614 ;
  assign n13616 = ( x32 & n13610 ) | ( x32 & ~n13615 ) | ( n13610 & ~n13615 ) ;
  assign n13617 = ( ~x32 & n13615 ) | ( ~x32 & n13616 ) | ( n13615 & n13616 ) ;
  assign n13618 = ( ~n13610 & n13616 ) | ( ~n13610 & n13617 ) | ( n13616 & n13617 ) ;
  assign n13619 = n2766 & n6201 ;
  assign n13620 = x116 & n2770 ;
  assign n13621 = x117 | n13620 ;
  assign n13622 = ( n2772 & n13620 ) | ( n2772 & n13621 ) | ( n13620 & n13621 ) ;
  assign n13623 = x115 & n2943 ;
  assign n13624 = n13622 | n13623 ;
  assign n13625 = ( x35 & n13619 ) | ( x35 & ~n13624 ) | ( n13619 & ~n13624 ) ;
  assign n13626 = ( ~x35 & n13624 ) | ( ~x35 & n13625 ) | ( n13624 & n13625 ) ;
  assign n13627 = ( ~n13619 & n13625 ) | ( ~n13619 & n13626 ) | ( n13625 & n13626 ) ;
  assign n13628 = n3224 & n5750 ;
  assign n13629 = x113 & n3228 ;
  assign n13630 = x114 | n13629 ;
  assign n13631 = ( n3230 & n13629 ) | ( n3230 & n13630 ) | ( n13629 & n13630 ) ;
  assign n13632 = x112 & n3413 ;
  assign n13633 = n13631 | n13632 ;
  assign n13634 = ( x38 & n13628 ) | ( x38 & ~n13633 ) | ( n13628 & ~n13633 ) ;
  assign n13635 = ( ~x38 & n13633 ) | ( ~x38 & n13634 ) | ( n13633 & n13634 ) ;
  assign n13636 = ( ~n13628 & n13634 ) | ( ~n13628 & n13635 ) | ( n13634 & n13635 ) ;
  assign n13637 = n3715 & n5130 ;
  assign n13638 = x110 & n3719 ;
  assign n13639 = x111 | n13638 ;
  assign n13640 = ( n3721 & n13638 ) | ( n3721 & n13639 ) | ( n13638 & n13639 ) ;
  assign n13641 = x109 & n3922 ;
  assign n13642 = n13640 | n13641 ;
  assign n13643 = ( x41 & n13637 ) | ( x41 & ~n13642 ) | ( n13637 & ~n13642 ) ;
  assign n13644 = ( ~x41 & n13642 ) | ( ~x41 & n13643 ) | ( n13642 & n13643 ) ;
  assign n13645 = ( ~n13637 & n13643 ) | ( ~n13637 & n13644 ) | ( n13643 & n13644 ) ;
  assign n13646 = n4227 & n4377 ;
  assign n13647 = x107 & n4231 ;
  assign n13648 = x108 | n13647 ;
  assign n13649 = ( n4233 & n13647 ) | ( n4233 & n13648 ) | ( n13647 & n13648 ) ;
  assign n13650 = x106 & n4470 ;
  assign n13651 = n13649 | n13650 ;
  assign n13652 = ( x44 & n13646 ) | ( x44 & ~n13651 ) | ( n13646 & ~n13651 ) ;
  assign n13653 = ( ~x44 & n13651 ) | ( ~x44 & n13652 ) | ( n13651 & n13652 ) ;
  assign n13654 = ( ~n13646 & n13652 ) | ( ~n13646 & n13653 ) | ( n13652 & n13653 ) ;
  assign n13655 = n3998 & n4787 ;
  assign n13656 = x104 & n4791 ;
  assign n13657 = x105 | n13656 ;
  assign n13658 = ( n4793 & n13656 ) | ( n4793 & n13657 ) | ( n13656 & n13657 ) ;
  assign n13659 = x103 & n5030 ;
  assign n13660 = n13658 | n13659 ;
  assign n13661 = ( x47 & n13655 ) | ( x47 & ~n13660 ) | ( n13655 & ~n13660 ) ;
  assign n13662 = ( ~x47 & n13660 ) | ( ~x47 & n13661 ) | ( n13660 & n13661 ) ;
  assign n13663 = ( ~n13655 & n13661 ) | ( ~n13655 & n13662 ) | ( n13661 & n13662 ) ;
  assign n13664 = n3486 & n5374 ;
  assign n13665 = x101 & n5378 ;
  assign n13666 = x102 | n13665 ;
  assign n13667 = ( n5380 & n13665 ) | ( n5380 & n13666 ) | ( n13665 & n13666 ) ;
  assign n13668 = x100 & n5638 ;
  assign n13669 = n13667 | n13668 ;
  assign n13670 = ( x50 & n13664 ) | ( x50 & ~n13669 ) | ( n13664 & ~n13669 ) ;
  assign n13671 = ( ~x50 & n13669 ) | ( ~x50 & n13670 ) | ( n13669 & n13670 ) ;
  assign n13672 = ( ~n13664 & n13670 ) | ( ~n13664 & n13671 ) | ( n13670 & n13671 ) ;
  assign n13673 = n2877 & n6027 ;
  assign n13674 = x98 & n6031 ;
  assign n13675 = x99 | n13674 ;
  assign n13676 = ( n6033 & n13674 ) | ( n6033 & n13675 ) | ( n13674 & n13675 ) ;
  assign n13677 = x97 & n6303 ;
  assign n13678 = n13676 | n13677 ;
  assign n13679 = ( x53 & n13673 ) | ( x53 & ~n13678 ) | ( n13673 & ~n13678 ) ;
  assign n13680 = ( ~x53 & n13678 ) | ( ~x53 & n13679 ) | ( n13678 & n13679 ) ;
  assign n13681 = ( ~n13673 & n13679 ) | ( ~n13673 & n13680 ) | ( n13679 & n13680 ) ;
  assign n13682 = n2449 & n6713 ;
  assign n13683 = x95 & n6717 ;
  assign n13684 = x96 | n13683 ;
  assign n13685 = ( n6719 & n13683 ) | ( n6719 & n13684 ) | ( n13683 & n13684 ) ;
  assign n13686 = x94 & n6980 ;
  assign n13687 = n13685 | n13686 ;
  assign n13688 = ( x56 & n13682 ) | ( x56 & ~n13687 ) | ( n13682 & ~n13687 ) ;
  assign n13689 = ( ~x56 & n13687 ) | ( ~x56 & n13688 ) | ( n13687 & n13688 ) ;
  assign n13690 = ( ~n13682 & n13688 ) | ( ~n13682 & n13689 ) | ( n13688 & n13689 ) ;
  assign n13691 = n2057 & n7423 ;
  assign n13692 = x92 & n7427 ;
  assign n13693 = x93 | n13692 ;
  assign n13694 = ( n7429 & n13692 ) | ( n7429 & n13693 ) | ( n13692 & n13693 ) ;
  assign n13695 = x91 & n7708 ;
  assign n13696 = n13694 | n13695 ;
  assign n13697 = ( x59 & n13691 ) | ( x59 & ~n13696 ) | ( n13691 & ~n13696 ) ;
  assign n13698 = ( ~x59 & n13696 ) | ( ~x59 & n13697 ) | ( n13696 & n13697 ) ;
  assign n13699 = ( ~n13691 & n13697 ) | ( ~n13691 & n13698 ) | ( n13697 & n13698 ) ;
  assign n13700 = n1701 & n8154 ;
  assign n13701 = x89 & n8158 ;
  assign n13702 = x90 | n13701 ;
  assign n13703 = ( n8160 & n13701 ) | ( n8160 & n13702 ) | ( n13701 & n13702 ) ;
  assign n13704 = x88 & n8439 ;
  assign n13705 = n13703 | n13704 ;
  assign n13706 = ( x62 & n13700 ) | ( x62 & ~n13705 ) | ( n13700 & ~n13705 ) ;
  assign n13707 = ( ~x62 & n13705 ) | ( ~x62 & n13706 ) | ( n13705 & n13706 ) ;
  assign n13708 = ( ~n13700 & n13706 ) | ( ~n13700 & n13707 ) | ( n13706 & n13707 ) ;
  assign n13709 = x86 & n8927 ;
  assign n13710 = ( ~x87 & n8693 ) | ( ~x87 & n8927 ) | ( n8693 & n8927 ) ;
  assign n13711 = ( n8693 & n13709 ) | ( n8693 & ~n13710 ) | ( n13709 & ~n13710 ) ;
  assign n13712 = ( n13523 & n13708 ) | ( n13523 & ~n13711 ) | ( n13708 & ~n13711 ) ;
  assign n13713 = ( ~n13523 & n13708 ) | ( ~n13523 & n13711 ) | ( n13708 & n13711 ) ;
  assign n13714 = ( ~n13708 & n13712 ) | ( ~n13708 & n13713 ) | ( n13712 & n13713 ) ;
  assign n13715 = ( n13533 & n13699 ) | ( n13533 & ~n13714 ) | ( n13699 & ~n13714 ) ;
  assign n13716 = ( ~n13533 & n13699 ) | ( ~n13533 & n13714 ) | ( n13699 & n13714 ) ;
  assign n13717 = ( ~n13699 & n13715 ) | ( ~n13699 & n13716 ) | ( n13715 & n13716 ) ;
  assign n13718 = ( n13536 & n13690 ) | ( n13536 & ~n13717 ) | ( n13690 & ~n13717 ) ;
  assign n13719 = ( ~n13536 & n13690 ) | ( ~n13536 & n13717 ) | ( n13690 & n13717 ) ;
  assign n13720 = ( ~n13690 & n13718 ) | ( ~n13690 & n13719 ) | ( n13718 & n13719 ) ;
  assign n13721 = ( n13539 & n13681 ) | ( n13539 & ~n13720 ) | ( n13681 & ~n13720 ) ;
  assign n13722 = ( ~n13539 & n13681 ) | ( ~n13539 & n13720 ) | ( n13681 & n13720 ) ;
  assign n13723 = ( ~n13681 & n13721 ) | ( ~n13681 & n13722 ) | ( n13721 & n13722 ) ;
  assign n13724 = ( n13542 & n13672 ) | ( n13542 & ~n13723 ) | ( n13672 & ~n13723 ) ;
  assign n13725 = ( ~n13542 & n13672 ) | ( ~n13542 & n13723 ) | ( n13672 & n13723 ) ;
  assign n13726 = ( ~n13672 & n13724 ) | ( ~n13672 & n13725 ) | ( n13724 & n13725 ) ;
  assign n13727 = ( n13545 & n13663 ) | ( n13545 & ~n13726 ) | ( n13663 & ~n13726 ) ;
  assign n13728 = ( ~n13545 & n13663 ) | ( ~n13545 & n13726 ) | ( n13663 & n13726 ) ;
  assign n13729 = ( ~n13663 & n13727 ) | ( ~n13663 & n13728 ) | ( n13727 & n13728 ) ;
  assign n13730 = ( n13548 & n13654 ) | ( n13548 & ~n13729 ) | ( n13654 & ~n13729 ) ;
  assign n13731 = ( ~n13548 & n13654 ) | ( ~n13548 & n13729 ) | ( n13654 & n13729 ) ;
  assign n13732 = ( ~n13654 & n13730 ) | ( ~n13654 & n13731 ) | ( n13730 & n13731 ) ;
  assign n13733 = ( n13551 & n13645 ) | ( n13551 & ~n13732 ) | ( n13645 & ~n13732 ) ;
  assign n13734 = ( ~n13551 & n13645 ) | ( ~n13551 & n13732 ) | ( n13645 & n13732 ) ;
  assign n13735 = ( ~n13645 & n13733 ) | ( ~n13645 & n13734 ) | ( n13733 & n13734 ) ;
  assign n13736 = ( n13554 & n13636 ) | ( n13554 & ~n13735 ) | ( n13636 & ~n13735 ) ;
  assign n13737 = ( ~n13554 & n13636 ) | ( ~n13554 & n13735 ) | ( n13636 & n13735 ) ;
  assign n13738 = ( ~n13636 & n13736 ) | ( ~n13636 & n13737 ) | ( n13736 & n13737 ) ;
  assign n13739 = ( n13557 & n13627 ) | ( n13557 & ~n13738 ) | ( n13627 & ~n13738 ) ;
  assign n13740 = ( ~n13557 & n13627 ) | ( ~n13557 & n13738 ) | ( n13627 & n13738 ) ;
  assign n13741 = ( ~n13627 & n13739 ) | ( ~n13627 & n13740 ) | ( n13739 & n13740 ) ;
  assign n13742 = ( n13569 & ~n13618 ) | ( n13569 & n13741 ) | ( ~n13618 & n13741 ) ;
  assign n13743 = ( n13569 & n13618 ) | ( n13569 & n13741 ) | ( n13618 & n13741 ) ;
  assign n13744 = ( n13618 & n13742 ) | ( n13618 & ~n13743 ) | ( n13742 & ~n13743 ) ;
  assign n13745 = ( n13572 & n13609 ) | ( n13572 & n13744 ) | ( n13609 & n13744 ) ;
  assign n13746 = ( n13572 & ~n13609 ) | ( n13572 & n13744 ) | ( ~n13609 & n13744 ) ;
  assign n13747 = ( n13609 & ~n13745 ) | ( n13609 & n13746 ) | ( ~n13745 & n13746 ) ;
  assign n13748 = ( n13575 & n13600 ) | ( n13575 & n13747 ) | ( n13600 & n13747 ) ;
  assign n13749 = ( n13575 & ~n13600 ) | ( n13575 & n13747 ) | ( ~n13600 & n13747 ) ;
  assign n13750 = ( n13600 & ~n13748 ) | ( n13600 & n13749 ) | ( ~n13748 & n13749 ) ;
  assign n13751 = ( n13578 & n13591 ) | ( n13578 & n13750 ) | ( n13591 & n13750 ) ;
  assign n13752 = ( ~n13578 & n13591 ) | ( ~n13578 & n13750 ) | ( n13591 & n13750 ) ;
  assign n13753 = ( n13578 & ~n13751 ) | ( n13578 & n13752 ) | ( ~n13751 & n13752 ) ;
  assign n13754 = ( n13581 & n13584 ) | ( n13581 & n13753 ) | ( n13584 & n13753 ) ;
  assign n13755 = ( n13581 & ~n13584 ) | ( n13581 & n13753 ) | ( ~n13584 & n13753 ) ;
  assign n13756 = ( n13584 & ~n13754 ) | ( n13584 & n13755 ) | ( ~n13754 & n13755 ) ;
  assign n13757 = n1949 & n7841 ;
  assign n13758 = x123 & n1953 ;
  assign n13759 = x124 | n13758 ;
  assign n13760 = ( n1955 & n13758 ) | ( n1955 & n13759 ) | ( n13758 & n13759 ) ;
  assign n13761 = x122 & n2114 ;
  assign n13762 = n13760 | n13761 ;
  assign n13763 = ( x29 & n13757 ) | ( x29 & ~n13762 ) | ( n13757 & ~n13762 ) ;
  assign n13764 = ( ~x29 & n13762 ) | ( ~x29 & n13763 ) | ( n13762 & n13763 ) ;
  assign n13765 = ( ~n13757 & n13763 ) | ( ~n13757 & n13764 ) | ( n13763 & n13764 ) ;
  assign n13766 = n2320 & n7113 ;
  assign n13767 = x120 & n2324 ;
  assign n13768 = x121 | n13767 ;
  assign n13769 = ( n2326 & n13767 ) | ( n2326 & n13768 ) | ( n13767 & n13768 ) ;
  assign n13770 = x119 & n2497 ;
  assign n13771 = n13769 | n13770 ;
  assign n13772 = ( x32 & n13766 ) | ( x32 & ~n13771 ) | ( n13766 & ~n13771 ) ;
  assign n13773 = ( ~x32 & n13771 ) | ( ~x32 & n13772 ) | ( n13771 & n13772 ) ;
  assign n13774 = ( ~n13766 & n13772 ) | ( ~n13766 & n13773 ) | ( n13772 & n13773 ) ;
  assign n13775 = n2766 & n6421 ;
  assign n13776 = x117 & n2770 ;
  assign n13777 = x118 | n13776 ;
  assign n13778 = ( n2772 & n13776 ) | ( n2772 & n13777 ) | ( n13776 & n13777 ) ;
  assign n13779 = x116 & n2943 ;
  assign n13780 = n13778 | n13779 ;
  assign n13781 = ( x35 & n13775 ) | ( x35 & ~n13780 ) | ( n13775 & ~n13780 ) ;
  assign n13782 = ( ~x35 & n13780 ) | ( ~x35 & n13781 ) | ( n13780 & n13781 ) ;
  assign n13783 = ( ~n13775 & n13781 ) | ( ~n13775 & n13782 ) | ( n13781 & n13782 ) ;
  assign n13784 = n3224 & n5765 ;
  assign n13785 = x114 & n3228 ;
  assign n13786 = x115 | n13785 ;
  assign n13787 = ( n3230 & n13785 ) | ( n3230 & n13786 ) | ( n13785 & n13786 ) ;
  assign n13788 = x113 & n3413 ;
  assign n13789 = n13787 | n13788 ;
  assign n13790 = ( x38 & n13784 ) | ( x38 & ~n13789 ) | ( n13784 & ~n13789 ) ;
  assign n13791 = ( ~x38 & n13789 ) | ( ~x38 & n13790 ) | ( n13789 & n13790 ) ;
  assign n13792 = ( ~n13784 & n13790 ) | ( ~n13784 & n13791 ) | ( n13790 & n13791 ) ;
  assign n13793 = n3715 & n5145 ;
  assign n13794 = x111 & n3719 ;
  assign n13795 = x112 | n13794 ;
  assign n13796 = ( n3721 & n13794 ) | ( n3721 & n13795 ) | ( n13794 & n13795 ) ;
  assign n13797 = x110 & n3922 ;
  assign n13798 = n13796 | n13797 ;
  assign n13799 = ( x41 & n13793 ) | ( x41 & ~n13798 ) | ( n13793 & ~n13798 ) ;
  assign n13800 = ( ~x41 & n13798 ) | ( ~x41 & n13799 ) | ( n13798 & n13799 ) ;
  assign n13801 = ( ~n13793 & n13799 ) | ( ~n13793 & n13800 ) | ( n13799 & n13800 ) ;
  assign n13802 = n4227 & n4734 ;
  assign n13803 = x108 & n4231 ;
  assign n13804 = x109 | n13803 ;
  assign n13805 = ( n4233 & n13803 ) | ( n4233 & n13804 ) | ( n13803 & n13804 ) ;
  assign n13806 = x107 & n4470 ;
  assign n13807 = n13805 | n13806 ;
  assign n13808 = ( x44 & n13802 ) | ( x44 & ~n13807 ) | ( n13802 & ~n13807 ) ;
  assign n13809 = ( ~x44 & n13807 ) | ( ~x44 & n13808 ) | ( n13807 & n13808 ) ;
  assign n13810 = ( ~n13802 & n13808 ) | ( ~n13802 & n13809 ) | ( n13808 & n13809 ) ;
  assign n13811 = n4013 & n4787 ;
  assign n13812 = x105 & n4791 ;
  assign n13813 = x106 | n13812 ;
  assign n13814 = ( n4793 & n13812 ) | ( n4793 & n13813 ) | ( n13812 & n13813 ) ;
  assign n13815 = x104 & n5030 ;
  assign n13816 = n13814 | n13815 ;
  assign n13817 = ( x47 & n13811 ) | ( x47 & ~n13816 ) | ( n13811 & ~n13816 ) ;
  assign n13818 = ( ~x47 & n13816 ) | ( ~x47 & n13817 ) | ( n13816 & n13817 ) ;
  assign n13819 = ( ~n13811 & n13817 ) | ( ~n13811 & n13818 ) | ( n13817 & n13818 ) ;
  assign n13820 = n3650 & n5374 ;
  assign n13821 = x102 & n5378 ;
  assign n13822 = x103 | n13821 ;
  assign n13823 = ( n5380 & n13821 ) | ( n5380 & n13822 ) | ( n13821 & n13822 ) ;
  assign n13824 = x101 & n5638 ;
  assign n13825 = n13823 | n13824 ;
  assign n13826 = ( x50 & n13820 ) | ( x50 & ~n13825 ) | ( n13820 & ~n13825 ) ;
  assign n13827 = ( ~x50 & n13825 ) | ( ~x50 & n13826 ) | ( n13825 & n13826 ) ;
  assign n13828 = ( ~n13820 & n13826 ) | ( ~n13820 & n13827 ) | ( n13826 & n13827 ) ;
  assign n13829 = n3162 & n6027 ;
  assign n13830 = x99 & n6031 ;
  assign n13831 = x100 | n13830 ;
  assign n13832 = ( n6033 & n13830 ) | ( n6033 & n13831 ) | ( n13830 & n13831 ) ;
  assign n13833 = x98 & n6303 ;
  assign n13834 = n13832 | n13833 ;
  assign n13835 = ( x53 & n13829 ) | ( x53 & ~n13834 ) | ( n13829 & ~n13834 ) ;
  assign n13836 = ( ~x53 & n13834 ) | ( ~x53 & n13835 ) | ( n13834 & n13835 ) ;
  assign n13837 = ( ~n13829 & n13835 ) | ( ~n13829 & n13836 ) | ( n13835 & n13836 ) ;
  assign n13838 = n2294 & n7423 ;
  assign n13839 = x93 & n7427 ;
  assign n13840 = x94 | n13839 ;
  assign n13841 = ( n7429 & n13839 ) | ( n7429 & n13840 ) | ( n13839 & n13840 ) ;
  assign n13842 = x92 & n7708 ;
  assign n13843 = n13841 | n13842 ;
  assign n13844 = ( x59 & n13838 ) | ( x59 & ~n13843 ) | ( n13838 & ~n13843 ) ;
  assign n13845 = ( ~x59 & n13843 ) | ( ~x59 & n13844 ) | ( n13843 & n13844 ) ;
  assign n13846 = ( ~n13838 & n13844 ) | ( ~n13838 & n13845 ) | ( n13844 & n13845 ) ;
  assign n13847 = n1914 & n8154 ;
  assign n13848 = x90 & n8158 ;
  assign n13849 = x91 | n13848 ;
  assign n13850 = ( n8160 & n13848 ) | ( n8160 & n13849 ) | ( n13848 & n13849 ) ;
  assign n13851 = x89 & n8439 ;
  assign n13852 = n13850 | n13851 ;
  assign n13853 = ( x62 & n13847 ) | ( x62 & ~n13852 ) | ( n13847 & ~n13852 ) ;
  assign n13854 = ( ~x62 & n13852 ) | ( ~x62 & n13853 ) | ( n13852 & n13853 ) ;
  assign n13855 = ( ~n13847 & n13853 ) | ( ~n13847 & n13854 ) | ( n13853 & n13854 ) ;
  assign n13856 = x87 & n8927 ;
  assign n13857 = ( ~x88 & n8693 ) | ( ~x88 & n8927 ) | ( n8693 & n8927 ) ;
  assign n13858 = ( n8693 & n13856 ) | ( n8693 & ~n13857 ) | ( n13856 & ~n13857 ) ;
  assign n13859 = ( ~x23 & n13711 ) | ( ~x23 & n13858 ) | ( n13711 & n13858 ) ;
  assign n13860 = ( n13711 & n13858 ) | ( n13711 & ~n13859 ) | ( n13858 & ~n13859 ) ;
  assign n13861 = ( x23 & n13859 ) | ( x23 & ~n13860 ) | ( n13859 & ~n13860 ) ;
  assign n13862 = ( n13712 & n13855 ) | ( n13712 & ~n13861 ) | ( n13855 & ~n13861 ) ;
  assign n13863 = ( ~n13712 & n13855 ) | ( ~n13712 & n13861 ) | ( n13855 & n13861 ) ;
  assign n13864 = ( ~n13855 & n13862 ) | ( ~n13855 & n13863 ) | ( n13862 & n13863 ) ;
  assign n13865 = ( n13715 & n13846 ) | ( n13715 & ~n13864 ) | ( n13846 & ~n13864 ) ;
  assign n13866 = ( ~n13715 & n13846 ) | ( ~n13715 & n13864 ) | ( n13846 & n13864 ) ;
  assign n13867 = ( ~n13846 & n13865 ) | ( ~n13846 & n13866 ) | ( n13865 & n13866 ) ;
  assign n13868 = n2585 & n6713 ;
  assign n13869 = x96 & n6717 ;
  assign n13870 = x97 | n13869 ;
  assign n13871 = ( n6719 & n13869 ) | ( n6719 & n13870 ) | ( n13869 & n13870 ) ;
  assign n13872 = x95 & n6980 ;
  assign n13873 = n13871 | n13872 ;
  assign n13874 = ( x56 & n13868 ) | ( x56 & ~n13873 ) | ( n13868 & ~n13873 ) ;
  assign n13875 = ( ~x56 & n13873 ) | ( ~x56 & n13874 ) | ( n13873 & n13874 ) ;
  assign n13876 = ( ~n13868 & n13874 ) | ( ~n13868 & n13875 ) | ( n13874 & n13875 ) ;
  assign n13877 = ( n13718 & ~n13867 ) | ( n13718 & n13876 ) | ( ~n13867 & n13876 ) ;
  assign n13878 = ( n13718 & n13867 ) | ( n13718 & n13876 ) | ( n13867 & n13876 ) ;
  assign n13879 = ( n13867 & n13877 ) | ( n13867 & ~n13878 ) | ( n13877 & ~n13878 ) ;
  assign n13880 = ( n13721 & n13837 ) | ( n13721 & ~n13879 ) | ( n13837 & ~n13879 ) ;
  assign n13881 = ( ~n13721 & n13837 ) | ( ~n13721 & n13879 ) | ( n13837 & n13879 ) ;
  assign n13882 = ( ~n13837 & n13880 ) | ( ~n13837 & n13881 ) | ( n13880 & n13881 ) ;
  assign n13883 = ( n13724 & n13828 ) | ( n13724 & ~n13882 ) | ( n13828 & ~n13882 ) ;
  assign n13884 = ( ~n13724 & n13828 ) | ( ~n13724 & n13882 ) | ( n13828 & n13882 ) ;
  assign n13885 = ( ~n13828 & n13883 ) | ( ~n13828 & n13884 ) | ( n13883 & n13884 ) ;
  assign n13886 = ( n13727 & n13819 ) | ( n13727 & ~n13885 ) | ( n13819 & ~n13885 ) ;
  assign n13887 = ( ~n13727 & n13819 ) | ( ~n13727 & n13885 ) | ( n13819 & n13885 ) ;
  assign n13888 = ( ~n13819 & n13886 ) | ( ~n13819 & n13887 ) | ( n13886 & n13887 ) ;
  assign n13889 = ( n13730 & n13810 ) | ( n13730 & ~n13888 ) | ( n13810 & ~n13888 ) ;
  assign n13890 = ( ~n13730 & n13810 ) | ( ~n13730 & n13888 ) | ( n13810 & n13888 ) ;
  assign n13891 = ( ~n13810 & n13889 ) | ( ~n13810 & n13890 ) | ( n13889 & n13890 ) ;
  assign n13892 = ( n13733 & n13801 ) | ( n13733 & ~n13891 ) | ( n13801 & ~n13891 ) ;
  assign n13893 = ( ~n13733 & n13801 ) | ( ~n13733 & n13891 ) | ( n13801 & n13891 ) ;
  assign n13894 = ( ~n13801 & n13892 ) | ( ~n13801 & n13893 ) | ( n13892 & n13893 ) ;
  assign n13895 = ( n13736 & n13792 ) | ( n13736 & ~n13894 ) | ( n13792 & ~n13894 ) ;
  assign n13896 = ( ~n13736 & n13792 ) | ( ~n13736 & n13894 ) | ( n13792 & n13894 ) ;
  assign n13897 = ( ~n13792 & n13895 ) | ( ~n13792 & n13896 ) | ( n13895 & n13896 ) ;
  assign n13898 = ( n13739 & n13783 ) | ( n13739 & ~n13897 ) | ( n13783 & ~n13897 ) ;
  assign n13899 = ( ~n13739 & n13783 ) | ( ~n13739 & n13897 ) | ( n13783 & n13897 ) ;
  assign n13900 = ( ~n13783 & n13898 ) | ( ~n13783 & n13899 ) | ( n13898 & n13899 ) ;
  assign n13901 = ( n13742 & ~n13774 ) | ( n13742 & n13900 ) | ( ~n13774 & n13900 ) ;
  assign n13902 = ( n13742 & n13774 ) | ( n13742 & n13900 ) | ( n13774 & n13900 ) ;
  assign n13903 = ( n13774 & n13901 ) | ( n13774 & ~n13902 ) | ( n13901 & ~n13902 ) ;
  assign n13904 = ( n13745 & n13765 ) | ( n13745 & n13903 ) | ( n13765 & n13903 ) ;
  assign n13905 = ( ~n13745 & n13765 ) | ( ~n13745 & n13903 ) | ( n13765 & n13903 ) ;
  assign n13906 = ( n13745 & ~n13904 ) | ( n13745 & n13905 ) | ( ~n13904 & n13905 ) ;
  assign n13907 = n1617 & n8846 ;
  assign n13908 = x126 & n1621 ;
  assign n13909 = x127 | n13908 ;
  assign n13910 = ( n1623 & n13908 ) | ( n1623 & n13909 ) | ( n13908 & n13909 ) ;
  assign n13911 = x125 & n1749 ;
  assign n13912 = n13910 | n13911 ;
  assign n13913 = ( x26 & n13907 ) | ( x26 & ~n13912 ) | ( n13907 & ~n13912 ) ;
  assign n13914 = ( ~x26 & n13912 ) | ( ~x26 & n13913 ) | ( n13912 & n13913 ) ;
  assign n13915 = ( ~n13907 & n13913 ) | ( ~n13907 & n13914 ) | ( n13913 & n13914 ) ;
  assign n13916 = ( n13748 & n13906 ) | ( n13748 & n13915 ) | ( n13906 & n13915 ) ;
  assign n13917 = ( n13748 & ~n13906 ) | ( n13748 & n13915 ) | ( ~n13906 & n13915 ) ;
  assign n13918 = ( n13906 & ~n13916 ) | ( n13906 & n13917 ) | ( ~n13916 & n13917 ) ;
  assign n13919 = ( n13751 & n13754 ) | ( n13751 & n13918 ) | ( n13754 & n13918 ) ;
  assign n13920 = ( n13751 & ~n13754 ) | ( n13751 & n13918 ) | ( ~n13754 & n13918 ) ;
  assign n13921 = ( n13754 & ~n13919 ) | ( n13754 & n13920 ) | ( ~n13919 & n13920 ) ;
  assign n13922 = n1617 & n8865 ;
  assign n13923 = x127 & n1621 ;
  assign n13924 = x126 | n13923 ;
  assign n13925 = ( n1749 & n13923 ) | ( n1749 & n13924 ) | ( n13923 & n13924 ) ;
  assign n13926 = ( x26 & n13922 ) | ( x26 & ~n13925 ) | ( n13922 & ~n13925 ) ;
  assign n13927 = ( ~x26 & n13925 ) | ( ~x26 & n13926 ) | ( n13925 & n13926 ) ;
  assign n13928 = ( ~n13922 & n13926 ) | ( ~n13922 & n13927 ) | ( n13926 & n13927 ) ;
  assign n13929 = n1949 & n8331 ;
  assign n13930 = x124 & n1953 ;
  assign n13931 = x125 | n13930 ;
  assign n13932 = ( n1955 & n13930 ) | ( n1955 & n13931 ) | ( n13930 & n13931 ) ;
  assign n13933 = x123 & n2114 ;
  assign n13934 = n13932 | n13933 ;
  assign n13935 = ( x29 & n13929 ) | ( x29 & ~n13934 ) | ( n13929 & ~n13934 ) ;
  assign n13936 = ( ~x29 & n13934 ) | ( ~x29 & n13935 ) | ( n13934 & n13935 ) ;
  assign n13937 = ( ~n13929 & n13935 ) | ( ~n13929 & n13936 ) | ( n13935 & n13936 ) ;
  assign n13938 = n2320 & n7582 ;
  assign n13939 = x121 & n2324 ;
  assign n13940 = x122 | n13939 ;
  assign n13941 = ( n2326 & n13939 ) | ( n2326 & n13940 ) | ( n13939 & n13940 ) ;
  assign n13942 = x120 & n2497 ;
  assign n13943 = n13941 | n13942 ;
  assign n13944 = ( x32 & n13938 ) | ( x32 & ~n13943 ) | ( n13938 & ~n13943 ) ;
  assign n13945 = ( ~x32 & n13943 ) | ( ~x32 & n13944 ) | ( n13943 & n13944 ) ;
  assign n13946 = ( ~n13938 & n13944 ) | ( ~n13938 & n13945 ) | ( n13944 & n13945 ) ;
  assign n13947 = n2766 & n6645 ;
  assign n13948 = x118 & n2770 ;
  assign n13949 = x119 | n13948 ;
  assign n13950 = ( n2772 & n13948 ) | ( n2772 & n13949 ) | ( n13948 & n13949 ) ;
  assign n13951 = x117 & n2943 ;
  assign n13952 = n13950 | n13951 ;
  assign n13953 = ( x35 & n13947 ) | ( x35 & ~n13952 ) | ( n13947 & ~n13952 ) ;
  assign n13954 = ( ~x35 & n13952 ) | ( ~x35 & n13953 ) | ( n13952 & n13953 ) ;
  assign n13955 = ( ~n13947 & n13953 ) | ( ~n13947 & n13954 ) | ( n13953 & n13954 ) ;
  assign n13956 = n3715 & n5542 ;
  assign n13957 = x112 & n3719 ;
  assign n13958 = x113 | n13957 ;
  assign n13959 = ( n3721 & n13957 ) | ( n3721 & n13958 ) | ( n13957 & n13958 ) ;
  assign n13960 = x111 & n3922 ;
  assign n13961 = n13959 | n13960 ;
  assign n13962 = ( x41 & n13956 ) | ( x41 & ~n13961 ) | ( n13956 & ~n13961 ) ;
  assign n13963 = ( ~x41 & n13961 ) | ( ~x41 & n13962 ) | ( n13961 & n13962 ) ;
  assign n13964 = ( ~n13956 & n13962 ) | ( ~n13956 & n13963 ) | ( n13962 & n13963 ) ;
  assign n13965 = n4362 & n4787 ;
  assign n13966 = x106 & n4791 ;
  assign n13967 = x107 | n13966 ;
  assign n13968 = ( n4793 & n13966 ) | ( n4793 & n13967 ) | ( n13966 & n13967 ) ;
  assign n13969 = x105 & n5030 ;
  assign n13970 = n13968 | n13969 ;
  assign n13971 = ( x47 & n13965 ) | ( x47 & ~n13970 ) | ( n13965 & ~n13970 ) ;
  assign n13972 = ( ~x47 & n13970 ) | ( ~x47 & n13971 ) | ( n13970 & n13971 ) ;
  assign n13973 = ( ~n13965 & n13971 ) | ( ~n13965 & n13972 ) | ( n13971 & n13972 ) ;
  assign n13974 = n3665 & n5374 ;
  assign n13975 = x103 & n5378 ;
  assign n13976 = x104 | n13975 ;
  assign n13977 = ( n5380 & n13975 ) | ( n5380 & n13976 ) | ( n13975 & n13976 ) ;
  assign n13978 = x102 & n5638 ;
  assign n13979 = n13977 | n13978 ;
  assign n13980 = ( x50 & n13974 ) | ( x50 & ~n13979 ) | ( n13974 & ~n13979 ) ;
  assign n13981 = ( ~x50 & n13979 ) | ( ~x50 & n13980 ) | ( n13979 & n13980 ) ;
  assign n13982 = ( ~n13974 & n13980 ) | ( ~n13974 & n13981 ) | ( n13980 & n13981 ) ;
  assign n13983 = n2725 & n6713 ;
  assign n13984 = x97 & n6717 ;
  assign n13985 = x98 | n13984 ;
  assign n13986 = ( n6719 & n13984 ) | ( n6719 & n13985 ) | ( n13984 & n13985 ) ;
  assign n13987 = x96 & n6980 ;
  assign n13988 = n13986 | n13987 ;
  assign n13989 = ( x56 & n13983 ) | ( x56 & ~n13988 ) | ( n13983 & ~n13988 ) ;
  assign n13990 = ( ~x56 & n13988 ) | ( ~x56 & n13989 ) | ( n13988 & n13989 ) ;
  assign n13991 = ( ~n13983 & n13989 ) | ( ~n13983 & n13990 ) | ( n13989 & n13990 ) ;
  assign n13992 = x88 & n8927 ;
  assign n13993 = ( ~x89 & n8693 ) | ( ~x89 & n8927 ) | ( n8693 & n8927 ) ;
  assign n13994 = ( n8693 & n13992 ) | ( n8693 & ~n13993 ) | ( n13992 & ~n13993 ) ;
  assign n13995 = n2042 & n8154 ;
  assign n13996 = x91 & n8158 ;
  assign n13997 = x92 | n13996 ;
  assign n13998 = ( n8160 & n13996 ) | ( n8160 & n13997 ) | ( n13996 & n13997 ) ;
  assign n13999 = x90 & n8439 ;
  assign n14000 = n13998 | n13999 ;
  assign n14001 = ( x62 & n13995 ) | ( x62 & ~n14000 ) | ( n13995 & ~n14000 ) ;
  assign n14002 = ( ~x62 & n14000 ) | ( ~x62 & n14001 ) | ( n14000 & n14001 ) ;
  assign n14003 = ( ~n13995 & n14001 ) | ( ~n13995 & n14002 ) | ( n14001 & n14002 ) ;
  assign n14004 = ( n13859 & ~n13994 ) | ( n13859 & n14003 ) | ( ~n13994 & n14003 ) ;
  assign n14005 = ( n13859 & n13994 ) | ( n13859 & n14003 ) | ( n13994 & n14003 ) ;
  assign n14006 = ( n13994 & n14004 ) | ( n13994 & ~n14005 ) | ( n14004 & ~n14005 ) ;
  assign n14007 = n2434 & n7423 ;
  assign n14008 = x94 & n7427 ;
  assign n14009 = x95 | n14008 ;
  assign n14010 = ( n7429 & n14008 ) | ( n7429 & n14009 ) | ( n14008 & n14009 ) ;
  assign n14011 = x93 & n7708 ;
  assign n14012 = n14010 | n14011 ;
  assign n14013 = ( x59 & n14007 ) | ( x59 & ~n14012 ) | ( n14007 & ~n14012 ) ;
  assign n14014 = ( ~x59 & n14012 ) | ( ~x59 & n14013 ) | ( n14012 & n14013 ) ;
  assign n14015 = ( ~n14007 & n14013 ) | ( ~n14007 & n14014 ) | ( n14013 & n14014 ) ;
  assign n14016 = ( n13862 & ~n14006 ) | ( n13862 & n14015 ) | ( ~n14006 & n14015 ) ;
  assign n14017 = ( n13862 & n14006 ) | ( n13862 & n14015 ) | ( n14006 & n14015 ) ;
  assign n14018 = ( n14006 & n14016 ) | ( n14006 & ~n14017 ) | ( n14016 & ~n14017 ) ;
  assign n14019 = ( n13865 & n13991 ) | ( n13865 & ~n14018 ) | ( n13991 & ~n14018 ) ;
  assign n14020 = ( ~n13865 & n13991 ) | ( ~n13865 & n14018 ) | ( n13991 & n14018 ) ;
  assign n14021 = ( ~n13991 & n14019 ) | ( ~n13991 & n14020 ) | ( n14019 & n14020 ) ;
  assign n14022 = n3326 & n6027 ;
  assign n14023 = x100 & n6031 ;
  assign n14024 = x101 | n14023 ;
  assign n14025 = ( n6033 & n14023 ) | ( n6033 & n14024 ) | ( n14023 & n14024 ) ;
  assign n14026 = x99 & n6303 ;
  assign n14027 = n14025 | n14026 ;
  assign n14028 = ( x53 & n14022 ) | ( x53 & ~n14027 ) | ( n14022 & ~n14027 ) ;
  assign n14029 = ( ~x53 & n14027 ) | ( ~x53 & n14028 ) | ( n14027 & n14028 ) ;
  assign n14030 = ( ~n14022 & n14028 ) | ( ~n14022 & n14029 ) | ( n14028 & n14029 ) ;
  assign n14031 = ( n13877 & ~n14021 ) | ( n13877 & n14030 ) | ( ~n14021 & n14030 ) ;
  assign n14032 = ( n13877 & n14021 ) | ( n13877 & n14030 ) | ( n14021 & n14030 ) ;
  assign n14033 = ( n14021 & n14031 ) | ( n14021 & ~n14032 ) | ( n14031 & ~n14032 ) ;
  assign n14034 = ( n13880 & n13982 ) | ( n13880 & ~n14033 ) | ( n13982 & ~n14033 ) ;
  assign n14035 = ( ~n13880 & n13982 ) | ( ~n13880 & n14033 ) | ( n13982 & n14033 ) ;
  assign n14036 = ( ~n13982 & n14034 ) | ( ~n13982 & n14035 ) | ( n14034 & n14035 ) ;
  assign n14037 = ( n13883 & n13973 ) | ( n13883 & ~n14036 ) | ( n13973 & ~n14036 ) ;
  assign n14038 = ( ~n13883 & n13973 ) | ( ~n13883 & n14036 ) | ( n13973 & n14036 ) ;
  assign n14039 = ( ~n13973 & n14037 ) | ( ~n13973 & n14038 ) | ( n14037 & n14038 ) ;
  assign n14040 = n4227 & n4934 ;
  assign n14041 = x109 & n4231 ;
  assign n14042 = x110 | n14041 ;
  assign n14043 = ( n4233 & n14041 ) | ( n4233 & n14042 ) | ( n14041 & n14042 ) ;
  assign n14044 = x108 & n4470 ;
  assign n14045 = n14043 | n14044 ;
  assign n14046 = ( x44 & n14040 ) | ( x44 & ~n14045 ) | ( n14040 & ~n14045 ) ;
  assign n14047 = ( ~x44 & n14045 ) | ( ~x44 & n14046 ) | ( n14045 & n14046 ) ;
  assign n14048 = ( ~n14040 & n14046 ) | ( ~n14040 & n14047 ) | ( n14046 & n14047 ) ;
  assign n14049 = ( n13886 & ~n14039 ) | ( n13886 & n14048 ) | ( ~n14039 & n14048 ) ;
  assign n14050 = ( n13886 & n14039 ) | ( n13886 & n14048 ) | ( n14039 & n14048 ) ;
  assign n14051 = ( n14039 & n14049 ) | ( n14039 & ~n14050 ) | ( n14049 & ~n14050 ) ;
  assign n14052 = ( n13889 & n13964 ) | ( n13889 & ~n14051 ) | ( n13964 & ~n14051 ) ;
  assign n14053 = ( ~n13889 & n13964 ) | ( ~n13889 & n14051 ) | ( n13964 & n14051 ) ;
  assign n14054 = ( ~n13964 & n14052 ) | ( ~n13964 & n14053 ) | ( n14052 & n14053 ) ;
  assign n14055 = n3224 & n5977 ;
  assign n14056 = x115 & n3228 ;
  assign n14057 = x116 | n14056 ;
  assign n14058 = ( n3230 & n14056 ) | ( n3230 & n14057 ) | ( n14056 & n14057 ) ;
  assign n14059 = x114 & n3413 ;
  assign n14060 = n14058 | n14059 ;
  assign n14061 = ( x38 & n14055 ) | ( x38 & ~n14060 ) | ( n14055 & ~n14060 ) ;
  assign n14062 = ( ~x38 & n14060 ) | ( ~x38 & n14061 ) | ( n14060 & n14061 ) ;
  assign n14063 = ( ~n14055 & n14061 ) | ( ~n14055 & n14062 ) | ( n14061 & n14062 ) ;
  assign n14064 = ( n13892 & ~n14054 ) | ( n13892 & n14063 ) | ( ~n14054 & n14063 ) ;
  assign n14065 = ( n13892 & n14054 ) | ( n13892 & n14063 ) | ( n14054 & n14063 ) ;
  assign n14066 = ( n14054 & n14064 ) | ( n14054 & ~n14065 ) | ( n14064 & ~n14065 ) ;
  assign n14067 = ( n13895 & n13955 ) | ( n13895 & ~n14066 ) | ( n13955 & ~n14066 ) ;
  assign n14068 = ( ~n13895 & n13955 ) | ( ~n13895 & n14066 ) | ( n13955 & n14066 ) ;
  assign n14069 = ( ~n13955 & n14067 ) | ( ~n13955 & n14068 ) | ( n14067 & n14068 ) ;
  assign n14070 = ( n13898 & n13946 ) | ( n13898 & ~n14069 ) | ( n13946 & ~n14069 ) ;
  assign n14071 = ( ~n13898 & n13946 ) | ( ~n13898 & n14069 ) | ( n13946 & n14069 ) ;
  assign n14072 = ( ~n13946 & n14070 ) | ( ~n13946 & n14071 ) | ( n14070 & n14071 ) ;
  assign n14073 = ( n13901 & ~n13937 ) | ( n13901 & n14072 ) | ( ~n13937 & n14072 ) ;
  assign n14074 = ( n13901 & n13937 ) | ( n13901 & n14072 ) | ( n13937 & n14072 ) ;
  assign n14075 = ( n13937 & n14073 ) | ( n13937 & ~n14074 ) | ( n14073 & ~n14074 ) ;
  assign n14076 = ( n13904 & n13928 ) | ( n13904 & n14075 ) | ( n13928 & n14075 ) ;
  assign n14077 = ( ~n13904 & n13928 ) | ( ~n13904 & n14075 ) | ( n13928 & n14075 ) ;
  assign n14078 = ( n13904 & ~n14076 ) | ( n13904 & n14077 ) | ( ~n14076 & n14077 ) ;
  assign n14079 = ( n13916 & n13919 ) | ( n13916 & n14078 ) | ( n13919 & n14078 ) ;
  assign n14080 = ( n13916 & ~n13919 ) | ( n13916 & n14078 ) | ( ~n13919 & n14078 ) ;
  assign n14081 = ( n13919 & ~n14079 ) | ( n13919 & n14080 ) | ( ~n14079 & n14080 ) ;
  assign n14082 = n1949 & n8587 ;
  assign n14083 = x125 & n1953 ;
  assign n14084 = x126 | n14083 ;
  assign n14085 = ( n1955 & n14083 ) | ( n1955 & n14084 ) | ( n14083 & n14084 ) ;
  assign n14086 = x124 & n2114 ;
  assign n14087 = n14085 | n14086 ;
  assign n14088 = ( x29 & n14082 ) | ( x29 & ~n14087 ) | ( n14082 & ~n14087 ) ;
  assign n14089 = ( ~x29 & n14087 ) | ( ~x29 & n14088 ) | ( n14087 & n14088 ) ;
  assign n14090 = ( ~n14082 & n14088 ) | ( ~n14082 & n14089 ) | ( n14088 & n14089 ) ;
  assign n14091 = n2320 & n7597 ;
  assign n14092 = x122 & n2324 ;
  assign n14093 = x123 | n14092 ;
  assign n14094 = ( n2326 & n14092 ) | ( n2326 & n14093 ) | ( n14092 & n14093 ) ;
  assign n14095 = x121 & n2497 ;
  assign n14096 = n14094 | n14095 ;
  assign n14097 = ( x32 & n14091 ) | ( x32 & ~n14096 ) | ( n14091 & ~n14096 ) ;
  assign n14098 = ( ~x32 & n14096 ) | ( ~x32 & n14097 ) | ( n14096 & n14097 ) ;
  assign n14099 = ( ~n14091 & n14097 ) | ( ~n14091 & n14098 ) | ( n14097 & n14098 ) ;
  assign n14100 = n2766 & n7098 ;
  assign n14101 = x119 & n2770 ;
  assign n14102 = x120 | n14101 ;
  assign n14103 = ( n2772 & n14101 ) | ( n2772 & n14102 ) | ( n14101 & n14102 ) ;
  assign n14104 = x118 & n2943 ;
  assign n14105 = n14103 | n14104 ;
  assign n14106 = ( x35 & n14100 ) | ( x35 & ~n14105 ) | ( n14100 & ~n14105 ) ;
  assign n14107 = ( ~x35 & n14105 ) | ( ~x35 & n14106 ) | ( n14105 & n14106 ) ;
  assign n14108 = ( ~n14100 & n14106 ) | ( ~n14100 & n14107 ) | ( n14106 & n14107 ) ;
  assign n14109 = n3224 & n6201 ;
  assign n14110 = x116 & n3228 ;
  assign n14111 = x117 | n14110 ;
  assign n14112 = ( n3230 & n14110 ) | ( n3230 & n14111 ) | ( n14110 & n14111 ) ;
  assign n14113 = x115 & n3413 ;
  assign n14114 = n14112 | n14113 ;
  assign n14115 = ( x38 & n14109 ) | ( x38 & ~n14114 ) | ( n14109 & ~n14114 ) ;
  assign n14116 = ( ~x38 & n14114 ) | ( ~x38 & n14115 ) | ( n14114 & n14115 ) ;
  assign n14117 = ( ~n14109 & n14115 ) | ( ~n14109 & n14116 ) | ( n14115 & n14116 ) ;
  assign n14118 = n3715 & n5750 ;
  assign n14119 = x113 & n3719 ;
  assign n14120 = x114 | n14119 ;
  assign n14121 = ( n3721 & n14119 ) | ( n3721 & n14120 ) | ( n14119 & n14120 ) ;
  assign n14122 = x112 & n3922 ;
  assign n14123 = n14121 | n14122 ;
  assign n14124 = ( x41 & n14118 ) | ( x41 & ~n14123 ) | ( n14118 & ~n14123 ) ;
  assign n14125 = ( ~x41 & n14123 ) | ( ~x41 & n14124 ) | ( n14123 & n14124 ) ;
  assign n14126 = ( ~n14118 & n14124 ) | ( ~n14118 & n14125 ) | ( n14124 & n14125 ) ;
  assign n14127 = n4227 & n5130 ;
  assign n14128 = x110 & n4231 ;
  assign n14129 = x111 | n14128 ;
  assign n14130 = ( n4233 & n14128 ) | ( n4233 & n14129 ) | ( n14128 & n14129 ) ;
  assign n14131 = x109 & n4470 ;
  assign n14132 = n14130 | n14131 ;
  assign n14133 = ( x44 & n14127 ) | ( x44 & ~n14132 ) | ( n14127 & ~n14132 ) ;
  assign n14134 = ( ~x44 & n14132 ) | ( ~x44 & n14133 ) | ( n14132 & n14133 ) ;
  assign n14135 = ( ~n14127 & n14133 ) | ( ~n14127 & n14134 ) | ( n14133 & n14134 ) ;
  assign n14136 = n4377 & n4787 ;
  assign n14137 = x107 & n4791 ;
  assign n14138 = x108 | n14137 ;
  assign n14139 = ( n4793 & n14137 ) | ( n4793 & n14138 ) | ( n14137 & n14138 ) ;
  assign n14140 = x106 & n5030 ;
  assign n14141 = n14139 | n14140 ;
  assign n14142 = ( x47 & n14136 ) | ( x47 & ~n14141 ) | ( n14136 & ~n14141 ) ;
  assign n14143 = ( ~x47 & n14141 ) | ( ~x47 & n14142 ) | ( n14141 & n14142 ) ;
  assign n14144 = ( ~n14136 & n14142 ) | ( ~n14136 & n14143 ) | ( n14142 & n14143 ) ;
  assign n14145 = n3998 & n5374 ;
  assign n14146 = x104 & n5378 ;
  assign n14147 = x105 | n14146 ;
  assign n14148 = ( n5380 & n14146 ) | ( n5380 & n14147 ) | ( n14146 & n14147 ) ;
  assign n14149 = x103 & n5638 ;
  assign n14150 = n14148 | n14149 ;
  assign n14151 = ( x50 & n14145 ) | ( x50 & ~n14150 ) | ( n14145 & ~n14150 ) ;
  assign n14152 = ( ~x50 & n14150 ) | ( ~x50 & n14151 ) | ( n14150 & n14151 ) ;
  assign n14153 = ( ~n14145 & n14151 ) | ( ~n14145 & n14152 ) | ( n14151 & n14152 ) ;
  assign n14154 = n2877 & n6713 ;
  assign n14155 = x98 & n6717 ;
  assign n14156 = x99 | n14155 ;
  assign n14157 = ( n6719 & n14155 ) | ( n6719 & n14156 ) | ( n14155 & n14156 ) ;
  assign n14158 = x97 & n6980 ;
  assign n14159 = n14157 | n14158 ;
  assign n14160 = ( x56 & n14154 ) | ( x56 & ~n14159 ) | ( n14154 & ~n14159 ) ;
  assign n14161 = ( ~x56 & n14159 ) | ( ~x56 & n14160 ) | ( n14159 & n14160 ) ;
  assign n14162 = ( ~n14154 & n14160 ) | ( ~n14154 & n14161 ) | ( n14160 & n14161 ) ;
  assign n14163 = n2449 & n7423 ;
  assign n14164 = x95 & n7427 ;
  assign n14165 = x96 | n14164 ;
  assign n14166 = ( n7429 & n14164 ) | ( n7429 & n14165 ) | ( n14164 & n14165 ) ;
  assign n14167 = x94 & n7708 ;
  assign n14168 = n14166 | n14167 ;
  assign n14169 = ( x59 & n14163 ) | ( x59 & ~n14168 ) | ( n14163 & ~n14168 ) ;
  assign n14170 = ( ~x59 & n14168 ) | ( ~x59 & n14169 ) | ( n14168 & n14169 ) ;
  assign n14171 = ( ~n14163 & n14169 ) | ( ~n14163 & n14170 ) | ( n14169 & n14170 ) ;
  assign n14172 = n2057 & n8154 ;
  assign n14173 = x92 & n8158 ;
  assign n14174 = x93 | n14173 ;
  assign n14175 = ( n8160 & n14173 ) | ( n8160 & n14174 ) | ( n14173 & n14174 ) ;
  assign n14176 = x91 & n8439 ;
  assign n14177 = n14175 | n14176 ;
  assign n14178 = ( x62 & n14172 ) | ( x62 & ~n14177 ) | ( n14172 & ~n14177 ) ;
  assign n14179 = ( ~x62 & n14177 ) | ( ~x62 & n14178 ) | ( n14177 & n14178 ) ;
  assign n14180 = ( ~n14172 & n14178 ) | ( ~n14172 & n14179 ) | ( n14178 & n14179 ) ;
  assign n14181 = x89 & n8927 ;
  assign n14182 = ( ~x90 & n8693 ) | ( ~x90 & n8927 ) | ( n8693 & n8927 ) ;
  assign n14183 = ( n8693 & n14181 ) | ( n8693 & ~n14182 ) | ( n14181 & ~n14182 ) ;
  assign n14184 = ( n13994 & n14180 ) | ( n13994 & ~n14183 ) | ( n14180 & ~n14183 ) ;
  assign n14185 = ( ~n13994 & n14180 ) | ( ~n13994 & n14183 ) | ( n14180 & n14183 ) ;
  assign n14186 = ( ~n14180 & n14184 ) | ( ~n14180 & n14185 ) | ( n14184 & n14185 ) ;
  assign n14187 = ( n14004 & n14171 ) | ( n14004 & ~n14186 ) | ( n14171 & ~n14186 ) ;
  assign n14188 = ( ~n14004 & n14171 ) | ( ~n14004 & n14186 ) | ( n14171 & n14186 ) ;
  assign n14189 = ( ~n14171 & n14187 ) | ( ~n14171 & n14188 ) | ( n14187 & n14188 ) ;
  assign n14190 = ( n14016 & n14162 ) | ( n14016 & ~n14189 ) | ( n14162 & ~n14189 ) ;
  assign n14191 = ( ~n14016 & n14162 ) | ( ~n14016 & n14189 ) | ( n14162 & n14189 ) ;
  assign n14192 = ( ~n14162 & n14190 ) | ( ~n14162 & n14191 ) | ( n14190 & n14191 ) ;
  assign n14193 = n3486 & n6027 ;
  assign n14194 = x101 & n6031 ;
  assign n14195 = x102 | n14194 ;
  assign n14196 = ( n6033 & n14194 ) | ( n6033 & n14195 ) | ( n14194 & n14195 ) ;
  assign n14197 = x100 & n6303 ;
  assign n14198 = n14196 | n14197 ;
  assign n14199 = ( x53 & n14193 ) | ( x53 & ~n14198 ) | ( n14193 & ~n14198 ) ;
  assign n14200 = ( ~x53 & n14198 ) | ( ~x53 & n14199 ) | ( n14198 & n14199 ) ;
  assign n14201 = ( ~n14193 & n14199 ) | ( ~n14193 & n14200 ) | ( n14199 & n14200 ) ;
  assign n14202 = ( n14019 & ~n14192 ) | ( n14019 & n14201 ) | ( ~n14192 & n14201 ) ;
  assign n14203 = ( n14019 & n14192 ) | ( n14019 & n14201 ) | ( n14192 & n14201 ) ;
  assign n14204 = ( n14192 & n14202 ) | ( n14192 & ~n14203 ) | ( n14202 & ~n14203 ) ;
  assign n14205 = ( n14031 & n14153 ) | ( n14031 & ~n14204 ) | ( n14153 & ~n14204 ) ;
  assign n14206 = ( ~n14031 & n14153 ) | ( ~n14031 & n14204 ) | ( n14153 & n14204 ) ;
  assign n14207 = ( ~n14153 & n14205 ) | ( ~n14153 & n14206 ) | ( n14205 & n14206 ) ;
  assign n14208 = ( n14034 & n14144 ) | ( n14034 & ~n14207 ) | ( n14144 & ~n14207 ) ;
  assign n14209 = ( ~n14034 & n14144 ) | ( ~n14034 & n14207 ) | ( n14144 & n14207 ) ;
  assign n14210 = ( ~n14144 & n14208 ) | ( ~n14144 & n14209 ) | ( n14208 & n14209 ) ;
  assign n14211 = ( n14037 & n14135 ) | ( n14037 & ~n14210 ) | ( n14135 & ~n14210 ) ;
  assign n14212 = ( ~n14037 & n14135 ) | ( ~n14037 & n14210 ) | ( n14135 & n14210 ) ;
  assign n14213 = ( ~n14135 & n14211 ) | ( ~n14135 & n14212 ) | ( n14211 & n14212 ) ;
  assign n14214 = ( n14049 & n14126 ) | ( n14049 & ~n14213 ) | ( n14126 & ~n14213 ) ;
  assign n14215 = ( ~n14049 & n14126 ) | ( ~n14049 & n14213 ) | ( n14126 & n14213 ) ;
  assign n14216 = ( ~n14126 & n14214 ) | ( ~n14126 & n14215 ) | ( n14214 & n14215 ) ;
  assign n14217 = ( n14052 & n14117 ) | ( n14052 & ~n14216 ) | ( n14117 & ~n14216 ) ;
  assign n14218 = ( ~n14052 & n14117 ) | ( ~n14052 & n14216 ) | ( n14117 & n14216 ) ;
  assign n14219 = ( ~n14117 & n14217 ) | ( ~n14117 & n14218 ) | ( n14217 & n14218 ) ;
  assign n14220 = ( n14064 & n14108 ) | ( n14064 & ~n14219 ) | ( n14108 & ~n14219 ) ;
  assign n14221 = ( ~n14064 & n14108 ) | ( ~n14064 & n14219 ) | ( n14108 & n14219 ) ;
  assign n14222 = ( ~n14108 & n14220 ) | ( ~n14108 & n14221 ) | ( n14220 & n14221 ) ;
  assign n14223 = ( n14067 & n14099 ) | ( n14067 & ~n14222 ) | ( n14099 & ~n14222 ) ;
  assign n14224 = ( ~n14067 & n14099 ) | ( ~n14067 & n14222 ) | ( n14099 & n14222 ) ;
  assign n14225 = ( ~n14099 & n14223 ) | ( ~n14099 & n14224 ) | ( n14223 & n14224 ) ;
  assign n14226 = ( n14070 & n14090 ) | ( n14070 & ~n14225 ) | ( n14090 & ~n14225 ) ;
  assign n14227 = ( ~n14070 & n14090 ) | ( ~n14070 & n14225 ) | ( n14090 & n14225 ) ;
  assign n14228 = ( ~n14090 & n14226 ) | ( ~n14090 & n14227 ) | ( n14226 & n14227 ) ;
  assign n14229 = n1617 & n8862 ;
  assign n14230 = ( x127 & n1749 ) | ( x127 & n14229 ) | ( n1749 & n14229 ) ;
  assign n14231 = x26 | n14230 ;
  assign n14232 = ~x26 & n14230 ;
  assign n14233 = ( ~n14230 & n14231 ) | ( ~n14230 & n14232 ) | ( n14231 & n14232 ) ;
  assign n14234 = ( n14073 & n14228 ) | ( n14073 & ~n14233 ) | ( n14228 & ~n14233 ) ;
  assign n14235 = ( ~n14073 & n14228 ) | ( ~n14073 & n14233 ) | ( n14228 & n14233 ) ;
  assign n14236 = ( ~n14228 & n14234 ) | ( ~n14228 & n14235 ) | ( n14234 & n14235 ) ;
  assign n14237 = ( n14076 & n14079 ) | ( n14076 & n14236 ) | ( n14079 & n14236 ) ;
  assign n14238 = ( n14076 & ~n14079 ) | ( n14076 & n14236 ) | ( ~n14079 & n14236 ) ;
  assign n14239 = ( n14079 & ~n14237 ) | ( n14079 & n14238 ) | ( ~n14237 & n14238 ) ;
  assign n14240 = n2766 & n7113 ;
  assign n14241 = x120 & n2770 ;
  assign n14242 = x121 | n14241 ;
  assign n14243 = ( n2772 & n14241 ) | ( n2772 & n14242 ) | ( n14241 & n14242 ) ;
  assign n14244 = x119 & n2943 ;
  assign n14245 = n14243 | n14244 ;
  assign n14246 = ( x35 & n14240 ) | ( x35 & ~n14245 ) | ( n14240 & ~n14245 ) ;
  assign n14247 = ( ~x35 & n14245 ) | ( ~x35 & n14246 ) | ( n14245 & n14246 ) ;
  assign n14248 = ( ~n14240 & n14246 ) | ( ~n14240 & n14247 ) | ( n14246 & n14247 ) ;
  assign n14249 = n3224 & n6421 ;
  assign n14250 = x117 & n3228 ;
  assign n14251 = x118 | n14250 ;
  assign n14252 = ( n3230 & n14250 ) | ( n3230 & n14251 ) | ( n14250 & n14251 ) ;
  assign n14253 = x116 & n3413 ;
  assign n14254 = n14252 | n14253 ;
  assign n14255 = ( x38 & n14249 ) | ( x38 & ~n14254 ) | ( n14249 & ~n14254 ) ;
  assign n14256 = ( ~x38 & n14254 ) | ( ~x38 & n14255 ) | ( n14254 & n14255 ) ;
  assign n14257 = ( ~n14249 & n14255 ) | ( ~n14249 & n14256 ) | ( n14255 & n14256 ) ;
  assign n14258 = n3715 & n5765 ;
  assign n14259 = x114 & n3719 ;
  assign n14260 = x115 | n14259 ;
  assign n14261 = ( n3721 & n14259 ) | ( n3721 & n14260 ) | ( n14259 & n14260 ) ;
  assign n14262 = x113 & n3922 ;
  assign n14263 = n14261 | n14262 ;
  assign n14264 = ( x41 & n14258 ) | ( x41 & ~n14263 ) | ( n14258 & ~n14263 ) ;
  assign n14265 = ( ~x41 & n14263 ) | ( ~x41 & n14264 ) | ( n14263 & n14264 ) ;
  assign n14266 = ( ~n14258 & n14264 ) | ( ~n14258 & n14265 ) | ( n14264 & n14265 ) ;
  assign n14267 = n4227 & n5145 ;
  assign n14268 = x111 & n4231 ;
  assign n14269 = x112 | n14268 ;
  assign n14270 = ( n4233 & n14268 ) | ( n4233 & n14269 ) | ( n14268 & n14269 ) ;
  assign n14271 = x110 & n4470 ;
  assign n14272 = n14270 | n14271 ;
  assign n14273 = ( x44 & n14267 ) | ( x44 & ~n14272 ) | ( n14267 & ~n14272 ) ;
  assign n14274 = ( ~x44 & n14272 ) | ( ~x44 & n14273 ) | ( n14272 & n14273 ) ;
  assign n14275 = ( ~n14267 & n14273 ) | ( ~n14267 & n14274 ) | ( n14273 & n14274 ) ;
  assign n14276 = n4734 & n4787 ;
  assign n14277 = x108 & n4791 ;
  assign n14278 = x109 | n14277 ;
  assign n14279 = ( n4793 & n14277 ) | ( n4793 & n14278 ) | ( n14277 & n14278 ) ;
  assign n14280 = x107 & n5030 ;
  assign n14281 = n14279 | n14280 ;
  assign n14282 = ( x47 & n14276 ) | ( x47 & ~n14281 ) | ( n14276 & ~n14281 ) ;
  assign n14283 = ( ~x47 & n14281 ) | ( ~x47 & n14282 ) | ( n14281 & n14282 ) ;
  assign n14284 = ( ~n14276 & n14282 ) | ( ~n14276 & n14283 ) | ( n14282 & n14283 ) ;
  assign n14285 = n4013 & n5374 ;
  assign n14286 = x105 & n5378 ;
  assign n14287 = x106 | n14286 ;
  assign n14288 = ( n5380 & n14286 ) | ( n5380 & n14287 ) | ( n14286 & n14287 ) ;
  assign n14289 = x104 & n5638 ;
  assign n14290 = n14288 | n14289 ;
  assign n14291 = ( x50 & n14285 ) | ( x50 & ~n14290 ) | ( n14285 & ~n14290 ) ;
  assign n14292 = ( ~x50 & n14290 ) | ( ~x50 & n14291 ) | ( n14290 & n14291 ) ;
  assign n14293 = ( ~n14285 & n14291 ) | ( ~n14285 & n14292 ) | ( n14291 & n14292 ) ;
  assign n14294 = n3650 & n6027 ;
  assign n14295 = x102 & n6031 ;
  assign n14296 = x103 | n14295 ;
  assign n14297 = ( n6033 & n14295 ) | ( n6033 & n14296 ) | ( n14295 & n14296 ) ;
  assign n14298 = x101 & n6303 ;
  assign n14299 = n14297 | n14298 ;
  assign n14300 = ( x53 & n14294 ) | ( x53 & ~n14299 ) | ( n14294 & ~n14299 ) ;
  assign n14301 = ( ~x53 & n14299 ) | ( ~x53 & n14300 ) | ( n14299 & n14300 ) ;
  assign n14302 = ( ~n14294 & n14300 ) | ( ~n14294 & n14301 ) | ( n14300 & n14301 ) ;
  assign n14303 = n3162 & n6713 ;
  assign n14304 = x99 & n6717 ;
  assign n14305 = x100 | n14304 ;
  assign n14306 = ( n6719 & n14304 ) | ( n6719 & n14305 ) | ( n14304 & n14305 ) ;
  assign n14307 = x98 & n6980 ;
  assign n14308 = n14306 | n14307 ;
  assign n14309 = ( x56 & n14303 ) | ( x56 & ~n14308 ) | ( n14303 & ~n14308 ) ;
  assign n14310 = ( ~x56 & n14308 ) | ( ~x56 & n14309 ) | ( n14308 & n14309 ) ;
  assign n14311 = ( ~n14303 & n14309 ) | ( ~n14303 & n14310 ) | ( n14309 & n14310 ) ;
  assign n14312 = n2585 & n7423 ;
  assign n14313 = x96 & n7427 ;
  assign n14314 = x97 | n14313 ;
  assign n14315 = ( n7429 & n14313 ) | ( n7429 & n14314 ) | ( n14313 & n14314 ) ;
  assign n14316 = x95 & n7708 ;
  assign n14317 = n14315 | n14316 ;
  assign n14318 = ( x59 & n14312 ) | ( x59 & ~n14317 ) | ( n14312 & ~n14317 ) ;
  assign n14319 = ( ~x59 & n14317 ) | ( ~x59 & n14318 ) | ( n14317 & n14318 ) ;
  assign n14320 = ( ~n14312 & n14318 ) | ( ~n14312 & n14319 ) | ( n14318 & n14319 ) ;
  assign n14321 = n2294 & n8154 ;
  assign n14322 = x93 & n8158 ;
  assign n14323 = x94 | n14322 ;
  assign n14324 = ( n8160 & n14322 ) | ( n8160 & n14323 ) | ( n14322 & n14323 ) ;
  assign n14325 = x92 & n8439 ;
  assign n14326 = n14324 | n14325 ;
  assign n14327 = ( x62 & n14321 ) | ( x62 & ~n14326 ) | ( n14321 & ~n14326 ) ;
  assign n14328 = ( ~x62 & n14326 ) | ( ~x62 & n14327 ) | ( n14326 & n14327 ) ;
  assign n14329 = ( ~n14321 & n14327 ) | ( ~n14321 & n14328 ) | ( n14327 & n14328 ) ;
  assign n14330 = x90 & n8927 ;
  assign n14331 = ( ~x91 & n8693 ) | ( ~x91 & n8927 ) | ( n8693 & n8927 ) ;
  assign n14332 = ( n8693 & n14330 ) | ( n8693 & ~n14331 ) | ( n14330 & ~n14331 ) ;
  assign n14333 = ( ~x26 & n14183 ) | ( ~x26 & n14332 ) | ( n14183 & n14332 ) ;
  assign n14334 = ( n14183 & n14332 ) | ( n14183 & ~n14333 ) | ( n14332 & ~n14333 ) ;
  assign n14335 = ( x26 & n14333 ) | ( x26 & ~n14334 ) | ( n14333 & ~n14334 ) ;
  assign n14336 = ( n14184 & n14329 ) | ( n14184 & ~n14335 ) | ( n14329 & ~n14335 ) ;
  assign n14337 = ( ~n14184 & n14329 ) | ( ~n14184 & n14335 ) | ( n14329 & n14335 ) ;
  assign n14338 = ( ~n14329 & n14336 ) | ( ~n14329 & n14337 ) | ( n14336 & n14337 ) ;
  assign n14339 = ( n14187 & n14320 ) | ( n14187 & ~n14338 ) | ( n14320 & ~n14338 ) ;
  assign n14340 = ( ~n14187 & n14320 ) | ( ~n14187 & n14338 ) | ( n14320 & n14338 ) ;
  assign n14341 = ( ~n14320 & n14339 ) | ( ~n14320 & n14340 ) | ( n14339 & n14340 ) ;
  assign n14342 = ( n14190 & n14311 ) | ( n14190 & ~n14341 ) | ( n14311 & ~n14341 ) ;
  assign n14343 = ( ~n14190 & n14311 ) | ( ~n14190 & n14341 ) | ( n14311 & n14341 ) ;
  assign n14344 = ( ~n14311 & n14342 ) | ( ~n14311 & n14343 ) | ( n14342 & n14343 ) ;
  assign n14345 = ( n14202 & n14302 ) | ( n14202 & ~n14344 ) | ( n14302 & ~n14344 ) ;
  assign n14346 = ( ~n14202 & n14302 ) | ( ~n14202 & n14344 ) | ( n14302 & n14344 ) ;
  assign n14347 = ( ~n14302 & n14345 ) | ( ~n14302 & n14346 ) | ( n14345 & n14346 ) ;
  assign n14348 = ( n14205 & n14293 ) | ( n14205 & ~n14347 ) | ( n14293 & ~n14347 ) ;
  assign n14349 = ( ~n14205 & n14293 ) | ( ~n14205 & n14347 ) | ( n14293 & n14347 ) ;
  assign n14350 = ( ~n14293 & n14348 ) | ( ~n14293 & n14349 ) | ( n14348 & n14349 ) ;
  assign n14351 = ( n14208 & n14284 ) | ( n14208 & ~n14350 ) | ( n14284 & ~n14350 ) ;
  assign n14352 = ( ~n14208 & n14284 ) | ( ~n14208 & n14350 ) | ( n14284 & n14350 ) ;
  assign n14353 = ( ~n14284 & n14351 ) | ( ~n14284 & n14352 ) | ( n14351 & n14352 ) ;
  assign n14354 = ( n14211 & n14275 ) | ( n14211 & ~n14353 ) | ( n14275 & ~n14353 ) ;
  assign n14355 = ( ~n14211 & n14275 ) | ( ~n14211 & n14353 ) | ( n14275 & n14353 ) ;
  assign n14356 = ( ~n14275 & n14354 ) | ( ~n14275 & n14355 ) | ( n14354 & n14355 ) ;
  assign n14357 = ( n14214 & n14266 ) | ( n14214 & ~n14356 ) | ( n14266 & ~n14356 ) ;
  assign n14358 = ( ~n14214 & n14266 ) | ( ~n14214 & n14356 ) | ( n14266 & n14356 ) ;
  assign n14359 = ( ~n14266 & n14357 ) | ( ~n14266 & n14358 ) | ( n14357 & n14358 ) ;
  assign n14360 = ( n14217 & n14257 ) | ( n14217 & ~n14359 ) | ( n14257 & ~n14359 ) ;
  assign n14361 = ( ~n14217 & n14257 ) | ( ~n14217 & n14359 ) | ( n14257 & n14359 ) ;
  assign n14362 = ( ~n14257 & n14360 ) | ( ~n14257 & n14361 ) | ( n14360 & n14361 ) ;
  assign n14363 = ( n14220 & n14248 ) | ( n14220 & ~n14362 ) | ( n14248 & ~n14362 ) ;
  assign n14364 = ( ~n14220 & n14248 ) | ( ~n14220 & n14362 ) | ( n14248 & n14362 ) ;
  assign n14365 = ( ~n14248 & n14363 ) | ( ~n14248 & n14364 ) | ( n14363 & n14364 ) ;
  assign n14366 = n2320 & n7841 ;
  assign n14367 = x123 & n2324 ;
  assign n14368 = x124 | n14367 ;
  assign n14369 = ( n2326 & n14367 ) | ( n2326 & n14368 ) | ( n14367 & n14368 ) ;
  assign n14370 = x122 & n2497 ;
  assign n14371 = n14369 | n14370 ;
  assign n14372 = ( x32 & n14366 ) | ( x32 & ~n14371 ) | ( n14366 & ~n14371 ) ;
  assign n14373 = ( ~x32 & n14371 ) | ( ~x32 & n14372 ) | ( n14371 & n14372 ) ;
  assign n14374 = ( ~n14366 & n14372 ) | ( ~n14366 & n14373 ) | ( n14372 & n14373 ) ;
  assign n14375 = ( n14223 & ~n14365 ) | ( n14223 & n14374 ) | ( ~n14365 & n14374 ) ;
  assign n14376 = ( n14223 & n14365 ) | ( n14223 & n14374 ) | ( n14365 & n14374 ) ;
  assign n14377 = ( n14365 & n14375 ) | ( n14365 & ~n14376 ) | ( n14375 & ~n14376 ) ;
  assign n14378 = n1949 & n8846 ;
  assign n14379 = x126 & n1953 ;
  assign n14380 = x127 | n14379 ;
  assign n14381 = ( n1955 & n14379 ) | ( n1955 & n14380 ) | ( n14379 & n14380 ) ;
  assign n14382 = x125 & n2114 ;
  assign n14383 = n14381 | n14382 ;
  assign n14384 = ( x29 & n14378 ) | ( x29 & ~n14383 ) | ( n14378 & ~n14383 ) ;
  assign n14385 = ( ~x29 & n14383 ) | ( ~x29 & n14384 ) | ( n14383 & n14384 ) ;
  assign n14386 = ( ~n14378 & n14384 ) | ( ~n14378 & n14385 ) | ( n14384 & n14385 ) ;
  assign n14387 = ( n14226 & ~n14377 ) | ( n14226 & n14386 ) | ( ~n14377 & n14386 ) ;
  assign n14388 = ( n14226 & n14377 ) | ( n14226 & n14386 ) | ( n14377 & n14386 ) ;
  assign n14389 = ( n14377 & n14387 ) | ( n14377 & ~n14388 ) | ( n14387 & ~n14388 ) ;
  assign n14390 = ( n14234 & ~n14237 ) | ( n14234 & n14389 ) | ( ~n14237 & n14389 ) ;
  assign n14391 = ( ~n14234 & n14237 ) | ( ~n14234 & n14389 ) | ( n14237 & n14389 ) ;
  assign n14392 = ( ~n14389 & n14390 ) | ( ~n14389 & n14391 ) | ( n14390 & n14391 ) ;
  assign n14393 = n1949 & n8865 ;
  assign n14394 = x127 & n1953 ;
  assign n14395 = x126 | n14394 ;
  assign n14396 = ( n2114 & n14394 ) | ( n2114 & n14395 ) | ( n14394 & n14395 ) ;
  assign n14397 = ( x29 & n14393 ) | ( x29 & ~n14396 ) | ( n14393 & ~n14396 ) ;
  assign n14398 = ( ~x29 & n14396 ) | ( ~x29 & n14397 ) | ( n14396 & n14397 ) ;
  assign n14399 = ( ~n14393 & n14397 ) | ( ~n14393 & n14398 ) | ( n14397 & n14398 ) ;
  assign n14400 = n2320 & n8331 ;
  assign n14401 = x124 & n2324 ;
  assign n14402 = x125 | n14401 ;
  assign n14403 = ( n2326 & n14401 ) | ( n2326 & n14402 ) | ( n14401 & n14402 ) ;
  assign n14404 = x123 & n2497 ;
  assign n14405 = n14403 | n14404 ;
  assign n14406 = ( x32 & n14400 ) | ( x32 & ~n14405 ) | ( n14400 & ~n14405 ) ;
  assign n14407 = ( ~x32 & n14405 ) | ( ~x32 & n14406 ) | ( n14405 & n14406 ) ;
  assign n14408 = ( ~n14400 & n14406 ) | ( ~n14400 & n14407 ) | ( n14406 & n14407 ) ;
  assign n14409 = n2766 & n7582 ;
  assign n14410 = x121 & n2770 ;
  assign n14411 = x122 | n14410 ;
  assign n14412 = ( n2772 & n14410 ) | ( n2772 & n14411 ) | ( n14410 & n14411 ) ;
  assign n14413 = x120 & n2943 ;
  assign n14414 = n14412 | n14413 ;
  assign n14415 = ( x35 & n14409 ) | ( x35 & ~n14414 ) | ( n14409 & ~n14414 ) ;
  assign n14416 = ( ~x35 & n14414 ) | ( ~x35 & n14415 ) | ( n14414 & n14415 ) ;
  assign n14417 = ( ~n14409 & n14415 ) | ( ~n14409 & n14416 ) | ( n14415 & n14416 ) ;
  assign n14418 = n3224 & n6645 ;
  assign n14419 = x118 & n3228 ;
  assign n14420 = x119 | n14419 ;
  assign n14421 = ( n3230 & n14419 ) | ( n3230 & n14420 ) | ( n14419 & n14420 ) ;
  assign n14422 = x117 & n3413 ;
  assign n14423 = n14421 | n14422 ;
  assign n14424 = ( x38 & n14418 ) | ( x38 & ~n14423 ) | ( n14418 & ~n14423 ) ;
  assign n14425 = ( ~x38 & n14423 ) | ( ~x38 & n14424 ) | ( n14423 & n14424 ) ;
  assign n14426 = ( ~n14418 & n14424 ) | ( ~n14418 & n14425 ) | ( n14424 & n14425 ) ;
  assign n14427 = n3715 & n5977 ;
  assign n14428 = x115 & n3719 ;
  assign n14429 = x116 | n14428 ;
  assign n14430 = ( n3721 & n14428 ) | ( n3721 & n14429 ) | ( n14428 & n14429 ) ;
  assign n14431 = x114 & n3922 ;
  assign n14432 = n14430 | n14431 ;
  assign n14433 = ( x41 & n14427 ) | ( x41 & ~n14432 ) | ( n14427 & ~n14432 ) ;
  assign n14434 = ( ~x41 & n14432 ) | ( ~x41 & n14433 ) | ( n14432 & n14433 ) ;
  assign n14435 = ( ~n14427 & n14433 ) | ( ~n14427 & n14434 ) | ( n14433 & n14434 ) ;
  assign n14436 = n4227 & n5542 ;
  assign n14437 = x112 & n4231 ;
  assign n14438 = x113 | n14437 ;
  assign n14439 = ( n4233 & n14437 ) | ( n4233 & n14438 ) | ( n14437 & n14438 ) ;
  assign n14440 = x111 & n4470 ;
  assign n14441 = n14439 | n14440 ;
  assign n14442 = ( x44 & n14436 ) | ( x44 & ~n14441 ) | ( n14436 & ~n14441 ) ;
  assign n14443 = ( ~x44 & n14441 ) | ( ~x44 & n14442 ) | ( n14441 & n14442 ) ;
  assign n14444 = ( ~n14436 & n14442 ) | ( ~n14436 & n14443 ) | ( n14442 & n14443 ) ;
  assign n14445 = n4787 & n4934 ;
  assign n14446 = x109 & n4791 ;
  assign n14447 = x110 | n14446 ;
  assign n14448 = ( n4793 & n14446 ) | ( n4793 & n14447 ) | ( n14446 & n14447 ) ;
  assign n14449 = x108 & n5030 ;
  assign n14450 = n14448 | n14449 ;
  assign n14451 = ( x47 & n14445 ) | ( x47 & ~n14450 ) | ( n14445 & ~n14450 ) ;
  assign n14452 = ( ~x47 & n14450 ) | ( ~x47 & n14451 ) | ( n14450 & n14451 ) ;
  assign n14453 = ( ~n14445 & n14451 ) | ( ~n14445 & n14452 ) | ( n14451 & n14452 ) ;
  assign n14454 = n4362 & n5374 ;
  assign n14455 = x106 & n5378 ;
  assign n14456 = x107 | n14455 ;
  assign n14457 = ( n5380 & n14455 ) | ( n5380 & n14456 ) | ( n14455 & n14456 ) ;
  assign n14458 = x105 & n5638 ;
  assign n14459 = n14457 | n14458 ;
  assign n14460 = ( x50 & n14454 ) | ( x50 & ~n14459 ) | ( n14454 & ~n14459 ) ;
  assign n14461 = ( ~x50 & n14459 ) | ( ~x50 & n14460 ) | ( n14459 & n14460 ) ;
  assign n14462 = ( ~n14454 & n14460 ) | ( ~n14454 & n14461 ) | ( n14460 & n14461 ) ;
  assign n14463 = n3665 & n6027 ;
  assign n14464 = x103 & n6031 ;
  assign n14465 = x104 | n14464 ;
  assign n14466 = ( n6033 & n14464 ) | ( n6033 & n14465 ) | ( n14464 & n14465 ) ;
  assign n14467 = x102 & n6303 ;
  assign n14468 = n14466 | n14467 ;
  assign n14469 = ( x53 & n14463 ) | ( x53 & ~n14468 ) | ( n14463 & ~n14468 ) ;
  assign n14470 = ( ~x53 & n14468 ) | ( ~x53 & n14469 ) | ( n14468 & n14469 ) ;
  assign n14471 = ( ~n14463 & n14469 ) | ( ~n14463 & n14470 ) | ( n14469 & n14470 ) ;
  assign n14472 = n3326 & n6713 ;
  assign n14473 = x100 & n6717 ;
  assign n14474 = x101 | n14473 ;
  assign n14475 = ( n6719 & n14473 ) | ( n6719 & n14474 ) | ( n14473 & n14474 ) ;
  assign n14476 = x99 & n6980 ;
  assign n14477 = n14475 | n14476 ;
  assign n14478 = ( x56 & n14472 ) | ( x56 & ~n14477 ) | ( n14472 & ~n14477 ) ;
  assign n14479 = ( ~x56 & n14477 ) | ( ~x56 & n14478 ) | ( n14477 & n14478 ) ;
  assign n14480 = ( ~n14472 & n14478 ) | ( ~n14472 & n14479 ) | ( n14478 & n14479 ) ;
  assign n14481 = n2434 & n8154 ;
  assign n14482 = x94 & n8158 ;
  assign n14483 = x95 | n14482 ;
  assign n14484 = ( n8160 & n14482 ) | ( n8160 & n14483 ) | ( n14482 & n14483 ) ;
  assign n14485 = x93 & n8439 ;
  assign n14486 = n14484 | n14485 ;
  assign n14487 = ( x62 & n14481 ) | ( x62 & ~n14486 ) | ( n14481 & ~n14486 ) ;
  assign n14488 = ( ~x62 & n14486 ) | ( ~x62 & n14487 ) | ( n14486 & n14487 ) ;
  assign n14489 = ( ~n14481 & n14487 ) | ( ~n14481 & n14488 ) | ( n14487 & n14488 ) ;
  assign n14490 = x91 & n8927 ;
  assign n14491 = ( ~x92 & n8693 ) | ( ~x92 & n8927 ) | ( n8693 & n8927 ) ;
  assign n14492 = ( n8693 & n14490 ) | ( n8693 & ~n14491 ) | ( n14490 & ~n14491 ) ;
  assign n14493 = ( ~n14333 & n14489 ) | ( ~n14333 & n14492 ) | ( n14489 & n14492 ) ;
  assign n14494 = ( n14489 & n14492 ) | ( n14489 & ~n14493 ) | ( n14492 & ~n14493 ) ;
  assign n14495 = ( n14333 & n14493 ) | ( n14333 & ~n14494 ) | ( n14493 & ~n14494 ) ;
  assign n14496 = n2725 & n7423 ;
  assign n14497 = x97 & n7427 ;
  assign n14498 = x98 | n14497 ;
  assign n14499 = ( n7429 & n14497 ) | ( n7429 & n14498 ) | ( n14497 & n14498 ) ;
  assign n14500 = x96 & n7708 ;
  assign n14501 = n14499 | n14500 ;
  assign n14502 = ( x59 & n14496 ) | ( x59 & ~n14501 ) | ( n14496 & ~n14501 ) ;
  assign n14503 = ( ~x59 & n14501 ) | ( ~x59 & n14502 ) | ( n14501 & n14502 ) ;
  assign n14504 = ( ~n14496 & n14502 ) | ( ~n14496 & n14503 ) | ( n14502 & n14503 ) ;
  assign n14505 = ( n14336 & ~n14495 ) | ( n14336 & n14504 ) | ( ~n14495 & n14504 ) ;
  assign n14506 = ( n14336 & n14495 ) | ( n14336 & n14504 ) | ( n14495 & n14504 ) ;
  assign n14507 = ( n14495 & n14505 ) | ( n14495 & ~n14506 ) | ( n14505 & ~n14506 ) ;
  assign n14508 = ( n14339 & n14480 ) | ( n14339 & ~n14507 ) | ( n14480 & ~n14507 ) ;
  assign n14509 = ( ~n14339 & n14480 ) | ( ~n14339 & n14507 ) | ( n14480 & n14507 ) ;
  assign n14510 = ( ~n14480 & n14508 ) | ( ~n14480 & n14509 ) | ( n14508 & n14509 ) ;
  assign n14511 = ( n14342 & n14471 ) | ( n14342 & ~n14510 ) | ( n14471 & ~n14510 ) ;
  assign n14512 = ( ~n14342 & n14471 ) | ( ~n14342 & n14510 ) | ( n14471 & n14510 ) ;
  assign n14513 = ( ~n14471 & n14511 ) | ( ~n14471 & n14512 ) | ( n14511 & n14512 ) ;
  assign n14514 = ( n14345 & n14462 ) | ( n14345 & ~n14513 ) | ( n14462 & ~n14513 ) ;
  assign n14515 = ( ~n14345 & n14462 ) | ( ~n14345 & n14513 ) | ( n14462 & n14513 ) ;
  assign n14516 = ( ~n14462 & n14514 ) | ( ~n14462 & n14515 ) | ( n14514 & n14515 ) ;
  assign n14517 = ( n14348 & n14453 ) | ( n14348 & ~n14516 ) | ( n14453 & ~n14516 ) ;
  assign n14518 = ( ~n14348 & n14453 ) | ( ~n14348 & n14516 ) | ( n14453 & n14516 ) ;
  assign n14519 = ( ~n14453 & n14517 ) | ( ~n14453 & n14518 ) | ( n14517 & n14518 ) ;
  assign n14520 = ( n14351 & n14444 ) | ( n14351 & ~n14519 ) | ( n14444 & ~n14519 ) ;
  assign n14521 = ( ~n14351 & n14444 ) | ( ~n14351 & n14519 ) | ( n14444 & n14519 ) ;
  assign n14522 = ( ~n14444 & n14520 ) | ( ~n14444 & n14521 ) | ( n14520 & n14521 ) ;
  assign n14523 = ( n14354 & n14435 ) | ( n14354 & ~n14522 ) | ( n14435 & ~n14522 ) ;
  assign n14524 = ( ~n14354 & n14435 ) | ( ~n14354 & n14522 ) | ( n14435 & n14522 ) ;
  assign n14525 = ( ~n14435 & n14523 ) | ( ~n14435 & n14524 ) | ( n14523 & n14524 ) ;
  assign n14526 = ( n14357 & n14426 ) | ( n14357 & ~n14525 ) | ( n14426 & ~n14525 ) ;
  assign n14527 = ( ~n14357 & n14426 ) | ( ~n14357 & n14525 ) | ( n14426 & n14525 ) ;
  assign n14528 = ( ~n14426 & n14526 ) | ( ~n14426 & n14527 ) | ( n14526 & n14527 ) ;
  assign n14529 = ( n14360 & n14417 ) | ( n14360 & ~n14528 ) | ( n14417 & ~n14528 ) ;
  assign n14530 = ( ~n14360 & n14417 ) | ( ~n14360 & n14528 ) | ( n14417 & n14528 ) ;
  assign n14531 = ( ~n14417 & n14529 ) | ( ~n14417 & n14530 ) | ( n14529 & n14530 ) ;
  assign n14532 = ( n14363 & n14408 ) | ( n14363 & ~n14531 ) | ( n14408 & ~n14531 ) ;
  assign n14533 = ( ~n14363 & n14408 ) | ( ~n14363 & n14531 ) | ( n14408 & n14531 ) ;
  assign n14534 = ( ~n14408 & n14532 ) | ( ~n14408 & n14533 ) | ( n14532 & n14533 ) ;
  assign n14535 = ( n14375 & n14399 ) | ( n14375 & ~n14534 ) | ( n14399 & ~n14534 ) ;
  assign n14536 = ( ~n14375 & n14399 ) | ( ~n14375 & n14534 ) | ( n14399 & n14534 ) ;
  assign n14537 = ( ~n14399 & n14535 ) | ( ~n14399 & n14536 ) | ( n14535 & n14536 ) ;
  assign n14538 = ( ~n14387 & n14390 ) | ( ~n14387 & n14537 ) | ( n14390 & n14537 ) ;
  assign n14539 = ( n14390 & n14537 ) | ( n14390 & ~n14538 ) | ( n14537 & ~n14538 ) ;
  assign n14540 = ( n14387 & n14538 ) | ( n14387 & ~n14539 ) | ( n14538 & ~n14539 ) ;
  assign n14541 = n2320 & n8587 ;
  assign n14542 = x125 & n2324 ;
  assign n14543 = x126 | n14542 ;
  assign n14544 = ( n2326 & n14542 ) | ( n2326 & n14543 ) | ( n14542 & n14543 ) ;
  assign n14545 = x124 & n2497 ;
  assign n14546 = n14544 | n14545 ;
  assign n14547 = ( x32 & n14541 ) | ( x32 & ~n14546 ) | ( n14541 & ~n14546 ) ;
  assign n14548 = ( ~x32 & n14546 ) | ( ~x32 & n14547 ) | ( n14546 & n14547 ) ;
  assign n14549 = ( ~n14541 & n14547 ) | ( ~n14541 & n14548 ) | ( n14547 & n14548 ) ;
  assign n14550 = n2766 & n7597 ;
  assign n14551 = x122 & n2770 ;
  assign n14552 = x123 | n14551 ;
  assign n14553 = ( n2772 & n14551 ) | ( n2772 & n14552 ) | ( n14551 & n14552 ) ;
  assign n14554 = x121 & n2943 ;
  assign n14555 = n14553 | n14554 ;
  assign n14556 = ( x35 & n14550 ) | ( x35 & ~n14555 ) | ( n14550 & ~n14555 ) ;
  assign n14557 = ( ~x35 & n14555 ) | ( ~x35 & n14556 ) | ( n14555 & n14556 ) ;
  assign n14558 = ( ~n14550 & n14556 ) | ( ~n14550 & n14557 ) | ( n14556 & n14557 ) ;
  assign n14559 = n3224 & n7098 ;
  assign n14560 = x119 & n3228 ;
  assign n14561 = x120 | n14560 ;
  assign n14562 = ( n3230 & n14560 ) | ( n3230 & n14561 ) | ( n14560 & n14561 ) ;
  assign n14563 = x118 & n3413 ;
  assign n14564 = n14562 | n14563 ;
  assign n14565 = ( x38 & n14559 ) | ( x38 & ~n14564 ) | ( n14559 & ~n14564 ) ;
  assign n14566 = ( ~x38 & n14564 ) | ( ~x38 & n14565 ) | ( n14564 & n14565 ) ;
  assign n14567 = ( ~n14559 & n14565 ) | ( ~n14559 & n14566 ) | ( n14565 & n14566 ) ;
  assign n14568 = n3715 & n6201 ;
  assign n14569 = x116 & n3719 ;
  assign n14570 = x117 | n14569 ;
  assign n14571 = ( n3721 & n14569 ) | ( n3721 & n14570 ) | ( n14569 & n14570 ) ;
  assign n14572 = x115 & n3922 ;
  assign n14573 = n14571 | n14572 ;
  assign n14574 = ( x41 & n14568 ) | ( x41 & ~n14573 ) | ( n14568 & ~n14573 ) ;
  assign n14575 = ( ~x41 & n14573 ) | ( ~x41 & n14574 ) | ( n14573 & n14574 ) ;
  assign n14576 = ( ~n14568 & n14574 ) | ( ~n14568 & n14575 ) | ( n14574 & n14575 ) ;
  assign n14577 = n4227 & n5750 ;
  assign n14578 = x113 & n4231 ;
  assign n14579 = x114 | n14578 ;
  assign n14580 = ( n4233 & n14578 ) | ( n4233 & n14579 ) | ( n14578 & n14579 ) ;
  assign n14581 = x112 & n4470 ;
  assign n14582 = n14580 | n14581 ;
  assign n14583 = ( x44 & n14577 ) | ( x44 & ~n14582 ) | ( n14577 & ~n14582 ) ;
  assign n14584 = ( ~x44 & n14582 ) | ( ~x44 & n14583 ) | ( n14582 & n14583 ) ;
  assign n14585 = ( ~n14577 & n14583 ) | ( ~n14577 & n14584 ) | ( n14583 & n14584 ) ;
  assign n14586 = n4787 & n5130 ;
  assign n14587 = x110 & n4791 ;
  assign n14588 = x111 | n14587 ;
  assign n14589 = ( n4793 & n14587 ) | ( n4793 & n14588 ) | ( n14587 & n14588 ) ;
  assign n14590 = x109 & n5030 ;
  assign n14591 = n14589 | n14590 ;
  assign n14592 = ( x47 & n14586 ) | ( x47 & ~n14591 ) | ( n14586 & ~n14591 ) ;
  assign n14593 = ( ~x47 & n14591 ) | ( ~x47 & n14592 ) | ( n14591 & n14592 ) ;
  assign n14594 = ( ~n14586 & n14592 ) | ( ~n14586 & n14593 ) | ( n14592 & n14593 ) ;
  assign n14595 = n4377 & n5374 ;
  assign n14596 = x107 & n5378 ;
  assign n14597 = x108 | n14596 ;
  assign n14598 = ( n5380 & n14596 ) | ( n5380 & n14597 ) | ( n14596 & n14597 ) ;
  assign n14599 = x106 & n5638 ;
  assign n14600 = n14598 | n14599 ;
  assign n14601 = ( x50 & n14595 ) | ( x50 & ~n14600 ) | ( n14595 & ~n14600 ) ;
  assign n14602 = ( ~x50 & n14600 ) | ( ~x50 & n14601 ) | ( n14600 & n14601 ) ;
  assign n14603 = ( ~n14595 & n14601 ) | ( ~n14595 & n14602 ) | ( n14601 & n14602 ) ;
  assign n14604 = n3998 & n6027 ;
  assign n14605 = x104 & n6031 ;
  assign n14606 = x105 | n14605 ;
  assign n14607 = ( n6033 & n14605 ) | ( n6033 & n14606 ) | ( n14605 & n14606 ) ;
  assign n14608 = x103 & n6303 ;
  assign n14609 = n14607 | n14608 ;
  assign n14610 = ( x53 & n14604 ) | ( x53 & ~n14609 ) | ( n14604 & ~n14609 ) ;
  assign n14611 = ( ~x53 & n14609 ) | ( ~x53 & n14610 ) | ( n14609 & n14610 ) ;
  assign n14612 = ( ~n14604 & n14610 ) | ( ~n14604 & n14611 ) | ( n14610 & n14611 ) ;
  assign n14613 = x92 & n8927 ;
  assign n14614 = ( ~x93 & n8693 ) | ( ~x93 & n8927 ) | ( n8693 & n8927 ) ;
  assign n14615 = ( n8693 & n14613 ) | ( n8693 & ~n14614 ) | ( n14613 & ~n14614 ) ;
  assign n14616 = ( n14333 & n14493 ) | ( n14333 & ~n14615 ) | ( n14493 & ~n14615 ) ;
  assign n14617 = ( n14333 & ~n14493 ) | ( n14333 & n14615 ) | ( ~n14493 & n14615 ) ;
  assign n14618 = ( ~n14333 & n14616 ) | ( ~n14333 & n14617 ) | ( n14616 & n14617 ) ;
  assign n14619 = n2877 & n7423 ;
  assign n14620 = x98 & n7427 ;
  assign n14621 = x99 | n14620 ;
  assign n14622 = ( n7429 & n14620 ) | ( n7429 & n14621 ) | ( n14620 & n14621 ) ;
  assign n14623 = x97 & n7708 ;
  assign n14624 = n14622 | n14623 ;
  assign n14625 = ( x59 & n14619 ) | ( x59 & ~n14624 ) | ( n14619 & ~n14624 ) ;
  assign n14626 = ( ~x59 & n14624 ) | ( ~x59 & n14625 ) | ( n14624 & n14625 ) ;
  assign n14627 = ( ~n14619 & n14625 ) | ( ~n14619 & n14626 ) | ( n14625 & n14626 ) ;
  assign n14628 = n2449 & n8154 ;
  assign n14629 = x95 & n8158 ;
  assign n14630 = x96 | n14629 ;
  assign n14631 = ( n8160 & n14629 ) | ( n8160 & n14630 ) | ( n14629 & n14630 ) ;
  assign n14632 = x94 & n8439 ;
  assign n14633 = n14631 | n14632 ;
  assign n14634 = ( x62 & n14628 ) | ( x62 & ~n14633 ) | ( n14628 & ~n14633 ) ;
  assign n14635 = ( ~x62 & n14633 ) | ( ~x62 & n14634 ) | ( n14633 & n14634 ) ;
  assign n14636 = ( ~n14628 & n14634 ) | ( ~n14628 & n14635 ) | ( n14634 & n14635 ) ;
  assign n14637 = ( ~n14618 & n14627 ) | ( ~n14618 & n14636 ) | ( n14627 & n14636 ) ;
  assign n14638 = ( n14627 & n14636 ) | ( n14627 & ~n14637 ) | ( n14636 & ~n14637 ) ;
  assign n14639 = ( n14618 & n14637 ) | ( n14618 & ~n14638 ) | ( n14637 & ~n14638 ) ;
  assign n14640 = n3486 & n6713 ;
  assign n14641 = x101 & n6717 ;
  assign n14642 = x102 | n14641 ;
  assign n14643 = ( n6719 & n14641 ) | ( n6719 & n14642 ) | ( n14641 & n14642 ) ;
  assign n14644 = x100 & n6980 ;
  assign n14645 = n14643 | n14644 ;
  assign n14646 = ( x56 & n14640 ) | ( x56 & ~n14645 ) | ( n14640 & ~n14645 ) ;
  assign n14647 = ( ~x56 & n14645 ) | ( ~x56 & n14646 ) | ( n14645 & n14646 ) ;
  assign n14648 = ( ~n14640 & n14646 ) | ( ~n14640 & n14647 ) | ( n14646 & n14647 ) ;
  assign n14649 = ( n14505 & ~n14639 ) | ( n14505 & n14648 ) | ( ~n14639 & n14648 ) ;
  assign n14650 = ( n14505 & n14639 ) | ( n14505 & n14648 ) | ( n14639 & n14648 ) ;
  assign n14651 = ( n14639 & n14649 ) | ( n14639 & ~n14650 ) | ( n14649 & ~n14650 ) ;
  assign n14652 = ( n14508 & n14612 ) | ( n14508 & ~n14651 ) | ( n14612 & ~n14651 ) ;
  assign n14653 = ( ~n14508 & n14612 ) | ( ~n14508 & n14651 ) | ( n14612 & n14651 ) ;
  assign n14654 = ( ~n14612 & n14652 ) | ( ~n14612 & n14653 ) | ( n14652 & n14653 ) ;
  assign n14655 = ( n14511 & n14603 ) | ( n14511 & ~n14654 ) | ( n14603 & ~n14654 ) ;
  assign n14656 = ( ~n14511 & n14603 ) | ( ~n14511 & n14654 ) | ( n14603 & n14654 ) ;
  assign n14657 = ( ~n14603 & n14655 ) | ( ~n14603 & n14656 ) | ( n14655 & n14656 ) ;
  assign n14658 = ( n14514 & n14594 ) | ( n14514 & ~n14657 ) | ( n14594 & ~n14657 ) ;
  assign n14659 = ( ~n14514 & n14594 ) | ( ~n14514 & n14657 ) | ( n14594 & n14657 ) ;
  assign n14660 = ( ~n14594 & n14658 ) | ( ~n14594 & n14659 ) | ( n14658 & n14659 ) ;
  assign n14661 = ( n14517 & n14585 ) | ( n14517 & ~n14660 ) | ( n14585 & ~n14660 ) ;
  assign n14662 = ( ~n14517 & n14585 ) | ( ~n14517 & n14660 ) | ( n14585 & n14660 ) ;
  assign n14663 = ( ~n14585 & n14661 ) | ( ~n14585 & n14662 ) | ( n14661 & n14662 ) ;
  assign n14664 = ( n14520 & n14576 ) | ( n14520 & ~n14663 ) | ( n14576 & ~n14663 ) ;
  assign n14665 = ( ~n14520 & n14576 ) | ( ~n14520 & n14663 ) | ( n14576 & n14663 ) ;
  assign n14666 = ( ~n14576 & n14664 ) | ( ~n14576 & n14665 ) | ( n14664 & n14665 ) ;
  assign n14667 = ( n14523 & n14567 ) | ( n14523 & ~n14666 ) | ( n14567 & ~n14666 ) ;
  assign n14668 = ( ~n14523 & n14567 ) | ( ~n14523 & n14666 ) | ( n14567 & n14666 ) ;
  assign n14669 = ( ~n14567 & n14667 ) | ( ~n14567 & n14668 ) | ( n14667 & n14668 ) ;
  assign n14670 = ( n14526 & n14558 ) | ( n14526 & ~n14669 ) | ( n14558 & ~n14669 ) ;
  assign n14671 = ( ~n14526 & n14558 ) | ( ~n14526 & n14669 ) | ( n14558 & n14669 ) ;
  assign n14672 = ( ~n14558 & n14670 ) | ( ~n14558 & n14671 ) | ( n14670 & n14671 ) ;
  assign n14673 = ( n14529 & n14549 ) | ( n14529 & ~n14672 ) | ( n14549 & ~n14672 ) ;
  assign n14674 = ( ~n14529 & n14549 ) | ( ~n14529 & n14672 ) | ( n14549 & n14672 ) ;
  assign n14675 = ( ~n14549 & n14673 ) | ( ~n14549 & n14674 ) | ( n14673 & n14674 ) ;
  assign n14676 = n1949 & n8862 ;
  assign n14677 = ( x127 & n2114 ) | ( x127 & n14676 ) | ( n2114 & n14676 ) ;
  assign n14678 = x29 | n14677 ;
  assign n14679 = ~x29 & n14677 ;
  assign n14680 = ( ~n14677 & n14678 ) | ( ~n14677 & n14679 ) | ( n14678 & n14679 ) ;
  assign n14681 = ( n14532 & ~n14675 ) | ( n14532 & n14680 ) | ( ~n14675 & n14680 ) ;
  assign n14682 = ( n14532 & n14675 ) | ( n14532 & n14680 ) | ( n14675 & n14680 ) ;
  assign n14683 = ( n14675 & n14681 ) | ( n14675 & ~n14682 ) | ( n14681 & ~n14682 ) ;
  assign n14684 = ( ~n14535 & n14538 ) | ( ~n14535 & n14683 ) | ( n14538 & n14683 ) ;
  assign n14685 = ( n14538 & n14683 ) | ( n14538 & ~n14684 ) | ( n14683 & ~n14684 ) ;
  assign n14686 = ( n14535 & n14684 ) | ( n14535 & ~n14685 ) | ( n14684 & ~n14685 ) ;
  assign n14687 = n2766 & n7841 ;
  assign n14688 = x123 & n2770 ;
  assign n14689 = x124 | n14688 ;
  assign n14690 = ( n2772 & n14688 ) | ( n2772 & n14689 ) | ( n14688 & n14689 ) ;
  assign n14691 = x122 & n2943 ;
  assign n14692 = n14690 | n14691 ;
  assign n14693 = ( x35 & n14687 ) | ( x35 & ~n14692 ) | ( n14687 & ~n14692 ) ;
  assign n14694 = ( ~x35 & n14692 ) | ( ~x35 & n14693 ) | ( n14692 & n14693 ) ;
  assign n14695 = ( ~n14687 & n14693 ) | ( ~n14687 & n14694 ) | ( n14693 & n14694 ) ;
  assign n14696 = n3224 & n7113 ;
  assign n14697 = x120 & n3228 ;
  assign n14698 = x121 | n14697 ;
  assign n14699 = ( n3230 & n14697 ) | ( n3230 & n14698 ) | ( n14697 & n14698 ) ;
  assign n14700 = x119 & n3413 ;
  assign n14701 = n14699 | n14700 ;
  assign n14702 = ( x38 & n14696 ) | ( x38 & ~n14701 ) | ( n14696 & ~n14701 ) ;
  assign n14703 = ( ~x38 & n14701 ) | ( ~x38 & n14702 ) | ( n14701 & n14702 ) ;
  assign n14704 = ( ~n14696 & n14702 ) | ( ~n14696 & n14703 ) | ( n14702 & n14703 ) ;
  assign n14705 = n3715 & n6421 ;
  assign n14706 = x117 & n3719 ;
  assign n14707 = x118 | n14706 ;
  assign n14708 = ( n3721 & n14706 ) | ( n3721 & n14707 ) | ( n14706 & n14707 ) ;
  assign n14709 = x116 & n3922 ;
  assign n14710 = n14708 | n14709 ;
  assign n14711 = ( x41 & n14705 ) | ( x41 & ~n14710 ) | ( n14705 & ~n14710 ) ;
  assign n14712 = ( ~x41 & n14710 ) | ( ~x41 & n14711 ) | ( n14710 & n14711 ) ;
  assign n14713 = ( ~n14705 & n14711 ) | ( ~n14705 & n14712 ) | ( n14711 & n14712 ) ;
  assign n14714 = n4227 & n5765 ;
  assign n14715 = x114 & n4231 ;
  assign n14716 = x115 | n14715 ;
  assign n14717 = ( n4233 & n14715 ) | ( n4233 & n14716 ) | ( n14715 & n14716 ) ;
  assign n14718 = x113 & n4470 ;
  assign n14719 = n14717 | n14718 ;
  assign n14720 = ( x44 & n14714 ) | ( x44 & ~n14719 ) | ( n14714 & ~n14719 ) ;
  assign n14721 = ( ~x44 & n14719 ) | ( ~x44 & n14720 ) | ( n14719 & n14720 ) ;
  assign n14722 = ( ~n14714 & n14720 ) | ( ~n14714 & n14721 ) | ( n14720 & n14721 ) ;
  assign n14723 = n4787 & n5145 ;
  assign n14724 = x111 & n4791 ;
  assign n14725 = x112 | n14724 ;
  assign n14726 = ( n4793 & n14724 ) | ( n4793 & n14725 ) | ( n14724 & n14725 ) ;
  assign n14727 = x110 & n5030 ;
  assign n14728 = n14726 | n14727 ;
  assign n14729 = ( x47 & n14723 ) | ( x47 & ~n14728 ) | ( n14723 & ~n14728 ) ;
  assign n14730 = ( ~x47 & n14728 ) | ( ~x47 & n14729 ) | ( n14728 & n14729 ) ;
  assign n14731 = ( ~n14723 & n14729 ) | ( ~n14723 & n14730 ) | ( n14729 & n14730 ) ;
  assign n14732 = n4734 & n5374 ;
  assign n14733 = x108 & n5378 ;
  assign n14734 = x109 | n14733 ;
  assign n14735 = ( n5380 & n14733 ) | ( n5380 & n14734 ) | ( n14733 & n14734 ) ;
  assign n14736 = x107 & n5638 ;
  assign n14737 = n14735 | n14736 ;
  assign n14738 = ( x50 & n14732 ) | ( x50 & ~n14737 ) | ( n14732 & ~n14737 ) ;
  assign n14739 = ( ~x50 & n14737 ) | ( ~x50 & n14738 ) | ( n14737 & n14738 ) ;
  assign n14740 = ( ~n14732 & n14738 ) | ( ~n14732 & n14739 ) | ( n14738 & n14739 ) ;
  assign n14741 = n4013 & n6027 ;
  assign n14742 = x105 & n6031 ;
  assign n14743 = x106 | n14742 ;
  assign n14744 = ( n6033 & n14742 ) | ( n6033 & n14743 ) | ( n14742 & n14743 ) ;
  assign n14745 = x104 & n6303 ;
  assign n14746 = n14744 | n14745 ;
  assign n14747 = ( x53 & n14741 ) | ( x53 & ~n14746 ) | ( n14741 & ~n14746 ) ;
  assign n14748 = ( ~x53 & n14746 ) | ( ~x53 & n14747 ) | ( n14746 & n14747 ) ;
  assign n14749 = ( ~n14741 & n14747 ) | ( ~n14741 & n14748 ) | ( n14747 & n14748 ) ;
  assign n14750 = n3650 & n6713 ;
  assign n14751 = x102 & n6717 ;
  assign n14752 = x103 | n14751 ;
  assign n14753 = ( n6719 & n14751 ) | ( n6719 & n14752 ) | ( n14751 & n14752 ) ;
  assign n14754 = x101 & n6980 ;
  assign n14755 = n14753 | n14754 ;
  assign n14756 = ( x56 & n14750 ) | ( x56 & ~n14755 ) | ( n14750 & ~n14755 ) ;
  assign n14757 = ( ~x56 & n14755 ) | ( ~x56 & n14756 ) | ( n14755 & n14756 ) ;
  assign n14758 = ( ~n14750 & n14756 ) | ( ~n14750 & n14757 ) | ( n14756 & n14757 ) ;
  assign n14759 = n3162 & n7423 ;
  assign n14760 = x99 & n7427 ;
  assign n14761 = x100 | n14760 ;
  assign n14762 = ( n7429 & n14760 ) | ( n7429 & n14761 ) | ( n14760 & n14761 ) ;
  assign n14763 = x98 & n7708 ;
  assign n14764 = n14762 | n14763 ;
  assign n14765 = ( x59 & n14759 ) | ( x59 & ~n14764 ) | ( n14759 & ~n14764 ) ;
  assign n14766 = ( ~x59 & n14764 ) | ( ~x59 & n14765 ) | ( n14764 & n14765 ) ;
  assign n14767 = ( ~n14759 & n14765 ) | ( ~n14759 & n14766 ) | ( n14765 & n14766 ) ;
  assign n14768 = n2585 & n8154 ;
  assign n14769 = x96 & n8158 ;
  assign n14770 = x97 | n14769 ;
  assign n14771 = ( n8160 & n14769 ) | ( n8160 & n14770 ) | ( n14769 & n14770 ) ;
  assign n14772 = x95 & n8439 ;
  assign n14773 = n14771 | n14772 ;
  assign n14774 = ( x62 & n14768 ) | ( x62 & ~n14773 ) | ( n14768 & ~n14773 ) ;
  assign n14775 = ( ~x62 & n14773 ) | ( ~x62 & n14774 ) | ( n14773 & n14774 ) ;
  assign n14776 = ( ~n14768 & n14774 ) | ( ~n14768 & n14775 ) | ( n14774 & n14775 ) ;
  assign n14777 = x93 & n8927 ;
  assign n14778 = ( ~x94 & n8693 ) | ( ~x94 & n8927 ) | ( n8693 & n8927 ) ;
  assign n14779 = ( n8693 & n14777 ) | ( n8693 & ~n14778 ) | ( n14777 & ~n14778 ) ;
  assign n14780 = ( ~x29 & n14615 ) | ( ~x29 & n14779 ) | ( n14615 & n14779 ) ;
  assign n14781 = ( n14615 & n14779 ) | ( n14615 & ~n14780 ) | ( n14779 & ~n14780 ) ;
  assign n14782 = ( x29 & n14780 ) | ( x29 & ~n14781 ) | ( n14780 & ~n14781 ) ;
  assign n14783 = ( n14616 & n14776 ) | ( n14616 & ~n14782 ) | ( n14776 & ~n14782 ) ;
  assign n14784 = ( ~n14616 & n14776 ) | ( ~n14616 & n14782 ) | ( n14776 & n14782 ) ;
  assign n14785 = ( ~n14776 & n14783 ) | ( ~n14776 & n14784 ) | ( n14783 & n14784 ) ;
  assign n14786 = ( n14637 & n14767 ) | ( n14637 & ~n14785 ) | ( n14767 & ~n14785 ) ;
  assign n14787 = ( ~n14637 & n14767 ) | ( ~n14637 & n14785 ) | ( n14767 & n14785 ) ;
  assign n14788 = ( ~n14767 & n14786 ) | ( ~n14767 & n14787 ) | ( n14786 & n14787 ) ;
  assign n14789 = ( n14649 & n14758 ) | ( n14649 & ~n14788 ) | ( n14758 & ~n14788 ) ;
  assign n14790 = ( ~n14649 & n14758 ) | ( ~n14649 & n14788 ) | ( n14758 & n14788 ) ;
  assign n14791 = ( ~n14758 & n14789 ) | ( ~n14758 & n14790 ) | ( n14789 & n14790 ) ;
  assign n14792 = ( n14652 & n14749 ) | ( n14652 & ~n14791 ) | ( n14749 & ~n14791 ) ;
  assign n14793 = ( ~n14652 & n14749 ) | ( ~n14652 & n14791 ) | ( n14749 & n14791 ) ;
  assign n14794 = ( ~n14749 & n14792 ) | ( ~n14749 & n14793 ) | ( n14792 & n14793 ) ;
  assign n14795 = ( n14655 & n14740 ) | ( n14655 & ~n14794 ) | ( n14740 & ~n14794 ) ;
  assign n14796 = ( ~n14655 & n14740 ) | ( ~n14655 & n14794 ) | ( n14740 & n14794 ) ;
  assign n14797 = ( ~n14740 & n14795 ) | ( ~n14740 & n14796 ) | ( n14795 & n14796 ) ;
  assign n14798 = ( n14658 & n14731 ) | ( n14658 & ~n14797 ) | ( n14731 & ~n14797 ) ;
  assign n14799 = ( ~n14658 & n14731 ) | ( ~n14658 & n14797 ) | ( n14731 & n14797 ) ;
  assign n14800 = ( ~n14731 & n14798 ) | ( ~n14731 & n14799 ) | ( n14798 & n14799 ) ;
  assign n14801 = ( n14661 & n14722 ) | ( n14661 & ~n14800 ) | ( n14722 & ~n14800 ) ;
  assign n14802 = ( ~n14661 & n14722 ) | ( ~n14661 & n14800 ) | ( n14722 & n14800 ) ;
  assign n14803 = ( ~n14722 & n14801 ) | ( ~n14722 & n14802 ) | ( n14801 & n14802 ) ;
  assign n14804 = ( n14664 & n14713 ) | ( n14664 & ~n14803 ) | ( n14713 & ~n14803 ) ;
  assign n14805 = ( ~n14664 & n14713 ) | ( ~n14664 & n14803 ) | ( n14713 & n14803 ) ;
  assign n14806 = ( ~n14713 & n14804 ) | ( ~n14713 & n14805 ) | ( n14804 & n14805 ) ;
  assign n14807 = ( n14667 & n14704 ) | ( n14667 & ~n14806 ) | ( n14704 & ~n14806 ) ;
  assign n14808 = ( ~n14667 & n14704 ) | ( ~n14667 & n14806 ) | ( n14704 & n14806 ) ;
  assign n14809 = ( ~n14704 & n14807 ) | ( ~n14704 & n14808 ) | ( n14807 & n14808 ) ;
  assign n14810 = ( n14670 & n14695 ) | ( n14670 & ~n14809 ) | ( n14695 & ~n14809 ) ;
  assign n14811 = ( ~n14670 & n14695 ) | ( ~n14670 & n14809 ) | ( n14695 & n14809 ) ;
  assign n14812 = ( ~n14695 & n14810 ) | ( ~n14695 & n14811 ) | ( n14810 & n14811 ) ;
  assign n14813 = n2320 & n8846 ;
  assign n14814 = x126 & n2324 ;
  assign n14815 = x127 | n14814 ;
  assign n14816 = ( n2326 & n14814 ) | ( n2326 & n14815 ) | ( n14814 & n14815 ) ;
  assign n14817 = x125 & n2497 ;
  assign n14818 = n14816 | n14817 ;
  assign n14819 = ( x32 & n14813 ) | ( x32 & ~n14818 ) | ( n14813 & ~n14818 ) ;
  assign n14820 = ( ~x32 & n14818 ) | ( ~x32 & n14819 ) | ( n14818 & n14819 ) ;
  assign n14821 = ( ~n14813 & n14819 ) | ( ~n14813 & n14820 ) | ( n14819 & n14820 ) ;
  assign n14822 = ( n14673 & ~n14812 ) | ( n14673 & n14821 ) | ( ~n14812 & n14821 ) ;
  assign n14823 = ( n14673 & n14812 ) | ( n14673 & n14821 ) | ( n14812 & n14821 ) ;
  assign n14824 = ( n14812 & n14822 ) | ( n14812 & ~n14823 ) | ( n14822 & ~n14823 ) ;
  assign n14825 = ( ~n14681 & n14684 ) | ( ~n14681 & n14824 ) | ( n14684 & n14824 ) ;
  assign n14826 = ( n14684 & n14824 ) | ( n14684 & ~n14825 ) | ( n14824 & ~n14825 ) ;
  assign n14827 = ( n14681 & n14825 ) | ( n14681 & ~n14826 ) | ( n14825 & ~n14826 ) ;
  assign n14828 = n2320 & n8865 ;
  assign n14829 = x127 & n2324 ;
  assign n14830 = x126 | n14829 ;
  assign n14831 = ( n2497 & n14829 ) | ( n2497 & n14830 ) | ( n14829 & n14830 ) ;
  assign n14832 = ( x32 & n14828 ) | ( x32 & ~n14831 ) | ( n14828 & ~n14831 ) ;
  assign n14833 = ( ~x32 & n14831 ) | ( ~x32 & n14832 ) | ( n14831 & n14832 ) ;
  assign n14834 = ( ~n14828 & n14832 ) | ( ~n14828 & n14833 ) | ( n14832 & n14833 ) ;
  assign n14835 = n3224 & n7582 ;
  assign n14836 = x121 & n3228 ;
  assign n14837 = x122 | n14836 ;
  assign n14838 = ( n3230 & n14836 ) | ( n3230 & n14837 ) | ( n14836 & n14837 ) ;
  assign n14839 = x120 & n3413 ;
  assign n14840 = n14838 | n14839 ;
  assign n14841 = ( x38 & n14835 ) | ( x38 & ~n14840 ) | ( n14835 & ~n14840 ) ;
  assign n14842 = ( ~x38 & n14840 ) | ( ~x38 & n14841 ) | ( n14840 & n14841 ) ;
  assign n14843 = ( ~n14835 & n14841 ) | ( ~n14835 & n14842 ) | ( n14841 & n14842 ) ;
  assign n14844 = n3715 & n6645 ;
  assign n14845 = x118 & n3719 ;
  assign n14846 = x119 | n14845 ;
  assign n14847 = ( n3721 & n14845 ) | ( n3721 & n14846 ) | ( n14845 & n14846 ) ;
  assign n14848 = x117 & n3922 ;
  assign n14849 = n14847 | n14848 ;
  assign n14850 = ( x41 & n14844 ) | ( x41 & ~n14849 ) | ( n14844 & ~n14849 ) ;
  assign n14851 = ( ~x41 & n14849 ) | ( ~x41 & n14850 ) | ( n14849 & n14850 ) ;
  assign n14852 = ( ~n14844 & n14850 ) | ( ~n14844 & n14851 ) | ( n14850 & n14851 ) ;
  assign n14853 = n4227 & n5977 ;
  assign n14854 = x115 & n4231 ;
  assign n14855 = x116 | n14854 ;
  assign n14856 = ( n4233 & n14854 ) | ( n4233 & n14855 ) | ( n14854 & n14855 ) ;
  assign n14857 = x114 & n4470 ;
  assign n14858 = n14856 | n14857 ;
  assign n14859 = ( x44 & n14853 ) | ( x44 & ~n14858 ) | ( n14853 & ~n14858 ) ;
  assign n14860 = ( ~x44 & n14858 ) | ( ~x44 & n14859 ) | ( n14858 & n14859 ) ;
  assign n14861 = ( ~n14853 & n14859 ) | ( ~n14853 & n14860 ) | ( n14859 & n14860 ) ;
  assign n14862 = n4787 & n5542 ;
  assign n14863 = x112 & n4791 ;
  assign n14864 = x113 | n14863 ;
  assign n14865 = ( n4793 & n14863 ) | ( n4793 & n14864 ) | ( n14863 & n14864 ) ;
  assign n14866 = x111 & n5030 ;
  assign n14867 = n14865 | n14866 ;
  assign n14868 = ( x47 & n14862 ) | ( x47 & ~n14867 ) | ( n14862 & ~n14867 ) ;
  assign n14869 = ( ~x47 & n14867 ) | ( ~x47 & n14868 ) | ( n14867 & n14868 ) ;
  assign n14870 = ( ~n14862 & n14868 ) | ( ~n14862 & n14869 ) | ( n14868 & n14869 ) ;
  assign n14871 = n4934 & n5374 ;
  assign n14872 = x109 & n5378 ;
  assign n14873 = x110 | n14872 ;
  assign n14874 = ( n5380 & n14872 ) | ( n5380 & n14873 ) | ( n14872 & n14873 ) ;
  assign n14875 = x108 & n5638 ;
  assign n14876 = n14874 | n14875 ;
  assign n14877 = ( x50 & n14871 ) | ( x50 & ~n14876 ) | ( n14871 & ~n14876 ) ;
  assign n14878 = ( ~x50 & n14876 ) | ( ~x50 & n14877 ) | ( n14876 & n14877 ) ;
  assign n14879 = ( ~n14871 & n14877 ) | ( ~n14871 & n14878 ) | ( n14877 & n14878 ) ;
  assign n14880 = n4362 & n6027 ;
  assign n14881 = x106 & n6031 ;
  assign n14882 = x107 | n14881 ;
  assign n14883 = ( n6033 & n14881 ) | ( n6033 & n14882 ) | ( n14881 & n14882 ) ;
  assign n14884 = x105 & n6303 ;
  assign n14885 = n14883 | n14884 ;
  assign n14886 = ( x53 & n14880 ) | ( x53 & ~n14885 ) | ( n14880 & ~n14885 ) ;
  assign n14887 = ( ~x53 & n14885 ) | ( ~x53 & n14886 ) | ( n14885 & n14886 ) ;
  assign n14888 = ( ~n14880 & n14886 ) | ( ~n14880 & n14887 ) | ( n14886 & n14887 ) ;
  assign n14889 = n3665 & n6713 ;
  assign n14890 = x103 & n6717 ;
  assign n14891 = x104 | n14890 ;
  assign n14892 = ( n6719 & n14890 ) | ( n6719 & n14891 ) | ( n14890 & n14891 ) ;
  assign n14893 = x102 & n6980 ;
  assign n14894 = n14892 | n14893 ;
  assign n14895 = ( x56 & n14889 ) | ( x56 & ~n14894 ) | ( n14889 & ~n14894 ) ;
  assign n14896 = ( ~x56 & n14894 ) | ( ~x56 & n14895 ) | ( n14894 & n14895 ) ;
  assign n14897 = ( ~n14889 & n14895 ) | ( ~n14889 & n14896 ) | ( n14895 & n14896 ) ;
  assign n14898 = n3326 & n7423 ;
  assign n14899 = x100 & n7427 ;
  assign n14900 = x101 | n14899 ;
  assign n14901 = ( n7429 & n14899 ) | ( n7429 & n14900 ) | ( n14899 & n14900 ) ;
  assign n14902 = x99 & n7708 ;
  assign n14903 = n14901 | n14902 ;
  assign n14904 = ( x59 & n14898 ) | ( x59 & ~n14903 ) | ( n14898 & ~n14903 ) ;
  assign n14905 = ( ~x59 & n14903 ) | ( ~x59 & n14904 ) | ( n14903 & n14904 ) ;
  assign n14906 = ( ~n14898 & n14904 ) | ( ~n14898 & n14905 ) | ( n14904 & n14905 ) ;
  assign n14907 = n2725 & n8154 ;
  assign n14908 = x97 & n8158 ;
  assign n14909 = x98 | n14908 ;
  assign n14910 = ( n8160 & n14908 ) | ( n8160 & n14909 ) | ( n14908 & n14909 ) ;
  assign n14911 = x96 & n8439 ;
  assign n14912 = n14910 | n14911 ;
  assign n14913 = ( x62 & n14907 ) | ( x62 & ~n14912 ) | ( n14907 & ~n14912 ) ;
  assign n14914 = ( ~x62 & n14912 ) | ( ~x62 & n14913 ) | ( n14912 & n14913 ) ;
  assign n14915 = ( ~n14907 & n14913 ) | ( ~n14907 & n14914 ) | ( n14913 & n14914 ) ;
  assign n14916 = x94 & n8927 ;
  assign n14917 = ( ~x95 & n8693 ) | ( ~x95 & n8927 ) | ( n8693 & n8927 ) ;
  assign n14918 = ( n8693 & n14916 ) | ( n8693 & ~n14917 ) | ( n14916 & ~n14917 ) ;
  assign n14919 = ( ~n14780 & n14915 ) | ( ~n14780 & n14918 ) | ( n14915 & n14918 ) ;
  assign n14920 = ( n14915 & n14918 ) | ( n14915 & ~n14919 ) | ( n14918 & ~n14919 ) ;
  assign n14921 = ( n14780 & n14919 ) | ( n14780 & ~n14920 ) | ( n14919 & ~n14920 ) ;
  assign n14922 = ( n14783 & n14906 ) | ( n14783 & ~n14921 ) | ( n14906 & ~n14921 ) ;
  assign n14923 = ( ~n14783 & n14906 ) | ( ~n14783 & n14921 ) | ( n14906 & n14921 ) ;
  assign n14924 = ( ~n14906 & n14922 ) | ( ~n14906 & n14923 ) | ( n14922 & n14923 ) ;
  assign n14925 = ( n14786 & n14897 ) | ( n14786 & ~n14924 ) | ( n14897 & ~n14924 ) ;
  assign n14926 = ( ~n14786 & n14897 ) | ( ~n14786 & n14924 ) | ( n14897 & n14924 ) ;
  assign n14927 = ( ~n14897 & n14925 ) | ( ~n14897 & n14926 ) | ( n14925 & n14926 ) ;
  assign n14928 = ( n14789 & n14888 ) | ( n14789 & ~n14927 ) | ( n14888 & ~n14927 ) ;
  assign n14929 = ( ~n14789 & n14888 ) | ( ~n14789 & n14927 ) | ( n14888 & n14927 ) ;
  assign n14930 = ( ~n14888 & n14928 ) | ( ~n14888 & n14929 ) | ( n14928 & n14929 ) ;
  assign n14931 = ( n14792 & n14879 ) | ( n14792 & ~n14930 ) | ( n14879 & ~n14930 ) ;
  assign n14932 = ( ~n14792 & n14879 ) | ( ~n14792 & n14930 ) | ( n14879 & n14930 ) ;
  assign n14933 = ( ~n14879 & n14931 ) | ( ~n14879 & n14932 ) | ( n14931 & n14932 ) ;
  assign n14934 = ( n14795 & n14870 ) | ( n14795 & ~n14933 ) | ( n14870 & ~n14933 ) ;
  assign n14935 = ( ~n14795 & n14870 ) | ( ~n14795 & n14933 ) | ( n14870 & n14933 ) ;
  assign n14936 = ( ~n14870 & n14934 ) | ( ~n14870 & n14935 ) | ( n14934 & n14935 ) ;
  assign n14937 = ( n14798 & n14861 ) | ( n14798 & ~n14936 ) | ( n14861 & ~n14936 ) ;
  assign n14938 = ( ~n14798 & n14861 ) | ( ~n14798 & n14936 ) | ( n14861 & n14936 ) ;
  assign n14939 = ( ~n14861 & n14937 ) | ( ~n14861 & n14938 ) | ( n14937 & n14938 ) ;
  assign n14940 = ( n14801 & n14852 ) | ( n14801 & ~n14939 ) | ( n14852 & ~n14939 ) ;
  assign n14941 = ( ~n14801 & n14852 ) | ( ~n14801 & n14939 ) | ( n14852 & n14939 ) ;
  assign n14942 = ( ~n14852 & n14940 ) | ( ~n14852 & n14941 ) | ( n14940 & n14941 ) ;
  assign n14943 = ( n14804 & n14843 ) | ( n14804 & ~n14942 ) | ( n14843 & ~n14942 ) ;
  assign n14944 = ( ~n14804 & n14843 ) | ( ~n14804 & n14942 ) | ( n14843 & n14942 ) ;
  assign n14945 = ( ~n14843 & n14943 ) | ( ~n14843 & n14944 ) | ( n14943 & n14944 ) ;
  assign n14946 = n2766 & n8331 ;
  assign n14947 = x124 & n2770 ;
  assign n14948 = x125 | n14947 ;
  assign n14949 = ( n2772 & n14947 ) | ( n2772 & n14948 ) | ( n14947 & n14948 ) ;
  assign n14950 = x123 & n2943 ;
  assign n14951 = n14949 | n14950 ;
  assign n14952 = ( x35 & n14946 ) | ( x35 & ~n14951 ) | ( n14946 & ~n14951 ) ;
  assign n14953 = ( ~x35 & n14951 ) | ( ~x35 & n14952 ) | ( n14951 & n14952 ) ;
  assign n14954 = ( ~n14946 & n14952 ) | ( ~n14946 & n14953 ) | ( n14952 & n14953 ) ;
  assign n14955 = ( n14807 & ~n14945 ) | ( n14807 & n14954 ) | ( ~n14945 & n14954 ) ;
  assign n14956 = ( n14807 & n14945 ) | ( n14807 & n14954 ) | ( n14945 & n14954 ) ;
  assign n14957 = ( n14945 & n14955 ) | ( n14945 & ~n14956 ) | ( n14955 & ~n14956 ) ;
  assign n14958 = ( n14810 & n14834 ) | ( n14810 & ~n14957 ) | ( n14834 & ~n14957 ) ;
  assign n14959 = ( ~n14810 & n14834 ) | ( ~n14810 & n14957 ) | ( n14834 & n14957 ) ;
  assign n14960 = ( ~n14834 & n14958 ) | ( ~n14834 & n14959 ) | ( n14958 & n14959 ) ;
  assign n14961 = ( ~n14822 & n14825 ) | ( ~n14822 & n14960 ) | ( n14825 & n14960 ) ;
  assign n14962 = ( n14825 & n14960 ) | ( n14825 & ~n14961 ) | ( n14960 & ~n14961 ) ;
  assign n14963 = ( n14822 & n14961 ) | ( n14822 & ~n14962 ) | ( n14961 & ~n14962 ) ;
  assign n14964 = n2320 & n8862 ;
  assign n14965 = ( x127 & n2497 ) | ( x127 & n14964 ) | ( n2497 & n14964 ) ;
  assign n14966 = x32 | n14965 ;
  assign n14967 = ~x32 & n14965 ;
  assign n14968 = ( ~n14965 & n14966 ) | ( ~n14965 & n14967 ) | ( n14966 & n14967 ) ;
  assign n14969 = n3224 & n7597 ;
  assign n14970 = x122 & n3228 ;
  assign n14971 = x123 | n14970 ;
  assign n14972 = ( n3230 & n14970 ) | ( n3230 & n14971 ) | ( n14970 & n14971 ) ;
  assign n14973 = x121 & n3413 ;
  assign n14974 = n14972 | n14973 ;
  assign n14975 = ( x38 & n14969 ) | ( x38 & ~n14974 ) | ( n14969 & ~n14974 ) ;
  assign n14976 = ( ~x38 & n14974 ) | ( ~x38 & n14975 ) | ( n14974 & n14975 ) ;
  assign n14977 = ( ~n14969 & n14975 ) | ( ~n14969 & n14976 ) | ( n14975 & n14976 ) ;
  assign n14978 = n3715 & n7098 ;
  assign n14979 = x119 & n3719 ;
  assign n14980 = x120 | n14979 ;
  assign n14981 = ( n3721 & n14979 ) | ( n3721 & n14980 ) | ( n14979 & n14980 ) ;
  assign n14982 = x118 & n3922 ;
  assign n14983 = n14981 | n14982 ;
  assign n14984 = ( x41 & n14978 ) | ( x41 & ~n14983 ) | ( n14978 & ~n14983 ) ;
  assign n14985 = ( ~x41 & n14983 ) | ( ~x41 & n14984 ) | ( n14983 & n14984 ) ;
  assign n14986 = ( ~n14978 & n14984 ) | ( ~n14978 & n14985 ) | ( n14984 & n14985 ) ;
  assign n14987 = n4227 & n6201 ;
  assign n14988 = x116 & n4231 ;
  assign n14989 = x117 | n14988 ;
  assign n14990 = ( n4233 & n14988 ) | ( n4233 & n14989 ) | ( n14988 & n14989 ) ;
  assign n14991 = x115 & n4470 ;
  assign n14992 = n14990 | n14991 ;
  assign n14993 = ( x44 & n14987 ) | ( x44 & ~n14992 ) | ( n14987 & ~n14992 ) ;
  assign n14994 = ( ~x44 & n14992 ) | ( ~x44 & n14993 ) | ( n14992 & n14993 ) ;
  assign n14995 = ( ~n14987 & n14993 ) | ( ~n14987 & n14994 ) | ( n14993 & n14994 ) ;
  assign n14996 = n4787 & n5750 ;
  assign n14997 = x113 & n4791 ;
  assign n14998 = x114 | n14997 ;
  assign n14999 = ( n4793 & n14997 ) | ( n4793 & n14998 ) | ( n14997 & n14998 ) ;
  assign n15000 = x112 & n5030 ;
  assign n15001 = n14999 | n15000 ;
  assign n15002 = ( x47 & n14996 ) | ( x47 & ~n15001 ) | ( n14996 & ~n15001 ) ;
  assign n15003 = ( ~x47 & n15001 ) | ( ~x47 & n15002 ) | ( n15001 & n15002 ) ;
  assign n15004 = ( ~n14996 & n15002 ) | ( ~n14996 & n15003 ) | ( n15002 & n15003 ) ;
  assign n15005 = n5130 & n5374 ;
  assign n15006 = x110 & n5378 ;
  assign n15007 = x111 | n15006 ;
  assign n15008 = ( n5380 & n15006 ) | ( n5380 & n15007 ) | ( n15006 & n15007 ) ;
  assign n15009 = x109 & n5638 ;
  assign n15010 = n15008 | n15009 ;
  assign n15011 = ( x50 & n15005 ) | ( x50 & ~n15010 ) | ( n15005 & ~n15010 ) ;
  assign n15012 = ( ~x50 & n15010 ) | ( ~x50 & n15011 ) | ( n15010 & n15011 ) ;
  assign n15013 = ( ~n15005 & n15011 ) | ( ~n15005 & n15012 ) | ( n15011 & n15012 ) ;
  assign n15014 = n4377 & n6027 ;
  assign n15015 = x107 & n6031 ;
  assign n15016 = x108 | n15015 ;
  assign n15017 = ( n6033 & n15015 ) | ( n6033 & n15016 ) | ( n15015 & n15016 ) ;
  assign n15018 = x106 & n6303 ;
  assign n15019 = n15017 | n15018 ;
  assign n15020 = ( x53 & n15014 ) | ( x53 & ~n15019 ) | ( n15014 & ~n15019 ) ;
  assign n15021 = ( ~x53 & n15019 ) | ( ~x53 & n15020 ) | ( n15019 & n15020 ) ;
  assign n15022 = ( ~n15014 & n15020 ) | ( ~n15014 & n15021 ) | ( n15020 & n15021 ) ;
  assign n15023 = n3998 & n6713 ;
  assign n15024 = x104 & n6717 ;
  assign n15025 = x105 | n15024 ;
  assign n15026 = ( n6719 & n15024 ) | ( n6719 & n15025 ) | ( n15024 & n15025 ) ;
  assign n15027 = x103 & n6980 ;
  assign n15028 = n15026 | n15027 ;
  assign n15029 = ( x56 & n15023 ) | ( x56 & ~n15028 ) | ( n15023 & ~n15028 ) ;
  assign n15030 = ( ~x56 & n15028 ) | ( ~x56 & n15029 ) | ( n15028 & n15029 ) ;
  assign n15031 = ( ~n15023 & n15029 ) | ( ~n15023 & n15030 ) | ( n15029 & n15030 ) ;
  assign n15032 = x95 & n8927 ;
  assign n15033 = ( ~x96 & n8693 ) | ( ~x96 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15034 = ( n8693 & n15032 ) | ( n8693 & ~n15033 ) | ( n15032 & ~n15033 ) ;
  assign n15035 = ( n14780 & n14919 ) | ( n14780 & ~n15034 ) | ( n14919 & ~n15034 ) ;
  assign n15036 = ( n14780 & ~n14919 ) | ( n14780 & n15034 ) | ( ~n14919 & n15034 ) ;
  assign n15037 = ( ~n14780 & n15035 ) | ( ~n14780 & n15036 ) | ( n15035 & n15036 ) ;
  assign n15038 = n3486 & n7423 ;
  assign n15039 = x101 & n7427 ;
  assign n15040 = x102 | n15039 ;
  assign n15041 = ( n7429 & n15039 ) | ( n7429 & n15040 ) | ( n15039 & n15040 ) ;
  assign n15042 = x100 & n7708 ;
  assign n15043 = n15041 | n15042 ;
  assign n15044 = ( x59 & n15038 ) | ( x59 & ~n15043 ) | ( n15038 & ~n15043 ) ;
  assign n15045 = ( ~x59 & n15043 ) | ( ~x59 & n15044 ) | ( n15043 & n15044 ) ;
  assign n15046 = ( ~n15038 & n15044 ) | ( ~n15038 & n15045 ) | ( n15044 & n15045 ) ;
  assign n15047 = n2877 & n8154 ;
  assign n15048 = x98 & n8158 ;
  assign n15049 = x99 | n15048 ;
  assign n15050 = ( n8160 & n15048 ) | ( n8160 & n15049 ) | ( n15048 & n15049 ) ;
  assign n15051 = x97 & n8439 ;
  assign n15052 = n15050 | n15051 ;
  assign n15053 = ( x62 & n15047 ) | ( x62 & ~n15052 ) | ( n15047 & ~n15052 ) ;
  assign n15054 = ( ~x62 & n15052 ) | ( ~x62 & n15053 ) | ( n15052 & n15053 ) ;
  assign n15055 = ( ~n15047 & n15053 ) | ( ~n15047 & n15054 ) | ( n15053 & n15054 ) ;
  assign n15056 = ( ~n15037 & n15046 ) | ( ~n15037 & n15055 ) | ( n15046 & n15055 ) ;
  assign n15057 = ( n15046 & n15055 ) | ( n15046 & ~n15056 ) | ( n15055 & ~n15056 ) ;
  assign n15058 = ( n15037 & n15056 ) | ( n15037 & ~n15057 ) | ( n15056 & ~n15057 ) ;
  assign n15059 = ( n14922 & n15031 ) | ( n14922 & ~n15058 ) | ( n15031 & ~n15058 ) ;
  assign n15060 = ( ~n14922 & n15031 ) | ( ~n14922 & n15058 ) | ( n15031 & n15058 ) ;
  assign n15061 = ( ~n15031 & n15059 ) | ( ~n15031 & n15060 ) | ( n15059 & n15060 ) ;
  assign n15062 = ( n14925 & n15022 ) | ( n14925 & ~n15061 ) | ( n15022 & ~n15061 ) ;
  assign n15063 = ( ~n14925 & n15022 ) | ( ~n14925 & n15061 ) | ( n15022 & n15061 ) ;
  assign n15064 = ( ~n15022 & n15062 ) | ( ~n15022 & n15063 ) | ( n15062 & n15063 ) ;
  assign n15065 = ( n14928 & n15013 ) | ( n14928 & ~n15064 ) | ( n15013 & ~n15064 ) ;
  assign n15066 = ( ~n14928 & n15013 ) | ( ~n14928 & n15064 ) | ( n15013 & n15064 ) ;
  assign n15067 = ( ~n15013 & n15065 ) | ( ~n15013 & n15066 ) | ( n15065 & n15066 ) ;
  assign n15068 = ( n14931 & n15004 ) | ( n14931 & ~n15067 ) | ( n15004 & ~n15067 ) ;
  assign n15069 = ( ~n14931 & n15004 ) | ( ~n14931 & n15067 ) | ( n15004 & n15067 ) ;
  assign n15070 = ( ~n15004 & n15068 ) | ( ~n15004 & n15069 ) | ( n15068 & n15069 ) ;
  assign n15071 = ( n14934 & n14995 ) | ( n14934 & ~n15070 ) | ( n14995 & ~n15070 ) ;
  assign n15072 = ( ~n14934 & n14995 ) | ( ~n14934 & n15070 ) | ( n14995 & n15070 ) ;
  assign n15073 = ( ~n14995 & n15071 ) | ( ~n14995 & n15072 ) | ( n15071 & n15072 ) ;
  assign n15074 = ( n14937 & n14986 ) | ( n14937 & ~n15073 ) | ( n14986 & ~n15073 ) ;
  assign n15075 = ( ~n14937 & n14986 ) | ( ~n14937 & n15073 ) | ( n14986 & n15073 ) ;
  assign n15076 = ( ~n14986 & n15074 ) | ( ~n14986 & n15075 ) | ( n15074 & n15075 ) ;
  assign n15077 = ( n14940 & n14977 ) | ( n14940 & ~n15076 ) | ( n14977 & ~n15076 ) ;
  assign n15078 = ( ~n14940 & n14977 ) | ( ~n14940 & n15076 ) | ( n14977 & n15076 ) ;
  assign n15079 = ( ~n14977 & n15077 ) | ( ~n14977 & n15078 ) | ( n15077 & n15078 ) ;
  assign n15080 = n2766 & n8587 ;
  assign n15081 = x125 & n2770 ;
  assign n15082 = x126 | n15081 ;
  assign n15083 = ( n2772 & n15081 ) | ( n2772 & n15082 ) | ( n15081 & n15082 ) ;
  assign n15084 = x124 & n2943 ;
  assign n15085 = n15083 | n15084 ;
  assign n15086 = ( x35 & n15080 ) | ( x35 & ~n15085 ) | ( n15080 & ~n15085 ) ;
  assign n15087 = ( ~x35 & n15085 ) | ( ~x35 & n15086 ) | ( n15085 & n15086 ) ;
  assign n15088 = ( ~n15080 & n15086 ) | ( ~n15080 & n15087 ) | ( n15086 & n15087 ) ;
  assign n15089 = ( n14943 & ~n15079 ) | ( n14943 & n15088 ) | ( ~n15079 & n15088 ) ;
  assign n15090 = ( n14943 & n15079 ) | ( n14943 & n15088 ) | ( n15079 & n15088 ) ;
  assign n15091 = ( n15079 & n15089 ) | ( n15079 & ~n15090 ) | ( n15089 & ~n15090 ) ;
  assign n15092 = ( n14955 & n14968 ) | ( n14955 & ~n15091 ) | ( n14968 & ~n15091 ) ;
  assign n15093 = ( ~n14955 & n14968 ) | ( ~n14955 & n15091 ) | ( n14968 & n15091 ) ;
  assign n15094 = ( ~n14968 & n15092 ) | ( ~n14968 & n15093 ) | ( n15092 & n15093 ) ;
  assign n15095 = ( ~n14958 & n14961 ) | ( ~n14958 & n15094 ) | ( n14961 & n15094 ) ;
  assign n15096 = ( n14961 & n15094 ) | ( n14961 & ~n15095 ) | ( n15094 & ~n15095 ) ;
  assign n15097 = ( n14958 & n15095 ) | ( n14958 & ~n15096 ) | ( n15095 & ~n15096 ) ;
  assign n15098 = n3224 & n7841 ;
  assign n15099 = x123 & n3228 ;
  assign n15100 = x124 | n15099 ;
  assign n15101 = ( n3230 & n15099 ) | ( n3230 & n15100 ) | ( n15099 & n15100 ) ;
  assign n15102 = x122 & n3413 ;
  assign n15103 = n15101 | n15102 ;
  assign n15104 = ( x38 & n15098 ) | ( x38 & ~n15103 ) | ( n15098 & ~n15103 ) ;
  assign n15105 = ( ~x38 & n15103 ) | ( ~x38 & n15104 ) | ( n15103 & n15104 ) ;
  assign n15106 = ( ~n15098 & n15104 ) | ( ~n15098 & n15105 ) | ( n15104 & n15105 ) ;
  assign n15107 = n3715 & n7113 ;
  assign n15108 = x120 & n3719 ;
  assign n15109 = x121 | n15108 ;
  assign n15110 = ( n3721 & n15108 ) | ( n3721 & n15109 ) | ( n15108 & n15109 ) ;
  assign n15111 = x119 & n3922 ;
  assign n15112 = n15110 | n15111 ;
  assign n15113 = ( x41 & n15107 ) | ( x41 & ~n15112 ) | ( n15107 & ~n15112 ) ;
  assign n15114 = ( ~x41 & n15112 ) | ( ~x41 & n15113 ) | ( n15112 & n15113 ) ;
  assign n15115 = ( ~n15107 & n15113 ) | ( ~n15107 & n15114 ) | ( n15113 & n15114 ) ;
  assign n15116 = n4227 & n6421 ;
  assign n15117 = x117 & n4231 ;
  assign n15118 = x118 | n15117 ;
  assign n15119 = ( n4233 & n15117 ) | ( n4233 & n15118 ) | ( n15117 & n15118 ) ;
  assign n15120 = x116 & n4470 ;
  assign n15121 = n15119 | n15120 ;
  assign n15122 = ( x44 & n15116 ) | ( x44 & ~n15121 ) | ( n15116 & ~n15121 ) ;
  assign n15123 = ( ~x44 & n15121 ) | ( ~x44 & n15122 ) | ( n15121 & n15122 ) ;
  assign n15124 = ( ~n15116 & n15122 ) | ( ~n15116 & n15123 ) | ( n15122 & n15123 ) ;
  assign n15125 = n4787 & n5765 ;
  assign n15126 = x114 & n4791 ;
  assign n15127 = x115 | n15126 ;
  assign n15128 = ( n4793 & n15126 ) | ( n4793 & n15127 ) | ( n15126 & n15127 ) ;
  assign n15129 = x113 & n5030 ;
  assign n15130 = n15128 | n15129 ;
  assign n15131 = ( x47 & n15125 ) | ( x47 & ~n15130 ) | ( n15125 & ~n15130 ) ;
  assign n15132 = ( ~x47 & n15130 ) | ( ~x47 & n15131 ) | ( n15130 & n15131 ) ;
  assign n15133 = ( ~n15125 & n15131 ) | ( ~n15125 & n15132 ) | ( n15131 & n15132 ) ;
  assign n15134 = n5145 & n5374 ;
  assign n15135 = x111 & n5378 ;
  assign n15136 = x112 | n15135 ;
  assign n15137 = ( n5380 & n15135 ) | ( n5380 & n15136 ) | ( n15135 & n15136 ) ;
  assign n15138 = x110 & n5638 ;
  assign n15139 = n15137 | n15138 ;
  assign n15140 = ( x50 & n15134 ) | ( x50 & ~n15139 ) | ( n15134 & ~n15139 ) ;
  assign n15141 = ( ~x50 & n15139 ) | ( ~x50 & n15140 ) | ( n15139 & n15140 ) ;
  assign n15142 = ( ~n15134 & n15140 ) | ( ~n15134 & n15141 ) | ( n15140 & n15141 ) ;
  assign n15143 = n4734 & n6027 ;
  assign n15144 = x108 & n6031 ;
  assign n15145 = x109 | n15144 ;
  assign n15146 = ( n6033 & n15144 ) | ( n6033 & n15145 ) | ( n15144 & n15145 ) ;
  assign n15147 = x107 & n6303 ;
  assign n15148 = n15146 | n15147 ;
  assign n15149 = ( x53 & n15143 ) | ( x53 & ~n15148 ) | ( n15143 & ~n15148 ) ;
  assign n15150 = ( ~x53 & n15148 ) | ( ~x53 & n15149 ) | ( n15148 & n15149 ) ;
  assign n15151 = ( ~n15143 & n15149 ) | ( ~n15143 & n15150 ) | ( n15149 & n15150 ) ;
  assign n15152 = n4013 & n6713 ;
  assign n15153 = x105 & n6717 ;
  assign n15154 = x106 | n15153 ;
  assign n15155 = ( n6719 & n15153 ) | ( n6719 & n15154 ) | ( n15153 & n15154 ) ;
  assign n15156 = x104 & n6980 ;
  assign n15157 = n15155 | n15156 ;
  assign n15158 = ( x56 & n15152 ) | ( x56 & ~n15157 ) | ( n15152 & ~n15157 ) ;
  assign n15159 = ( ~x56 & n15157 ) | ( ~x56 & n15158 ) | ( n15157 & n15158 ) ;
  assign n15160 = ( ~n15152 & n15158 ) | ( ~n15152 & n15159 ) | ( n15158 & n15159 ) ;
  assign n15161 = n3650 & n7423 ;
  assign n15162 = x102 & n7427 ;
  assign n15163 = x103 | n15162 ;
  assign n15164 = ( n7429 & n15162 ) | ( n7429 & n15163 ) | ( n15162 & n15163 ) ;
  assign n15165 = x101 & n7708 ;
  assign n15166 = n15164 | n15165 ;
  assign n15167 = ( x59 & n15161 ) | ( x59 & ~n15166 ) | ( n15161 & ~n15166 ) ;
  assign n15168 = ( ~x59 & n15166 ) | ( ~x59 & n15167 ) | ( n15166 & n15167 ) ;
  assign n15169 = ( ~n15161 & n15167 ) | ( ~n15161 & n15168 ) | ( n15167 & n15168 ) ;
  assign n15170 = n3162 & n8154 ;
  assign n15171 = x99 & n8158 ;
  assign n15172 = x100 | n15171 ;
  assign n15173 = ( n8160 & n15171 ) | ( n8160 & n15172 ) | ( n15171 & n15172 ) ;
  assign n15174 = x98 & n8439 ;
  assign n15175 = n15173 | n15174 ;
  assign n15176 = ( x62 & n15170 ) | ( x62 & ~n15175 ) | ( n15170 & ~n15175 ) ;
  assign n15177 = ( ~x62 & n15175 ) | ( ~x62 & n15176 ) | ( n15175 & n15176 ) ;
  assign n15178 = ( ~n15170 & n15176 ) | ( ~n15170 & n15177 ) | ( n15176 & n15177 ) ;
  assign n15179 = x96 & n8927 ;
  assign n15180 = ( ~x97 & n8693 ) | ( ~x97 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15181 = ( n8693 & n15179 ) | ( n8693 & ~n15180 ) | ( n15179 & ~n15180 ) ;
  assign n15182 = ( ~x32 & n15034 ) | ( ~x32 & n15181 ) | ( n15034 & n15181 ) ;
  assign n15183 = ( n15034 & n15181 ) | ( n15034 & ~n15182 ) | ( n15181 & ~n15182 ) ;
  assign n15184 = ( x32 & n15182 ) | ( x32 & ~n15183 ) | ( n15182 & ~n15183 ) ;
  assign n15185 = ( n15035 & n15178 ) | ( n15035 & ~n15184 ) | ( n15178 & ~n15184 ) ;
  assign n15186 = ( ~n15035 & n15178 ) | ( ~n15035 & n15184 ) | ( n15178 & n15184 ) ;
  assign n15187 = ( ~n15178 & n15185 ) | ( ~n15178 & n15186 ) | ( n15185 & n15186 ) ;
  assign n15188 = ( n15056 & n15169 ) | ( n15056 & ~n15187 ) | ( n15169 & ~n15187 ) ;
  assign n15189 = ( ~n15056 & n15169 ) | ( ~n15056 & n15187 ) | ( n15169 & n15187 ) ;
  assign n15190 = ( ~n15169 & n15188 ) | ( ~n15169 & n15189 ) | ( n15188 & n15189 ) ;
  assign n15191 = ( n15059 & n15160 ) | ( n15059 & ~n15190 ) | ( n15160 & ~n15190 ) ;
  assign n15192 = ( ~n15059 & n15160 ) | ( ~n15059 & n15190 ) | ( n15160 & n15190 ) ;
  assign n15193 = ( ~n15160 & n15191 ) | ( ~n15160 & n15192 ) | ( n15191 & n15192 ) ;
  assign n15194 = ( n15062 & n15151 ) | ( n15062 & ~n15193 ) | ( n15151 & ~n15193 ) ;
  assign n15195 = ( ~n15062 & n15151 ) | ( ~n15062 & n15193 ) | ( n15151 & n15193 ) ;
  assign n15196 = ( ~n15151 & n15194 ) | ( ~n15151 & n15195 ) | ( n15194 & n15195 ) ;
  assign n15197 = ( n15065 & n15142 ) | ( n15065 & ~n15196 ) | ( n15142 & ~n15196 ) ;
  assign n15198 = ( ~n15065 & n15142 ) | ( ~n15065 & n15196 ) | ( n15142 & n15196 ) ;
  assign n15199 = ( ~n15142 & n15197 ) | ( ~n15142 & n15198 ) | ( n15197 & n15198 ) ;
  assign n15200 = ( n15068 & n15133 ) | ( n15068 & ~n15199 ) | ( n15133 & ~n15199 ) ;
  assign n15201 = ( ~n15068 & n15133 ) | ( ~n15068 & n15199 ) | ( n15133 & n15199 ) ;
  assign n15202 = ( ~n15133 & n15200 ) | ( ~n15133 & n15201 ) | ( n15200 & n15201 ) ;
  assign n15203 = ( n15071 & n15124 ) | ( n15071 & ~n15202 ) | ( n15124 & ~n15202 ) ;
  assign n15204 = ( ~n15071 & n15124 ) | ( ~n15071 & n15202 ) | ( n15124 & n15202 ) ;
  assign n15205 = ( ~n15124 & n15203 ) | ( ~n15124 & n15204 ) | ( n15203 & n15204 ) ;
  assign n15206 = ( n15074 & n15115 ) | ( n15074 & ~n15205 ) | ( n15115 & ~n15205 ) ;
  assign n15207 = ( ~n15074 & n15115 ) | ( ~n15074 & n15205 ) | ( n15115 & n15205 ) ;
  assign n15208 = ( ~n15115 & n15206 ) | ( ~n15115 & n15207 ) | ( n15206 & n15207 ) ;
  assign n15209 = ( n15077 & n15106 ) | ( n15077 & ~n15208 ) | ( n15106 & ~n15208 ) ;
  assign n15210 = ( ~n15077 & n15106 ) | ( ~n15077 & n15208 ) | ( n15106 & n15208 ) ;
  assign n15211 = ( ~n15106 & n15209 ) | ( ~n15106 & n15210 ) | ( n15209 & n15210 ) ;
  assign n15212 = n2766 & n8846 ;
  assign n15213 = x126 & n2770 ;
  assign n15214 = x127 | n15213 ;
  assign n15215 = ( n2772 & n15213 ) | ( n2772 & n15214 ) | ( n15213 & n15214 ) ;
  assign n15216 = x125 & n2943 ;
  assign n15217 = n15215 | n15216 ;
  assign n15218 = ( x35 & n15212 ) | ( x35 & ~n15217 ) | ( n15212 & ~n15217 ) ;
  assign n15219 = ( ~x35 & n15217 ) | ( ~x35 & n15218 ) | ( n15217 & n15218 ) ;
  assign n15220 = ( ~n15212 & n15218 ) | ( ~n15212 & n15219 ) | ( n15218 & n15219 ) ;
  assign n15221 = ( n15089 & ~n15211 ) | ( n15089 & n15220 ) | ( ~n15211 & n15220 ) ;
  assign n15222 = ( n15089 & n15211 ) | ( n15089 & n15220 ) | ( n15211 & n15220 ) ;
  assign n15223 = ( n15211 & n15221 ) | ( n15211 & ~n15222 ) | ( n15221 & ~n15222 ) ;
  assign n15224 = ( ~n15092 & n15095 ) | ( ~n15092 & n15223 ) | ( n15095 & n15223 ) ;
  assign n15225 = ( n15095 & n15223 ) | ( n15095 & ~n15224 ) | ( n15223 & ~n15224 ) ;
  assign n15226 = ( n15092 & n15224 ) | ( n15092 & ~n15225 ) | ( n15224 & ~n15225 ) ;
  assign n15227 = n2766 & n8865 ;
  assign n15228 = x127 & n2770 ;
  assign n15229 = x126 | n15228 ;
  assign n15230 = ( n2943 & n15228 ) | ( n2943 & n15229 ) | ( n15228 & n15229 ) ;
  assign n15231 = ( x35 & n15227 ) | ( x35 & ~n15230 ) | ( n15227 & ~n15230 ) ;
  assign n15232 = ( ~x35 & n15230 ) | ( ~x35 & n15231 ) | ( n15230 & n15231 ) ;
  assign n15233 = ( ~n15227 & n15231 ) | ( ~n15227 & n15232 ) | ( n15231 & n15232 ) ;
  assign n15234 = n3715 & n7582 ;
  assign n15235 = x121 & n3719 ;
  assign n15236 = x122 | n15235 ;
  assign n15237 = ( n3721 & n15235 ) | ( n3721 & n15236 ) | ( n15235 & n15236 ) ;
  assign n15238 = x120 & n3922 ;
  assign n15239 = n15237 | n15238 ;
  assign n15240 = ( x41 & n15234 ) | ( x41 & ~n15239 ) | ( n15234 & ~n15239 ) ;
  assign n15241 = ( ~x41 & n15239 ) | ( ~x41 & n15240 ) | ( n15239 & n15240 ) ;
  assign n15242 = ( ~n15234 & n15240 ) | ( ~n15234 & n15241 ) | ( n15240 & n15241 ) ;
  assign n15243 = n4227 & n6645 ;
  assign n15244 = x118 & n4231 ;
  assign n15245 = x119 | n15244 ;
  assign n15246 = ( n4233 & n15244 ) | ( n4233 & n15245 ) | ( n15244 & n15245 ) ;
  assign n15247 = x117 & n4470 ;
  assign n15248 = n15246 | n15247 ;
  assign n15249 = ( x44 & n15243 ) | ( x44 & ~n15248 ) | ( n15243 & ~n15248 ) ;
  assign n15250 = ( ~x44 & n15248 ) | ( ~x44 & n15249 ) | ( n15248 & n15249 ) ;
  assign n15251 = ( ~n15243 & n15249 ) | ( ~n15243 & n15250 ) | ( n15249 & n15250 ) ;
  assign n15252 = n5374 & n5542 ;
  assign n15253 = x112 & n5378 ;
  assign n15254 = x113 | n15253 ;
  assign n15255 = ( n5380 & n15253 ) | ( n5380 & n15254 ) | ( n15253 & n15254 ) ;
  assign n15256 = x111 & n5638 ;
  assign n15257 = n15255 | n15256 ;
  assign n15258 = ( x50 & n15252 ) | ( x50 & ~n15257 ) | ( n15252 & ~n15257 ) ;
  assign n15259 = ( ~x50 & n15257 ) | ( ~x50 & n15258 ) | ( n15257 & n15258 ) ;
  assign n15260 = ( ~n15252 & n15258 ) | ( ~n15252 & n15259 ) | ( n15258 & n15259 ) ;
  assign n15261 = n4362 & n6713 ;
  assign n15262 = x106 & n6717 ;
  assign n15263 = x107 | n15262 ;
  assign n15264 = ( n6719 & n15262 ) | ( n6719 & n15263 ) | ( n15262 & n15263 ) ;
  assign n15265 = x105 & n6980 ;
  assign n15266 = n15264 | n15265 ;
  assign n15267 = ( x56 & n15261 ) | ( x56 & ~n15266 ) | ( n15261 & ~n15266 ) ;
  assign n15268 = ( ~x56 & n15266 ) | ( ~x56 & n15267 ) | ( n15266 & n15267 ) ;
  assign n15269 = ( ~n15261 & n15267 ) | ( ~n15261 & n15268 ) | ( n15267 & n15268 ) ;
  assign n15270 = n3665 & n7423 ;
  assign n15271 = x103 & n7427 ;
  assign n15272 = x104 | n15271 ;
  assign n15273 = ( n7429 & n15271 ) | ( n7429 & n15272 ) | ( n15271 & n15272 ) ;
  assign n15274 = x102 & n7708 ;
  assign n15275 = n15273 | n15274 ;
  assign n15276 = ( x59 & n15270 ) | ( x59 & ~n15275 ) | ( n15270 & ~n15275 ) ;
  assign n15277 = ( ~x59 & n15275 ) | ( ~x59 & n15276 ) | ( n15275 & n15276 ) ;
  assign n15278 = ( ~n15270 & n15276 ) | ( ~n15270 & n15277 ) | ( n15276 & n15277 ) ;
  assign n15279 = n3326 & n8154 ;
  assign n15280 = x100 & n8158 ;
  assign n15281 = x101 | n15280 ;
  assign n15282 = ( n8160 & n15280 ) | ( n8160 & n15281 ) | ( n15280 & n15281 ) ;
  assign n15283 = x99 & n8439 ;
  assign n15284 = n15282 | n15283 ;
  assign n15285 = ( x62 & n15279 ) | ( x62 & ~n15284 ) | ( n15279 & ~n15284 ) ;
  assign n15286 = ( ~x62 & n15284 ) | ( ~x62 & n15285 ) | ( n15284 & n15285 ) ;
  assign n15287 = ( ~n15279 & n15285 ) | ( ~n15279 & n15286 ) | ( n15285 & n15286 ) ;
  assign n15288 = x97 & n8927 ;
  assign n15289 = ( ~x98 & n8693 ) | ( ~x98 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15290 = ( n8693 & n15288 ) | ( n8693 & ~n15289 ) | ( n15288 & ~n15289 ) ;
  assign n15291 = ( ~n15182 & n15287 ) | ( ~n15182 & n15290 ) | ( n15287 & n15290 ) ;
  assign n15292 = ( n15287 & n15290 ) | ( n15287 & ~n15291 ) | ( n15290 & ~n15291 ) ;
  assign n15293 = ( n15182 & n15291 ) | ( n15182 & ~n15292 ) | ( n15291 & ~n15292 ) ;
  assign n15294 = ( n15185 & n15278 ) | ( n15185 & ~n15293 ) | ( n15278 & ~n15293 ) ;
  assign n15295 = ( ~n15185 & n15278 ) | ( ~n15185 & n15293 ) | ( n15278 & n15293 ) ;
  assign n15296 = ( ~n15278 & n15294 ) | ( ~n15278 & n15295 ) | ( n15294 & n15295 ) ;
  assign n15297 = ( n15188 & n15269 ) | ( n15188 & ~n15296 ) | ( n15269 & ~n15296 ) ;
  assign n15298 = ( ~n15188 & n15269 ) | ( ~n15188 & n15296 ) | ( n15269 & n15296 ) ;
  assign n15299 = ( ~n15269 & n15297 ) | ( ~n15269 & n15298 ) | ( n15297 & n15298 ) ;
  assign n15300 = n4934 & n6027 ;
  assign n15301 = x109 & n6031 ;
  assign n15302 = x110 | n15301 ;
  assign n15303 = ( n6033 & n15301 ) | ( n6033 & n15302 ) | ( n15301 & n15302 ) ;
  assign n15304 = x108 & n6303 ;
  assign n15305 = n15303 | n15304 ;
  assign n15306 = ( x53 & n15300 ) | ( x53 & ~n15305 ) | ( n15300 & ~n15305 ) ;
  assign n15307 = ( ~x53 & n15305 ) | ( ~x53 & n15306 ) | ( n15305 & n15306 ) ;
  assign n15308 = ( ~n15300 & n15306 ) | ( ~n15300 & n15307 ) | ( n15306 & n15307 ) ;
  assign n15309 = ( n15191 & ~n15299 ) | ( n15191 & n15308 ) | ( ~n15299 & n15308 ) ;
  assign n15310 = ( n15191 & n15299 ) | ( n15191 & n15308 ) | ( n15299 & n15308 ) ;
  assign n15311 = ( n15299 & n15309 ) | ( n15299 & ~n15310 ) | ( n15309 & ~n15310 ) ;
  assign n15312 = ( n15194 & n15260 ) | ( n15194 & ~n15311 ) | ( n15260 & ~n15311 ) ;
  assign n15313 = ( ~n15194 & n15260 ) | ( ~n15194 & n15311 ) | ( n15260 & n15311 ) ;
  assign n15314 = ( ~n15260 & n15312 ) | ( ~n15260 & n15313 ) | ( n15312 & n15313 ) ;
  assign n15315 = n4787 & n5977 ;
  assign n15316 = x115 & n4791 ;
  assign n15317 = x116 | n15316 ;
  assign n15318 = ( n4793 & n15316 ) | ( n4793 & n15317 ) | ( n15316 & n15317 ) ;
  assign n15319 = x114 & n5030 ;
  assign n15320 = n15318 | n15319 ;
  assign n15321 = ( x47 & n15315 ) | ( x47 & ~n15320 ) | ( n15315 & ~n15320 ) ;
  assign n15322 = ( ~x47 & n15320 ) | ( ~x47 & n15321 ) | ( n15320 & n15321 ) ;
  assign n15323 = ( ~n15315 & n15321 ) | ( ~n15315 & n15322 ) | ( n15321 & n15322 ) ;
  assign n15324 = ( n15197 & ~n15314 ) | ( n15197 & n15323 ) | ( ~n15314 & n15323 ) ;
  assign n15325 = ( n15197 & n15314 ) | ( n15197 & n15323 ) | ( n15314 & n15323 ) ;
  assign n15326 = ( n15314 & n15324 ) | ( n15314 & ~n15325 ) | ( n15324 & ~n15325 ) ;
  assign n15327 = ( n15200 & n15251 ) | ( n15200 & ~n15326 ) | ( n15251 & ~n15326 ) ;
  assign n15328 = ( ~n15200 & n15251 ) | ( ~n15200 & n15326 ) | ( n15251 & n15326 ) ;
  assign n15329 = ( ~n15251 & n15327 ) | ( ~n15251 & n15328 ) | ( n15327 & n15328 ) ;
  assign n15330 = ( n15203 & n15242 ) | ( n15203 & ~n15329 ) | ( n15242 & ~n15329 ) ;
  assign n15331 = ( ~n15203 & n15242 ) | ( ~n15203 & n15329 ) | ( n15242 & n15329 ) ;
  assign n15332 = ( ~n15242 & n15330 ) | ( ~n15242 & n15331 ) | ( n15330 & n15331 ) ;
  assign n15333 = n3224 & n8331 ;
  assign n15334 = x124 & n3228 ;
  assign n15335 = x125 | n15334 ;
  assign n15336 = ( n3230 & n15334 ) | ( n3230 & n15335 ) | ( n15334 & n15335 ) ;
  assign n15337 = x123 & n3413 ;
  assign n15338 = n15336 | n15337 ;
  assign n15339 = ( x38 & n15333 ) | ( x38 & ~n15338 ) | ( n15333 & ~n15338 ) ;
  assign n15340 = ( ~x38 & n15338 ) | ( ~x38 & n15339 ) | ( n15338 & n15339 ) ;
  assign n15341 = ( ~n15333 & n15339 ) | ( ~n15333 & n15340 ) | ( n15339 & n15340 ) ;
  assign n15342 = ( n15206 & ~n15332 ) | ( n15206 & n15341 ) | ( ~n15332 & n15341 ) ;
  assign n15343 = ( n15206 & n15332 ) | ( n15206 & n15341 ) | ( n15332 & n15341 ) ;
  assign n15344 = ( n15332 & n15342 ) | ( n15332 & ~n15343 ) | ( n15342 & ~n15343 ) ;
  assign n15345 = ( n15209 & n15233 ) | ( n15209 & ~n15344 ) | ( n15233 & ~n15344 ) ;
  assign n15346 = ( ~n15209 & n15233 ) | ( ~n15209 & n15344 ) | ( n15233 & n15344 ) ;
  assign n15347 = ( ~n15233 & n15345 ) | ( ~n15233 & n15346 ) | ( n15345 & n15346 ) ;
  assign n15348 = ( ~n15221 & n15224 ) | ( ~n15221 & n15347 ) | ( n15224 & n15347 ) ;
  assign n15349 = ( n15224 & n15347 ) | ( n15224 & ~n15348 ) | ( n15347 & ~n15348 ) ;
  assign n15350 = ( n15221 & n15348 ) | ( n15221 & ~n15349 ) | ( n15348 & ~n15349 ) ;
  assign n15351 = n2766 & n8862 ;
  assign n15352 = ( x127 & n2943 ) | ( x127 & n15351 ) | ( n2943 & n15351 ) ;
  assign n15353 = x35 | n15352 ;
  assign n15354 = ~x35 & n15352 ;
  assign n15355 = ( ~n15352 & n15353 ) | ( ~n15352 & n15354 ) | ( n15353 & n15354 ) ;
  assign n15356 = n3715 & n7597 ;
  assign n15357 = x122 & n3719 ;
  assign n15358 = x123 | n15357 ;
  assign n15359 = ( n3721 & n15357 ) | ( n3721 & n15358 ) | ( n15357 & n15358 ) ;
  assign n15360 = x121 & n3922 ;
  assign n15361 = n15359 | n15360 ;
  assign n15362 = ( x41 & n15356 ) | ( x41 & ~n15361 ) | ( n15356 & ~n15361 ) ;
  assign n15363 = ( ~x41 & n15361 ) | ( ~x41 & n15362 ) | ( n15361 & n15362 ) ;
  assign n15364 = ( ~n15356 & n15362 ) | ( ~n15356 & n15363 ) | ( n15362 & n15363 ) ;
  assign n15365 = n4227 & n7098 ;
  assign n15366 = x119 & n4231 ;
  assign n15367 = x120 | n15366 ;
  assign n15368 = ( n4233 & n15366 ) | ( n4233 & n15367 ) | ( n15366 & n15367 ) ;
  assign n15369 = x118 & n4470 ;
  assign n15370 = n15368 | n15369 ;
  assign n15371 = ( x44 & n15365 ) | ( x44 & ~n15370 ) | ( n15365 & ~n15370 ) ;
  assign n15372 = ( ~x44 & n15370 ) | ( ~x44 & n15371 ) | ( n15370 & n15371 ) ;
  assign n15373 = ( ~n15365 & n15371 ) | ( ~n15365 & n15372 ) | ( n15371 & n15372 ) ;
  assign n15374 = n4787 & n6201 ;
  assign n15375 = x116 & n4791 ;
  assign n15376 = x117 | n15375 ;
  assign n15377 = ( n4793 & n15375 ) | ( n4793 & n15376 ) | ( n15375 & n15376 ) ;
  assign n15378 = x115 & n5030 ;
  assign n15379 = n15377 | n15378 ;
  assign n15380 = ( x47 & n15374 ) | ( x47 & ~n15379 ) | ( n15374 & ~n15379 ) ;
  assign n15381 = ( ~x47 & n15379 ) | ( ~x47 & n15380 ) | ( n15379 & n15380 ) ;
  assign n15382 = ( ~n15374 & n15380 ) | ( ~n15374 & n15381 ) | ( n15380 & n15381 ) ;
  assign n15383 = n5374 & n5750 ;
  assign n15384 = x113 & n5378 ;
  assign n15385 = x114 | n15384 ;
  assign n15386 = ( n5380 & n15384 ) | ( n5380 & n15385 ) | ( n15384 & n15385 ) ;
  assign n15387 = x112 & n5638 ;
  assign n15388 = n15386 | n15387 ;
  assign n15389 = ( x50 & n15383 ) | ( x50 & ~n15388 ) | ( n15383 & ~n15388 ) ;
  assign n15390 = ( ~x50 & n15388 ) | ( ~x50 & n15389 ) | ( n15388 & n15389 ) ;
  assign n15391 = ( ~n15383 & n15389 ) | ( ~n15383 & n15390 ) | ( n15389 & n15390 ) ;
  assign n15392 = n4377 & n6713 ;
  assign n15393 = x107 & n6717 ;
  assign n15394 = x108 | n15393 ;
  assign n15395 = ( n6719 & n15393 ) | ( n6719 & n15394 ) | ( n15393 & n15394 ) ;
  assign n15396 = x106 & n6980 ;
  assign n15397 = n15395 | n15396 ;
  assign n15398 = ( x56 & n15392 ) | ( x56 & ~n15397 ) | ( n15392 & ~n15397 ) ;
  assign n15399 = ( ~x56 & n15397 ) | ( ~x56 & n15398 ) | ( n15397 & n15398 ) ;
  assign n15400 = ( ~n15392 & n15398 ) | ( ~n15392 & n15399 ) | ( n15398 & n15399 ) ;
  assign n15401 = x98 & n8927 ;
  assign n15402 = ( ~x99 & n8693 ) | ( ~x99 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15403 = ( n8693 & n15401 ) | ( n8693 & ~n15402 ) | ( n15401 & ~n15402 ) ;
  assign n15404 = ( n15182 & n15291 ) | ( n15182 & ~n15403 ) | ( n15291 & ~n15403 ) ;
  assign n15405 = ( n15182 & ~n15291 ) | ( n15182 & n15403 ) | ( ~n15291 & n15403 ) ;
  assign n15406 = ( ~n15182 & n15404 ) | ( ~n15182 & n15405 ) | ( n15404 & n15405 ) ;
  assign n15407 = n3998 & n7423 ;
  assign n15408 = x104 & n7427 ;
  assign n15409 = x105 | n15408 ;
  assign n15410 = ( n7429 & n15408 ) | ( n7429 & n15409 ) | ( n15408 & n15409 ) ;
  assign n15411 = x103 & n7708 ;
  assign n15412 = n15410 | n15411 ;
  assign n15413 = ( x59 & n15407 ) | ( x59 & ~n15412 ) | ( n15407 & ~n15412 ) ;
  assign n15414 = ( ~x59 & n15412 ) | ( ~x59 & n15413 ) | ( n15412 & n15413 ) ;
  assign n15415 = ( ~n15407 & n15413 ) | ( ~n15407 & n15414 ) | ( n15413 & n15414 ) ;
  assign n15416 = n3486 & n8154 ;
  assign n15417 = x101 & n8158 ;
  assign n15418 = x102 | n15417 ;
  assign n15419 = ( n8160 & n15417 ) | ( n8160 & n15418 ) | ( n15417 & n15418 ) ;
  assign n15420 = x100 & n8439 ;
  assign n15421 = n15419 | n15420 ;
  assign n15422 = ( x62 & n15416 ) | ( x62 & ~n15421 ) | ( n15416 & ~n15421 ) ;
  assign n15423 = ( ~x62 & n15421 ) | ( ~x62 & n15422 ) | ( n15421 & n15422 ) ;
  assign n15424 = ( ~n15416 & n15422 ) | ( ~n15416 & n15423 ) | ( n15422 & n15423 ) ;
  assign n15425 = ( ~n15406 & n15415 ) | ( ~n15406 & n15424 ) | ( n15415 & n15424 ) ;
  assign n15426 = ( n15415 & n15424 ) | ( n15415 & ~n15425 ) | ( n15424 & ~n15425 ) ;
  assign n15427 = ( n15406 & n15425 ) | ( n15406 & ~n15426 ) | ( n15425 & ~n15426 ) ;
  assign n15428 = ( n15294 & n15400 ) | ( n15294 & ~n15427 ) | ( n15400 & ~n15427 ) ;
  assign n15429 = ( ~n15294 & n15400 ) | ( ~n15294 & n15427 ) | ( n15400 & n15427 ) ;
  assign n15430 = ( ~n15400 & n15428 ) | ( ~n15400 & n15429 ) | ( n15428 & n15429 ) ;
  assign n15431 = n5130 & n6027 ;
  assign n15432 = x110 & n6031 ;
  assign n15433 = x111 | n15432 ;
  assign n15434 = ( n6033 & n15432 ) | ( n6033 & n15433 ) | ( n15432 & n15433 ) ;
  assign n15435 = x109 & n6303 ;
  assign n15436 = n15434 | n15435 ;
  assign n15437 = ( x53 & n15431 ) | ( x53 & ~n15436 ) | ( n15431 & ~n15436 ) ;
  assign n15438 = ( ~x53 & n15436 ) | ( ~x53 & n15437 ) | ( n15436 & n15437 ) ;
  assign n15439 = ( ~n15431 & n15437 ) | ( ~n15431 & n15438 ) | ( n15437 & n15438 ) ;
  assign n15440 = ( n15297 & ~n15430 ) | ( n15297 & n15439 ) | ( ~n15430 & n15439 ) ;
  assign n15441 = ( n15297 & n15430 ) | ( n15297 & n15439 ) | ( n15430 & n15439 ) ;
  assign n15442 = ( n15430 & n15440 ) | ( n15430 & ~n15441 ) | ( n15440 & ~n15441 ) ;
  assign n15443 = ( n15309 & n15391 ) | ( n15309 & ~n15442 ) | ( n15391 & ~n15442 ) ;
  assign n15444 = ( ~n15309 & n15391 ) | ( ~n15309 & n15442 ) | ( n15391 & n15442 ) ;
  assign n15445 = ( ~n15391 & n15443 ) | ( ~n15391 & n15444 ) | ( n15443 & n15444 ) ;
  assign n15446 = ( n15312 & n15382 ) | ( n15312 & ~n15445 ) | ( n15382 & ~n15445 ) ;
  assign n15447 = ( ~n15312 & n15382 ) | ( ~n15312 & n15445 ) | ( n15382 & n15445 ) ;
  assign n15448 = ( ~n15382 & n15446 ) | ( ~n15382 & n15447 ) | ( n15446 & n15447 ) ;
  assign n15449 = ( n15324 & n15373 ) | ( n15324 & ~n15448 ) | ( n15373 & ~n15448 ) ;
  assign n15450 = ( ~n15324 & n15373 ) | ( ~n15324 & n15448 ) | ( n15373 & n15448 ) ;
  assign n15451 = ( ~n15373 & n15449 ) | ( ~n15373 & n15450 ) | ( n15449 & n15450 ) ;
  assign n15452 = ( n15327 & n15364 ) | ( n15327 & ~n15451 ) | ( n15364 & ~n15451 ) ;
  assign n15453 = ( ~n15327 & n15364 ) | ( ~n15327 & n15451 ) | ( n15364 & n15451 ) ;
  assign n15454 = ( ~n15364 & n15452 ) | ( ~n15364 & n15453 ) | ( n15452 & n15453 ) ;
  assign n15455 = n3224 & n8587 ;
  assign n15456 = x125 & n3228 ;
  assign n15457 = x126 | n15456 ;
  assign n15458 = ( n3230 & n15456 ) | ( n3230 & n15457 ) | ( n15456 & n15457 ) ;
  assign n15459 = x124 & n3413 ;
  assign n15460 = n15458 | n15459 ;
  assign n15461 = ( x38 & n15455 ) | ( x38 & ~n15460 ) | ( n15455 & ~n15460 ) ;
  assign n15462 = ( ~x38 & n15460 ) | ( ~x38 & n15461 ) | ( n15460 & n15461 ) ;
  assign n15463 = ( ~n15455 & n15461 ) | ( ~n15455 & n15462 ) | ( n15461 & n15462 ) ;
  assign n15464 = ( n15330 & ~n15454 ) | ( n15330 & n15463 ) | ( ~n15454 & n15463 ) ;
  assign n15465 = ( n15330 & n15454 ) | ( n15330 & n15463 ) | ( n15454 & n15463 ) ;
  assign n15466 = ( n15454 & n15464 ) | ( n15454 & ~n15465 ) | ( n15464 & ~n15465 ) ;
  assign n15467 = ( n15342 & n15355 ) | ( n15342 & ~n15466 ) | ( n15355 & ~n15466 ) ;
  assign n15468 = ( ~n15342 & n15355 ) | ( ~n15342 & n15466 ) | ( n15355 & n15466 ) ;
  assign n15469 = ( ~n15355 & n15467 ) | ( ~n15355 & n15468 ) | ( n15467 & n15468 ) ;
  assign n15470 = ( ~n15345 & n15348 ) | ( ~n15345 & n15469 ) | ( n15348 & n15469 ) ;
  assign n15471 = ( n15348 & n15469 ) | ( n15348 & ~n15470 ) | ( n15469 & ~n15470 ) ;
  assign n15472 = ( n15345 & n15470 ) | ( n15345 & ~n15471 ) | ( n15470 & ~n15471 ) ;
  assign n15473 = n3224 & n8846 ;
  assign n15474 = x126 & n3228 ;
  assign n15475 = x127 | n15474 ;
  assign n15476 = ( n3230 & n15474 ) | ( n3230 & n15475 ) | ( n15474 & n15475 ) ;
  assign n15477 = x125 & n3413 ;
  assign n15478 = n15476 | n15477 ;
  assign n15479 = ( x38 & n15473 ) | ( x38 & ~n15478 ) | ( n15473 & ~n15478 ) ;
  assign n15480 = ( ~x38 & n15478 ) | ( ~x38 & n15479 ) | ( n15478 & n15479 ) ;
  assign n15481 = ( ~n15473 & n15479 ) | ( ~n15473 & n15480 ) | ( n15479 & n15480 ) ;
  assign n15482 = n3715 & n7841 ;
  assign n15483 = x123 & n3719 ;
  assign n15484 = x124 | n15483 ;
  assign n15485 = ( n3721 & n15483 ) | ( n3721 & n15484 ) | ( n15483 & n15484 ) ;
  assign n15486 = x122 & n3922 ;
  assign n15487 = n15485 | n15486 ;
  assign n15488 = ( x41 & n15482 ) | ( x41 & ~n15487 ) | ( n15482 & ~n15487 ) ;
  assign n15489 = ( ~x41 & n15487 ) | ( ~x41 & n15488 ) | ( n15487 & n15488 ) ;
  assign n15490 = ( ~n15482 & n15488 ) | ( ~n15482 & n15489 ) | ( n15488 & n15489 ) ;
  assign n15491 = n4227 & n7113 ;
  assign n15492 = x120 & n4231 ;
  assign n15493 = x121 | n15492 ;
  assign n15494 = ( n4233 & n15492 ) | ( n4233 & n15493 ) | ( n15492 & n15493 ) ;
  assign n15495 = x119 & n4470 ;
  assign n15496 = n15494 | n15495 ;
  assign n15497 = ( x44 & n15491 ) | ( x44 & ~n15496 ) | ( n15491 & ~n15496 ) ;
  assign n15498 = ( ~x44 & n15496 ) | ( ~x44 & n15497 ) | ( n15496 & n15497 ) ;
  assign n15499 = ( ~n15491 & n15497 ) | ( ~n15491 & n15498 ) | ( n15497 & n15498 ) ;
  assign n15500 = n4787 & n6421 ;
  assign n15501 = x117 & n4791 ;
  assign n15502 = x118 | n15501 ;
  assign n15503 = ( n4793 & n15501 ) | ( n4793 & n15502 ) | ( n15501 & n15502 ) ;
  assign n15504 = x116 & n5030 ;
  assign n15505 = n15503 | n15504 ;
  assign n15506 = ( x47 & n15500 ) | ( x47 & ~n15505 ) | ( n15500 & ~n15505 ) ;
  assign n15507 = ( ~x47 & n15505 ) | ( ~x47 & n15506 ) | ( n15505 & n15506 ) ;
  assign n15508 = ( ~n15500 & n15506 ) | ( ~n15500 & n15507 ) | ( n15506 & n15507 ) ;
  assign n15509 = n5374 & n5765 ;
  assign n15510 = x114 & n5378 ;
  assign n15511 = x115 | n15510 ;
  assign n15512 = ( n5380 & n15510 ) | ( n5380 & n15511 ) | ( n15510 & n15511 ) ;
  assign n15513 = x113 & n5638 ;
  assign n15514 = n15512 | n15513 ;
  assign n15515 = ( x50 & n15509 ) | ( x50 & ~n15514 ) | ( n15509 & ~n15514 ) ;
  assign n15516 = ( ~x50 & n15514 ) | ( ~x50 & n15515 ) | ( n15514 & n15515 ) ;
  assign n15517 = ( ~n15509 & n15515 ) | ( ~n15509 & n15516 ) | ( n15515 & n15516 ) ;
  assign n15518 = n5145 & n6027 ;
  assign n15519 = x111 & n6031 ;
  assign n15520 = x112 | n15519 ;
  assign n15521 = ( n6033 & n15519 ) | ( n6033 & n15520 ) | ( n15519 & n15520 ) ;
  assign n15522 = x110 & n6303 ;
  assign n15523 = n15521 | n15522 ;
  assign n15524 = ( x53 & n15518 ) | ( x53 & ~n15523 ) | ( n15518 & ~n15523 ) ;
  assign n15525 = ( ~x53 & n15523 ) | ( ~x53 & n15524 ) | ( n15523 & n15524 ) ;
  assign n15526 = ( ~n15518 & n15524 ) | ( ~n15518 & n15525 ) | ( n15524 & n15525 ) ;
  assign n15527 = n4734 & n6713 ;
  assign n15528 = x108 & n6717 ;
  assign n15529 = x109 | n15528 ;
  assign n15530 = ( n6719 & n15528 ) | ( n6719 & n15529 ) | ( n15528 & n15529 ) ;
  assign n15531 = x107 & n6980 ;
  assign n15532 = n15530 | n15531 ;
  assign n15533 = ( x56 & n15527 ) | ( x56 & ~n15532 ) | ( n15527 & ~n15532 ) ;
  assign n15534 = ( ~x56 & n15532 ) | ( ~x56 & n15533 ) | ( n15532 & n15533 ) ;
  assign n15535 = ( ~n15527 & n15533 ) | ( ~n15527 & n15534 ) | ( n15533 & n15534 ) ;
  assign n15536 = n4013 & n7423 ;
  assign n15537 = x105 & n7427 ;
  assign n15538 = x106 | n15537 ;
  assign n15539 = ( n7429 & n15537 ) | ( n7429 & n15538 ) | ( n15537 & n15538 ) ;
  assign n15540 = x104 & n7708 ;
  assign n15541 = n15539 | n15540 ;
  assign n15542 = ( x59 & n15536 ) | ( x59 & ~n15541 ) | ( n15536 & ~n15541 ) ;
  assign n15543 = ( ~x59 & n15541 ) | ( ~x59 & n15542 ) | ( n15541 & n15542 ) ;
  assign n15544 = ( ~n15536 & n15542 ) | ( ~n15536 & n15543 ) | ( n15542 & n15543 ) ;
  assign n15545 = n3650 & n8154 ;
  assign n15546 = x102 & n8158 ;
  assign n15547 = x103 | n15546 ;
  assign n15548 = ( n8160 & n15546 ) | ( n8160 & n15547 ) | ( n15546 & n15547 ) ;
  assign n15549 = x101 & n8439 ;
  assign n15550 = n15548 | n15549 ;
  assign n15551 = ( x62 & n15545 ) | ( x62 & ~n15550 ) | ( n15545 & ~n15550 ) ;
  assign n15552 = ( ~x62 & n15550 ) | ( ~x62 & n15551 ) | ( n15550 & n15551 ) ;
  assign n15553 = ( ~n15545 & n15551 ) | ( ~n15545 & n15552 ) | ( n15551 & n15552 ) ;
  assign n15554 = x99 & n8927 ;
  assign n15555 = ( ~x100 & n8693 ) | ( ~x100 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15556 = ( n8693 & n15554 ) | ( n8693 & ~n15555 ) | ( n15554 & ~n15555 ) ;
  assign n15557 = ( ~x35 & n15403 ) | ( ~x35 & n15556 ) | ( n15403 & n15556 ) ;
  assign n15558 = ( n15403 & n15556 ) | ( n15403 & ~n15557 ) | ( n15556 & ~n15557 ) ;
  assign n15559 = ( x35 & n15557 ) | ( x35 & ~n15558 ) | ( n15557 & ~n15558 ) ;
  assign n15560 = ( n15404 & n15553 ) | ( n15404 & ~n15559 ) | ( n15553 & ~n15559 ) ;
  assign n15561 = ( ~n15404 & n15553 ) | ( ~n15404 & n15559 ) | ( n15553 & n15559 ) ;
  assign n15562 = ( ~n15553 & n15560 ) | ( ~n15553 & n15561 ) | ( n15560 & n15561 ) ;
  assign n15563 = ( n15425 & n15544 ) | ( n15425 & ~n15562 ) | ( n15544 & ~n15562 ) ;
  assign n15564 = ( ~n15425 & n15544 ) | ( ~n15425 & n15562 ) | ( n15544 & n15562 ) ;
  assign n15565 = ( ~n15544 & n15563 ) | ( ~n15544 & n15564 ) | ( n15563 & n15564 ) ;
  assign n15566 = ( n15428 & n15535 ) | ( n15428 & ~n15565 ) | ( n15535 & ~n15565 ) ;
  assign n15567 = ( ~n15428 & n15535 ) | ( ~n15428 & n15565 ) | ( n15535 & n15565 ) ;
  assign n15568 = ( ~n15535 & n15566 ) | ( ~n15535 & n15567 ) | ( n15566 & n15567 ) ;
  assign n15569 = ( n15440 & n15526 ) | ( n15440 & ~n15568 ) | ( n15526 & ~n15568 ) ;
  assign n15570 = ( ~n15440 & n15526 ) | ( ~n15440 & n15568 ) | ( n15526 & n15568 ) ;
  assign n15571 = ( ~n15526 & n15569 ) | ( ~n15526 & n15570 ) | ( n15569 & n15570 ) ;
  assign n15572 = ( n15443 & n15517 ) | ( n15443 & ~n15571 ) | ( n15517 & ~n15571 ) ;
  assign n15573 = ( ~n15443 & n15517 ) | ( ~n15443 & n15571 ) | ( n15517 & n15571 ) ;
  assign n15574 = ( ~n15517 & n15572 ) | ( ~n15517 & n15573 ) | ( n15572 & n15573 ) ;
  assign n15575 = ( n15446 & n15508 ) | ( n15446 & ~n15574 ) | ( n15508 & ~n15574 ) ;
  assign n15576 = ( ~n15446 & n15508 ) | ( ~n15446 & n15574 ) | ( n15508 & n15574 ) ;
  assign n15577 = ( ~n15508 & n15575 ) | ( ~n15508 & n15576 ) | ( n15575 & n15576 ) ;
  assign n15578 = ( n15449 & n15499 ) | ( n15449 & ~n15577 ) | ( n15499 & ~n15577 ) ;
  assign n15579 = ( ~n15449 & n15499 ) | ( ~n15449 & n15577 ) | ( n15499 & n15577 ) ;
  assign n15580 = ( ~n15499 & n15578 ) | ( ~n15499 & n15579 ) | ( n15578 & n15579 ) ;
  assign n15581 = ( n15452 & n15490 ) | ( n15452 & ~n15580 ) | ( n15490 & ~n15580 ) ;
  assign n15582 = ( ~n15452 & n15490 ) | ( ~n15452 & n15580 ) | ( n15490 & n15580 ) ;
  assign n15583 = ( ~n15490 & n15581 ) | ( ~n15490 & n15582 ) | ( n15581 & n15582 ) ;
  assign n15584 = ( n15464 & n15481 ) | ( n15464 & ~n15583 ) | ( n15481 & ~n15583 ) ;
  assign n15585 = ( ~n15464 & n15481 ) | ( ~n15464 & n15583 ) | ( n15481 & n15583 ) ;
  assign n15586 = ( ~n15481 & n15584 ) | ( ~n15481 & n15585 ) | ( n15584 & n15585 ) ;
  assign n15587 = ( ~n15467 & n15470 ) | ( ~n15467 & n15586 ) | ( n15470 & n15586 ) ;
  assign n15588 = ( n15470 & n15586 ) | ( n15470 & ~n15587 ) | ( n15586 & ~n15587 ) ;
  assign n15589 = ( n15467 & n15587 ) | ( n15467 & ~n15588 ) | ( n15587 & ~n15588 ) ;
  assign n15590 = n3224 & n8865 ;
  assign n15591 = x127 & n3228 ;
  assign n15592 = x126 | n15591 ;
  assign n15593 = ( n3413 & n15591 ) | ( n3413 & n15592 ) | ( n15591 & n15592 ) ;
  assign n15594 = ( x38 & n15590 ) | ( x38 & ~n15593 ) | ( n15590 & ~n15593 ) ;
  assign n15595 = ( ~x38 & n15593 ) | ( ~x38 & n15594 ) | ( n15593 & n15594 ) ;
  assign n15596 = ( ~n15590 & n15594 ) | ( ~n15590 & n15595 ) | ( n15594 & n15595 ) ;
  assign n15597 = n3715 & n8331 ;
  assign n15598 = x124 & n3719 ;
  assign n15599 = x125 | n15598 ;
  assign n15600 = ( n3721 & n15598 ) | ( n3721 & n15599 ) | ( n15598 & n15599 ) ;
  assign n15601 = x123 & n3922 ;
  assign n15602 = n15600 | n15601 ;
  assign n15603 = ( x41 & n15597 ) | ( x41 & ~n15602 ) | ( n15597 & ~n15602 ) ;
  assign n15604 = ( ~x41 & n15602 ) | ( ~x41 & n15603 ) | ( n15602 & n15603 ) ;
  assign n15605 = ( ~n15597 & n15603 ) | ( ~n15597 & n15604 ) | ( n15603 & n15604 ) ;
  assign n15606 = n4787 & n6645 ;
  assign n15607 = x118 & n4791 ;
  assign n15608 = x119 | n15607 ;
  assign n15609 = ( n4793 & n15607 ) | ( n4793 & n15608 ) | ( n15607 & n15608 ) ;
  assign n15610 = x117 & n5030 ;
  assign n15611 = n15609 | n15610 ;
  assign n15612 = ( x47 & n15606 ) | ( x47 & ~n15611 ) | ( n15606 & ~n15611 ) ;
  assign n15613 = ( ~x47 & n15611 ) | ( ~x47 & n15612 ) | ( n15611 & n15612 ) ;
  assign n15614 = ( ~n15606 & n15612 ) | ( ~n15606 & n15613 ) | ( n15612 & n15613 ) ;
  assign n15615 = n5542 & n6027 ;
  assign n15616 = x112 & n6031 ;
  assign n15617 = x113 | n15616 ;
  assign n15618 = ( n6033 & n15616 ) | ( n6033 & n15617 ) | ( n15616 & n15617 ) ;
  assign n15619 = x111 & n6303 ;
  assign n15620 = n15618 | n15619 ;
  assign n15621 = ( x53 & n15615 ) | ( x53 & ~n15620 ) | ( n15615 & ~n15620 ) ;
  assign n15622 = ( ~x53 & n15620 ) | ( ~x53 & n15621 ) | ( n15620 & n15621 ) ;
  assign n15623 = ( ~n15615 & n15621 ) | ( ~n15615 & n15622 ) | ( n15621 & n15622 ) ;
  assign n15624 = n4362 & n7423 ;
  assign n15625 = x106 & n7427 ;
  assign n15626 = x107 | n15625 ;
  assign n15627 = ( n7429 & n15625 ) | ( n7429 & n15626 ) | ( n15625 & n15626 ) ;
  assign n15628 = x105 & n7708 ;
  assign n15629 = n15627 | n15628 ;
  assign n15630 = ( x59 & n15624 ) | ( x59 & ~n15629 ) | ( n15624 & ~n15629 ) ;
  assign n15631 = ( ~x59 & n15629 ) | ( ~x59 & n15630 ) | ( n15629 & n15630 ) ;
  assign n15632 = ( ~n15624 & n15630 ) | ( ~n15624 & n15631 ) | ( n15630 & n15631 ) ;
  assign n15633 = n3665 & n8154 ;
  assign n15634 = x103 & n8158 ;
  assign n15635 = x104 | n15634 ;
  assign n15636 = ( n8160 & n15634 ) | ( n8160 & n15635 ) | ( n15634 & n15635 ) ;
  assign n15637 = x102 & n8439 ;
  assign n15638 = n15636 | n15637 ;
  assign n15639 = ( x62 & n15633 ) | ( x62 & ~n15638 ) | ( n15633 & ~n15638 ) ;
  assign n15640 = ( ~x62 & n15638 ) | ( ~x62 & n15639 ) | ( n15638 & n15639 ) ;
  assign n15641 = ( ~n15633 & n15639 ) | ( ~n15633 & n15640 ) | ( n15639 & n15640 ) ;
  assign n15642 = x100 & n8927 ;
  assign n15643 = ( ~x101 & n8693 ) | ( ~x101 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15644 = ( n8693 & n15642 ) | ( n8693 & ~n15643 ) | ( n15642 & ~n15643 ) ;
  assign n15645 = ( n15557 & n15641 ) | ( n15557 & ~n15644 ) | ( n15641 & ~n15644 ) ;
  assign n15646 = ( ~n15557 & n15641 ) | ( ~n15557 & n15644 ) | ( n15641 & n15644 ) ;
  assign n15647 = ( ~n15641 & n15645 ) | ( ~n15641 & n15646 ) | ( n15645 & n15646 ) ;
  assign n15648 = ( n15560 & n15632 ) | ( n15560 & ~n15647 ) | ( n15632 & ~n15647 ) ;
  assign n15649 = ( ~n15560 & n15632 ) | ( ~n15560 & n15647 ) | ( n15632 & n15647 ) ;
  assign n15650 = ( ~n15632 & n15648 ) | ( ~n15632 & n15649 ) | ( n15648 & n15649 ) ;
  assign n15651 = n4934 & n6713 ;
  assign n15652 = x109 & n6717 ;
  assign n15653 = x110 | n15652 ;
  assign n15654 = ( n6719 & n15652 ) | ( n6719 & n15653 ) | ( n15652 & n15653 ) ;
  assign n15655 = x108 & n6980 ;
  assign n15656 = n15654 | n15655 ;
  assign n15657 = ( x56 & n15651 ) | ( x56 & ~n15656 ) | ( n15651 & ~n15656 ) ;
  assign n15658 = ( ~x56 & n15656 ) | ( ~x56 & n15657 ) | ( n15656 & n15657 ) ;
  assign n15659 = ( ~n15651 & n15657 ) | ( ~n15651 & n15658 ) | ( n15657 & n15658 ) ;
  assign n15660 = ( n15563 & ~n15650 ) | ( n15563 & n15659 ) | ( ~n15650 & n15659 ) ;
  assign n15661 = ( n15563 & n15650 ) | ( n15563 & n15659 ) | ( n15650 & n15659 ) ;
  assign n15662 = ( n15650 & n15660 ) | ( n15650 & ~n15661 ) | ( n15660 & ~n15661 ) ;
  assign n15663 = ( n15566 & n15623 ) | ( n15566 & ~n15662 ) | ( n15623 & ~n15662 ) ;
  assign n15664 = ( ~n15566 & n15623 ) | ( ~n15566 & n15662 ) | ( n15623 & n15662 ) ;
  assign n15665 = ( ~n15623 & n15663 ) | ( ~n15623 & n15664 ) | ( n15663 & n15664 ) ;
  assign n15666 = n5374 & n5977 ;
  assign n15667 = x115 & n5378 ;
  assign n15668 = x116 | n15667 ;
  assign n15669 = ( n5380 & n15667 ) | ( n5380 & n15668 ) | ( n15667 & n15668 ) ;
  assign n15670 = x114 & n5638 ;
  assign n15671 = n15669 | n15670 ;
  assign n15672 = ( x50 & n15666 ) | ( x50 & ~n15671 ) | ( n15666 & ~n15671 ) ;
  assign n15673 = ( ~x50 & n15671 ) | ( ~x50 & n15672 ) | ( n15671 & n15672 ) ;
  assign n15674 = ( ~n15666 & n15672 ) | ( ~n15666 & n15673 ) | ( n15672 & n15673 ) ;
  assign n15675 = ( n15569 & ~n15665 ) | ( n15569 & n15674 ) | ( ~n15665 & n15674 ) ;
  assign n15676 = ( n15569 & n15665 ) | ( n15569 & n15674 ) | ( n15665 & n15674 ) ;
  assign n15677 = ( n15665 & n15675 ) | ( n15665 & ~n15676 ) | ( n15675 & ~n15676 ) ;
  assign n15678 = ( n15572 & n15614 ) | ( n15572 & ~n15677 ) | ( n15614 & ~n15677 ) ;
  assign n15679 = ( ~n15572 & n15614 ) | ( ~n15572 & n15677 ) | ( n15614 & n15677 ) ;
  assign n15680 = ( ~n15614 & n15678 ) | ( ~n15614 & n15679 ) | ( n15678 & n15679 ) ;
  assign n15681 = n4227 & n7582 ;
  assign n15682 = x121 & n4231 ;
  assign n15683 = x122 | n15682 ;
  assign n15684 = ( n4233 & n15682 ) | ( n4233 & n15683 ) | ( n15682 & n15683 ) ;
  assign n15685 = x120 & n4470 ;
  assign n15686 = n15684 | n15685 ;
  assign n15687 = ( x44 & n15681 ) | ( x44 & ~n15686 ) | ( n15681 & ~n15686 ) ;
  assign n15688 = ( ~x44 & n15686 ) | ( ~x44 & n15687 ) | ( n15686 & n15687 ) ;
  assign n15689 = ( ~n15681 & n15687 ) | ( ~n15681 & n15688 ) | ( n15687 & n15688 ) ;
  assign n15690 = ( n15575 & ~n15680 ) | ( n15575 & n15689 ) | ( ~n15680 & n15689 ) ;
  assign n15691 = ( n15575 & n15680 ) | ( n15575 & n15689 ) | ( n15680 & n15689 ) ;
  assign n15692 = ( n15680 & n15690 ) | ( n15680 & ~n15691 ) | ( n15690 & ~n15691 ) ;
  assign n15693 = ( n15578 & n15605 ) | ( n15578 & ~n15692 ) | ( n15605 & ~n15692 ) ;
  assign n15694 = ( ~n15578 & n15605 ) | ( ~n15578 & n15692 ) | ( n15605 & n15692 ) ;
  assign n15695 = ( ~n15605 & n15693 ) | ( ~n15605 & n15694 ) | ( n15693 & n15694 ) ;
  assign n15696 = ( n15581 & n15596 ) | ( n15581 & ~n15695 ) | ( n15596 & ~n15695 ) ;
  assign n15697 = ( ~n15581 & n15596 ) | ( ~n15581 & n15695 ) | ( n15596 & n15695 ) ;
  assign n15698 = ( ~n15596 & n15696 ) | ( ~n15596 & n15697 ) | ( n15696 & n15697 ) ;
  assign n15699 = ( ~n15584 & n15587 ) | ( ~n15584 & n15698 ) | ( n15587 & n15698 ) ;
  assign n15700 = ( n15587 & n15698 ) | ( n15587 & ~n15699 ) | ( n15698 & ~n15699 ) ;
  assign n15701 = ( n15584 & n15699 ) | ( n15584 & ~n15700 ) | ( n15699 & ~n15700 ) ;
  assign n15702 = n3224 & n8862 ;
  assign n15703 = ( x127 & n3413 ) | ( x127 & n15702 ) | ( n3413 & n15702 ) ;
  assign n15704 = x38 | n15703 ;
  assign n15705 = ~x38 & n15703 ;
  assign n15706 = ( ~n15703 & n15704 ) | ( ~n15703 & n15705 ) | ( n15704 & n15705 ) ;
  assign n15707 = n3715 & n8587 ;
  assign n15708 = x125 & n3719 ;
  assign n15709 = x126 | n15708 ;
  assign n15710 = ( n3721 & n15708 ) | ( n3721 & n15709 ) | ( n15708 & n15709 ) ;
  assign n15711 = x124 & n3922 ;
  assign n15712 = n15710 | n15711 ;
  assign n15713 = ( x41 & n15707 ) | ( x41 & ~n15712 ) | ( n15707 & ~n15712 ) ;
  assign n15714 = ( ~x41 & n15712 ) | ( ~x41 & n15713 ) | ( n15712 & n15713 ) ;
  assign n15715 = ( ~n15707 & n15713 ) | ( ~n15707 & n15714 ) | ( n15713 & n15714 ) ;
  assign n15716 = n4787 & n7098 ;
  assign n15717 = x119 & n4791 ;
  assign n15718 = x120 | n15717 ;
  assign n15719 = ( n4793 & n15717 ) | ( n4793 & n15718 ) | ( n15717 & n15718 ) ;
  assign n15720 = x118 & n5030 ;
  assign n15721 = n15719 | n15720 ;
  assign n15722 = ( x47 & n15716 ) | ( x47 & ~n15721 ) | ( n15716 & ~n15721 ) ;
  assign n15723 = ( ~x47 & n15721 ) | ( ~x47 & n15722 ) | ( n15721 & n15722 ) ;
  assign n15724 = ( ~n15716 & n15722 ) | ( ~n15716 & n15723 ) | ( n15722 & n15723 ) ;
  assign n15725 = n5374 & n6201 ;
  assign n15726 = x116 & n5378 ;
  assign n15727 = x117 | n15726 ;
  assign n15728 = ( n5380 & n15726 ) | ( n5380 & n15727 ) | ( n15726 & n15727 ) ;
  assign n15729 = x115 & n5638 ;
  assign n15730 = n15728 | n15729 ;
  assign n15731 = ( x50 & n15725 ) | ( x50 & ~n15730 ) | ( n15725 & ~n15730 ) ;
  assign n15732 = ( ~x50 & n15730 ) | ( ~x50 & n15731 ) | ( n15730 & n15731 ) ;
  assign n15733 = ( ~n15725 & n15731 ) | ( ~n15725 & n15732 ) | ( n15731 & n15732 ) ;
  assign n15734 = n5750 & n6027 ;
  assign n15735 = x113 & n6031 ;
  assign n15736 = x114 | n15735 ;
  assign n15737 = ( n6033 & n15735 ) | ( n6033 & n15736 ) | ( n15735 & n15736 ) ;
  assign n15738 = x112 & n6303 ;
  assign n15739 = n15737 | n15738 ;
  assign n15740 = ( x53 & n15734 ) | ( x53 & ~n15739 ) | ( n15734 & ~n15739 ) ;
  assign n15741 = ( ~x53 & n15739 ) | ( ~x53 & n15740 ) | ( n15739 & n15740 ) ;
  assign n15742 = ( ~n15734 & n15740 ) | ( ~n15734 & n15741 ) | ( n15740 & n15741 ) ;
  assign n15743 = x101 & n8927 ;
  assign n15744 = ( ~x102 & n8693 ) | ( ~x102 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15745 = ( n8693 & n15743 ) | ( n8693 & ~n15744 ) | ( n15743 & ~n15744 ) ;
  assign n15746 = ( ~n15644 & n15645 ) | ( ~n15644 & n15745 ) | ( n15645 & n15745 ) ;
  assign n15747 = ( n15644 & n15645 ) | ( n15644 & n15745 ) | ( n15645 & n15745 ) ;
  assign n15748 = ( n15644 & n15746 ) | ( n15644 & ~n15747 ) | ( n15746 & ~n15747 ) ;
  assign n15749 = n4377 & n7423 ;
  assign n15750 = x107 & n7427 ;
  assign n15751 = x108 | n15750 ;
  assign n15752 = ( n7429 & n15750 ) | ( n7429 & n15751 ) | ( n15750 & n15751 ) ;
  assign n15753 = x106 & n7708 ;
  assign n15754 = n15752 | n15753 ;
  assign n15755 = ( x59 & n15749 ) | ( x59 & ~n15754 ) | ( n15749 & ~n15754 ) ;
  assign n15756 = ( ~x59 & n15754 ) | ( ~x59 & n15755 ) | ( n15754 & n15755 ) ;
  assign n15757 = ( ~n15749 & n15755 ) | ( ~n15749 & n15756 ) | ( n15755 & n15756 ) ;
  assign n15758 = n3998 & n8154 ;
  assign n15759 = x104 & n8158 ;
  assign n15760 = x105 | n15759 ;
  assign n15761 = ( n8160 & n15759 ) | ( n8160 & n15760 ) | ( n15759 & n15760 ) ;
  assign n15762 = x103 & n8439 ;
  assign n15763 = n15761 | n15762 ;
  assign n15764 = ( x62 & n15758 ) | ( x62 & ~n15763 ) | ( n15758 & ~n15763 ) ;
  assign n15765 = ( ~x62 & n15763 ) | ( ~x62 & n15764 ) | ( n15763 & n15764 ) ;
  assign n15766 = ( ~n15758 & n15764 ) | ( ~n15758 & n15765 ) | ( n15764 & n15765 ) ;
  assign n15767 = ( ~n15748 & n15757 ) | ( ~n15748 & n15766 ) | ( n15757 & n15766 ) ;
  assign n15768 = ( n15757 & n15766 ) | ( n15757 & ~n15767 ) | ( n15766 & ~n15767 ) ;
  assign n15769 = ( n15748 & n15767 ) | ( n15748 & ~n15768 ) | ( n15767 & ~n15768 ) ;
  assign n15770 = n5130 & n6713 ;
  assign n15771 = x110 & n6717 ;
  assign n15772 = x111 | n15771 ;
  assign n15773 = ( n6719 & n15771 ) | ( n6719 & n15772 ) | ( n15771 & n15772 ) ;
  assign n15774 = x109 & n6980 ;
  assign n15775 = n15773 | n15774 ;
  assign n15776 = ( x56 & n15770 ) | ( x56 & ~n15775 ) | ( n15770 & ~n15775 ) ;
  assign n15777 = ( ~x56 & n15775 ) | ( ~x56 & n15776 ) | ( n15775 & n15776 ) ;
  assign n15778 = ( ~n15770 & n15776 ) | ( ~n15770 & n15777 ) | ( n15776 & n15777 ) ;
  assign n15779 = ( n15648 & ~n15769 ) | ( n15648 & n15778 ) | ( ~n15769 & n15778 ) ;
  assign n15780 = ( n15648 & n15769 ) | ( n15648 & n15778 ) | ( n15769 & n15778 ) ;
  assign n15781 = ( n15769 & n15779 ) | ( n15769 & ~n15780 ) | ( n15779 & ~n15780 ) ;
  assign n15782 = ( n15660 & n15742 ) | ( n15660 & ~n15781 ) | ( n15742 & ~n15781 ) ;
  assign n15783 = ( ~n15660 & n15742 ) | ( ~n15660 & n15781 ) | ( n15742 & n15781 ) ;
  assign n15784 = ( ~n15742 & n15782 ) | ( ~n15742 & n15783 ) | ( n15782 & n15783 ) ;
  assign n15785 = ( n15663 & n15733 ) | ( n15663 & ~n15784 ) | ( n15733 & ~n15784 ) ;
  assign n15786 = ( ~n15663 & n15733 ) | ( ~n15663 & n15784 ) | ( n15733 & n15784 ) ;
  assign n15787 = ( ~n15733 & n15785 ) | ( ~n15733 & n15786 ) | ( n15785 & n15786 ) ;
  assign n15788 = ( n15675 & n15724 ) | ( n15675 & ~n15787 ) | ( n15724 & ~n15787 ) ;
  assign n15789 = ( ~n15675 & n15724 ) | ( ~n15675 & n15787 ) | ( n15724 & n15787 ) ;
  assign n15790 = ( ~n15724 & n15788 ) | ( ~n15724 & n15789 ) | ( n15788 & n15789 ) ;
  assign n15791 = n4227 & n7597 ;
  assign n15792 = x122 & n4231 ;
  assign n15793 = x123 | n15792 ;
  assign n15794 = ( n4233 & n15792 ) | ( n4233 & n15793 ) | ( n15792 & n15793 ) ;
  assign n15795 = x121 & n4470 ;
  assign n15796 = n15794 | n15795 ;
  assign n15797 = ( x44 & n15791 ) | ( x44 & ~n15796 ) | ( n15791 & ~n15796 ) ;
  assign n15798 = ( ~x44 & n15796 ) | ( ~x44 & n15797 ) | ( n15796 & n15797 ) ;
  assign n15799 = ( ~n15791 & n15797 ) | ( ~n15791 & n15798 ) | ( n15797 & n15798 ) ;
  assign n15800 = ( n15678 & ~n15790 ) | ( n15678 & n15799 ) | ( ~n15790 & n15799 ) ;
  assign n15801 = ( n15678 & n15790 ) | ( n15678 & n15799 ) | ( n15790 & n15799 ) ;
  assign n15802 = ( n15790 & n15800 ) | ( n15790 & ~n15801 ) | ( n15800 & ~n15801 ) ;
  assign n15803 = ( n15690 & n15715 ) | ( n15690 & ~n15802 ) | ( n15715 & ~n15802 ) ;
  assign n15804 = ( ~n15690 & n15715 ) | ( ~n15690 & n15802 ) | ( n15715 & n15802 ) ;
  assign n15805 = ( ~n15715 & n15803 ) | ( ~n15715 & n15804 ) | ( n15803 & n15804 ) ;
  assign n15806 = ( n15693 & n15706 ) | ( n15693 & ~n15805 ) | ( n15706 & ~n15805 ) ;
  assign n15807 = ( ~n15693 & n15706 ) | ( ~n15693 & n15805 ) | ( n15706 & n15805 ) ;
  assign n15808 = ( ~n15706 & n15806 ) | ( ~n15706 & n15807 ) | ( n15806 & n15807 ) ;
  assign n15809 = ( ~n15696 & n15699 ) | ( ~n15696 & n15808 ) | ( n15699 & n15808 ) ;
  assign n15810 = ( n15699 & n15808 ) | ( n15699 & ~n15809 ) | ( n15808 & ~n15809 ) ;
  assign n15811 = ( n15696 & n15809 ) | ( n15696 & ~n15810 ) | ( n15809 & ~n15810 ) ;
  assign n15812 = n3715 & n8846 ;
  assign n15813 = x126 & n3719 ;
  assign n15814 = x127 | n15813 ;
  assign n15815 = ( n3721 & n15813 ) | ( n3721 & n15814 ) | ( n15813 & n15814 ) ;
  assign n15816 = x125 & n3922 ;
  assign n15817 = n15815 | n15816 ;
  assign n15818 = ( x41 & n15812 ) | ( x41 & ~n15817 ) | ( n15812 & ~n15817 ) ;
  assign n15819 = ( ~x41 & n15817 ) | ( ~x41 & n15818 ) | ( n15817 & n15818 ) ;
  assign n15820 = ( ~n15812 & n15818 ) | ( ~n15812 & n15819 ) | ( n15818 & n15819 ) ;
  assign n15821 = n4227 & n7841 ;
  assign n15822 = x123 & n4231 ;
  assign n15823 = x124 | n15822 ;
  assign n15824 = ( n4233 & n15822 ) | ( n4233 & n15823 ) | ( n15822 & n15823 ) ;
  assign n15825 = x122 & n4470 ;
  assign n15826 = n15824 | n15825 ;
  assign n15827 = ( x44 & n15821 ) | ( x44 & ~n15826 ) | ( n15821 & ~n15826 ) ;
  assign n15828 = ( ~x44 & n15826 ) | ( ~x44 & n15827 ) | ( n15826 & n15827 ) ;
  assign n15829 = ( ~n15821 & n15827 ) | ( ~n15821 & n15828 ) | ( n15827 & n15828 ) ;
  assign n15830 = n4787 & n7113 ;
  assign n15831 = x120 & n4791 ;
  assign n15832 = x121 | n15831 ;
  assign n15833 = ( n4793 & n15831 ) | ( n4793 & n15832 ) | ( n15831 & n15832 ) ;
  assign n15834 = x119 & n5030 ;
  assign n15835 = n15833 | n15834 ;
  assign n15836 = ( x47 & n15830 ) | ( x47 & ~n15835 ) | ( n15830 & ~n15835 ) ;
  assign n15837 = ( ~x47 & n15835 ) | ( ~x47 & n15836 ) | ( n15835 & n15836 ) ;
  assign n15838 = ( ~n15830 & n15836 ) | ( ~n15830 & n15837 ) | ( n15836 & n15837 ) ;
  assign n15839 = n5374 & n6421 ;
  assign n15840 = x117 & n5378 ;
  assign n15841 = x118 | n15840 ;
  assign n15842 = ( n5380 & n15840 ) | ( n5380 & n15841 ) | ( n15840 & n15841 ) ;
  assign n15843 = x116 & n5638 ;
  assign n15844 = n15842 | n15843 ;
  assign n15845 = ( x50 & n15839 ) | ( x50 & ~n15844 ) | ( n15839 & ~n15844 ) ;
  assign n15846 = ( ~x50 & n15844 ) | ( ~x50 & n15845 ) | ( n15844 & n15845 ) ;
  assign n15847 = ( ~n15839 & n15845 ) | ( ~n15839 & n15846 ) | ( n15845 & n15846 ) ;
  assign n15848 = n5765 & n6027 ;
  assign n15849 = x114 & n6031 ;
  assign n15850 = x115 | n15849 ;
  assign n15851 = ( n6033 & n15849 ) | ( n6033 & n15850 ) | ( n15849 & n15850 ) ;
  assign n15852 = x113 & n6303 ;
  assign n15853 = n15851 | n15852 ;
  assign n15854 = ( x53 & n15848 ) | ( x53 & ~n15853 ) | ( n15848 & ~n15853 ) ;
  assign n15855 = ( ~x53 & n15853 ) | ( ~x53 & n15854 ) | ( n15853 & n15854 ) ;
  assign n15856 = ( ~n15848 & n15854 ) | ( ~n15848 & n15855 ) | ( n15854 & n15855 ) ;
  assign n15857 = n5145 & n6713 ;
  assign n15858 = x111 & n6717 ;
  assign n15859 = x112 | n15858 ;
  assign n15860 = ( n6719 & n15858 ) | ( n6719 & n15859 ) | ( n15858 & n15859 ) ;
  assign n15861 = x110 & n6980 ;
  assign n15862 = n15860 | n15861 ;
  assign n15863 = ( x56 & n15857 ) | ( x56 & ~n15862 ) | ( n15857 & ~n15862 ) ;
  assign n15864 = ( ~x56 & n15862 ) | ( ~x56 & n15863 ) | ( n15862 & n15863 ) ;
  assign n15865 = ( ~n15857 & n15863 ) | ( ~n15857 & n15864 ) | ( n15863 & n15864 ) ;
  assign n15866 = n4734 & n7423 ;
  assign n15867 = x108 & n7427 ;
  assign n15868 = x109 | n15867 ;
  assign n15869 = ( n7429 & n15867 ) | ( n7429 & n15868 ) | ( n15867 & n15868 ) ;
  assign n15870 = x107 & n7708 ;
  assign n15871 = n15869 | n15870 ;
  assign n15872 = ( x59 & n15866 ) | ( x59 & ~n15871 ) | ( n15866 & ~n15871 ) ;
  assign n15873 = ( ~x59 & n15871 ) | ( ~x59 & n15872 ) | ( n15871 & n15872 ) ;
  assign n15874 = ( ~n15866 & n15872 ) | ( ~n15866 & n15873 ) | ( n15872 & n15873 ) ;
  assign n15875 = n4013 & n8154 ;
  assign n15876 = x105 & n8158 ;
  assign n15877 = x106 | n15876 ;
  assign n15878 = ( n8160 & n15876 ) | ( n8160 & n15877 ) | ( n15876 & n15877 ) ;
  assign n15879 = x104 & n8439 ;
  assign n15880 = n15878 | n15879 ;
  assign n15881 = ( x62 & n15875 ) | ( x62 & ~n15880 ) | ( n15875 & ~n15880 ) ;
  assign n15882 = ( ~x62 & n15880 ) | ( ~x62 & n15881 ) | ( n15880 & n15881 ) ;
  assign n15883 = ( ~n15875 & n15881 ) | ( ~n15875 & n15882 ) | ( n15881 & n15882 ) ;
  assign n15884 = x102 & n8927 ;
  assign n15885 = ( ~x103 & n8693 ) | ( ~x103 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15886 = ( n8693 & n15884 ) | ( n8693 & ~n15885 ) | ( n15884 & ~n15885 ) ;
  assign n15887 = ( ~x38 & n15644 ) | ( ~x38 & n15886 ) | ( n15644 & n15886 ) ;
  assign n15888 = ( n15644 & n15886 ) | ( n15644 & ~n15887 ) | ( n15886 & ~n15887 ) ;
  assign n15889 = ( x38 & n15887 ) | ( x38 & ~n15888 ) | ( n15887 & ~n15888 ) ;
  assign n15890 = ( n15746 & n15883 ) | ( n15746 & ~n15889 ) | ( n15883 & ~n15889 ) ;
  assign n15891 = ( ~n15746 & n15883 ) | ( ~n15746 & n15889 ) | ( n15883 & n15889 ) ;
  assign n15892 = ( ~n15883 & n15890 ) | ( ~n15883 & n15891 ) | ( n15890 & n15891 ) ;
  assign n15893 = ( n15767 & n15874 ) | ( n15767 & ~n15892 ) | ( n15874 & ~n15892 ) ;
  assign n15894 = ( ~n15767 & n15874 ) | ( ~n15767 & n15892 ) | ( n15874 & n15892 ) ;
  assign n15895 = ( ~n15874 & n15893 ) | ( ~n15874 & n15894 ) | ( n15893 & n15894 ) ;
  assign n15896 = ( n15779 & n15865 ) | ( n15779 & ~n15895 ) | ( n15865 & ~n15895 ) ;
  assign n15897 = ( ~n15779 & n15865 ) | ( ~n15779 & n15895 ) | ( n15865 & n15895 ) ;
  assign n15898 = ( ~n15865 & n15896 ) | ( ~n15865 & n15897 ) | ( n15896 & n15897 ) ;
  assign n15899 = ( n15782 & n15856 ) | ( n15782 & ~n15898 ) | ( n15856 & ~n15898 ) ;
  assign n15900 = ( ~n15782 & n15856 ) | ( ~n15782 & n15898 ) | ( n15856 & n15898 ) ;
  assign n15901 = ( ~n15856 & n15899 ) | ( ~n15856 & n15900 ) | ( n15899 & n15900 ) ;
  assign n15902 = ( n15785 & n15847 ) | ( n15785 & ~n15901 ) | ( n15847 & ~n15901 ) ;
  assign n15903 = ( ~n15785 & n15847 ) | ( ~n15785 & n15901 ) | ( n15847 & n15901 ) ;
  assign n15904 = ( ~n15847 & n15902 ) | ( ~n15847 & n15903 ) | ( n15902 & n15903 ) ;
  assign n15905 = ( n15788 & n15838 ) | ( n15788 & ~n15904 ) | ( n15838 & ~n15904 ) ;
  assign n15906 = ( ~n15788 & n15838 ) | ( ~n15788 & n15904 ) | ( n15838 & n15904 ) ;
  assign n15907 = ( ~n15838 & n15905 ) | ( ~n15838 & n15906 ) | ( n15905 & n15906 ) ;
  assign n15908 = ( n15800 & n15829 ) | ( n15800 & ~n15907 ) | ( n15829 & ~n15907 ) ;
  assign n15909 = ( ~n15800 & n15829 ) | ( ~n15800 & n15907 ) | ( n15829 & n15907 ) ;
  assign n15910 = ( ~n15829 & n15908 ) | ( ~n15829 & n15909 ) | ( n15908 & n15909 ) ;
  assign n15911 = ( n15803 & n15820 ) | ( n15803 & ~n15910 ) | ( n15820 & ~n15910 ) ;
  assign n15912 = ( ~n15803 & n15820 ) | ( ~n15803 & n15910 ) | ( n15820 & n15910 ) ;
  assign n15913 = ( ~n15820 & n15911 ) | ( ~n15820 & n15912 ) | ( n15911 & n15912 ) ;
  assign n15914 = ( ~n15806 & n15809 ) | ( ~n15806 & n15913 ) | ( n15809 & n15913 ) ;
  assign n15915 = ( n15809 & n15913 ) | ( n15809 & ~n15914 ) | ( n15913 & ~n15914 ) ;
  assign n15916 = ( n15806 & n15914 ) | ( n15806 & ~n15915 ) | ( n15914 & ~n15915 ) ;
  assign n15917 = n3715 & n8865 ;
  assign n15918 = x127 & n3719 ;
  assign n15919 = x126 | n15918 ;
  assign n15920 = ( n3922 & n15918 ) | ( n3922 & n15919 ) | ( n15918 & n15919 ) ;
  assign n15921 = ( x41 & n15917 ) | ( x41 & ~n15920 ) | ( n15917 & ~n15920 ) ;
  assign n15922 = ( ~x41 & n15920 ) | ( ~x41 & n15921 ) | ( n15920 & n15921 ) ;
  assign n15923 = ( ~n15917 & n15921 ) | ( ~n15917 & n15922 ) | ( n15921 & n15922 ) ;
  assign n15924 = n4787 & n7582 ;
  assign n15925 = x121 & n4791 ;
  assign n15926 = x122 | n15925 ;
  assign n15927 = ( n4793 & n15925 ) | ( n4793 & n15926 ) | ( n15925 & n15926 ) ;
  assign n15928 = x120 & n5030 ;
  assign n15929 = n15927 | n15928 ;
  assign n15930 = ( x47 & n15924 ) | ( x47 & ~n15929 ) | ( n15924 & ~n15929 ) ;
  assign n15931 = ( ~x47 & n15929 ) | ( ~x47 & n15930 ) | ( n15929 & n15930 ) ;
  assign n15932 = ( ~n15924 & n15930 ) | ( ~n15924 & n15931 ) | ( n15930 & n15931 ) ;
  assign n15933 = n5977 & n6027 ;
  assign n15934 = x115 & n6031 ;
  assign n15935 = x116 | n15934 ;
  assign n15936 = ( n6033 & n15934 ) | ( n6033 & n15935 ) | ( n15934 & n15935 ) ;
  assign n15937 = x114 & n6303 ;
  assign n15938 = n15936 | n15937 ;
  assign n15939 = ( x53 & n15933 ) | ( x53 & ~n15938 ) | ( n15933 & ~n15938 ) ;
  assign n15940 = ( ~x53 & n15938 ) | ( ~x53 & n15939 ) | ( n15938 & n15939 ) ;
  assign n15941 = ( ~n15933 & n15939 ) | ( ~n15933 & n15940 ) | ( n15939 & n15940 ) ;
  assign n15942 = n4934 & n7423 ;
  assign n15943 = x109 & n7427 ;
  assign n15944 = x110 | n15943 ;
  assign n15945 = ( n7429 & n15943 ) | ( n7429 & n15944 ) | ( n15943 & n15944 ) ;
  assign n15946 = x108 & n7708 ;
  assign n15947 = n15945 | n15946 ;
  assign n15948 = ( x59 & n15942 ) | ( x59 & ~n15947 ) | ( n15942 & ~n15947 ) ;
  assign n15949 = ( ~x59 & n15947 ) | ( ~x59 & n15948 ) | ( n15947 & n15948 ) ;
  assign n15950 = ( ~n15942 & n15948 ) | ( ~n15942 & n15949 ) | ( n15948 & n15949 ) ;
  assign n15951 = n4362 & n8154 ;
  assign n15952 = x106 & n8158 ;
  assign n15953 = x107 | n15952 ;
  assign n15954 = ( n8160 & n15952 ) | ( n8160 & n15953 ) | ( n15952 & n15953 ) ;
  assign n15955 = x105 & n8439 ;
  assign n15956 = n15954 | n15955 ;
  assign n15957 = ( x62 & n15951 ) | ( x62 & ~n15956 ) | ( n15951 & ~n15956 ) ;
  assign n15958 = ( ~x62 & n15956 ) | ( ~x62 & n15957 ) | ( n15956 & n15957 ) ;
  assign n15959 = ( ~n15951 & n15957 ) | ( ~n15951 & n15958 ) | ( n15957 & n15958 ) ;
  assign n15960 = x103 & n8927 ;
  assign n15961 = ( ~x104 & n8693 ) | ( ~x104 & n8927 ) | ( n8693 & n8927 ) ;
  assign n15962 = ( n8693 & n15960 ) | ( n8693 & ~n15961 ) | ( n15960 & ~n15961 ) ;
  assign n15963 = ( n15887 & n15959 ) | ( n15887 & ~n15962 ) | ( n15959 & ~n15962 ) ;
  assign n15964 = ( ~n15887 & n15959 ) | ( ~n15887 & n15962 ) | ( n15959 & n15962 ) ;
  assign n15965 = ( ~n15959 & n15963 ) | ( ~n15959 & n15964 ) | ( n15963 & n15964 ) ;
  assign n15966 = ( n15890 & n15950 ) | ( n15890 & ~n15965 ) | ( n15950 & ~n15965 ) ;
  assign n15967 = ( ~n15890 & n15950 ) | ( ~n15890 & n15965 ) | ( n15950 & n15965 ) ;
  assign n15968 = ( ~n15950 & n15966 ) | ( ~n15950 & n15967 ) | ( n15966 & n15967 ) ;
  assign n15969 = n5542 & n6713 ;
  assign n15970 = x112 & n6717 ;
  assign n15971 = x113 | n15970 ;
  assign n15972 = ( n6719 & n15970 ) | ( n6719 & n15971 ) | ( n15970 & n15971 ) ;
  assign n15973 = x111 & n6980 ;
  assign n15974 = n15972 | n15973 ;
  assign n15975 = ( x56 & n15969 ) | ( x56 & ~n15974 ) | ( n15969 & ~n15974 ) ;
  assign n15976 = ( ~x56 & n15974 ) | ( ~x56 & n15975 ) | ( n15974 & n15975 ) ;
  assign n15977 = ( ~n15969 & n15975 ) | ( ~n15969 & n15976 ) | ( n15975 & n15976 ) ;
  assign n15978 = ( n15893 & ~n15968 ) | ( n15893 & n15977 ) | ( ~n15968 & n15977 ) ;
  assign n15979 = ( n15893 & n15968 ) | ( n15893 & n15977 ) | ( n15968 & n15977 ) ;
  assign n15980 = ( n15968 & n15978 ) | ( n15968 & ~n15979 ) | ( n15978 & ~n15979 ) ;
  assign n15981 = ( n15896 & n15941 ) | ( n15896 & ~n15980 ) | ( n15941 & ~n15980 ) ;
  assign n15982 = ( ~n15896 & n15941 ) | ( ~n15896 & n15980 ) | ( n15941 & n15980 ) ;
  assign n15983 = ( ~n15941 & n15981 ) | ( ~n15941 & n15982 ) | ( n15981 & n15982 ) ;
  assign n15984 = n5374 & n6645 ;
  assign n15985 = x118 & n5378 ;
  assign n15986 = x119 | n15985 ;
  assign n15987 = ( n5380 & n15985 ) | ( n5380 & n15986 ) | ( n15985 & n15986 ) ;
  assign n15988 = x117 & n5638 ;
  assign n15989 = n15987 | n15988 ;
  assign n15990 = ( x50 & n15984 ) | ( x50 & ~n15989 ) | ( n15984 & ~n15989 ) ;
  assign n15991 = ( ~x50 & n15989 ) | ( ~x50 & n15990 ) | ( n15989 & n15990 ) ;
  assign n15992 = ( ~n15984 & n15990 ) | ( ~n15984 & n15991 ) | ( n15990 & n15991 ) ;
  assign n15993 = ( n15899 & ~n15983 ) | ( n15899 & n15992 ) | ( ~n15983 & n15992 ) ;
  assign n15994 = ( n15899 & n15983 ) | ( n15899 & n15992 ) | ( n15983 & n15992 ) ;
  assign n15995 = ( n15983 & n15993 ) | ( n15983 & ~n15994 ) | ( n15993 & ~n15994 ) ;
  assign n15996 = ( n15902 & n15932 ) | ( n15902 & ~n15995 ) | ( n15932 & ~n15995 ) ;
  assign n15997 = ( ~n15902 & n15932 ) | ( ~n15902 & n15995 ) | ( n15932 & n15995 ) ;
  assign n15998 = ( ~n15932 & n15996 ) | ( ~n15932 & n15997 ) | ( n15996 & n15997 ) ;
  assign n15999 = n4227 & n8331 ;
  assign n16000 = x124 & n4231 ;
  assign n16001 = x125 | n16000 ;
  assign n16002 = ( n4233 & n16000 ) | ( n4233 & n16001 ) | ( n16000 & n16001 ) ;
  assign n16003 = x123 & n4470 ;
  assign n16004 = n16002 | n16003 ;
  assign n16005 = ( x44 & n15999 ) | ( x44 & ~n16004 ) | ( n15999 & ~n16004 ) ;
  assign n16006 = ( ~x44 & n16004 ) | ( ~x44 & n16005 ) | ( n16004 & n16005 ) ;
  assign n16007 = ( ~n15999 & n16005 ) | ( ~n15999 & n16006 ) | ( n16005 & n16006 ) ;
  assign n16008 = ( n15905 & ~n15998 ) | ( n15905 & n16007 ) | ( ~n15998 & n16007 ) ;
  assign n16009 = ( n15905 & n15998 ) | ( n15905 & n16007 ) | ( n15998 & n16007 ) ;
  assign n16010 = ( n15998 & n16008 ) | ( n15998 & ~n16009 ) | ( n16008 & ~n16009 ) ;
  assign n16011 = ( n15908 & n15923 ) | ( n15908 & ~n16010 ) | ( n15923 & ~n16010 ) ;
  assign n16012 = ( ~n15908 & n15923 ) | ( ~n15908 & n16010 ) | ( n15923 & n16010 ) ;
  assign n16013 = ( ~n15923 & n16011 ) | ( ~n15923 & n16012 ) | ( n16011 & n16012 ) ;
  assign n16014 = ( ~n15911 & n15914 ) | ( ~n15911 & n16013 ) | ( n15914 & n16013 ) ;
  assign n16015 = ( n15914 & n16013 ) | ( n15914 & ~n16014 ) | ( n16013 & ~n16014 ) ;
  assign n16016 = ( n15911 & n16014 ) | ( n15911 & ~n16015 ) | ( n16014 & ~n16015 ) ;
  assign n16017 = n3715 & n8862 ;
  assign n16018 = ( x127 & n3922 ) | ( x127 & n16017 ) | ( n3922 & n16017 ) ;
  assign n16019 = x41 | n16018 ;
  assign n16020 = ~x41 & n16018 ;
  assign n16021 = ( ~n16018 & n16019 ) | ( ~n16018 & n16020 ) | ( n16019 & n16020 ) ;
  assign n16022 = n4787 & n7597 ;
  assign n16023 = x122 & n4791 ;
  assign n16024 = x123 | n16023 ;
  assign n16025 = ( n4793 & n16023 ) | ( n4793 & n16024 ) | ( n16023 & n16024 ) ;
  assign n16026 = x121 & n5030 ;
  assign n16027 = n16025 | n16026 ;
  assign n16028 = ( x47 & n16022 ) | ( x47 & ~n16027 ) | ( n16022 & ~n16027 ) ;
  assign n16029 = ( ~x47 & n16027 ) | ( ~x47 & n16028 ) | ( n16027 & n16028 ) ;
  assign n16030 = ( ~n16022 & n16028 ) | ( ~n16022 & n16029 ) | ( n16028 & n16029 ) ;
  assign n16031 = n5374 & n7098 ;
  assign n16032 = x119 & n5378 ;
  assign n16033 = x120 | n16032 ;
  assign n16034 = ( n5380 & n16032 ) | ( n5380 & n16033 ) | ( n16032 & n16033 ) ;
  assign n16035 = x118 & n5638 ;
  assign n16036 = n16034 | n16035 ;
  assign n16037 = ( x50 & n16031 ) | ( x50 & ~n16036 ) | ( n16031 & ~n16036 ) ;
  assign n16038 = ( ~x50 & n16036 ) | ( ~x50 & n16037 ) | ( n16036 & n16037 ) ;
  assign n16039 = ( ~n16031 & n16037 ) | ( ~n16031 & n16038 ) | ( n16037 & n16038 ) ;
  assign n16040 = n6027 & n6201 ;
  assign n16041 = x116 & n6031 ;
  assign n16042 = x117 | n16041 ;
  assign n16043 = ( n6033 & n16041 ) | ( n6033 & n16042 ) | ( n16041 & n16042 ) ;
  assign n16044 = x115 & n6303 ;
  assign n16045 = n16043 | n16044 ;
  assign n16046 = ( x53 & n16040 ) | ( x53 & ~n16045 ) | ( n16040 & ~n16045 ) ;
  assign n16047 = ( ~x53 & n16045 ) | ( ~x53 & n16046 ) | ( n16045 & n16046 ) ;
  assign n16048 = ( ~n16040 & n16046 ) | ( ~n16040 & n16047 ) | ( n16046 & n16047 ) ;
  assign n16049 = x104 & n8927 ;
  assign n16050 = ( ~x105 & n8693 ) | ( ~x105 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16051 = ( n8693 & n16049 ) | ( n8693 & ~n16050 ) | ( n16049 & ~n16050 ) ;
  assign n16052 = ( ~n15962 & n15963 ) | ( ~n15962 & n16051 ) | ( n15963 & n16051 ) ;
  assign n16053 = ( n15962 & n15963 ) | ( n15962 & ~n16051 ) | ( n15963 & ~n16051 ) ;
  assign n16054 = ( ~n15963 & n16052 ) | ( ~n15963 & n16053 ) | ( n16052 & n16053 ) ;
  assign n16055 = n5130 & n7423 ;
  assign n16056 = x110 & n7427 ;
  assign n16057 = x111 | n16056 ;
  assign n16058 = ( n7429 & n16056 ) | ( n7429 & n16057 ) | ( n16056 & n16057 ) ;
  assign n16059 = x109 & n7708 ;
  assign n16060 = n16058 | n16059 ;
  assign n16061 = ( x59 & n16055 ) | ( x59 & ~n16060 ) | ( n16055 & ~n16060 ) ;
  assign n16062 = ( ~x59 & n16060 ) | ( ~x59 & n16061 ) | ( n16060 & n16061 ) ;
  assign n16063 = ( ~n16055 & n16061 ) | ( ~n16055 & n16062 ) | ( n16061 & n16062 ) ;
  assign n16064 = n4377 & n8154 ;
  assign n16065 = x107 & n8158 ;
  assign n16066 = x108 | n16065 ;
  assign n16067 = ( n8160 & n16065 ) | ( n8160 & n16066 ) | ( n16065 & n16066 ) ;
  assign n16068 = x106 & n8439 ;
  assign n16069 = n16067 | n16068 ;
  assign n16070 = ( x62 & n16064 ) | ( x62 & ~n16069 ) | ( n16064 & ~n16069 ) ;
  assign n16071 = ( ~x62 & n16069 ) | ( ~x62 & n16070 ) | ( n16069 & n16070 ) ;
  assign n16072 = ( ~n16064 & n16070 ) | ( ~n16064 & n16071 ) | ( n16070 & n16071 ) ;
  assign n16073 = ( ~n16054 & n16063 ) | ( ~n16054 & n16072 ) | ( n16063 & n16072 ) ;
  assign n16074 = ( n16063 & n16072 ) | ( n16063 & ~n16073 ) | ( n16072 & ~n16073 ) ;
  assign n16075 = ( n16054 & n16073 ) | ( n16054 & ~n16074 ) | ( n16073 & ~n16074 ) ;
  assign n16076 = n5750 & n6713 ;
  assign n16077 = x113 & n6717 ;
  assign n16078 = x114 | n16077 ;
  assign n16079 = ( n6719 & n16077 ) | ( n6719 & n16078 ) | ( n16077 & n16078 ) ;
  assign n16080 = x112 & n6980 ;
  assign n16081 = n16079 | n16080 ;
  assign n16082 = ( x56 & n16076 ) | ( x56 & ~n16081 ) | ( n16076 & ~n16081 ) ;
  assign n16083 = ( ~x56 & n16081 ) | ( ~x56 & n16082 ) | ( n16081 & n16082 ) ;
  assign n16084 = ( ~n16076 & n16082 ) | ( ~n16076 & n16083 ) | ( n16082 & n16083 ) ;
  assign n16085 = ( n15966 & ~n16075 ) | ( n15966 & n16084 ) | ( ~n16075 & n16084 ) ;
  assign n16086 = ( n15966 & n16075 ) | ( n15966 & n16084 ) | ( n16075 & n16084 ) ;
  assign n16087 = ( n16075 & n16085 ) | ( n16075 & ~n16086 ) | ( n16085 & ~n16086 ) ;
  assign n16088 = ( n15978 & n16048 ) | ( n15978 & ~n16087 ) | ( n16048 & ~n16087 ) ;
  assign n16089 = ( ~n15978 & n16048 ) | ( ~n15978 & n16087 ) | ( n16048 & n16087 ) ;
  assign n16090 = ( ~n16048 & n16088 ) | ( ~n16048 & n16089 ) | ( n16088 & n16089 ) ;
  assign n16091 = ( n15981 & n16039 ) | ( n15981 & ~n16090 ) | ( n16039 & ~n16090 ) ;
  assign n16092 = ( ~n15981 & n16039 ) | ( ~n15981 & n16090 ) | ( n16039 & n16090 ) ;
  assign n16093 = ( ~n16039 & n16091 ) | ( ~n16039 & n16092 ) | ( n16091 & n16092 ) ;
  assign n16094 = ( n15993 & n16030 ) | ( n15993 & ~n16093 ) | ( n16030 & ~n16093 ) ;
  assign n16095 = ( ~n15993 & n16030 ) | ( ~n15993 & n16093 ) | ( n16030 & n16093 ) ;
  assign n16096 = ( ~n16030 & n16094 ) | ( ~n16030 & n16095 ) | ( n16094 & n16095 ) ;
  assign n16097 = n4227 & n8587 ;
  assign n16098 = x125 & n4231 ;
  assign n16099 = x126 | n16098 ;
  assign n16100 = ( n4233 & n16098 ) | ( n4233 & n16099 ) | ( n16098 & n16099 ) ;
  assign n16101 = x124 & n4470 ;
  assign n16102 = n16100 | n16101 ;
  assign n16103 = ( x44 & n16097 ) | ( x44 & ~n16102 ) | ( n16097 & ~n16102 ) ;
  assign n16104 = ( ~x44 & n16102 ) | ( ~x44 & n16103 ) | ( n16102 & n16103 ) ;
  assign n16105 = ( ~n16097 & n16103 ) | ( ~n16097 & n16104 ) | ( n16103 & n16104 ) ;
  assign n16106 = ( n15996 & ~n16096 ) | ( n15996 & n16105 ) | ( ~n16096 & n16105 ) ;
  assign n16107 = ( n15996 & n16096 ) | ( n15996 & n16105 ) | ( n16096 & n16105 ) ;
  assign n16108 = ( n16096 & n16106 ) | ( n16096 & ~n16107 ) | ( n16106 & ~n16107 ) ;
  assign n16109 = ( n16008 & n16021 ) | ( n16008 & ~n16108 ) | ( n16021 & ~n16108 ) ;
  assign n16110 = ( ~n16008 & n16021 ) | ( ~n16008 & n16108 ) | ( n16021 & n16108 ) ;
  assign n16111 = ( ~n16021 & n16109 ) | ( ~n16021 & n16110 ) | ( n16109 & n16110 ) ;
  assign n16112 = ( ~n16011 & n16014 ) | ( ~n16011 & n16111 ) | ( n16014 & n16111 ) ;
  assign n16113 = ( n16014 & n16111 ) | ( n16014 & ~n16112 ) | ( n16111 & ~n16112 ) ;
  assign n16114 = ( n16011 & n16112 ) | ( n16011 & ~n16113 ) | ( n16112 & ~n16113 ) ;
  assign n16115 = n4227 & n8846 ;
  assign n16116 = x126 & n4231 ;
  assign n16117 = x127 | n16116 ;
  assign n16118 = ( n4233 & n16116 ) | ( n4233 & n16117 ) | ( n16116 & n16117 ) ;
  assign n16119 = x125 & n4470 ;
  assign n16120 = n16118 | n16119 ;
  assign n16121 = ( x44 & n16115 ) | ( x44 & ~n16120 ) | ( n16115 & ~n16120 ) ;
  assign n16122 = ( ~x44 & n16120 ) | ( ~x44 & n16121 ) | ( n16120 & n16121 ) ;
  assign n16123 = ( ~n16115 & n16121 ) | ( ~n16115 & n16122 ) | ( n16121 & n16122 ) ;
  assign n16124 = n4787 & n7841 ;
  assign n16125 = x123 & n4791 ;
  assign n16126 = x124 | n16125 ;
  assign n16127 = ( n4793 & n16125 ) | ( n4793 & n16126 ) | ( n16125 & n16126 ) ;
  assign n16128 = x122 & n5030 ;
  assign n16129 = n16127 | n16128 ;
  assign n16130 = ( x47 & n16124 ) | ( x47 & ~n16129 ) | ( n16124 & ~n16129 ) ;
  assign n16131 = ( ~x47 & n16129 ) | ( ~x47 & n16130 ) | ( n16129 & n16130 ) ;
  assign n16132 = ( ~n16124 & n16130 ) | ( ~n16124 & n16131 ) | ( n16130 & n16131 ) ;
  assign n16133 = n5374 & n7113 ;
  assign n16134 = x120 & n5378 ;
  assign n16135 = x121 | n16134 ;
  assign n16136 = ( n5380 & n16134 ) | ( n5380 & n16135 ) | ( n16134 & n16135 ) ;
  assign n16137 = x119 & n5638 ;
  assign n16138 = n16136 | n16137 ;
  assign n16139 = ( x50 & n16133 ) | ( x50 & ~n16138 ) | ( n16133 & ~n16138 ) ;
  assign n16140 = ( ~x50 & n16138 ) | ( ~x50 & n16139 ) | ( n16138 & n16139 ) ;
  assign n16141 = ( ~n16133 & n16139 ) | ( ~n16133 & n16140 ) | ( n16139 & n16140 ) ;
  assign n16142 = n6027 & n6421 ;
  assign n16143 = x117 & n6031 ;
  assign n16144 = x118 | n16143 ;
  assign n16145 = ( n6033 & n16143 ) | ( n6033 & n16144 ) | ( n16143 & n16144 ) ;
  assign n16146 = x116 & n6303 ;
  assign n16147 = n16145 | n16146 ;
  assign n16148 = ( x53 & n16142 ) | ( x53 & ~n16147 ) | ( n16142 & ~n16147 ) ;
  assign n16149 = ( ~x53 & n16147 ) | ( ~x53 & n16148 ) | ( n16147 & n16148 ) ;
  assign n16150 = ( ~n16142 & n16148 ) | ( ~n16142 & n16149 ) | ( n16148 & n16149 ) ;
  assign n16151 = n5765 & n6713 ;
  assign n16152 = x114 & n6717 ;
  assign n16153 = x115 | n16152 ;
  assign n16154 = ( n6719 & n16152 ) | ( n6719 & n16153 ) | ( n16152 & n16153 ) ;
  assign n16155 = x113 & n6980 ;
  assign n16156 = n16154 | n16155 ;
  assign n16157 = ( x56 & n16151 ) | ( x56 & ~n16156 ) | ( n16151 & ~n16156 ) ;
  assign n16158 = ( ~x56 & n16156 ) | ( ~x56 & n16157 ) | ( n16156 & n16157 ) ;
  assign n16159 = ( ~n16151 & n16157 ) | ( ~n16151 & n16158 ) | ( n16157 & n16158 ) ;
  assign n16160 = n5145 & n7423 ;
  assign n16161 = x111 & n7427 ;
  assign n16162 = x112 | n16161 ;
  assign n16163 = ( n7429 & n16161 ) | ( n7429 & n16162 ) | ( n16161 & n16162 ) ;
  assign n16164 = x110 & n7708 ;
  assign n16165 = n16163 | n16164 ;
  assign n16166 = ( x59 & n16160 ) | ( x59 & ~n16165 ) | ( n16160 & ~n16165 ) ;
  assign n16167 = ( ~x59 & n16165 ) | ( ~x59 & n16166 ) | ( n16165 & n16166 ) ;
  assign n16168 = ( ~n16160 & n16166 ) | ( ~n16160 & n16167 ) | ( n16166 & n16167 ) ;
  assign n16169 = n4734 & n8154 ;
  assign n16170 = x108 & n8158 ;
  assign n16171 = x109 | n16170 ;
  assign n16172 = ( n8160 & n16170 ) | ( n8160 & n16171 ) | ( n16170 & n16171 ) ;
  assign n16173 = x107 & n8439 ;
  assign n16174 = n16172 | n16173 ;
  assign n16175 = ( x62 & n16169 ) | ( x62 & ~n16174 ) | ( n16169 & ~n16174 ) ;
  assign n16176 = ( ~x62 & n16174 ) | ( ~x62 & n16175 ) | ( n16174 & n16175 ) ;
  assign n16177 = ( ~n16169 & n16175 ) | ( ~n16169 & n16176 ) | ( n16175 & n16176 ) ;
  assign n16178 = x105 & n8927 ;
  assign n16179 = ( ~x106 & n8693 ) | ( ~x106 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16180 = ( n8693 & n16178 ) | ( n8693 & ~n16179 ) | ( n16178 & ~n16179 ) ;
  assign n16181 = ( ~x41 & n15962 ) | ( ~x41 & n16180 ) | ( n15962 & n16180 ) ;
  assign n16182 = ( n15962 & n16180 ) | ( n15962 & ~n16181 ) | ( n16180 & ~n16181 ) ;
  assign n16183 = ( x41 & n16181 ) | ( x41 & ~n16182 ) | ( n16181 & ~n16182 ) ;
  assign n16184 = ( n16052 & n16177 ) | ( n16052 & ~n16183 ) | ( n16177 & ~n16183 ) ;
  assign n16185 = ( ~n16052 & n16177 ) | ( ~n16052 & n16183 ) | ( n16177 & n16183 ) ;
  assign n16186 = ( ~n16177 & n16184 ) | ( ~n16177 & n16185 ) | ( n16184 & n16185 ) ;
  assign n16187 = ( n16073 & n16168 ) | ( n16073 & ~n16186 ) | ( n16168 & ~n16186 ) ;
  assign n16188 = ( ~n16073 & n16168 ) | ( ~n16073 & n16186 ) | ( n16168 & n16186 ) ;
  assign n16189 = ( ~n16168 & n16187 ) | ( ~n16168 & n16188 ) | ( n16187 & n16188 ) ;
  assign n16190 = ( n16085 & n16159 ) | ( n16085 & ~n16189 ) | ( n16159 & ~n16189 ) ;
  assign n16191 = ( ~n16085 & n16159 ) | ( ~n16085 & n16189 ) | ( n16159 & n16189 ) ;
  assign n16192 = ( ~n16159 & n16190 ) | ( ~n16159 & n16191 ) | ( n16190 & n16191 ) ;
  assign n16193 = ( n16088 & n16150 ) | ( n16088 & ~n16192 ) | ( n16150 & ~n16192 ) ;
  assign n16194 = ( ~n16088 & n16150 ) | ( ~n16088 & n16192 ) | ( n16150 & n16192 ) ;
  assign n16195 = ( ~n16150 & n16193 ) | ( ~n16150 & n16194 ) | ( n16193 & n16194 ) ;
  assign n16196 = ( n16091 & n16141 ) | ( n16091 & ~n16195 ) | ( n16141 & ~n16195 ) ;
  assign n16197 = ( ~n16091 & n16141 ) | ( ~n16091 & n16195 ) | ( n16141 & n16195 ) ;
  assign n16198 = ( ~n16141 & n16196 ) | ( ~n16141 & n16197 ) | ( n16196 & n16197 ) ;
  assign n16199 = ( n16094 & n16132 ) | ( n16094 & ~n16198 ) | ( n16132 & ~n16198 ) ;
  assign n16200 = ( ~n16094 & n16132 ) | ( ~n16094 & n16198 ) | ( n16132 & n16198 ) ;
  assign n16201 = ( ~n16132 & n16199 ) | ( ~n16132 & n16200 ) | ( n16199 & n16200 ) ;
  assign n16202 = ( n16106 & n16123 ) | ( n16106 & ~n16201 ) | ( n16123 & ~n16201 ) ;
  assign n16203 = ( ~n16106 & n16123 ) | ( ~n16106 & n16201 ) | ( n16123 & n16201 ) ;
  assign n16204 = ( ~n16123 & n16202 ) | ( ~n16123 & n16203 ) | ( n16202 & n16203 ) ;
  assign n16205 = ( ~n16109 & n16112 ) | ( ~n16109 & n16204 ) | ( n16112 & n16204 ) ;
  assign n16206 = ( n16112 & n16204 ) | ( n16112 & ~n16205 ) | ( n16204 & ~n16205 ) ;
  assign n16207 = ( n16109 & n16205 ) | ( n16109 & ~n16206 ) | ( n16205 & ~n16206 ) ;
  assign n16208 = n4227 & n8865 ;
  assign n16209 = x127 & n4231 ;
  assign n16210 = x126 | n16209 ;
  assign n16211 = ( n4470 & n16209 ) | ( n4470 & n16210 ) | ( n16209 & n16210 ) ;
  assign n16212 = ( x44 & n16208 ) | ( x44 & ~n16211 ) | ( n16208 & ~n16211 ) ;
  assign n16213 = ( ~x44 & n16211 ) | ( ~x44 & n16212 ) | ( n16211 & n16212 ) ;
  assign n16214 = ( ~n16208 & n16212 ) | ( ~n16208 & n16213 ) | ( n16212 & n16213 ) ;
  assign n16215 = n4787 & n8331 ;
  assign n16216 = x124 & n4791 ;
  assign n16217 = x125 | n16216 ;
  assign n16218 = ( n4793 & n16216 ) | ( n4793 & n16217 ) | ( n16216 & n16217 ) ;
  assign n16219 = x123 & n5030 ;
  assign n16220 = n16218 | n16219 ;
  assign n16221 = ( x47 & n16215 ) | ( x47 & ~n16220 ) | ( n16215 & ~n16220 ) ;
  assign n16222 = ( ~x47 & n16220 ) | ( ~x47 & n16221 ) | ( n16220 & n16221 ) ;
  assign n16223 = ( ~n16215 & n16221 ) | ( ~n16215 & n16222 ) | ( n16221 & n16222 ) ;
  assign n16224 = n5374 & n7582 ;
  assign n16225 = x121 & n5378 ;
  assign n16226 = x122 | n16225 ;
  assign n16227 = ( n5380 & n16225 ) | ( n5380 & n16226 ) | ( n16225 & n16226 ) ;
  assign n16228 = x120 & n5638 ;
  assign n16229 = n16227 | n16228 ;
  assign n16230 = ( x50 & n16224 ) | ( x50 & ~n16229 ) | ( n16224 & ~n16229 ) ;
  assign n16231 = ( ~x50 & n16229 ) | ( ~x50 & n16230 ) | ( n16229 & n16230 ) ;
  assign n16232 = ( ~n16224 & n16230 ) | ( ~n16224 & n16231 ) | ( n16230 & n16231 ) ;
  assign n16233 = n6027 & n6645 ;
  assign n16234 = x118 & n6031 ;
  assign n16235 = x119 | n16234 ;
  assign n16236 = ( n6033 & n16234 ) | ( n6033 & n16235 ) | ( n16234 & n16235 ) ;
  assign n16237 = x117 & n6303 ;
  assign n16238 = n16236 | n16237 ;
  assign n16239 = ( x53 & n16233 ) | ( x53 & ~n16238 ) | ( n16233 & ~n16238 ) ;
  assign n16240 = ( ~x53 & n16238 ) | ( ~x53 & n16239 ) | ( n16238 & n16239 ) ;
  assign n16241 = ( ~n16233 & n16239 ) | ( ~n16233 & n16240 ) | ( n16239 & n16240 ) ;
  assign n16242 = n5977 & n6713 ;
  assign n16243 = x115 & n6717 ;
  assign n16244 = x116 | n16243 ;
  assign n16245 = ( n6719 & n16243 ) | ( n6719 & n16244 ) | ( n16243 & n16244 ) ;
  assign n16246 = x114 & n6980 ;
  assign n16247 = n16245 | n16246 ;
  assign n16248 = ( x56 & n16242 ) | ( x56 & ~n16247 ) | ( n16242 & ~n16247 ) ;
  assign n16249 = ( ~x56 & n16247 ) | ( ~x56 & n16248 ) | ( n16247 & n16248 ) ;
  assign n16250 = ( ~n16242 & n16248 ) | ( ~n16242 & n16249 ) | ( n16248 & n16249 ) ;
  assign n16251 = n5542 & n7423 ;
  assign n16252 = x112 & n7427 ;
  assign n16253 = x113 | n16252 ;
  assign n16254 = ( n7429 & n16252 ) | ( n7429 & n16253 ) | ( n16252 & n16253 ) ;
  assign n16255 = x111 & n7708 ;
  assign n16256 = n16254 | n16255 ;
  assign n16257 = ( x59 & n16251 ) | ( x59 & ~n16256 ) | ( n16251 & ~n16256 ) ;
  assign n16258 = ( ~x59 & n16256 ) | ( ~x59 & n16257 ) | ( n16256 & n16257 ) ;
  assign n16259 = ( ~n16251 & n16257 ) | ( ~n16251 & n16258 ) | ( n16257 & n16258 ) ;
  assign n16260 = n4934 & n8154 ;
  assign n16261 = x109 & n8158 ;
  assign n16262 = x110 | n16261 ;
  assign n16263 = ( n8160 & n16261 ) | ( n8160 & n16262 ) | ( n16261 & n16262 ) ;
  assign n16264 = x108 & n8439 ;
  assign n16265 = n16263 | n16264 ;
  assign n16266 = ( x62 & n16260 ) | ( x62 & ~n16265 ) | ( n16260 & ~n16265 ) ;
  assign n16267 = ( ~x62 & n16265 ) | ( ~x62 & n16266 ) | ( n16265 & n16266 ) ;
  assign n16268 = ( ~n16260 & n16266 ) | ( ~n16260 & n16267 ) | ( n16266 & n16267 ) ;
  assign n16269 = x106 & n8927 ;
  assign n16270 = ( ~x107 & n8693 ) | ( ~x107 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16271 = ( n8693 & n16269 ) | ( n8693 & ~n16270 ) | ( n16269 & ~n16270 ) ;
  assign n16272 = ( n16181 & n16268 ) | ( n16181 & ~n16271 ) | ( n16268 & ~n16271 ) ;
  assign n16273 = ( ~n16181 & n16268 ) | ( ~n16181 & n16271 ) | ( n16268 & n16271 ) ;
  assign n16274 = ( ~n16268 & n16272 ) | ( ~n16268 & n16273 ) | ( n16272 & n16273 ) ;
  assign n16275 = ( n16184 & n16259 ) | ( n16184 & ~n16274 ) | ( n16259 & ~n16274 ) ;
  assign n16276 = ( ~n16184 & n16259 ) | ( ~n16184 & n16274 ) | ( n16259 & n16274 ) ;
  assign n16277 = ( ~n16259 & n16275 ) | ( ~n16259 & n16276 ) | ( n16275 & n16276 ) ;
  assign n16278 = ( n16187 & n16250 ) | ( n16187 & ~n16277 ) | ( n16250 & ~n16277 ) ;
  assign n16279 = ( ~n16187 & n16250 ) | ( ~n16187 & n16277 ) | ( n16250 & n16277 ) ;
  assign n16280 = ( ~n16250 & n16278 ) | ( ~n16250 & n16279 ) | ( n16278 & n16279 ) ;
  assign n16281 = ( n16190 & n16241 ) | ( n16190 & ~n16280 ) | ( n16241 & ~n16280 ) ;
  assign n16282 = ( ~n16190 & n16241 ) | ( ~n16190 & n16280 ) | ( n16241 & n16280 ) ;
  assign n16283 = ( ~n16241 & n16281 ) | ( ~n16241 & n16282 ) | ( n16281 & n16282 ) ;
  assign n16284 = ( n16193 & n16232 ) | ( n16193 & ~n16283 ) | ( n16232 & ~n16283 ) ;
  assign n16285 = ( ~n16193 & n16232 ) | ( ~n16193 & n16283 ) | ( n16232 & n16283 ) ;
  assign n16286 = ( ~n16232 & n16284 ) | ( ~n16232 & n16285 ) | ( n16284 & n16285 ) ;
  assign n16287 = ( n16196 & n16223 ) | ( n16196 & ~n16286 ) | ( n16223 & ~n16286 ) ;
  assign n16288 = ( ~n16196 & n16223 ) | ( ~n16196 & n16286 ) | ( n16223 & n16286 ) ;
  assign n16289 = ( ~n16223 & n16287 ) | ( ~n16223 & n16288 ) | ( n16287 & n16288 ) ;
  assign n16290 = ( n16199 & n16214 ) | ( n16199 & ~n16289 ) | ( n16214 & ~n16289 ) ;
  assign n16291 = ( ~n16199 & n16214 ) | ( ~n16199 & n16289 ) | ( n16214 & n16289 ) ;
  assign n16292 = ( ~n16214 & n16290 ) | ( ~n16214 & n16291 ) | ( n16290 & n16291 ) ;
  assign n16293 = ( ~n16202 & n16205 ) | ( ~n16202 & n16292 ) | ( n16205 & n16292 ) ;
  assign n16294 = ( n16205 & n16292 ) | ( n16205 & ~n16293 ) | ( n16292 & ~n16293 ) ;
  assign n16295 = ( n16202 & n16293 ) | ( n16202 & ~n16294 ) | ( n16293 & ~n16294 ) ;
  assign n16296 = n4227 & n8862 ;
  assign n16297 = ( x127 & n4470 ) | ( x127 & n16296 ) | ( n4470 & n16296 ) ;
  assign n16298 = x44 | n16297 ;
  assign n16299 = ~x44 & n16297 ;
  assign n16300 = ( ~n16297 & n16298 ) | ( ~n16297 & n16299 ) | ( n16298 & n16299 ) ;
  assign n16301 = n4787 & n8587 ;
  assign n16302 = x125 & n4791 ;
  assign n16303 = x126 | n16302 ;
  assign n16304 = ( n4793 & n16302 ) | ( n4793 & n16303 ) | ( n16302 & n16303 ) ;
  assign n16305 = x124 & n5030 ;
  assign n16306 = n16304 | n16305 ;
  assign n16307 = ( x47 & n16301 ) | ( x47 & ~n16306 ) | ( n16301 & ~n16306 ) ;
  assign n16308 = ( ~x47 & n16306 ) | ( ~x47 & n16307 ) | ( n16306 & n16307 ) ;
  assign n16309 = ( ~n16301 & n16307 ) | ( ~n16301 & n16308 ) | ( n16307 & n16308 ) ;
  assign n16310 = n5374 & n7597 ;
  assign n16311 = x122 & n5378 ;
  assign n16312 = x123 | n16311 ;
  assign n16313 = ( n5380 & n16311 ) | ( n5380 & n16312 ) | ( n16311 & n16312 ) ;
  assign n16314 = x121 & n5638 ;
  assign n16315 = n16313 | n16314 ;
  assign n16316 = ( x50 & n16310 ) | ( x50 & ~n16315 ) | ( n16310 & ~n16315 ) ;
  assign n16317 = ( ~x50 & n16315 ) | ( ~x50 & n16316 ) | ( n16315 & n16316 ) ;
  assign n16318 = ( ~n16310 & n16316 ) | ( ~n16310 & n16317 ) | ( n16316 & n16317 ) ;
  assign n16319 = n6027 & n7098 ;
  assign n16320 = x119 & n6031 ;
  assign n16321 = x120 | n16320 ;
  assign n16322 = ( n6033 & n16320 ) | ( n6033 & n16321 ) | ( n16320 & n16321 ) ;
  assign n16323 = x118 & n6303 ;
  assign n16324 = n16322 | n16323 ;
  assign n16325 = ( x53 & n16319 ) | ( x53 & ~n16324 ) | ( n16319 & ~n16324 ) ;
  assign n16326 = ( ~x53 & n16324 ) | ( ~x53 & n16325 ) | ( n16324 & n16325 ) ;
  assign n16327 = ( ~n16319 & n16325 ) | ( ~n16319 & n16326 ) | ( n16325 & n16326 ) ;
  assign n16328 = n6201 & n6713 ;
  assign n16329 = x116 & n6717 ;
  assign n16330 = x117 | n16329 ;
  assign n16331 = ( n6719 & n16329 ) | ( n6719 & n16330 ) | ( n16329 & n16330 ) ;
  assign n16332 = x115 & n6980 ;
  assign n16333 = n16331 | n16332 ;
  assign n16334 = ( x56 & n16328 ) | ( x56 & ~n16333 ) | ( n16328 & ~n16333 ) ;
  assign n16335 = ( ~x56 & n16333 ) | ( ~x56 & n16334 ) | ( n16333 & n16334 ) ;
  assign n16336 = ( ~n16328 & n16334 ) | ( ~n16328 & n16335 ) | ( n16334 & n16335 ) ;
  assign n16337 = n5750 & n7423 ;
  assign n16338 = x113 & n7427 ;
  assign n16339 = x114 | n16338 ;
  assign n16340 = ( n7429 & n16338 ) | ( n7429 & n16339 ) | ( n16338 & n16339 ) ;
  assign n16341 = x112 & n7708 ;
  assign n16342 = n16340 | n16341 ;
  assign n16343 = ( x59 & n16337 ) | ( x59 & ~n16342 ) | ( n16337 & ~n16342 ) ;
  assign n16344 = ( ~x59 & n16342 ) | ( ~x59 & n16343 ) | ( n16342 & n16343 ) ;
  assign n16345 = ( ~n16337 & n16343 ) | ( ~n16337 & n16344 ) | ( n16343 & n16344 ) ;
  assign n16346 = x107 & n8927 ;
  assign n16347 = ( ~x108 & n8693 ) | ( ~x108 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16348 = ( n8693 & n16346 ) | ( n8693 & ~n16347 ) | ( n16346 & ~n16347 ) ;
  assign n16349 = n5130 & n8154 ;
  assign n16350 = x110 & n8158 ;
  assign n16351 = x111 | n16350 ;
  assign n16352 = ( n8160 & n16350 ) | ( n8160 & n16351 ) | ( n16350 & n16351 ) ;
  assign n16353 = x109 & n8439 ;
  assign n16354 = n16352 | n16353 ;
  assign n16355 = ( x62 & n16349 ) | ( x62 & ~n16354 ) | ( n16349 & ~n16354 ) ;
  assign n16356 = ( ~x62 & n16354 ) | ( ~x62 & n16355 ) | ( n16354 & n16355 ) ;
  assign n16357 = ( ~n16349 & n16355 ) | ( ~n16349 & n16356 ) | ( n16355 & n16356 ) ;
  assign n16358 = ( ~n16271 & n16348 ) | ( ~n16271 & n16357 ) | ( n16348 & n16357 ) ;
  assign n16359 = ( n16348 & n16357 ) | ( n16348 & ~n16358 ) | ( n16357 & ~n16358 ) ;
  assign n16360 = ( n16271 & n16358 ) | ( n16271 & ~n16359 ) | ( n16358 & ~n16359 ) ;
  assign n16361 = ( n16272 & n16345 ) | ( n16272 & ~n16360 ) | ( n16345 & ~n16360 ) ;
  assign n16362 = ( ~n16272 & n16345 ) | ( ~n16272 & n16360 ) | ( n16345 & n16360 ) ;
  assign n16363 = ( ~n16345 & n16361 ) | ( ~n16345 & n16362 ) | ( n16361 & n16362 ) ;
  assign n16364 = ( n16275 & n16336 ) | ( n16275 & ~n16363 ) | ( n16336 & ~n16363 ) ;
  assign n16365 = ( ~n16275 & n16336 ) | ( ~n16275 & n16363 ) | ( n16336 & n16363 ) ;
  assign n16366 = ( ~n16336 & n16364 ) | ( ~n16336 & n16365 ) | ( n16364 & n16365 ) ;
  assign n16367 = ( n16278 & n16327 ) | ( n16278 & ~n16366 ) | ( n16327 & ~n16366 ) ;
  assign n16368 = ( ~n16278 & n16327 ) | ( ~n16278 & n16366 ) | ( n16327 & n16366 ) ;
  assign n16369 = ( ~n16327 & n16367 ) | ( ~n16327 & n16368 ) | ( n16367 & n16368 ) ;
  assign n16370 = ( n16281 & n16318 ) | ( n16281 & ~n16369 ) | ( n16318 & ~n16369 ) ;
  assign n16371 = ( ~n16281 & n16318 ) | ( ~n16281 & n16369 ) | ( n16318 & n16369 ) ;
  assign n16372 = ( ~n16318 & n16370 ) | ( ~n16318 & n16371 ) | ( n16370 & n16371 ) ;
  assign n16373 = ( n16284 & n16309 ) | ( n16284 & ~n16372 ) | ( n16309 & ~n16372 ) ;
  assign n16374 = ( ~n16284 & n16309 ) | ( ~n16284 & n16372 ) | ( n16309 & n16372 ) ;
  assign n16375 = ( ~n16309 & n16373 ) | ( ~n16309 & n16374 ) | ( n16373 & n16374 ) ;
  assign n16376 = ( n16287 & n16300 ) | ( n16287 & ~n16375 ) | ( n16300 & ~n16375 ) ;
  assign n16377 = ( ~n16287 & n16300 ) | ( ~n16287 & n16375 ) | ( n16300 & n16375 ) ;
  assign n16378 = ( ~n16300 & n16376 ) | ( ~n16300 & n16377 ) | ( n16376 & n16377 ) ;
  assign n16379 = ( ~n16290 & n16293 ) | ( ~n16290 & n16378 ) | ( n16293 & n16378 ) ;
  assign n16380 = ( n16293 & n16378 ) | ( n16293 & ~n16379 ) | ( n16378 & ~n16379 ) ;
  assign n16381 = ( n16290 & n16379 ) | ( n16290 & ~n16380 ) | ( n16379 & ~n16380 ) ;
  assign n16382 = n4787 & n8846 ;
  assign n16383 = x126 & n4791 ;
  assign n16384 = x127 | n16383 ;
  assign n16385 = ( n4793 & n16383 ) | ( n4793 & n16384 ) | ( n16383 & n16384 ) ;
  assign n16386 = x125 & n5030 ;
  assign n16387 = n16385 | n16386 ;
  assign n16388 = ( x47 & n16382 ) | ( x47 & ~n16387 ) | ( n16382 & ~n16387 ) ;
  assign n16389 = ( ~x47 & n16387 ) | ( ~x47 & n16388 ) | ( n16387 & n16388 ) ;
  assign n16390 = ( ~n16382 & n16388 ) | ( ~n16382 & n16389 ) | ( n16388 & n16389 ) ;
  assign n16391 = n5374 & n7841 ;
  assign n16392 = x123 & n5378 ;
  assign n16393 = x124 | n16392 ;
  assign n16394 = ( n5380 & n16392 ) | ( n5380 & n16393 ) | ( n16392 & n16393 ) ;
  assign n16395 = x122 & n5638 ;
  assign n16396 = n16394 | n16395 ;
  assign n16397 = ( x50 & n16391 ) | ( x50 & ~n16396 ) | ( n16391 & ~n16396 ) ;
  assign n16398 = ( ~x50 & n16396 ) | ( ~x50 & n16397 ) | ( n16396 & n16397 ) ;
  assign n16399 = ( ~n16391 & n16397 ) | ( ~n16391 & n16398 ) | ( n16397 & n16398 ) ;
  assign n16400 = n6027 & n7113 ;
  assign n16401 = x120 & n6031 ;
  assign n16402 = x121 | n16401 ;
  assign n16403 = ( n6033 & n16401 ) | ( n6033 & n16402 ) | ( n16401 & n16402 ) ;
  assign n16404 = x119 & n6303 ;
  assign n16405 = n16403 | n16404 ;
  assign n16406 = ( x53 & n16400 ) | ( x53 & ~n16405 ) | ( n16400 & ~n16405 ) ;
  assign n16407 = ( ~x53 & n16405 ) | ( ~x53 & n16406 ) | ( n16405 & n16406 ) ;
  assign n16408 = ( ~n16400 & n16406 ) | ( ~n16400 & n16407 ) | ( n16406 & n16407 ) ;
  assign n16409 = n6421 & n6713 ;
  assign n16410 = x117 & n6717 ;
  assign n16411 = x118 | n16410 ;
  assign n16412 = ( n6719 & n16410 ) | ( n6719 & n16411 ) | ( n16410 & n16411 ) ;
  assign n16413 = x116 & n6980 ;
  assign n16414 = n16412 | n16413 ;
  assign n16415 = ( x56 & n16409 ) | ( x56 & ~n16414 ) | ( n16409 & ~n16414 ) ;
  assign n16416 = ( ~x56 & n16414 ) | ( ~x56 & n16415 ) | ( n16414 & n16415 ) ;
  assign n16417 = ( ~n16409 & n16415 ) | ( ~n16409 & n16416 ) | ( n16415 & n16416 ) ;
  assign n16418 = n5765 & n7423 ;
  assign n16419 = x114 & n7427 ;
  assign n16420 = x115 | n16419 ;
  assign n16421 = ( n7429 & n16419 ) | ( n7429 & n16420 ) | ( n16419 & n16420 ) ;
  assign n16422 = x113 & n7708 ;
  assign n16423 = n16421 | n16422 ;
  assign n16424 = ( x59 & n16418 ) | ( x59 & ~n16423 ) | ( n16418 & ~n16423 ) ;
  assign n16425 = ( ~x59 & n16423 ) | ( ~x59 & n16424 ) | ( n16423 & n16424 ) ;
  assign n16426 = ( ~n16418 & n16424 ) | ( ~n16418 & n16425 ) | ( n16424 & n16425 ) ;
  assign n16427 = n5145 & n8154 ;
  assign n16428 = x111 & n8158 ;
  assign n16429 = x112 | n16428 ;
  assign n16430 = ( n8160 & n16428 ) | ( n8160 & n16429 ) | ( n16428 & n16429 ) ;
  assign n16431 = x110 & n8439 ;
  assign n16432 = n16430 | n16431 ;
  assign n16433 = ( x62 & n16427 ) | ( x62 & ~n16432 ) | ( n16427 & ~n16432 ) ;
  assign n16434 = ( ~x62 & n16432 ) | ( ~x62 & n16433 ) | ( n16432 & n16433 ) ;
  assign n16435 = ( ~n16427 & n16433 ) | ( ~n16427 & n16434 ) | ( n16433 & n16434 ) ;
  assign n16436 = x108 & n8927 ;
  assign n16437 = ( ~x109 & n8693 ) | ( ~x109 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16438 = ( n8693 & n16436 ) | ( n8693 & ~n16437 ) | ( n16436 & ~n16437 ) ;
  assign n16439 = ( ~x44 & n16271 ) | ( ~x44 & n16438 ) | ( n16271 & n16438 ) ;
  assign n16440 = ( n16271 & n16438 ) | ( n16271 & ~n16439 ) | ( n16438 & ~n16439 ) ;
  assign n16441 = ( x44 & n16439 ) | ( x44 & ~n16440 ) | ( n16439 & ~n16440 ) ;
  assign n16442 = ( n16358 & n16435 ) | ( n16358 & ~n16441 ) | ( n16435 & ~n16441 ) ;
  assign n16443 = ( ~n16358 & n16435 ) | ( ~n16358 & n16441 ) | ( n16435 & n16441 ) ;
  assign n16444 = ( ~n16435 & n16442 ) | ( ~n16435 & n16443 ) | ( n16442 & n16443 ) ;
  assign n16445 = ( n16361 & n16426 ) | ( n16361 & ~n16444 ) | ( n16426 & ~n16444 ) ;
  assign n16446 = ( ~n16361 & n16426 ) | ( ~n16361 & n16444 ) | ( n16426 & n16444 ) ;
  assign n16447 = ( ~n16426 & n16445 ) | ( ~n16426 & n16446 ) | ( n16445 & n16446 ) ;
  assign n16448 = ( n16364 & n16417 ) | ( n16364 & ~n16447 ) | ( n16417 & ~n16447 ) ;
  assign n16449 = ( ~n16364 & n16417 ) | ( ~n16364 & n16447 ) | ( n16417 & n16447 ) ;
  assign n16450 = ( ~n16417 & n16448 ) | ( ~n16417 & n16449 ) | ( n16448 & n16449 ) ;
  assign n16451 = ( n16367 & n16408 ) | ( n16367 & ~n16450 ) | ( n16408 & ~n16450 ) ;
  assign n16452 = ( ~n16367 & n16408 ) | ( ~n16367 & n16450 ) | ( n16408 & n16450 ) ;
  assign n16453 = ( ~n16408 & n16451 ) | ( ~n16408 & n16452 ) | ( n16451 & n16452 ) ;
  assign n16454 = ( n16370 & n16399 ) | ( n16370 & ~n16453 ) | ( n16399 & ~n16453 ) ;
  assign n16455 = ( ~n16370 & n16399 ) | ( ~n16370 & n16453 ) | ( n16399 & n16453 ) ;
  assign n16456 = ( ~n16399 & n16454 ) | ( ~n16399 & n16455 ) | ( n16454 & n16455 ) ;
  assign n16457 = ( n16373 & n16390 ) | ( n16373 & ~n16456 ) | ( n16390 & ~n16456 ) ;
  assign n16458 = ( ~n16373 & n16390 ) | ( ~n16373 & n16456 ) | ( n16390 & n16456 ) ;
  assign n16459 = ( ~n16390 & n16457 ) | ( ~n16390 & n16458 ) | ( n16457 & n16458 ) ;
  assign n16460 = ( ~n16376 & n16379 ) | ( ~n16376 & n16459 ) | ( n16379 & n16459 ) ;
  assign n16461 = ( n16379 & n16459 ) | ( n16379 & ~n16460 ) | ( n16459 & ~n16460 ) ;
  assign n16462 = ( n16376 & n16460 ) | ( n16376 & ~n16461 ) | ( n16460 & ~n16461 ) ;
  assign n16463 = n4787 & n8865 ;
  assign n16464 = x127 & n4791 ;
  assign n16465 = x126 | n16464 ;
  assign n16466 = ( n5030 & n16464 ) | ( n5030 & n16465 ) | ( n16464 & n16465 ) ;
  assign n16467 = ( x47 & n16463 ) | ( x47 & ~n16466 ) | ( n16463 & ~n16466 ) ;
  assign n16468 = ( ~x47 & n16466 ) | ( ~x47 & n16467 ) | ( n16466 & n16467 ) ;
  assign n16469 = ( ~n16463 & n16467 ) | ( ~n16463 & n16468 ) | ( n16467 & n16468 ) ;
  assign n16470 = n5374 & n8331 ;
  assign n16471 = x124 & n5378 ;
  assign n16472 = x125 | n16471 ;
  assign n16473 = ( n5380 & n16471 ) | ( n5380 & n16472 ) | ( n16471 & n16472 ) ;
  assign n16474 = x123 & n5638 ;
  assign n16475 = n16473 | n16474 ;
  assign n16476 = ( x50 & n16470 ) | ( x50 & ~n16475 ) | ( n16470 & ~n16475 ) ;
  assign n16477 = ( ~x50 & n16475 ) | ( ~x50 & n16476 ) | ( n16475 & n16476 ) ;
  assign n16478 = ( ~n16470 & n16476 ) | ( ~n16470 & n16477 ) | ( n16476 & n16477 ) ;
  assign n16479 = n6027 & n7582 ;
  assign n16480 = x121 & n6031 ;
  assign n16481 = x122 | n16480 ;
  assign n16482 = ( n6033 & n16480 ) | ( n6033 & n16481 ) | ( n16480 & n16481 ) ;
  assign n16483 = x120 & n6303 ;
  assign n16484 = n16482 | n16483 ;
  assign n16485 = ( x53 & n16479 ) | ( x53 & ~n16484 ) | ( n16479 & ~n16484 ) ;
  assign n16486 = ( ~x53 & n16484 ) | ( ~x53 & n16485 ) | ( n16484 & n16485 ) ;
  assign n16487 = ( ~n16479 & n16485 ) | ( ~n16479 & n16486 ) | ( n16485 & n16486 ) ;
  assign n16488 = n6645 & n6713 ;
  assign n16489 = x118 & n6717 ;
  assign n16490 = x119 | n16489 ;
  assign n16491 = ( n6719 & n16489 ) | ( n6719 & n16490 ) | ( n16489 & n16490 ) ;
  assign n16492 = x117 & n6980 ;
  assign n16493 = n16491 | n16492 ;
  assign n16494 = ( x56 & n16488 ) | ( x56 & ~n16493 ) | ( n16488 & ~n16493 ) ;
  assign n16495 = ( ~x56 & n16493 ) | ( ~x56 & n16494 ) | ( n16493 & n16494 ) ;
  assign n16496 = ( ~n16488 & n16494 ) | ( ~n16488 & n16495 ) | ( n16494 & n16495 ) ;
  assign n16497 = n5977 & n7423 ;
  assign n16498 = x115 & n7427 ;
  assign n16499 = x116 | n16498 ;
  assign n16500 = ( n7429 & n16498 ) | ( n7429 & n16499 ) | ( n16498 & n16499 ) ;
  assign n16501 = x114 & n7708 ;
  assign n16502 = n16500 | n16501 ;
  assign n16503 = ( x59 & n16497 ) | ( x59 & ~n16502 ) | ( n16497 & ~n16502 ) ;
  assign n16504 = ( ~x59 & n16502 ) | ( ~x59 & n16503 ) | ( n16502 & n16503 ) ;
  assign n16505 = ( ~n16497 & n16503 ) | ( ~n16497 & n16504 ) | ( n16503 & n16504 ) ;
  assign n16506 = n5542 & n8154 ;
  assign n16507 = x112 & n8158 ;
  assign n16508 = x113 | n16507 ;
  assign n16509 = ( n8160 & n16507 ) | ( n8160 & n16508 ) | ( n16507 & n16508 ) ;
  assign n16510 = x111 & n8439 ;
  assign n16511 = n16509 | n16510 ;
  assign n16512 = ( x62 & n16506 ) | ( x62 & ~n16511 ) | ( n16506 & ~n16511 ) ;
  assign n16513 = ( ~x62 & n16511 ) | ( ~x62 & n16512 ) | ( n16511 & n16512 ) ;
  assign n16514 = ( ~n16506 & n16512 ) | ( ~n16506 & n16513 ) | ( n16512 & n16513 ) ;
  assign n16515 = x109 & n8927 ;
  assign n16516 = ( ~x110 & n8693 ) | ( ~x110 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16517 = ( n8693 & n16515 ) | ( n8693 & ~n16516 ) | ( n16515 & ~n16516 ) ;
  assign n16518 = ( ~n16439 & n16514 ) | ( ~n16439 & n16517 ) | ( n16514 & n16517 ) ;
  assign n16519 = ( n16514 & n16517 ) | ( n16514 & ~n16518 ) | ( n16517 & ~n16518 ) ;
  assign n16520 = ( n16439 & n16518 ) | ( n16439 & ~n16519 ) | ( n16518 & ~n16519 ) ;
  assign n16521 = ( n16442 & n16505 ) | ( n16442 & ~n16520 ) | ( n16505 & ~n16520 ) ;
  assign n16522 = ( ~n16442 & n16505 ) | ( ~n16442 & n16520 ) | ( n16505 & n16520 ) ;
  assign n16523 = ( ~n16505 & n16521 ) | ( ~n16505 & n16522 ) | ( n16521 & n16522 ) ;
  assign n16524 = ( n16445 & n16496 ) | ( n16445 & ~n16523 ) | ( n16496 & ~n16523 ) ;
  assign n16525 = ( ~n16445 & n16496 ) | ( ~n16445 & n16523 ) | ( n16496 & n16523 ) ;
  assign n16526 = ( ~n16496 & n16524 ) | ( ~n16496 & n16525 ) | ( n16524 & n16525 ) ;
  assign n16527 = ( n16448 & n16487 ) | ( n16448 & ~n16526 ) | ( n16487 & ~n16526 ) ;
  assign n16528 = ( ~n16448 & n16487 ) | ( ~n16448 & n16526 ) | ( n16487 & n16526 ) ;
  assign n16529 = ( ~n16487 & n16527 ) | ( ~n16487 & n16528 ) | ( n16527 & n16528 ) ;
  assign n16530 = ( n16451 & n16478 ) | ( n16451 & ~n16529 ) | ( n16478 & ~n16529 ) ;
  assign n16531 = ( ~n16451 & n16478 ) | ( ~n16451 & n16529 ) | ( n16478 & n16529 ) ;
  assign n16532 = ( ~n16478 & n16530 ) | ( ~n16478 & n16531 ) | ( n16530 & n16531 ) ;
  assign n16533 = ( n16454 & n16469 ) | ( n16454 & ~n16532 ) | ( n16469 & ~n16532 ) ;
  assign n16534 = ( ~n16454 & n16469 ) | ( ~n16454 & n16532 ) | ( n16469 & n16532 ) ;
  assign n16535 = ( ~n16469 & n16533 ) | ( ~n16469 & n16534 ) | ( n16533 & n16534 ) ;
  assign n16536 = ( ~n16457 & n16460 ) | ( ~n16457 & n16535 ) | ( n16460 & n16535 ) ;
  assign n16537 = ( n16460 & n16535 ) | ( n16460 & ~n16536 ) | ( n16535 & ~n16536 ) ;
  assign n16538 = ( n16457 & n16536 ) | ( n16457 & ~n16537 ) | ( n16536 & ~n16537 ) ;
  assign n16539 = n4787 & n8862 ;
  assign n16540 = ( x127 & n5030 ) | ( x127 & n16539 ) | ( n5030 & n16539 ) ;
  assign n16541 = x47 | n16540 ;
  assign n16542 = ~x47 & n16540 ;
  assign n16543 = ( ~n16540 & n16541 ) | ( ~n16540 & n16542 ) | ( n16541 & n16542 ) ;
  assign n16544 = n5374 & n8587 ;
  assign n16545 = x125 & n5378 ;
  assign n16546 = x126 | n16545 ;
  assign n16547 = ( n5380 & n16545 ) | ( n5380 & n16546 ) | ( n16545 & n16546 ) ;
  assign n16548 = x124 & n5638 ;
  assign n16549 = n16547 | n16548 ;
  assign n16550 = ( x50 & n16544 ) | ( x50 & ~n16549 ) | ( n16544 & ~n16549 ) ;
  assign n16551 = ( ~x50 & n16549 ) | ( ~x50 & n16550 ) | ( n16549 & n16550 ) ;
  assign n16552 = ( ~n16544 & n16550 ) | ( ~n16544 & n16551 ) | ( n16550 & n16551 ) ;
  assign n16553 = n6713 & n7098 ;
  assign n16554 = x119 & n6717 ;
  assign n16555 = x120 | n16554 ;
  assign n16556 = ( n6719 & n16554 ) | ( n6719 & n16555 ) | ( n16554 & n16555 ) ;
  assign n16557 = x118 & n6980 ;
  assign n16558 = n16556 | n16557 ;
  assign n16559 = ( x56 & n16553 ) | ( x56 & ~n16558 ) | ( n16553 & ~n16558 ) ;
  assign n16560 = ( ~x56 & n16558 ) | ( ~x56 & n16559 ) | ( n16558 & n16559 ) ;
  assign n16561 = ( ~n16553 & n16559 ) | ( ~n16553 & n16560 ) | ( n16559 & n16560 ) ;
  assign n16562 = x110 & n8927 ;
  assign n16563 = ( ~x111 & n8693 ) | ( ~x111 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16564 = ( n8693 & n16562 ) | ( n8693 & ~n16563 ) | ( n16562 & ~n16563 ) ;
  assign n16565 = ( n16439 & n16518 ) | ( n16439 & ~n16564 ) | ( n16518 & ~n16564 ) ;
  assign n16566 = ( n16439 & ~n16518 ) | ( n16439 & n16564 ) | ( ~n16518 & n16564 ) ;
  assign n16567 = ( ~n16439 & n16565 ) | ( ~n16439 & n16566 ) | ( n16565 & n16566 ) ;
  assign n16568 = n6201 & n7423 ;
  assign n16569 = x116 & n7427 ;
  assign n16570 = x117 | n16569 ;
  assign n16571 = ( n7429 & n16569 ) | ( n7429 & n16570 ) | ( n16569 & n16570 ) ;
  assign n16572 = x115 & n7708 ;
  assign n16573 = n16571 | n16572 ;
  assign n16574 = ( x59 & n16568 ) | ( x59 & ~n16573 ) | ( n16568 & ~n16573 ) ;
  assign n16575 = ( ~x59 & n16573 ) | ( ~x59 & n16574 ) | ( n16573 & n16574 ) ;
  assign n16576 = ( ~n16568 & n16574 ) | ( ~n16568 & n16575 ) | ( n16574 & n16575 ) ;
  assign n16577 = n5750 & n8154 ;
  assign n16578 = x113 & n8158 ;
  assign n16579 = x114 | n16578 ;
  assign n16580 = ( n8160 & n16578 ) | ( n8160 & n16579 ) | ( n16578 & n16579 ) ;
  assign n16581 = x112 & n8439 ;
  assign n16582 = n16580 | n16581 ;
  assign n16583 = ( x62 & n16577 ) | ( x62 & ~n16582 ) | ( n16577 & ~n16582 ) ;
  assign n16584 = ( ~x62 & n16582 ) | ( ~x62 & n16583 ) | ( n16582 & n16583 ) ;
  assign n16585 = ( ~n16577 & n16583 ) | ( ~n16577 & n16584 ) | ( n16583 & n16584 ) ;
  assign n16586 = ( ~n16567 & n16576 ) | ( ~n16567 & n16585 ) | ( n16576 & n16585 ) ;
  assign n16587 = ( n16576 & n16585 ) | ( n16576 & ~n16586 ) | ( n16585 & ~n16586 ) ;
  assign n16588 = ( n16567 & n16586 ) | ( n16567 & ~n16587 ) | ( n16586 & ~n16587 ) ;
  assign n16589 = ( n16521 & n16561 ) | ( n16521 & ~n16588 ) | ( n16561 & ~n16588 ) ;
  assign n16590 = ( ~n16521 & n16561 ) | ( ~n16521 & n16588 ) | ( n16561 & n16588 ) ;
  assign n16591 = ( ~n16561 & n16589 ) | ( ~n16561 & n16590 ) | ( n16589 & n16590 ) ;
  assign n16592 = n6027 & n7597 ;
  assign n16593 = x122 & n6031 ;
  assign n16594 = x123 | n16593 ;
  assign n16595 = ( n6033 & n16593 ) | ( n6033 & n16594 ) | ( n16593 & n16594 ) ;
  assign n16596 = x121 & n6303 ;
  assign n16597 = n16595 | n16596 ;
  assign n16598 = ( x53 & n16592 ) | ( x53 & ~n16597 ) | ( n16592 & ~n16597 ) ;
  assign n16599 = ( ~x53 & n16597 ) | ( ~x53 & n16598 ) | ( n16597 & n16598 ) ;
  assign n16600 = ( ~n16592 & n16598 ) | ( ~n16592 & n16599 ) | ( n16598 & n16599 ) ;
  assign n16601 = ( n16524 & ~n16591 ) | ( n16524 & n16600 ) | ( ~n16591 & n16600 ) ;
  assign n16602 = ( n16524 & n16591 ) | ( n16524 & n16600 ) | ( n16591 & n16600 ) ;
  assign n16603 = ( n16591 & n16601 ) | ( n16591 & ~n16602 ) | ( n16601 & ~n16602 ) ;
  assign n16604 = ( n16527 & n16552 ) | ( n16527 & ~n16603 ) | ( n16552 & ~n16603 ) ;
  assign n16605 = ( ~n16527 & n16552 ) | ( ~n16527 & n16603 ) | ( n16552 & n16603 ) ;
  assign n16606 = ( ~n16552 & n16604 ) | ( ~n16552 & n16605 ) | ( n16604 & n16605 ) ;
  assign n16607 = ( n16530 & n16543 ) | ( n16530 & ~n16606 ) | ( n16543 & ~n16606 ) ;
  assign n16608 = ( ~n16530 & n16543 ) | ( ~n16530 & n16606 ) | ( n16543 & n16606 ) ;
  assign n16609 = ( ~n16543 & n16607 ) | ( ~n16543 & n16608 ) | ( n16607 & n16608 ) ;
  assign n16610 = ( ~n16533 & n16536 ) | ( ~n16533 & n16609 ) | ( n16536 & n16609 ) ;
  assign n16611 = ( n16536 & n16609 ) | ( n16536 & ~n16610 ) | ( n16609 & ~n16610 ) ;
  assign n16612 = ( n16533 & n16610 ) | ( n16533 & ~n16611 ) | ( n16610 & ~n16611 ) ;
  assign n16613 = n5374 & n8846 ;
  assign n16614 = x126 & n5378 ;
  assign n16615 = x127 | n16614 ;
  assign n16616 = ( n5380 & n16614 ) | ( n5380 & n16615 ) | ( n16614 & n16615 ) ;
  assign n16617 = x125 & n5638 ;
  assign n16618 = n16616 | n16617 ;
  assign n16619 = ( x50 & n16613 ) | ( x50 & ~n16618 ) | ( n16613 & ~n16618 ) ;
  assign n16620 = ( ~x50 & n16618 ) | ( ~x50 & n16619 ) | ( n16618 & n16619 ) ;
  assign n16621 = ( ~n16613 & n16619 ) | ( ~n16613 & n16620 ) | ( n16619 & n16620 ) ;
  assign n16622 = n6027 & n7841 ;
  assign n16623 = x123 & n6031 ;
  assign n16624 = x124 | n16623 ;
  assign n16625 = ( n6033 & n16623 ) | ( n6033 & n16624 ) | ( n16623 & n16624 ) ;
  assign n16626 = x122 & n6303 ;
  assign n16627 = n16625 | n16626 ;
  assign n16628 = ( x53 & n16622 ) | ( x53 & ~n16627 ) | ( n16622 & ~n16627 ) ;
  assign n16629 = ( ~x53 & n16627 ) | ( ~x53 & n16628 ) | ( n16627 & n16628 ) ;
  assign n16630 = ( ~n16622 & n16628 ) | ( ~n16622 & n16629 ) | ( n16628 & n16629 ) ;
  assign n16631 = n6713 & n7113 ;
  assign n16632 = x120 & n6717 ;
  assign n16633 = x121 | n16632 ;
  assign n16634 = ( n6719 & n16632 ) | ( n6719 & n16633 ) | ( n16632 & n16633 ) ;
  assign n16635 = x119 & n6980 ;
  assign n16636 = n16634 | n16635 ;
  assign n16637 = ( x56 & n16631 ) | ( x56 & ~n16636 ) | ( n16631 & ~n16636 ) ;
  assign n16638 = ( ~x56 & n16636 ) | ( ~x56 & n16637 ) | ( n16636 & n16637 ) ;
  assign n16639 = ( ~n16631 & n16637 ) | ( ~n16631 & n16638 ) | ( n16637 & n16638 ) ;
  assign n16640 = n6421 & n7423 ;
  assign n16641 = x117 & n7427 ;
  assign n16642 = x118 | n16641 ;
  assign n16643 = ( n7429 & n16641 ) | ( n7429 & n16642 ) | ( n16641 & n16642 ) ;
  assign n16644 = x116 & n7708 ;
  assign n16645 = n16643 | n16644 ;
  assign n16646 = ( x59 & n16640 ) | ( x59 & ~n16645 ) | ( n16640 & ~n16645 ) ;
  assign n16647 = ( ~x59 & n16645 ) | ( ~x59 & n16646 ) | ( n16645 & n16646 ) ;
  assign n16648 = ( ~n16640 & n16646 ) | ( ~n16640 & n16647 ) | ( n16646 & n16647 ) ;
  assign n16649 = n5765 & n8154 ;
  assign n16650 = x114 & n8158 ;
  assign n16651 = x115 | n16650 ;
  assign n16652 = ( n8160 & n16650 ) | ( n8160 & n16651 ) | ( n16650 & n16651 ) ;
  assign n16653 = x113 & n8439 ;
  assign n16654 = n16652 | n16653 ;
  assign n16655 = ( x62 & n16649 ) | ( x62 & ~n16654 ) | ( n16649 & ~n16654 ) ;
  assign n16656 = ( ~x62 & n16654 ) | ( ~x62 & n16655 ) | ( n16654 & n16655 ) ;
  assign n16657 = ( ~n16649 & n16655 ) | ( ~n16649 & n16656 ) | ( n16655 & n16656 ) ;
  assign n16658 = x111 & n8927 ;
  assign n16659 = ( ~x112 & n8693 ) | ( ~x112 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16660 = ( n8693 & n16658 ) | ( n8693 & ~n16659 ) | ( n16658 & ~n16659 ) ;
  assign n16661 = ( ~x47 & n16564 ) | ( ~x47 & n16660 ) | ( n16564 & n16660 ) ;
  assign n16662 = ( n16564 & n16660 ) | ( n16564 & ~n16661 ) | ( n16660 & ~n16661 ) ;
  assign n16663 = ( x47 & n16661 ) | ( x47 & ~n16662 ) | ( n16661 & ~n16662 ) ;
  assign n16664 = ( n16565 & n16657 ) | ( n16565 & ~n16663 ) | ( n16657 & ~n16663 ) ;
  assign n16665 = ( ~n16565 & n16657 ) | ( ~n16565 & n16663 ) | ( n16657 & n16663 ) ;
  assign n16666 = ( ~n16657 & n16664 ) | ( ~n16657 & n16665 ) | ( n16664 & n16665 ) ;
  assign n16667 = ( n16586 & n16648 ) | ( n16586 & ~n16666 ) | ( n16648 & ~n16666 ) ;
  assign n16668 = ( ~n16586 & n16648 ) | ( ~n16586 & n16666 ) | ( n16648 & n16666 ) ;
  assign n16669 = ( ~n16648 & n16667 ) | ( ~n16648 & n16668 ) | ( n16667 & n16668 ) ;
  assign n16670 = ( n16589 & n16639 ) | ( n16589 & ~n16669 ) | ( n16639 & ~n16669 ) ;
  assign n16671 = ( ~n16589 & n16639 ) | ( ~n16589 & n16669 ) | ( n16639 & n16669 ) ;
  assign n16672 = ( ~n16639 & n16670 ) | ( ~n16639 & n16671 ) | ( n16670 & n16671 ) ;
  assign n16673 = ( n16601 & n16630 ) | ( n16601 & ~n16672 ) | ( n16630 & ~n16672 ) ;
  assign n16674 = ( ~n16601 & n16630 ) | ( ~n16601 & n16672 ) | ( n16630 & n16672 ) ;
  assign n16675 = ( ~n16630 & n16673 ) | ( ~n16630 & n16674 ) | ( n16673 & n16674 ) ;
  assign n16676 = ( n16604 & n16621 ) | ( n16604 & ~n16675 ) | ( n16621 & ~n16675 ) ;
  assign n16677 = ( ~n16604 & n16621 ) | ( ~n16604 & n16675 ) | ( n16621 & n16675 ) ;
  assign n16678 = ( ~n16621 & n16676 ) | ( ~n16621 & n16677 ) | ( n16676 & n16677 ) ;
  assign n16679 = ( ~n16607 & n16610 ) | ( ~n16607 & n16678 ) | ( n16610 & n16678 ) ;
  assign n16680 = ( n16610 & n16678 ) | ( n16610 & ~n16679 ) | ( n16678 & ~n16679 ) ;
  assign n16681 = ( n16607 & n16679 ) | ( n16607 & ~n16680 ) | ( n16679 & ~n16680 ) ;
  assign n16682 = n5374 & n8865 ;
  assign n16683 = x127 & n5378 ;
  assign n16684 = x126 | n16683 ;
  assign n16685 = ( n5638 & n16683 ) | ( n5638 & n16684 ) | ( n16683 & n16684 ) ;
  assign n16686 = ( x50 & n16682 ) | ( x50 & ~n16685 ) | ( n16682 & ~n16685 ) ;
  assign n16687 = ( ~x50 & n16685 ) | ( ~x50 & n16686 ) | ( n16685 & n16686 ) ;
  assign n16688 = ( ~n16682 & n16686 ) | ( ~n16682 & n16687 ) | ( n16686 & n16687 ) ;
  assign n16689 = n6027 & n8331 ;
  assign n16690 = x124 & n6031 ;
  assign n16691 = x125 | n16690 ;
  assign n16692 = ( n6033 & n16690 ) | ( n6033 & n16691 ) | ( n16690 & n16691 ) ;
  assign n16693 = x123 & n6303 ;
  assign n16694 = n16692 | n16693 ;
  assign n16695 = ( x53 & n16689 ) | ( x53 & ~n16694 ) | ( n16689 & ~n16694 ) ;
  assign n16696 = ( ~x53 & n16694 ) | ( ~x53 & n16695 ) | ( n16694 & n16695 ) ;
  assign n16697 = ( ~n16689 & n16695 ) | ( ~n16689 & n16696 ) | ( n16695 & n16696 ) ;
  assign n16698 = n6713 & n7582 ;
  assign n16699 = x121 & n6717 ;
  assign n16700 = x122 | n16699 ;
  assign n16701 = ( n6719 & n16699 ) | ( n6719 & n16700 ) | ( n16699 & n16700 ) ;
  assign n16702 = x120 & n6980 ;
  assign n16703 = n16701 | n16702 ;
  assign n16704 = ( x56 & n16698 ) | ( x56 & ~n16703 ) | ( n16698 & ~n16703 ) ;
  assign n16705 = ( ~x56 & n16703 ) | ( ~x56 & n16704 ) | ( n16703 & n16704 ) ;
  assign n16706 = ( ~n16698 & n16704 ) | ( ~n16698 & n16705 ) | ( n16704 & n16705 ) ;
  assign n16707 = n6645 & n7423 ;
  assign n16708 = x118 & n7427 ;
  assign n16709 = x119 | n16708 ;
  assign n16710 = ( n7429 & n16708 ) | ( n7429 & n16709 ) | ( n16708 & n16709 ) ;
  assign n16711 = x117 & n7708 ;
  assign n16712 = n16710 | n16711 ;
  assign n16713 = ( x59 & n16707 ) | ( x59 & ~n16712 ) | ( n16707 & ~n16712 ) ;
  assign n16714 = ( ~x59 & n16712 ) | ( ~x59 & n16713 ) | ( n16712 & n16713 ) ;
  assign n16715 = ( ~n16707 & n16713 ) | ( ~n16707 & n16714 ) | ( n16713 & n16714 ) ;
  assign n16716 = x112 & n8927 ;
  assign n16717 = ( ~x113 & n8693 ) | ( ~x113 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16718 = ( n8693 & n16716 ) | ( n8693 & ~n16717 ) | ( n16716 & ~n16717 ) ;
  assign n16719 = n5977 & n8154 ;
  assign n16720 = x115 & n8158 ;
  assign n16721 = x116 | n16720 ;
  assign n16722 = ( n8160 & n16720 ) | ( n8160 & n16721 ) | ( n16720 & n16721 ) ;
  assign n16723 = x114 & n8439 ;
  assign n16724 = n16722 | n16723 ;
  assign n16725 = ( x62 & n16719 ) | ( x62 & ~n16724 ) | ( n16719 & ~n16724 ) ;
  assign n16726 = ( ~x62 & n16724 ) | ( ~x62 & n16725 ) | ( n16724 & n16725 ) ;
  assign n16727 = ( ~n16719 & n16725 ) | ( ~n16719 & n16726 ) | ( n16725 & n16726 ) ;
  assign n16728 = ( n16661 & ~n16718 ) | ( n16661 & n16727 ) | ( ~n16718 & n16727 ) ;
  assign n16729 = ( n16661 & n16718 ) | ( n16661 & n16727 ) | ( n16718 & n16727 ) ;
  assign n16730 = ( n16718 & n16728 ) | ( n16718 & ~n16729 ) | ( n16728 & ~n16729 ) ;
  assign n16731 = ( n16664 & n16715 ) | ( n16664 & ~n16730 ) | ( n16715 & ~n16730 ) ;
  assign n16732 = ( ~n16664 & n16715 ) | ( ~n16664 & n16730 ) | ( n16715 & n16730 ) ;
  assign n16733 = ( ~n16715 & n16731 ) | ( ~n16715 & n16732 ) | ( n16731 & n16732 ) ;
  assign n16734 = ( n16667 & n16706 ) | ( n16667 & ~n16733 ) | ( n16706 & ~n16733 ) ;
  assign n16735 = ( ~n16667 & n16706 ) | ( ~n16667 & n16733 ) | ( n16706 & n16733 ) ;
  assign n16736 = ( ~n16706 & n16734 ) | ( ~n16706 & n16735 ) | ( n16734 & n16735 ) ;
  assign n16737 = ( n16670 & n16697 ) | ( n16670 & ~n16736 ) | ( n16697 & ~n16736 ) ;
  assign n16738 = ( ~n16670 & n16697 ) | ( ~n16670 & n16736 ) | ( n16697 & n16736 ) ;
  assign n16739 = ( ~n16697 & n16737 ) | ( ~n16697 & n16738 ) | ( n16737 & n16738 ) ;
  assign n16740 = ( n16673 & n16688 ) | ( n16673 & ~n16739 ) | ( n16688 & ~n16739 ) ;
  assign n16741 = ( ~n16673 & n16688 ) | ( ~n16673 & n16739 ) | ( n16688 & n16739 ) ;
  assign n16742 = ( ~n16688 & n16740 ) | ( ~n16688 & n16741 ) | ( n16740 & n16741 ) ;
  assign n16743 = ( ~n16676 & n16679 ) | ( ~n16676 & n16742 ) | ( n16679 & n16742 ) ;
  assign n16744 = ( n16679 & n16742 ) | ( n16679 & ~n16743 ) | ( n16742 & ~n16743 ) ;
  assign n16745 = ( n16676 & n16743 ) | ( n16676 & ~n16744 ) | ( n16743 & ~n16744 ) ;
  assign n16746 = n5374 & n8862 ;
  assign n16747 = ( x127 & n5638 ) | ( x127 & n16746 ) | ( n5638 & n16746 ) ;
  assign n16748 = x50 | n16747 ;
  assign n16749 = ~x50 & n16747 ;
  assign n16750 = ( ~n16747 & n16748 ) | ( ~n16747 & n16749 ) | ( n16748 & n16749 ) ;
  assign n16751 = n6027 & n8587 ;
  assign n16752 = x125 & n6031 ;
  assign n16753 = x126 | n16752 ;
  assign n16754 = ( n6033 & n16752 ) | ( n6033 & n16753 ) | ( n16752 & n16753 ) ;
  assign n16755 = x124 & n6303 ;
  assign n16756 = n16754 | n16755 ;
  assign n16757 = ( x53 & n16751 ) | ( x53 & ~n16756 ) | ( n16751 & ~n16756 ) ;
  assign n16758 = ( ~x53 & n16756 ) | ( ~x53 & n16757 ) | ( n16756 & n16757 ) ;
  assign n16759 = ( ~n16751 & n16757 ) | ( ~n16751 & n16758 ) | ( n16757 & n16758 ) ;
  assign n16760 = n6713 & n7597 ;
  assign n16761 = x122 & n6717 ;
  assign n16762 = x123 | n16761 ;
  assign n16763 = ( n6719 & n16761 ) | ( n6719 & n16762 ) | ( n16761 & n16762 ) ;
  assign n16764 = x121 & n6980 ;
  assign n16765 = n16763 | n16764 ;
  assign n16766 = ( x56 & n16760 ) | ( x56 & ~n16765 ) | ( n16760 & ~n16765 ) ;
  assign n16767 = ( ~x56 & n16765 ) | ( ~x56 & n16766 ) | ( n16765 & n16766 ) ;
  assign n16768 = ( ~n16760 & n16766 ) | ( ~n16760 & n16767 ) | ( n16766 & n16767 ) ;
  assign n16769 = n7098 & n7423 ;
  assign n16770 = x119 & n7427 ;
  assign n16771 = x120 | n16770 ;
  assign n16772 = ( n7429 & n16770 ) | ( n7429 & n16771 ) | ( n16770 & n16771 ) ;
  assign n16773 = x118 & n7708 ;
  assign n16774 = n16772 | n16773 ;
  assign n16775 = ( x59 & n16769 ) | ( x59 & ~n16774 ) | ( n16769 & ~n16774 ) ;
  assign n16776 = ( ~x59 & n16774 ) | ( ~x59 & n16775 ) | ( n16774 & n16775 ) ;
  assign n16777 = ( ~n16769 & n16775 ) | ( ~n16769 & n16776 ) | ( n16775 & n16776 ) ;
  assign n16778 = n6201 & n8154 ;
  assign n16779 = x116 & n8158 ;
  assign n16780 = x117 | n16779 ;
  assign n16781 = ( n8160 & n16779 ) | ( n8160 & n16780 ) | ( n16779 & n16780 ) ;
  assign n16782 = x115 & n8439 ;
  assign n16783 = n16781 | n16782 ;
  assign n16784 = ( x62 & n16778 ) | ( x62 & ~n16783 ) | ( n16778 & ~n16783 ) ;
  assign n16785 = ( ~x62 & n16783 ) | ( ~x62 & n16784 ) | ( n16783 & n16784 ) ;
  assign n16786 = ( ~n16778 & n16784 ) | ( ~n16778 & n16785 ) | ( n16784 & n16785 ) ;
  assign n16787 = x113 & n8927 ;
  assign n16788 = ( ~x114 & n8693 ) | ( ~x114 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16789 = ( n8693 & n16787 ) | ( n8693 & ~n16788 ) | ( n16787 & ~n16788 ) ;
  assign n16790 = ( ~n16718 & n16786 ) | ( ~n16718 & n16789 ) | ( n16786 & n16789 ) ;
  assign n16791 = ( n16786 & n16789 ) | ( n16786 & ~n16790 ) | ( n16789 & ~n16790 ) ;
  assign n16792 = ( n16718 & n16790 ) | ( n16718 & ~n16791 ) | ( n16790 & ~n16791 ) ;
  assign n16793 = ( n16728 & n16777 ) | ( n16728 & ~n16792 ) | ( n16777 & ~n16792 ) ;
  assign n16794 = ( ~n16728 & n16777 ) | ( ~n16728 & n16792 ) | ( n16777 & n16792 ) ;
  assign n16795 = ( ~n16777 & n16793 ) | ( ~n16777 & n16794 ) | ( n16793 & n16794 ) ;
  assign n16796 = ( n16731 & n16768 ) | ( n16731 & ~n16795 ) | ( n16768 & ~n16795 ) ;
  assign n16797 = ( ~n16731 & n16768 ) | ( ~n16731 & n16795 ) | ( n16768 & n16795 ) ;
  assign n16798 = ( ~n16768 & n16796 ) | ( ~n16768 & n16797 ) | ( n16796 & n16797 ) ;
  assign n16799 = ( n16734 & n16759 ) | ( n16734 & ~n16798 ) | ( n16759 & ~n16798 ) ;
  assign n16800 = ( ~n16734 & n16759 ) | ( ~n16734 & n16798 ) | ( n16759 & n16798 ) ;
  assign n16801 = ( ~n16759 & n16799 ) | ( ~n16759 & n16800 ) | ( n16799 & n16800 ) ;
  assign n16802 = ( n16737 & n16750 ) | ( n16737 & ~n16801 ) | ( n16750 & ~n16801 ) ;
  assign n16803 = ( ~n16737 & n16750 ) | ( ~n16737 & n16801 ) | ( n16750 & n16801 ) ;
  assign n16804 = ( ~n16750 & n16802 ) | ( ~n16750 & n16803 ) | ( n16802 & n16803 ) ;
  assign n16805 = ( ~n16740 & n16743 ) | ( ~n16740 & n16804 ) | ( n16743 & n16804 ) ;
  assign n16806 = ( n16743 & n16804 ) | ( n16743 & ~n16805 ) | ( n16804 & ~n16805 ) ;
  assign n16807 = ( n16740 & n16805 ) | ( n16740 & ~n16806 ) | ( n16805 & ~n16806 ) ;
  assign n16808 = n6027 & n8846 ;
  assign n16809 = x126 & n6031 ;
  assign n16810 = x127 | n16809 ;
  assign n16811 = ( n6033 & n16809 ) | ( n6033 & n16810 ) | ( n16809 & n16810 ) ;
  assign n16812 = x125 & n6303 ;
  assign n16813 = n16811 | n16812 ;
  assign n16814 = ( x53 & n16808 ) | ( x53 & ~n16813 ) | ( n16808 & ~n16813 ) ;
  assign n16815 = ( ~x53 & n16813 ) | ( ~x53 & n16814 ) | ( n16813 & n16814 ) ;
  assign n16816 = ( ~n16808 & n16814 ) | ( ~n16808 & n16815 ) | ( n16814 & n16815 ) ;
  assign n16817 = n6713 & n7841 ;
  assign n16818 = x123 & n6717 ;
  assign n16819 = x124 | n16818 ;
  assign n16820 = ( n6719 & n16818 ) | ( n6719 & n16819 ) | ( n16818 & n16819 ) ;
  assign n16821 = x122 & n6980 ;
  assign n16822 = n16820 | n16821 ;
  assign n16823 = ( x56 & n16817 ) | ( x56 & ~n16822 ) | ( n16817 & ~n16822 ) ;
  assign n16824 = ( ~x56 & n16822 ) | ( ~x56 & n16823 ) | ( n16822 & n16823 ) ;
  assign n16825 = ( ~n16817 & n16823 ) | ( ~n16817 & n16824 ) | ( n16823 & n16824 ) ;
  assign n16826 = n7113 & n7423 ;
  assign n16827 = x120 & n7427 ;
  assign n16828 = x121 | n16827 ;
  assign n16829 = ( n7429 & n16827 ) | ( n7429 & n16828 ) | ( n16827 & n16828 ) ;
  assign n16830 = x119 & n7708 ;
  assign n16831 = n16829 | n16830 ;
  assign n16832 = ( x59 & n16826 ) | ( x59 & ~n16831 ) | ( n16826 & ~n16831 ) ;
  assign n16833 = ( ~x59 & n16831 ) | ( ~x59 & n16832 ) | ( n16831 & n16832 ) ;
  assign n16834 = ( ~n16826 & n16832 ) | ( ~n16826 & n16833 ) | ( n16832 & n16833 ) ;
  assign n16835 = n6421 & n8154 ;
  assign n16836 = x117 & n8158 ;
  assign n16837 = x118 | n16836 ;
  assign n16838 = ( n8160 & n16836 ) | ( n8160 & n16837 ) | ( n16836 & n16837 ) ;
  assign n16839 = x116 & n8439 ;
  assign n16840 = n16838 | n16839 ;
  assign n16841 = ( x62 & n16835 ) | ( x62 & ~n16840 ) | ( n16835 & ~n16840 ) ;
  assign n16842 = ( ~x62 & n16840 ) | ( ~x62 & n16841 ) | ( n16840 & n16841 ) ;
  assign n16843 = ( ~n16835 & n16841 ) | ( ~n16835 & n16842 ) | ( n16841 & n16842 ) ;
  assign n16844 = x114 & n8927 ;
  assign n16845 = ( ~x115 & n8693 ) | ( ~x115 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16846 = ( n8693 & n16844 ) | ( n8693 & ~n16845 ) | ( n16844 & ~n16845 ) ;
  assign n16847 = ( ~x50 & n16718 ) | ( ~x50 & n16846 ) | ( n16718 & n16846 ) ;
  assign n16848 = ( n16718 & n16846 ) | ( n16718 & ~n16847 ) | ( n16846 & ~n16847 ) ;
  assign n16849 = ( x50 & n16847 ) | ( x50 & ~n16848 ) | ( n16847 & ~n16848 ) ;
  assign n16850 = ( n16790 & n16843 ) | ( n16790 & ~n16849 ) | ( n16843 & ~n16849 ) ;
  assign n16851 = ( ~n16790 & n16843 ) | ( ~n16790 & n16849 ) | ( n16843 & n16849 ) ;
  assign n16852 = ( ~n16843 & n16850 ) | ( ~n16843 & n16851 ) | ( n16850 & n16851 ) ;
  assign n16853 = ( n16793 & n16834 ) | ( n16793 & ~n16852 ) | ( n16834 & ~n16852 ) ;
  assign n16854 = ( ~n16793 & n16834 ) | ( ~n16793 & n16852 ) | ( n16834 & n16852 ) ;
  assign n16855 = ( ~n16834 & n16853 ) | ( ~n16834 & n16854 ) | ( n16853 & n16854 ) ;
  assign n16856 = ( n16796 & n16825 ) | ( n16796 & ~n16855 ) | ( n16825 & ~n16855 ) ;
  assign n16857 = ( ~n16796 & n16825 ) | ( ~n16796 & n16855 ) | ( n16825 & n16855 ) ;
  assign n16858 = ( ~n16825 & n16856 ) | ( ~n16825 & n16857 ) | ( n16856 & n16857 ) ;
  assign n16859 = ( n16799 & n16816 ) | ( n16799 & ~n16858 ) | ( n16816 & ~n16858 ) ;
  assign n16860 = ( ~n16799 & n16816 ) | ( ~n16799 & n16858 ) | ( n16816 & n16858 ) ;
  assign n16861 = ( ~n16816 & n16859 ) | ( ~n16816 & n16860 ) | ( n16859 & n16860 ) ;
  assign n16862 = ( ~n16802 & n16805 ) | ( ~n16802 & n16861 ) | ( n16805 & n16861 ) ;
  assign n16863 = ( n16805 & n16861 ) | ( n16805 & ~n16862 ) | ( n16861 & ~n16862 ) ;
  assign n16864 = ( n16802 & n16862 ) | ( n16802 & ~n16863 ) | ( n16862 & ~n16863 ) ;
  assign n16865 = n6027 & n8865 ;
  assign n16866 = x127 & n6031 ;
  assign n16867 = x126 | n16866 ;
  assign n16868 = ( n6303 & n16866 ) | ( n6303 & n16867 ) | ( n16866 & n16867 ) ;
  assign n16869 = ( x53 & n16865 ) | ( x53 & ~n16868 ) | ( n16865 & ~n16868 ) ;
  assign n16870 = ( ~x53 & n16868 ) | ( ~x53 & n16869 ) | ( n16868 & n16869 ) ;
  assign n16871 = ( ~n16865 & n16869 ) | ( ~n16865 & n16870 ) | ( n16869 & n16870 ) ;
  assign n16872 = n6713 & n8331 ;
  assign n16873 = x124 & n6717 ;
  assign n16874 = x125 | n16873 ;
  assign n16875 = ( n6719 & n16873 ) | ( n6719 & n16874 ) | ( n16873 & n16874 ) ;
  assign n16876 = x123 & n6980 ;
  assign n16877 = n16875 | n16876 ;
  assign n16878 = ( x56 & n16872 ) | ( x56 & ~n16877 ) | ( n16872 & ~n16877 ) ;
  assign n16879 = ( ~x56 & n16877 ) | ( ~x56 & n16878 ) | ( n16877 & n16878 ) ;
  assign n16880 = ( ~n16872 & n16878 ) | ( ~n16872 & n16879 ) | ( n16878 & n16879 ) ;
  assign n16881 = n7423 & n7582 ;
  assign n16882 = x121 & n7427 ;
  assign n16883 = x122 | n16882 ;
  assign n16884 = ( n7429 & n16882 ) | ( n7429 & n16883 ) | ( n16882 & n16883 ) ;
  assign n16885 = x120 & n7708 ;
  assign n16886 = n16884 | n16885 ;
  assign n16887 = ( x59 & n16881 ) | ( x59 & ~n16886 ) | ( n16881 & ~n16886 ) ;
  assign n16888 = ( ~x59 & n16886 ) | ( ~x59 & n16887 ) | ( n16886 & n16887 ) ;
  assign n16889 = ( ~n16881 & n16887 ) | ( ~n16881 & n16888 ) | ( n16887 & n16888 ) ;
  assign n16890 = n6645 & n8154 ;
  assign n16891 = x118 & n8158 ;
  assign n16892 = x119 | n16891 ;
  assign n16893 = ( n8160 & n16891 ) | ( n8160 & n16892 ) | ( n16891 & n16892 ) ;
  assign n16894 = x117 & n8439 ;
  assign n16895 = n16893 | n16894 ;
  assign n16896 = ( x62 & n16890 ) | ( x62 & ~n16895 ) | ( n16890 & ~n16895 ) ;
  assign n16897 = ( ~x62 & n16895 ) | ( ~x62 & n16896 ) | ( n16895 & n16896 ) ;
  assign n16898 = ( ~n16890 & n16896 ) | ( ~n16890 & n16897 ) | ( n16896 & n16897 ) ;
  assign n16899 = x115 & n8927 ;
  assign n16900 = ( ~x116 & n8693 ) | ( ~x116 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16901 = ( n8693 & n16899 ) | ( n8693 & ~n16900 ) | ( n16899 & ~n16900 ) ;
  assign n16902 = ( ~n16847 & n16898 ) | ( ~n16847 & n16901 ) | ( n16898 & n16901 ) ;
  assign n16903 = ( n16898 & n16901 ) | ( n16898 & ~n16902 ) | ( n16901 & ~n16902 ) ;
  assign n16904 = ( n16847 & n16902 ) | ( n16847 & ~n16903 ) | ( n16902 & ~n16903 ) ;
  assign n16905 = ( n16850 & n16889 ) | ( n16850 & ~n16904 ) | ( n16889 & ~n16904 ) ;
  assign n16906 = ( ~n16850 & n16889 ) | ( ~n16850 & n16904 ) | ( n16889 & n16904 ) ;
  assign n16907 = ( ~n16889 & n16905 ) | ( ~n16889 & n16906 ) | ( n16905 & n16906 ) ;
  assign n16908 = ( n16853 & n16880 ) | ( n16853 & ~n16907 ) | ( n16880 & ~n16907 ) ;
  assign n16909 = ( ~n16853 & n16880 ) | ( ~n16853 & n16907 ) | ( n16880 & n16907 ) ;
  assign n16910 = ( ~n16880 & n16908 ) | ( ~n16880 & n16909 ) | ( n16908 & n16909 ) ;
  assign n16911 = ( n16856 & n16871 ) | ( n16856 & ~n16910 ) | ( n16871 & ~n16910 ) ;
  assign n16912 = ( ~n16856 & n16871 ) | ( ~n16856 & n16910 ) | ( n16871 & n16910 ) ;
  assign n16913 = ( ~n16871 & n16911 ) | ( ~n16871 & n16912 ) | ( n16911 & n16912 ) ;
  assign n16914 = ( ~n16859 & n16862 ) | ( ~n16859 & n16913 ) | ( n16862 & n16913 ) ;
  assign n16915 = ( n16862 & n16913 ) | ( n16862 & ~n16914 ) | ( n16913 & ~n16914 ) ;
  assign n16916 = ( n16859 & n16914 ) | ( n16859 & ~n16915 ) | ( n16914 & ~n16915 ) ;
  assign n16917 = n6027 & n8862 ;
  assign n16918 = ( x127 & n6303 ) | ( x127 & n16917 ) | ( n6303 & n16917 ) ;
  assign n16919 = x53 | n16918 ;
  assign n16920 = ~x53 & n16918 ;
  assign n16921 = ( ~n16918 & n16919 ) | ( ~n16918 & n16920 ) | ( n16919 & n16920 ) ;
  assign n16922 = n6713 & n8587 ;
  assign n16923 = x125 & n6717 ;
  assign n16924 = x126 | n16923 ;
  assign n16925 = ( n6719 & n16923 ) | ( n6719 & n16924 ) | ( n16923 & n16924 ) ;
  assign n16926 = x124 & n6980 ;
  assign n16927 = n16925 | n16926 ;
  assign n16928 = ( x56 & n16922 ) | ( x56 & ~n16927 ) | ( n16922 & ~n16927 ) ;
  assign n16929 = ( ~x56 & n16927 ) | ( ~x56 & n16928 ) | ( n16927 & n16928 ) ;
  assign n16930 = ( ~n16922 & n16928 ) | ( ~n16922 & n16929 ) | ( n16928 & n16929 ) ;
  assign n16931 = x116 & n8927 ;
  assign n16932 = ( ~x117 & n8693 ) | ( ~x117 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16933 = ( n8693 & n16931 ) | ( n8693 & ~n16932 ) | ( n16931 & ~n16932 ) ;
  assign n16934 = ( n16847 & n16902 ) | ( n16847 & ~n16933 ) | ( n16902 & ~n16933 ) ;
  assign n16935 = ( n16847 & ~n16902 ) | ( n16847 & n16933 ) | ( ~n16902 & n16933 ) ;
  assign n16936 = ( ~n16847 & n16934 ) | ( ~n16847 & n16935 ) | ( n16934 & n16935 ) ;
  assign n16937 = n7423 & n7597 ;
  assign n16938 = x122 & n7427 ;
  assign n16939 = x123 | n16938 ;
  assign n16940 = ( n7429 & n16938 ) | ( n7429 & n16939 ) | ( n16938 & n16939 ) ;
  assign n16941 = x121 & n7708 ;
  assign n16942 = n16940 | n16941 ;
  assign n16943 = ( x59 & n16937 ) | ( x59 & ~n16942 ) | ( n16937 & ~n16942 ) ;
  assign n16944 = ( ~x59 & n16942 ) | ( ~x59 & n16943 ) | ( n16942 & n16943 ) ;
  assign n16945 = ( ~n16937 & n16943 ) | ( ~n16937 & n16944 ) | ( n16943 & n16944 ) ;
  assign n16946 = n7098 & n8154 ;
  assign n16947 = x119 & n8158 ;
  assign n16948 = x120 | n16947 ;
  assign n16949 = ( n8160 & n16947 ) | ( n8160 & n16948 ) | ( n16947 & n16948 ) ;
  assign n16950 = x118 & n8439 ;
  assign n16951 = n16949 | n16950 ;
  assign n16952 = ( x62 & n16946 ) | ( x62 & ~n16951 ) | ( n16946 & ~n16951 ) ;
  assign n16953 = ( ~x62 & n16951 ) | ( ~x62 & n16952 ) | ( n16951 & n16952 ) ;
  assign n16954 = ( ~n16946 & n16952 ) | ( ~n16946 & n16953 ) | ( n16952 & n16953 ) ;
  assign n16955 = ( ~n16936 & n16945 ) | ( ~n16936 & n16954 ) | ( n16945 & n16954 ) ;
  assign n16956 = ( n16945 & n16954 ) | ( n16945 & ~n16955 ) | ( n16954 & ~n16955 ) ;
  assign n16957 = ( n16936 & n16955 ) | ( n16936 & ~n16956 ) | ( n16955 & ~n16956 ) ;
  assign n16958 = ( n16905 & n16930 ) | ( n16905 & ~n16957 ) | ( n16930 & ~n16957 ) ;
  assign n16959 = ( ~n16905 & n16930 ) | ( ~n16905 & n16957 ) | ( n16930 & n16957 ) ;
  assign n16960 = ( ~n16930 & n16958 ) | ( ~n16930 & n16959 ) | ( n16958 & n16959 ) ;
  assign n16961 = ( n16908 & n16921 ) | ( n16908 & ~n16960 ) | ( n16921 & ~n16960 ) ;
  assign n16962 = ( ~n16908 & n16921 ) | ( ~n16908 & n16960 ) | ( n16921 & n16960 ) ;
  assign n16963 = ( ~n16921 & n16961 ) | ( ~n16921 & n16962 ) | ( n16961 & n16962 ) ;
  assign n16964 = ( ~n16911 & n16914 ) | ( ~n16911 & n16963 ) | ( n16914 & n16963 ) ;
  assign n16965 = ( n16914 & n16963 ) | ( n16914 & ~n16964 ) | ( n16963 & ~n16964 ) ;
  assign n16966 = ( n16911 & n16964 ) | ( n16911 & ~n16965 ) | ( n16964 & ~n16965 ) ;
  assign n16967 = n7423 & n7841 ;
  assign n16968 = x123 & n7427 ;
  assign n16969 = x124 | n16968 ;
  assign n16970 = ( n7429 & n16968 ) | ( n7429 & n16969 ) | ( n16968 & n16969 ) ;
  assign n16971 = x122 & n7708 ;
  assign n16972 = n16970 | n16971 ;
  assign n16973 = ( x59 & n16967 ) | ( x59 & ~n16972 ) | ( n16967 & ~n16972 ) ;
  assign n16974 = ( ~x59 & n16972 ) | ( ~x59 & n16973 ) | ( n16972 & n16973 ) ;
  assign n16975 = ( ~n16967 & n16973 ) | ( ~n16967 & n16974 ) | ( n16973 & n16974 ) ;
  assign n16976 = n7113 & n8154 ;
  assign n16977 = x120 & n8158 ;
  assign n16978 = x121 | n16977 ;
  assign n16979 = ( n8160 & n16977 ) | ( n8160 & n16978 ) | ( n16977 & n16978 ) ;
  assign n16980 = x119 & n8439 ;
  assign n16981 = n16979 | n16980 ;
  assign n16982 = ( x62 & n16976 ) | ( x62 & ~n16981 ) | ( n16976 & ~n16981 ) ;
  assign n16983 = ( ~x62 & n16981 ) | ( ~x62 & n16982 ) | ( n16981 & n16982 ) ;
  assign n16984 = ( ~n16976 & n16982 ) | ( ~n16976 & n16983 ) | ( n16982 & n16983 ) ;
  assign n16985 = x117 & n8927 ;
  assign n16986 = ( ~x118 & n8693 ) | ( ~x118 & n8927 ) | ( n8693 & n8927 ) ;
  assign n16987 = ( n8693 & n16985 ) | ( n8693 & ~n16986 ) | ( n16985 & ~n16986 ) ;
  assign n16988 = ( ~x53 & n16933 ) | ( ~x53 & n16987 ) | ( n16933 & n16987 ) ;
  assign n16989 = ( n16933 & n16987 ) | ( n16933 & ~n16988 ) | ( n16987 & ~n16988 ) ;
  assign n16990 = ( x53 & n16988 ) | ( x53 & ~n16989 ) | ( n16988 & ~n16989 ) ;
  assign n16991 = ( n16934 & n16984 ) | ( n16934 & ~n16990 ) | ( n16984 & ~n16990 ) ;
  assign n16992 = ( ~n16934 & n16984 ) | ( ~n16934 & n16990 ) | ( n16984 & n16990 ) ;
  assign n16993 = ( ~n16984 & n16991 ) | ( ~n16984 & n16992 ) | ( n16991 & n16992 ) ;
  assign n16994 = ( n16955 & n16975 ) | ( n16955 & ~n16993 ) | ( n16975 & ~n16993 ) ;
  assign n16995 = ( ~n16955 & n16975 ) | ( ~n16955 & n16993 ) | ( n16975 & n16993 ) ;
  assign n16996 = ( ~n16975 & n16994 ) | ( ~n16975 & n16995 ) | ( n16994 & n16995 ) ;
  assign n16997 = n6713 & n8846 ;
  assign n16998 = x126 & n6717 ;
  assign n16999 = x127 | n16998 ;
  assign n17000 = ( n6719 & n16998 ) | ( n6719 & n16999 ) | ( n16998 & n16999 ) ;
  assign n17001 = x125 & n6980 ;
  assign n17002 = n17000 | n17001 ;
  assign n17003 = ( x56 & n16997 ) | ( x56 & ~n17002 ) | ( n16997 & ~n17002 ) ;
  assign n17004 = ( ~x56 & n17002 ) | ( ~x56 & n17003 ) | ( n17002 & n17003 ) ;
  assign n17005 = ( ~n16997 & n17003 ) | ( ~n16997 & n17004 ) | ( n17003 & n17004 ) ;
  assign n17006 = ( n16958 & ~n16996 ) | ( n16958 & n17005 ) | ( ~n16996 & n17005 ) ;
  assign n17007 = ( n16958 & n16996 ) | ( n16958 & n17005 ) | ( n16996 & n17005 ) ;
  assign n17008 = ( n16996 & n17006 ) | ( n16996 & ~n17007 ) | ( n17006 & ~n17007 ) ;
  assign n17009 = ( ~n16961 & n16964 ) | ( ~n16961 & n17008 ) | ( n16964 & n17008 ) ;
  assign n17010 = ( n16964 & n17008 ) | ( n16964 & ~n17009 ) | ( n17008 & ~n17009 ) ;
  assign n17011 = ( n16961 & n17009 ) | ( n16961 & ~n17010 ) | ( n17009 & ~n17010 ) ;
  assign n17012 = n6713 & n8865 ;
  assign n17013 = x127 & n6717 ;
  assign n17014 = x126 | n17013 ;
  assign n17015 = ( n6980 & n17013 ) | ( n6980 & n17014 ) | ( n17013 & n17014 ) ;
  assign n17016 = ( x56 & n17012 ) | ( x56 & ~n17015 ) | ( n17012 & ~n17015 ) ;
  assign n17017 = ( ~x56 & n17015 ) | ( ~x56 & n17016 ) | ( n17015 & n17016 ) ;
  assign n17018 = ( ~n17012 & n17016 ) | ( ~n17012 & n17017 ) | ( n17016 & n17017 ) ;
  assign n17019 = n7423 & n8331 ;
  assign n17020 = x124 & n7427 ;
  assign n17021 = x125 | n17020 ;
  assign n17022 = ( n7429 & n17020 ) | ( n7429 & n17021 ) | ( n17020 & n17021 ) ;
  assign n17023 = x123 & n7708 ;
  assign n17024 = n17022 | n17023 ;
  assign n17025 = ( x59 & n17019 ) | ( x59 & ~n17024 ) | ( n17019 & ~n17024 ) ;
  assign n17026 = ( ~x59 & n17024 ) | ( ~x59 & n17025 ) | ( n17024 & n17025 ) ;
  assign n17027 = ( ~n17019 & n17025 ) | ( ~n17019 & n17026 ) | ( n17025 & n17026 ) ;
  assign n17028 = x118 & n8927 ;
  assign n17029 = ( ~x119 & n8693 ) | ( ~x119 & n8927 ) | ( n8693 & n8927 ) ;
  assign n17030 = ( n8693 & n17028 ) | ( n8693 & ~n17029 ) | ( n17028 & ~n17029 ) ;
  assign n17031 = n7582 & n8154 ;
  assign n17032 = x121 & n8158 ;
  assign n17033 = x122 | n17032 ;
  assign n17034 = ( n8160 & n17032 ) | ( n8160 & n17033 ) | ( n17032 & n17033 ) ;
  assign n17035 = x120 & n8439 ;
  assign n17036 = n17034 | n17035 ;
  assign n17037 = ( x62 & n17031 ) | ( x62 & ~n17036 ) | ( n17031 & ~n17036 ) ;
  assign n17038 = ( ~x62 & n17036 ) | ( ~x62 & n17037 ) | ( n17036 & n17037 ) ;
  assign n17039 = ( ~n17031 & n17037 ) | ( ~n17031 & n17038 ) | ( n17037 & n17038 ) ;
  assign n17040 = ( n16988 & ~n17030 ) | ( n16988 & n17039 ) | ( ~n17030 & n17039 ) ;
  assign n17041 = ( n16988 & n17030 ) | ( n16988 & n17039 ) | ( n17030 & n17039 ) ;
  assign n17042 = ( n17030 & n17040 ) | ( n17030 & ~n17041 ) | ( n17040 & ~n17041 ) ;
  assign n17043 = ( n16991 & n17027 ) | ( n16991 & ~n17042 ) | ( n17027 & ~n17042 ) ;
  assign n17044 = ( ~n16991 & n17027 ) | ( ~n16991 & n17042 ) | ( n17027 & n17042 ) ;
  assign n17045 = ( ~n17027 & n17043 ) | ( ~n17027 & n17044 ) | ( n17043 & n17044 ) ;
  assign n17046 = ( n16994 & n17018 ) | ( n16994 & ~n17045 ) | ( n17018 & ~n17045 ) ;
  assign n17047 = ( ~n16994 & n17018 ) | ( ~n16994 & n17045 ) | ( n17018 & n17045 ) ;
  assign n17048 = ( ~n17018 & n17046 ) | ( ~n17018 & n17047 ) | ( n17046 & n17047 ) ;
  assign n17049 = ( ~n17006 & n17009 ) | ( ~n17006 & n17048 ) | ( n17009 & n17048 ) ;
  assign n17050 = ( n17009 & n17048 ) | ( n17009 & ~n17049 ) | ( n17048 & ~n17049 ) ;
  assign n17051 = ( n17006 & n17049 ) | ( n17006 & ~n17050 ) | ( n17049 & ~n17050 ) ;
  assign n17052 = n7423 & n8587 ;
  assign n17053 = x125 & n7427 ;
  assign n17054 = x126 | n17053 ;
  assign n17055 = ( n7429 & n17053 ) | ( n7429 & n17054 ) | ( n17053 & n17054 ) ;
  assign n17056 = x124 & n7708 ;
  assign n17057 = n17055 | n17056 ;
  assign n17058 = ( x59 & n17052 ) | ( x59 & ~n17057 ) | ( n17052 & ~n17057 ) ;
  assign n17059 = ( ~x59 & n17057 ) | ( ~x59 & n17058 ) | ( n17057 & n17058 ) ;
  assign n17060 = ( ~n17052 & n17058 ) | ( ~n17052 & n17059 ) | ( n17058 & n17059 ) ;
  assign n17061 = n7597 & n8154 ;
  assign n17062 = x122 & n8158 ;
  assign n17063 = x123 | n17062 ;
  assign n17064 = ( n8160 & n17062 ) | ( n8160 & n17063 ) | ( n17062 & n17063 ) ;
  assign n17065 = x121 & n8439 ;
  assign n17066 = n17064 | n17065 ;
  assign n17067 = ( x62 & n17061 ) | ( x62 & ~n17066 ) | ( n17061 & ~n17066 ) ;
  assign n17068 = ( ~x62 & n17066 ) | ( ~x62 & n17067 ) | ( n17066 & n17067 ) ;
  assign n17069 = ( ~n17061 & n17067 ) | ( ~n17061 & n17068 ) | ( n17067 & n17068 ) ;
  assign n17070 = x119 & n8927 ;
  assign n17071 = ( ~x120 & n8693 ) | ( ~x120 & n8927 ) | ( n8693 & n8927 ) ;
  assign n17072 = ( n8693 & n17070 ) | ( n8693 & ~n17071 ) | ( n17070 & ~n17071 ) ;
  assign n17073 = ( ~n17030 & n17069 ) | ( ~n17030 & n17072 ) | ( n17069 & n17072 ) ;
  assign n17074 = ( n17069 & n17072 ) | ( n17069 & ~n17073 ) | ( n17072 & ~n17073 ) ;
  assign n17075 = ( n17030 & n17073 ) | ( n17030 & ~n17074 ) | ( n17073 & ~n17074 ) ;
  assign n17076 = ( n17040 & n17060 ) | ( n17040 & ~n17075 ) | ( n17060 & ~n17075 ) ;
  assign n17077 = ( ~n17040 & n17060 ) | ( ~n17040 & n17075 ) | ( n17060 & n17075 ) ;
  assign n17078 = ( ~n17060 & n17076 ) | ( ~n17060 & n17077 ) | ( n17076 & n17077 ) ;
  assign n17079 = n6713 & n8862 ;
  assign n17080 = ( x127 & n6980 ) | ( x127 & n17079 ) | ( n6980 & n17079 ) ;
  assign n17081 = x56 | n17080 ;
  assign n17082 = ~x56 & n17080 ;
  assign n17083 = ( ~n17080 & n17081 ) | ( ~n17080 & n17082 ) | ( n17081 & n17082 ) ;
  assign n17084 = ( n17043 & ~n17078 ) | ( n17043 & n17083 ) | ( ~n17078 & n17083 ) ;
  assign n17085 = ( n17043 & n17078 ) | ( n17043 & n17083 ) | ( n17078 & n17083 ) ;
  assign n17086 = ( n17078 & n17084 ) | ( n17078 & ~n17085 ) | ( n17084 & ~n17085 ) ;
  assign n17087 = ( ~n17046 & n17049 ) | ( ~n17046 & n17086 ) | ( n17049 & n17086 ) ;
  assign n17088 = ( n17049 & n17086 ) | ( n17049 & ~n17087 ) | ( n17086 & ~n17087 ) ;
  assign n17089 = ( n17046 & n17087 ) | ( n17046 & ~n17088 ) | ( n17087 & ~n17088 ) ;
  assign n17090 = n7841 & n8154 ;
  assign n17091 = x123 & n8158 ;
  assign n17092 = x124 | n17091 ;
  assign n17093 = ( n8160 & n17091 ) | ( n8160 & n17092 ) | ( n17091 & n17092 ) ;
  assign n17094 = x122 & n8439 ;
  assign n17095 = n17093 | n17094 ;
  assign n17096 = ( x62 & n17090 ) | ( x62 & ~n17095 ) | ( n17090 & ~n17095 ) ;
  assign n17097 = ( ~x62 & n17095 ) | ( ~x62 & n17096 ) | ( n17095 & n17096 ) ;
  assign n17098 = ( ~n17090 & n17096 ) | ( ~n17090 & n17097 ) | ( n17096 & n17097 ) ;
  assign n17099 = x120 & n8927 ;
  assign n17100 = ( ~x121 & n8693 ) | ( ~x121 & n8927 ) | ( n8693 & n8927 ) ;
  assign n17101 = ( n8693 & n17099 ) | ( n8693 & ~n17100 ) | ( n17099 & ~n17100 ) ;
  assign n17102 = ( ~x56 & n17030 ) | ( ~x56 & n17101 ) | ( n17030 & n17101 ) ;
  assign n17103 = ( n17030 & n17101 ) | ( n17030 & ~n17102 ) | ( n17101 & ~n17102 ) ;
  assign n17104 = ( x56 & n17102 ) | ( x56 & ~n17103 ) | ( n17102 & ~n17103 ) ;
  assign n17105 = ( n17073 & n17098 ) | ( n17073 & ~n17104 ) | ( n17098 & ~n17104 ) ;
  assign n17106 = ( ~n17073 & n17098 ) | ( ~n17073 & n17104 ) | ( n17098 & n17104 ) ;
  assign n17107 = ( ~n17098 & n17105 ) | ( ~n17098 & n17106 ) | ( n17105 & n17106 ) ;
  assign n17108 = n7423 & n8846 ;
  assign n17109 = x126 & n7427 ;
  assign n17110 = x127 | n17109 ;
  assign n17111 = ( n7429 & n17109 ) | ( n7429 & n17110 ) | ( n17109 & n17110 ) ;
  assign n17112 = x125 & n7708 ;
  assign n17113 = n17111 | n17112 ;
  assign n17114 = ( x59 & n17108 ) | ( x59 & ~n17113 ) | ( n17108 & ~n17113 ) ;
  assign n17115 = ( ~x59 & n17113 ) | ( ~x59 & n17114 ) | ( n17113 & n17114 ) ;
  assign n17116 = ( ~n17108 & n17114 ) | ( ~n17108 & n17115 ) | ( n17114 & n17115 ) ;
  assign n17117 = ( n17076 & ~n17107 ) | ( n17076 & n17116 ) | ( ~n17107 & n17116 ) ;
  assign n17118 = ( n17076 & n17107 ) | ( n17076 & n17116 ) | ( n17107 & n17116 ) ;
  assign n17119 = ( n17107 & n17117 ) | ( n17107 & ~n17118 ) | ( n17117 & ~n17118 ) ;
  assign n17120 = ( ~n17084 & n17087 ) | ( ~n17084 & n17119 ) | ( n17087 & n17119 ) ;
  assign n17121 = ( n17087 & n17119 ) | ( n17087 & ~n17120 ) | ( n17119 & ~n17120 ) ;
  assign n17122 = ( n17084 & n17120 ) | ( n17084 & ~n17121 ) | ( n17120 & ~n17121 ) ;
  assign n17123 = n7423 & n8865 ;
  assign n17124 = x127 & n7427 ;
  assign n17125 = x126 | n17124 ;
  assign n17126 = ( n7708 & n17124 ) | ( n7708 & n17125 ) | ( n17124 & n17125 ) ;
  assign n17127 = ( x59 & n17123 ) | ( x59 & ~n17126 ) | ( n17123 & ~n17126 ) ;
  assign n17128 = ( ~x59 & n17126 ) | ( ~x59 & n17127 ) | ( n17126 & n17127 ) ;
  assign n17129 = ( ~n17123 & n17127 ) | ( ~n17123 & n17128 ) | ( n17127 & n17128 ) ;
  assign n17130 = n8154 & n8331 ;
  assign n17131 = x124 & n8158 ;
  assign n17132 = x125 | n17131 ;
  assign n17133 = ( n8160 & n17131 ) | ( n8160 & n17132 ) | ( n17131 & n17132 ) ;
  assign n17134 = x123 & n8439 ;
  assign n17135 = n17133 | n17134 ;
  assign n17136 = ( x62 & n17130 ) | ( x62 & ~n17135 ) | ( n17130 & ~n17135 ) ;
  assign n17137 = ( ~x62 & n17135 ) | ( ~x62 & n17136 ) | ( n17135 & n17136 ) ;
  assign n17138 = ( ~n17130 & n17136 ) | ( ~n17130 & n17137 ) | ( n17136 & n17137 ) ;
  assign n17139 = x121 & n8927 ;
  assign n17140 = ( ~x122 & n8693 ) | ( ~x122 & n8927 ) | ( n8693 & n8927 ) ;
  assign n17141 = ( n8693 & n17139 ) | ( n8693 & ~n17140 ) | ( n17139 & ~n17140 ) ;
  assign n17142 = ( ~n17102 & n17138 ) | ( ~n17102 & n17141 ) | ( n17138 & n17141 ) ;
  assign n17143 = ( n17138 & n17141 ) | ( n17138 & ~n17142 ) | ( n17141 & ~n17142 ) ;
  assign n17144 = ( n17102 & n17142 ) | ( n17102 & ~n17143 ) | ( n17142 & ~n17143 ) ;
  assign n17145 = ( n17105 & n17129 ) | ( n17105 & ~n17144 ) | ( n17129 & ~n17144 ) ;
  assign n17146 = ( ~n17105 & n17129 ) | ( ~n17105 & n17144 ) | ( n17129 & n17144 ) ;
  assign n17147 = ( ~n17129 & n17145 ) | ( ~n17129 & n17146 ) | ( n17145 & n17146 ) ;
  assign n17148 = ( ~n17117 & n17120 ) | ( ~n17117 & n17147 ) | ( n17120 & n17147 ) ;
  assign n17149 = ( n17120 & n17147 ) | ( n17120 & ~n17148 ) | ( n17147 & ~n17148 ) ;
  assign n17150 = ( n17117 & n17148 ) | ( n17117 & ~n17149 ) | ( n17148 & ~n17149 ) ;
  assign n17151 = x122 & n8927 ;
  assign n17152 = ( ~x123 & n8693 ) | ( ~x123 & n8927 ) | ( n8693 & n8927 ) ;
  assign n17153 = ( n8693 & n17151 ) | ( n8693 & ~n17152 ) | ( n17151 & ~n17152 ) ;
  assign n17154 = ( n17102 & n17142 ) | ( n17102 & ~n17153 ) | ( n17142 & ~n17153 ) ;
  assign n17155 = ( n17102 & ~n17142 ) | ( n17102 & n17153 ) | ( ~n17142 & n17153 ) ;
  assign n17156 = ( ~n17102 & n17154 ) | ( ~n17102 & n17155 ) | ( n17154 & n17155 ) ;
  assign n17157 = n8154 & n8587 ;
  assign n17158 = x125 & n8158 ;
  assign n17159 = x126 | n17158 ;
  assign n17160 = ( n8160 & n17158 ) | ( n8160 & n17159 ) | ( n17158 & n17159 ) ;
  assign n17161 = x124 & n8439 ;
  assign n17162 = n17160 | n17161 ;
  assign n17163 = ( x62 & n17157 ) | ( x62 & ~n17162 ) | ( n17157 & ~n17162 ) ;
  assign n17164 = ( ~x62 & n17162 ) | ( ~x62 & n17163 ) | ( n17162 & n17163 ) ;
  assign n17165 = ( ~n17157 & n17163 ) | ( ~n17157 & n17164 ) | ( n17163 & n17164 ) ;
  assign n17166 = n7423 & n8862 ;
  assign n17167 = ( x127 & n7708 ) | ( x127 & n17166 ) | ( n7708 & n17166 ) ;
  assign n17168 = x59 | n17167 ;
  assign n17169 = ~x59 & n17167 ;
  assign n17170 = ( ~n17167 & n17168 ) | ( ~n17167 & n17169 ) | ( n17168 & n17169 ) ;
  assign n17171 = ( ~n17156 & n17165 ) | ( ~n17156 & n17170 ) | ( n17165 & n17170 ) ;
  assign n17172 = ( n17165 & n17170 ) | ( n17165 & ~n17171 ) | ( n17170 & ~n17171 ) ;
  assign n17173 = ( n17156 & n17171 ) | ( n17156 & ~n17172 ) | ( n17171 & ~n17172 ) ;
  assign n17174 = ( ~n17145 & n17148 ) | ( ~n17145 & n17173 ) | ( n17148 & n17173 ) ;
  assign n17175 = ( n17148 & n17173 ) | ( n17148 & ~n17174 ) | ( n17173 & ~n17174 ) ;
  assign n17176 = ( n17145 & n17174 ) | ( n17145 & ~n17175 ) | ( n17174 & ~n17175 ) ;
  assign n17177 = n8154 & n8846 ;
  assign n17178 = x126 & n8158 ;
  assign n17179 = x127 | n17178 ;
  assign n17180 = ( n8160 & n17178 ) | ( n8160 & n17179 ) | ( n17178 & n17179 ) ;
  assign n17181 = x125 & n8439 ;
  assign n17182 = n17180 | n17181 ;
  assign n17183 = ( x62 & n17177 ) | ( x62 & ~n17182 ) | ( n17177 & ~n17182 ) ;
  assign n17184 = ( ~x62 & n17182 ) | ( ~x62 & n17183 ) | ( n17182 & n17183 ) ;
  assign n17185 = ( ~n17177 & n17183 ) | ( ~n17177 & n17184 ) | ( n17183 & n17184 ) ;
  assign n17186 = x123 & n8927 ;
  assign n17187 = ( ~x124 & n8693 ) | ( ~x124 & n8927 ) | ( n8693 & n8927 ) ;
  assign n17188 = ( n8693 & n17186 ) | ( n8693 & ~n17187 ) | ( n17186 & ~n17187 ) ;
  assign n17189 = ( ~x59 & n17153 ) | ( ~x59 & n17188 ) | ( n17153 & n17188 ) ;
  assign n17190 = ( n17153 & n17188 ) | ( n17153 & ~n17189 ) | ( n17188 & ~n17189 ) ;
  assign n17191 = ( x59 & n17189 ) | ( x59 & ~n17190 ) | ( n17189 & ~n17190 ) ;
  assign n17192 = ( n17154 & n17185 ) | ( n17154 & ~n17191 ) | ( n17185 & ~n17191 ) ;
  assign n17193 = ( ~n17154 & n17185 ) | ( ~n17154 & n17191 ) | ( n17185 & n17191 ) ;
  assign n17194 = ( ~n17185 & n17192 ) | ( ~n17185 & n17193 ) | ( n17192 & n17193 ) ;
  assign n17195 = ( ~n17171 & n17174 ) | ( ~n17171 & n17194 ) | ( n17174 & n17194 ) ;
  assign n17196 = ( n17174 & n17194 ) | ( n17174 & ~n17195 ) | ( n17194 & ~n17195 ) ;
  assign n17197 = ( n17171 & n17195 ) | ( n17171 & ~n17196 ) | ( n17195 & ~n17196 ) ;
  assign n17198 = x124 & n8927 ;
  assign n17199 = ( ~x125 & n8693 ) | ( ~x125 & n8927 ) | ( n8693 & n8927 ) ;
  assign n17200 = ( n8693 & n17198 ) | ( n8693 & ~n17199 ) | ( n17198 & ~n17199 ) ;
  assign n17201 = n8154 & n8865 ;
  assign n17202 = x127 & n8158 ;
  assign n17203 = x126 | n17202 ;
  assign n17204 = ( n8439 & n17202 ) | ( n8439 & n17203 ) | ( n17202 & n17203 ) ;
  assign n17205 = ( x62 & n17201 ) | ( x62 & ~n17204 ) | ( n17201 & ~n17204 ) ;
  assign n17206 = ( ~x62 & n17204 ) | ( ~x62 & n17205 ) | ( n17204 & n17205 ) ;
  assign n17207 = ( ~n17201 & n17205 ) | ( ~n17201 & n17206 ) | ( n17205 & n17206 ) ;
  assign n17208 = ( n17189 & ~n17200 ) | ( n17189 & n17207 ) | ( ~n17200 & n17207 ) ;
  assign n17209 = ( n17189 & n17200 ) | ( n17189 & n17207 ) | ( n17200 & n17207 ) ;
  assign n17210 = ( n17200 & n17208 ) | ( n17200 & ~n17209 ) | ( n17208 & ~n17209 ) ;
  assign n17211 = ( ~n17192 & n17195 ) | ( ~n17192 & n17210 ) | ( n17195 & n17210 ) ;
  assign n17212 = ( n17195 & n17210 ) | ( n17195 & ~n17211 ) | ( n17210 & ~n17211 ) ;
  assign n17213 = ( n17192 & n17211 ) | ( n17192 & ~n17212 ) | ( n17211 & ~n17212 ) ;
  assign n17214 = x125 & n8927 ;
  assign n17215 = ( ~x126 & n8693 ) | ( ~x126 & n8927 ) | ( n8693 & n8927 ) ;
  assign n17216 = ( n8693 & n17214 ) | ( n8693 & ~n17215 ) | ( n17214 & ~n17215 ) ;
  assign n17217 = n8154 & n8862 ;
  assign n17218 = ( x127 & n8439 ) | ( x127 & n17217 ) | ( n8439 & n17217 ) ;
  assign n17219 = x62 | n17218 ;
  assign n17220 = ~x62 & n17218 ;
  assign n17221 = ( ~n17218 & n17219 ) | ( ~n17218 & n17220 ) | ( n17219 & n17220 ) ;
  assign n17222 = ( ~n17200 & n17216 ) | ( ~n17200 & n17221 ) | ( n17216 & n17221 ) ;
  assign n17223 = ( n17216 & n17221 ) | ( n17216 & ~n17222 ) | ( n17221 & ~n17222 ) ;
  assign n17224 = ( n17200 & n17222 ) | ( n17200 & ~n17223 ) | ( n17222 & ~n17223 ) ;
  assign n17225 = ( ~n17208 & n17211 ) | ( ~n17208 & n17224 ) | ( n17211 & n17224 ) ;
  assign n17226 = ( n17211 & n17224 ) | ( n17211 & ~n17225 ) | ( n17224 & ~n17225 ) ;
  assign n17227 = ( n17208 & n17225 ) | ( n17208 & ~n17226 ) | ( n17225 & ~n17226 ) ;
  assign n17228 = x63 & x127 ;
  assign n17229 = x62 & ~x127 ;
  assign n17230 = x126 & n8927 ;
  assign n17231 = ( n17228 & n17229 ) | ( n17228 & ~n17230 ) | ( n17229 & ~n17230 ) ;
  assign n17232 = n17200 & ~n17231 ;
  assign n17233 = ~n17200 & n17231 ;
  assign n17234 = n17232 | n17233 ;
  assign n17235 = ( ~n17222 & n17225 ) | ( ~n17222 & n17234 ) | ( n17225 & n17234 ) ;
  assign n17236 = ( n17225 & n17234 ) | ( n17225 & ~n17235 ) | ( n17234 & ~n17235 ) ;
  assign n17237 = ( n17222 & n17235 ) | ( n17222 & ~n17236 ) | ( n17235 & ~n17236 ) ;
  assign n17238 = ( ~n17228 & n17232 ) | ( ~n17228 & n17235 ) | ( n17232 & n17235 ) ;
  assign n17239 = ( n17232 & n17235 ) | ( n17232 & ~n17238 ) | ( n17235 & ~n17238 ) ;
  assign n17240 = ( n17228 & n17238 ) | ( n17228 & ~n17239 ) | ( n17238 & ~n17239 ) ;
  assign y0 = n129 ;
  assign y1 = n146 ;
  assign y2 = n160 ;
  assign y3 = n181 ;
  assign y4 = n213 ;
  assign y5 = n242 ;
  assign y6 = n274 ;
  assign y7 = n318 ;
  assign y8 = n358 ;
  assign y9 = n402 ;
  assign y10 = n458 ;
  assign y11 = n510 ;
  assign y12 = n566 ;
  assign y13 = n634 ;
  assign y14 = n698 ;
  assign y15 = n766 ;
  assign y16 = n846 ;
  assign y17 = n922 ;
  assign y18 = n1002 ;
  assign y19 = n1094 ;
  assign y20 = n1182 ;
  assign y21 = n1274 ;
  assign y22 = n1378 ;
  assign y23 = n1478 ;
  assign y24 = n1582 ;
  assign y25 = n1698 ;
  assign y26 = n1810 ;
  assign y27 = n1926 ;
  assign y28 = n2054 ;
  assign y29 = n2178 ;
  assign y30 = n2306 ;
  assign y31 = n2446 ;
  assign y32 = n2582 ;
  assign y33 = n2722 ;
  assign y34 = n2874 ;
  assign y35 = n3022 ;
  assign y36 = n3174 ;
  assign y37 = n3338 ;
  assign y38 = n3498 ;
  assign y39 = n3662 ;
  assign y40 = n3838 ;
  assign y41 = n4010 ;
  assign y42 = n4186 ;
  assign y43 = n4374 ;
  assign y44 = n4558 ;
  assign y45 = n4746 ;
  assign y46 = n4946 ;
  assign y47 = n5142 ;
  assign y48 = n5342 ;
  assign y49 = n5554 ;
  assign y50 = n5762 ;
  assign y51 = n5974 ;
  assign y52 = n6198 ;
  assign y53 = n6418 ;
  assign y54 = n6642 ;
  assign y55 = n6878 ;
  assign y56 = n7110 ;
  assign y57 = n7346 ;
  assign y58 = n7594 ;
  assign y59 = n7838 ;
  assign y60 = n8086 ;
  assign y61 = n8346 ;
  assign y62 = n8602 ;
  assign y63 = n8861 ;
  assign y64 = n9118 ;
  assign y65 = n9370 ;
  assign y66 = n9616 ;
  assign y67 = n9860 ;
  assign y68 = n10102 ;
  assign y69 = n10339 ;
  assign y70 = n10571 ;
  assign y71 = n10801 ;
  assign y72 = n11026 ;
  assign y73 = n11246 ;
  assign y74 = n11464 ;
  assign y75 = n11677 ;
  assign y76 = n11885 ;
  assign y77 = n12091 ;
  assign y78 = n12292 ;
  assign y79 = n12488 ;
  assign y80 = n12682 ;
  assign y81 = n12871 ;
  assign y82 = n13055 ;
  assign y83 = n13237 ;
  assign y84 = n13414 ;
  assign y85 = n13586 ;
  assign y86 = n13756 ;
  assign y87 = n13921 ;
  assign y88 = n14081 ;
  assign y89 = n14239 ;
  assign y90 = n14392 ;
  assign y91 = n14540 ;
  assign y92 = n14686 ;
  assign y93 = n14827 ;
  assign y94 = n14963 ;
  assign y95 = n15097 ;
  assign y96 = n15226 ;
  assign y97 = n15350 ;
  assign y98 = n15472 ;
  assign y99 = n15589 ;
  assign y100 = n15701 ;
  assign y101 = n15811 ;
  assign y102 = n15916 ;
  assign y103 = n16016 ;
  assign y104 = n16114 ;
  assign y105 = n16207 ;
  assign y106 = n16295 ;
  assign y107 = n16381 ;
  assign y108 = n16462 ;
  assign y109 = n16538 ;
  assign y110 = n16612 ;
  assign y111 = n16681 ;
  assign y112 = n16745 ;
  assign y113 = n16807 ;
  assign y114 = n16864 ;
  assign y115 = n16916 ;
  assign y116 = n16966 ;
  assign y117 = n17011 ;
  assign y118 = n17051 ;
  assign y119 = n17089 ;
  assign y120 = n17122 ;
  assign y121 = n17150 ;
  assign y122 = n17176 ;
  assign y123 = n17197 ;
  assign y124 = n17213 ;
  assign y125 = n17227 ;
  assign y126 = n17237 ;
  assign y127 = n17240 ;
endmodule
