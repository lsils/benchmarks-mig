module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 ;
  assign n129 = x124 | x125 ;
  assign n130 = x126 | n129 ;
  assign n131 = x126 | x127 ;
  assign n132 = ( x127 & n130 ) | ( x127 & ~n131 ) | ( n130 & ~n131 ) ;
  assign n133 = x126 & x127 ;
  assign n134 = x125 & ~x127 ;
  assign n135 = n133 | n134 ;
  assign n136 = ~x126 & x127 ;
  assign n137 = x122 | x123 ;
  assign n138 = n136 | n137 ;
  assign n139 = x125 & x127 ;
  assign n140 = x124 | n139 ;
  assign n141 = n138 | n140 ;
  assign n142 = ( ~n130 & n135 ) | ( ~n130 & n141 ) | ( n135 & n141 ) ;
  assign n143 = ~x126 & n139 ;
  assign n144 = x125 | x127 ;
  assign n145 = ~n137 & n144 ;
  assign n146 = ~n143 & n145 ;
  assign n147 = ( ~x124 & n143 ) | ( ~x124 & n146 ) | ( n143 & n146 ) ;
  assign n148 = n139 & ~n147 ;
  assign n149 = ( n136 & ~n137 ) | ( n136 & n144 ) | ( ~n137 & n144 ) ;
  assign n150 = ( x126 & n137 ) | ( x126 & ~n140 ) | ( n137 & ~n140 ) ;
  assign n151 = ( n148 & n149 ) | ( n148 & n150 ) | ( n149 & n150 ) ;
  assign n152 = ~x126 & n134 ;
  assign n153 = x120 | x121 ;
  assign n154 = ~n132 & n153 ;
  assign n155 = ( x122 & ~n152 ) | ( x122 & n154 ) | ( ~n152 & n154 ) ;
  assign n156 = x123 & n129 ;
  assign n157 = ~n135 & n156 ;
  assign n158 = n132 & ~n153 ;
  assign n159 = ( n146 & n157 ) | ( n146 & ~n158 ) | ( n157 & ~n158 ) ;
  assign n160 = x122 & n133 ;
  assign n161 = ~x125 & x126 ;
  assign n162 = x123 | n161 ;
  assign n163 = ( x122 & n160 ) | ( x122 & ~n162 ) | ( n160 & ~n162 ) ;
  assign n164 = ( n155 & n159 ) | ( n155 & ~n163 ) | ( n159 & ~n163 ) ;
  assign n165 = x126 | n134 ;
  assign n166 = x124 & ~n145 ;
  assign n167 = n165 & n166 ;
  assign n168 = n147 | n167 ;
  assign n169 = ( ~n131 & n164 ) | ( ~n131 & n168 ) | ( n164 & n168 ) ;
  assign n170 = n151 | n169 ;
  assign n171 = ( n131 & n147 ) | ( n131 & n167 ) | ( n147 & n167 ) ;
  assign n172 = ~n164 & n171 ;
  assign n173 = ~n151 & n164 ;
  assign n174 = ( n164 & n172 ) | ( n164 & ~n173 ) | ( n172 & ~n173 ) ;
  assign n175 = x118 | x119 ;
  assign n176 = x120 | n175 ;
  assign n177 = ~n142 & n176 ;
  assign n178 = n153 & n170 ;
  assign n179 = ( x121 & n170 ) | ( x121 & ~n177 ) | ( n170 & ~n177 ) ;
  assign n180 = n142 & ~n176 ;
  assign n181 = n179 & ~n180 ;
  assign n182 = ( n177 & ~n178 ) | ( n177 & n181 ) | ( ~n178 & n181 ) ;
  assign n183 = n142 | n170 ;
  assign n184 = ( ~x122 & n178 ) | ( ~x122 & n183 ) | ( n178 & n183 ) ;
  assign n185 = ( x122 & n178 ) | ( x122 & n183 ) | ( n178 & n183 ) ;
  assign n186 = ( x122 & n184 ) | ( x122 & ~n185 ) | ( n184 & ~n185 ) ;
  assign n187 = ( ~n132 & n182 ) | ( ~n132 & n186 ) | ( n182 & n186 ) ;
  assign n188 = ~x122 & n142 ;
  assign n189 = ( ~x122 & n154 ) | ( ~x122 & n158 ) | ( n154 & n158 ) ;
  assign n190 = ( ~x122 & x126 ) | ( ~x122 & n134 ) | ( x126 & n134 ) ;
  assign n191 = ( n165 & n189 ) | ( n165 & ~n190 ) | ( n189 & ~n190 ) ;
  assign n192 = n170 & ~n191 ;
  assign n193 = ( ~x123 & n188 ) | ( ~x123 & n192 ) | ( n188 & n192 ) ;
  assign n194 = ( x123 & n188 ) | ( x123 & n192 ) | ( n188 & n192 ) ;
  assign n195 = ( x123 & n193 ) | ( x123 & ~n194 ) | ( n193 & ~n194 ) ;
  assign n196 = ( ~n131 & n187 ) | ( ~n131 & n195 ) | ( n187 & n195 ) ;
  assign n197 = n174 | n196 ;
  assign n198 = ( n132 & ~n182 ) | ( n132 & n197 ) | ( ~n182 & n197 ) ;
  assign n199 = n132 & ~n182 ;
  assign n200 = ( n186 & ~n198 ) | ( n186 & n199 ) | ( ~n198 & n199 ) ;
  assign n201 = ( n186 & n198 ) | ( n186 & n199 ) | ( n198 & n199 ) ;
  assign n202 = ( n198 & n200 ) | ( n198 & ~n201 ) | ( n200 & ~n201 ) ;
  assign n203 = ~n175 & n197 ;
  assign n204 = x116 | x117 ;
  assign n205 = x118 | n204 ;
  assign n206 = n170 & ~n205 ;
  assign n207 = ~n170 & n205 ;
  assign n208 = ( x119 & ~n197 ) | ( x119 & n207 ) | ( ~n197 & n207 ) ;
  assign n209 = ( n203 & ~n206 ) | ( n203 & n208 ) | ( ~n206 & n208 ) ;
  assign n210 = n170 & ~n197 ;
  assign n211 = ( x120 & n203 ) | ( x120 & n210 ) | ( n203 & n210 ) ;
  assign n212 = ( ~x120 & n203 ) | ( ~x120 & n210 ) | ( n203 & n210 ) ;
  assign n213 = ( x120 & ~n211 ) | ( x120 & n212 ) | ( ~n211 & n212 ) ;
  assign n214 = ( ~n142 & n209 ) | ( ~n142 & n213 ) | ( n209 & n213 ) ;
  assign n215 = ( n142 & n170 ) | ( n142 & ~n197 ) | ( n170 & ~n197 ) ;
  assign n216 = n183 & ~n215 ;
  assign n217 = ( ~x121 & n212 ) | ( ~x121 & n216 ) | ( n212 & n216 ) ;
  assign n218 = ( x121 & n212 ) | ( x121 & n216 ) | ( n212 & n216 ) ;
  assign n219 = ( x121 & n217 ) | ( x121 & ~n218 ) | ( n217 & ~n218 ) ;
  assign n220 = ( ~n132 & n214 ) | ( ~n132 & n219 ) | ( n214 & n219 ) ;
  assign n221 = ( ~n131 & n202 ) | ( ~n131 & n220 ) | ( n202 & n220 ) ;
  assign n222 = n174 & ~n195 ;
  assign n223 = n187 & n222 ;
  assign n224 = ( n195 & ~n196 ) | ( n195 & n223 ) | ( ~n196 & n223 ) ;
  assign n225 = n221 | n224 ;
  assign n226 = n220 & n224 ;
  assign n227 = ( n202 & ~n221 ) | ( n202 & n226 ) | ( ~n221 & n226 ) ;
  assign n228 = ( n132 & ~n214 ) | ( n132 & n225 ) | ( ~n214 & n225 ) ;
  assign n229 = n132 & ~n214 ;
  assign n230 = ( n219 & n228 ) | ( n219 & n229 ) | ( n228 & n229 ) ;
  assign n231 = ( n219 & ~n228 ) | ( n219 & n229 ) | ( ~n228 & n229 ) ;
  assign n232 = ( n228 & ~n230 ) | ( n228 & n231 ) | ( ~n230 & n231 ) ;
  assign n233 = ~n204 & n225 ;
  assign n234 = x114 | x115 ;
  assign n235 = x116 | n234 ;
  assign n236 = n197 & ~n235 ;
  assign n237 = ~n197 & n235 ;
  assign n238 = ( x117 & ~n225 ) | ( x117 & n237 ) | ( ~n225 & n237 ) ;
  assign n239 = ( n233 & ~n236 ) | ( n233 & n238 ) | ( ~n236 & n238 ) ;
  assign n240 = n197 & ~n225 ;
  assign n241 = ( x118 & n233 ) | ( x118 & n240 ) | ( n233 & n240 ) ;
  assign n242 = ( ~x118 & n233 ) | ( ~x118 & n240 ) | ( n233 & n240 ) ;
  assign n243 = ( x118 & ~n241 ) | ( x118 & n242 ) | ( ~n241 & n242 ) ;
  assign n244 = ( ~n170 & n239 ) | ( ~n170 & n243 ) | ( n239 & n243 ) ;
  assign n245 = ~n170 & n197 ;
  assign n246 = ( n210 & n225 ) | ( n210 & n245 ) | ( n225 & n245 ) ;
  assign n247 = ( x119 & n242 ) | ( x119 & n246 ) | ( n242 & n246 ) ;
  assign n248 = ( ~x119 & n242 ) | ( ~x119 & n246 ) | ( n242 & n246 ) ;
  assign n249 = ( x119 & ~n247 ) | ( x119 & n248 ) | ( ~n247 & n248 ) ;
  assign n250 = ( ~n142 & n244 ) | ( ~n142 & n249 ) | ( n244 & n249 ) ;
  assign n251 = n142 & ~n209 ;
  assign n252 = ( n142 & ~n209 ) | ( n142 & n225 ) | ( ~n209 & n225 ) ;
  assign n253 = ( ~n213 & n251 ) | ( ~n213 & n252 ) | ( n251 & n252 ) ;
  assign n254 = ( n213 & n251 ) | ( n213 & n252 ) | ( n251 & n252 ) ;
  assign n255 = ( n213 & n253 ) | ( n213 & ~n254 ) | ( n253 & ~n254 ) ;
  assign n256 = ( ~n132 & n250 ) | ( ~n132 & n255 ) | ( n250 & n255 ) ;
  assign n257 = ( ~n131 & n232 ) | ( ~n131 & n256 ) | ( n232 & n256 ) ;
  assign n258 = n227 | n257 ;
  assign n259 = ( n132 & ~n250 ) | ( n132 & n258 ) | ( ~n250 & n258 ) ;
  assign n260 = n132 & ~n250 ;
  assign n261 = ( n255 & ~n259 ) | ( n255 & n260 ) | ( ~n259 & n260 ) ;
  assign n262 = ( n255 & n259 ) | ( n255 & n260 ) | ( n259 & n260 ) ;
  assign n263 = ( n259 & n261 ) | ( n259 & ~n262 ) | ( n261 & ~n262 ) ;
  assign n264 = ~n234 & n258 ;
  assign n265 = x112 | x113 ;
  assign n266 = x114 | n265 ;
  assign n267 = n225 & ~n266 ;
  assign n268 = ~n225 & n266 ;
  assign n269 = ( x115 & ~n258 ) | ( x115 & n268 ) | ( ~n258 & n268 ) ;
  assign n270 = ( n264 & ~n267 ) | ( n264 & n269 ) | ( ~n267 & n269 ) ;
  assign n271 = n225 & ~n258 ;
  assign n272 = ( x116 & n264 ) | ( x116 & n271 ) | ( n264 & n271 ) ;
  assign n273 = ( ~x116 & n264 ) | ( ~x116 & n271 ) | ( n264 & n271 ) ;
  assign n274 = ( x116 & ~n272 ) | ( x116 & n273 ) | ( ~n272 & n273 ) ;
  assign n275 = ( ~n197 & n270 ) | ( ~n197 & n274 ) | ( n270 & n274 ) ;
  assign n276 = ~n197 & n225 ;
  assign n277 = ( n240 & n258 ) | ( n240 & n276 ) | ( n258 & n276 ) ;
  assign n278 = ( x117 & n273 ) | ( x117 & n277 ) | ( n273 & n277 ) ;
  assign n279 = ( ~x117 & n273 ) | ( ~x117 & n277 ) | ( n273 & n277 ) ;
  assign n280 = ( x117 & ~n278 ) | ( x117 & n279 ) | ( ~n278 & n279 ) ;
  assign n281 = ( ~n170 & n275 ) | ( ~n170 & n280 ) | ( n275 & n280 ) ;
  assign n282 = n170 & ~n239 ;
  assign n283 = ( n170 & ~n239 ) | ( n170 & n258 ) | ( ~n239 & n258 ) ;
  assign n284 = ( ~n243 & n282 ) | ( ~n243 & n283 ) | ( n282 & n283 ) ;
  assign n285 = ( n243 & n282 ) | ( n243 & n283 ) | ( n282 & n283 ) ;
  assign n286 = ( n243 & n284 ) | ( n243 & ~n285 ) | ( n284 & ~n285 ) ;
  assign n287 = ( ~n142 & n281 ) | ( ~n142 & n286 ) | ( n281 & n286 ) ;
  assign n288 = ( n142 & ~n244 ) | ( n142 & n258 ) | ( ~n244 & n258 ) ;
  assign n289 = n142 & ~n244 ;
  assign n290 = ( n249 & n288 ) | ( n249 & n289 ) | ( n288 & n289 ) ;
  assign n291 = ( ~n249 & n288 ) | ( ~n249 & n289 ) | ( n288 & n289 ) ;
  assign n292 = ( n249 & ~n290 ) | ( n249 & n291 ) | ( ~n290 & n291 ) ;
  assign n293 = ( ~n132 & n287 ) | ( ~n132 & n292 ) | ( n287 & n292 ) ;
  assign n294 = ( ~n131 & n263 ) | ( ~n131 & n293 ) | ( n263 & n293 ) ;
  assign n295 = n232 & ~n257 ;
  assign n296 = n227 & n256 ;
  assign n297 = n295 | n296 ;
  assign n298 = n294 | n297 ;
  assign n299 = n263 & ~n294 ;
  assign n300 = n293 & n297 ;
  assign n301 = n299 | n300 ;
  assign n302 = x110 | x111 ;
  assign n303 = x112 | n302 ;
  assign n304 = ~n258 & n303 ;
  assign n305 = ( x113 & ~n298 ) | ( x113 & n304 ) | ( ~n298 & n304 ) ;
  assign n306 = ~n265 & n298 ;
  assign n307 = n258 & ~n303 ;
  assign n308 = ( n305 & n306 ) | ( n305 & ~n307 ) | ( n306 & ~n307 ) ;
  assign n309 = n258 & ~n298 ;
  assign n310 = ( x114 & n306 ) | ( x114 & n309 ) | ( n306 & n309 ) ;
  assign n311 = ( ~x114 & n306 ) | ( ~x114 & n309 ) | ( n306 & n309 ) ;
  assign n312 = ( x114 & ~n310 ) | ( x114 & n311 ) | ( ~n310 & n311 ) ;
  assign n313 = ( ~n225 & n308 ) | ( ~n225 & n312 ) | ( n308 & n312 ) ;
  assign n314 = ~n225 & n258 ;
  assign n315 = ( n271 & n298 ) | ( n271 & n314 ) | ( n298 & n314 ) ;
  assign n316 = ( ~x115 & n311 ) | ( ~x115 & n315 ) | ( n311 & n315 ) ;
  assign n317 = ( x115 & n311 ) | ( x115 & n315 ) | ( n311 & n315 ) ;
  assign n318 = ( x115 & n316 ) | ( x115 & ~n317 ) | ( n316 & ~n317 ) ;
  assign n319 = ( ~n197 & n313 ) | ( ~n197 & n318 ) | ( n313 & n318 ) ;
  assign n320 = n197 & ~n270 ;
  assign n321 = ( n197 & ~n270 ) | ( n197 & n298 ) | ( ~n270 & n298 ) ;
  assign n322 = ( ~n274 & n320 ) | ( ~n274 & n321 ) | ( n320 & n321 ) ;
  assign n323 = ( n274 & n320 ) | ( n274 & n321 ) | ( n320 & n321 ) ;
  assign n324 = ( n274 & n322 ) | ( n274 & ~n323 ) | ( n322 & ~n323 ) ;
  assign n325 = ( ~n170 & n319 ) | ( ~n170 & n324 ) | ( n319 & n324 ) ;
  assign n326 = ( n170 & ~n275 ) | ( n170 & n298 ) | ( ~n275 & n298 ) ;
  assign n327 = n170 & ~n275 ;
  assign n328 = ( n280 & n326 ) | ( n280 & n327 ) | ( n326 & n327 ) ;
  assign n329 = ( ~n280 & n326 ) | ( ~n280 & n327 ) | ( n326 & n327 ) ;
  assign n330 = ( n280 & ~n328 ) | ( n280 & n329 ) | ( ~n328 & n329 ) ;
  assign n331 = ( ~n142 & n325 ) | ( ~n142 & n330 ) | ( n325 & n330 ) ;
  assign n332 = n142 & ~n281 ;
  assign n333 = ( n142 & ~n281 ) | ( n142 & n298 ) | ( ~n281 & n298 ) ;
  assign n334 = ( n286 & n332 ) | ( n286 & n333 ) | ( n332 & n333 ) ;
  assign n335 = ( ~n286 & n332 ) | ( ~n286 & n333 ) | ( n332 & n333 ) ;
  assign n336 = ( n286 & ~n334 ) | ( n286 & n335 ) | ( ~n334 & n335 ) ;
  assign n337 = ( ~n132 & n331 ) | ( ~n132 & n336 ) | ( n331 & n336 ) ;
  assign n338 = ( n132 & ~n287 ) | ( n132 & n298 ) | ( ~n287 & n298 ) ;
  assign n339 = n132 & ~n287 ;
  assign n340 = ( n292 & n338 ) | ( n292 & n339 ) | ( n338 & n339 ) ;
  assign n341 = ( ~n292 & n338 ) | ( ~n292 & n339 ) | ( n338 & n339 ) ;
  assign n342 = ( n292 & ~n340 ) | ( n292 & n341 ) | ( ~n340 & n341 ) ;
  assign n343 = ( ~n131 & n337 ) | ( ~n131 & n342 ) | ( n337 & n342 ) ;
  assign n344 = n301 | n343 ;
  assign n345 = n342 & ~n343 ;
  assign n346 = n301 & n337 ;
  assign n347 = n345 | n346 ;
  assign n348 = ( n132 & ~n331 ) | ( n132 & n344 ) | ( ~n331 & n344 ) ;
  assign n349 = n132 & ~n331 ;
  assign n350 = ( n336 & n348 ) | ( n336 & n349 ) | ( n348 & n349 ) ;
  assign n351 = ( n336 & ~n348 ) | ( n336 & n349 ) | ( ~n348 & n349 ) ;
  assign n352 = ( n348 & ~n350 ) | ( n348 & n351 ) | ( ~n350 & n351 ) ;
  assign n353 = x108 | x109 ;
  assign n354 = x110 | n353 ;
  assign n355 = n298 & ~n354 ;
  assign n356 = ~n302 & n344 ;
  assign n357 = ~n298 & n354 ;
  assign n358 = ( x111 & ~n344 ) | ( x111 & n357 ) | ( ~n344 & n357 ) ;
  assign n359 = ( ~n355 & n356 ) | ( ~n355 & n358 ) | ( n356 & n358 ) ;
  assign n360 = n298 & ~n344 ;
  assign n361 = ( ~x112 & n356 ) | ( ~x112 & n360 ) | ( n356 & n360 ) ;
  assign n362 = ( x112 & n356 ) | ( x112 & n360 ) | ( n356 & n360 ) ;
  assign n363 = ( x112 & n361 ) | ( x112 & ~n362 ) | ( n361 & ~n362 ) ;
  assign n364 = ( ~n258 & n359 ) | ( ~n258 & n363 ) | ( n359 & n363 ) ;
  assign n365 = ~n258 & n298 ;
  assign n366 = ( n309 & n344 ) | ( n309 & n365 ) | ( n344 & n365 ) ;
  assign n367 = ( x113 & n361 ) | ( x113 & n366 ) | ( n361 & n366 ) ;
  assign n368 = ( ~x113 & n361 ) | ( ~x113 & n366 ) | ( n361 & n366 ) ;
  assign n369 = ( x113 & ~n367 ) | ( x113 & n368 ) | ( ~n367 & n368 ) ;
  assign n370 = ( ~n225 & n364 ) | ( ~n225 & n369 ) | ( n364 & n369 ) ;
  assign n371 = ( n225 & ~n308 ) | ( n225 & n344 ) | ( ~n308 & n344 ) ;
  assign n372 = n225 & ~n308 ;
  assign n373 = ( n312 & n371 ) | ( n312 & n372 ) | ( n371 & n372 ) ;
  assign n374 = ( ~n312 & n371 ) | ( ~n312 & n372 ) | ( n371 & n372 ) ;
  assign n375 = ( n312 & ~n373 ) | ( n312 & n374 ) | ( ~n373 & n374 ) ;
  assign n376 = ( ~n197 & n370 ) | ( ~n197 & n375 ) | ( n370 & n375 ) ;
  assign n377 = ( n197 & ~n313 ) | ( n197 & n344 ) | ( ~n313 & n344 ) ;
  assign n378 = n197 & ~n313 ;
  assign n379 = ( n318 & n377 ) | ( n318 & n378 ) | ( n377 & n378 ) ;
  assign n380 = ( ~n318 & n377 ) | ( ~n318 & n378 ) | ( n377 & n378 ) ;
  assign n381 = ( n318 & ~n379 ) | ( n318 & n380 ) | ( ~n379 & n380 ) ;
  assign n382 = ( ~n170 & n376 ) | ( ~n170 & n381 ) | ( n376 & n381 ) ;
  assign n383 = ( n170 & ~n319 ) | ( n170 & n344 ) | ( ~n319 & n344 ) ;
  assign n384 = n170 & ~n319 ;
  assign n385 = ( n324 & n383 ) | ( n324 & n384 ) | ( n383 & n384 ) ;
  assign n386 = ( ~n324 & n383 ) | ( ~n324 & n384 ) | ( n383 & n384 ) ;
  assign n387 = ( n324 & ~n385 ) | ( n324 & n386 ) | ( ~n385 & n386 ) ;
  assign n388 = ( ~n142 & n382 ) | ( ~n142 & n387 ) | ( n382 & n387 ) ;
  assign n389 = ~n142 & n325 ;
  assign n390 = ( ~n142 & n325 ) | ( ~n142 & n344 ) | ( n325 & n344 ) ;
  assign n391 = ( ~n330 & n389 ) | ( ~n330 & n390 ) | ( n389 & n390 ) ;
  assign n392 = ( n330 & n389 ) | ( n330 & n390 ) | ( n389 & n390 ) ;
  assign n393 = ( n330 & n391 ) | ( n330 & ~n392 ) | ( n391 & ~n392 ) ;
  assign n394 = ( ~n132 & n388 ) | ( ~n132 & n393 ) | ( n388 & n393 ) ;
  assign n395 = ( ~n131 & n352 ) | ( ~n131 & n394 ) | ( n352 & n394 ) ;
  assign n396 = n347 | n395 ;
  assign n397 = n352 & ~n395 ;
  assign n398 = n347 & n394 ;
  assign n399 = n397 | n398 ;
  assign n400 = ( n132 & ~n388 ) | ( n132 & n396 ) | ( ~n388 & n396 ) ;
  assign n401 = n132 & ~n388 ;
  assign n402 = ( n393 & n400 ) | ( n393 & n401 ) | ( n400 & n401 ) ;
  assign n403 = ( n393 & ~n400 ) | ( n393 & n401 ) | ( ~n400 & n401 ) ;
  assign n404 = ( n400 & ~n402 ) | ( n400 & n403 ) | ( ~n402 & n403 ) ;
  assign n405 = ~n353 & n396 ;
  assign n406 = x106 | x107 ;
  assign n407 = x108 | n406 ;
  assign n408 = n344 & ~n407 ;
  assign n409 = ~n344 & n407 ;
  assign n410 = ( x109 & ~n396 ) | ( x109 & n409 ) | ( ~n396 & n409 ) ;
  assign n411 = ( n405 & ~n408 ) | ( n405 & n410 ) | ( ~n408 & n410 ) ;
  assign n412 = n344 & ~n396 ;
  assign n413 = ( x110 & n405 ) | ( x110 & n412 ) | ( n405 & n412 ) ;
  assign n414 = ( ~x110 & n405 ) | ( ~x110 & n412 ) | ( n405 & n412 ) ;
  assign n415 = ( x110 & ~n413 ) | ( x110 & n414 ) | ( ~n413 & n414 ) ;
  assign n416 = ( ~n298 & n411 ) | ( ~n298 & n415 ) | ( n411 & n415 ) ;
  assign n417 = ~n298 & n344 ;
  assign n418 = ( n360 & n396 ) | ( n360 & n417 ) | ( n396 & n417 ) ;
  assign n419 = ( ~x111 & n414 ) | ( ~x111 & n418 ) | ( n414 & n418 ) ;
  assign n420 = ( x111 & n414 ) | ( x111 & n418 ) | ( n414 & n418 ) ;
  assign n421 = ( x111 & n419 ) | ( x111 & ~n420 ) | ( n419 & ~n420 ) ;
  assign n422 = ( ~n258 & n416 ) | ( ~n258 & n421 ) | ( n416 & n421 ) ;
  assign n423 = ( n258 & ~n359 ) | ( n258 & n396 ) | ( ~n359 & n396 ) ;
  assign n424 = n258 & ~n359 ;
  assign n425 = ( n363 & n423 ) | ( n363 & n424 ) | ( n423 & n424 ) ;
  assign n426 = ( ~n363 & n423 ) | ( ~n363 & n424 ) | ( n423 & n424 ) ;
  assign n427 = ( n363 & ~n425 ) | ( n363 & n426 ) | ( ~n425 & n426 ) ;
  assign n428 = ( ~n225 & n422 ) | ( ~n225 & n427 ) | ( n422 & n427 ) ;
  assign n429 = n225 & ~n364 ;
  assign n430 = ( n225 & ~n364 ) | ( n225 & n396 ) | ( ~n364 & n396 ) ;
  assign n431 = ( n369 & n429 ) | ( n369 & n430 ) | ( n429 & n430 ) ;
  assign n432 = ( ~n369 & n429 ) | ( ~n369 & n430 ) | ( n429 & n430 ) ;
  assign n433 = ( n369 & ~n431 ) | ( n369 & n432 ) | ( ~n431 & n432 ) ;
  assign n434 = ( ~n197 & n428 ) | ( ~n197 & n433 ) | ( n428 & n433 ) ;
  assign n435 = ~n197 & n370 ;
  assign n436 = ( ~n197 & n370 ) | ( ~n197 & n396 ) | ( n370 & n396 ) ;
  assign n437 = ( n375 & n435 ) | ( n375 & n436 ) | ( n435 & n436 ) ;
  assign n438 = ( ~n375 & n435 ) | ( ~n375 & n436 ) | ( n435 & n436 ) ;
  assign n439 = ( n375 & ~n437 ) | ( n375 & n438 ) | ( ~n437 & n438 ) ;
  assign n440 = ( ~n170 & n434 ) | ( ~n170 & n439 ) | ( n434 & n439 ) ;
  assign n441 = ( n170 & ~n376 ) | ( n170 & n396 ) | ( ~n376 & n396 ) ;
  assign n442 = n170 & ~n376 ;
  assign n443 = ( n381 & n441 ) | ( n381 & n442 ) | ( n441 & n442 ) ;
  assign n444 = ( ~n381 & n441 ) | ( ~n381 & n442 ) | ( n441 & n442 ) ;
  assign n445 = ( n381 & ~n443 ) | ( n381 & n444 ) | ( ~n443 & n444 ) ;
  assign n446 = ( ~n142 & n440 ) | ( ~n142 & n445 ) | ( n440 & n445 ) ;
  assign n447 = ( n142 & ~n382 ) | ( n142 & n396 ) | ( ~n382 & n396 ) ;
  assign n448 = n142 & ~n382 ;
  assign n449 = ( n387 & n447 ) | ( n387 & n448 ) | ( n447 & n448 ) ;
  assign n450 = ( ~n387 & n447 ) | ( ~n387 & n448 ) | ( n447 & n448 ) ;
  assign n451 = ( n387 & ~n449 ) | ( n387 & n450 ) | ( ~n449 & n450 ) ;
  assign n452 = ( ~n132 & n446 ) | ( ~n132 & n451 ) | ( n446 & n451 ) ;
  assign n453 = ( ~n131 & n404 ) | ( ~n131 & n452 ) | ( n404 & n452 ) ;
  assign n454 = n399 | n453 ;
  assign n455 = n404 & ~n453 ;
  assign n456 = n399 & n452 ;
  assign n457 = n455 | n456 ;
  assign n458 = ( n132 & ~n446 ) | ( n132 & n454 ) | ( ~n446 & n454 ) ;
  assign n459 = n132 & ~n446 ;
  assign n460 = ( n451 & ~n458 ) | ( n451 & n459 ) | ( ~n458 & n459 ) ;
  assign n461 = ( n451 & n458 ) | ( n451 & n459 ) | ( n458 & n459 ) ;
  assign n462 = ( n458 & n460 ) | ( n458 & ~n461 ) | ( n460 & ~n461 ) ;
  assign n463 = x104 | x105 ;
  assign n464 = x106 | n463 ;
  assign n465 = n396 & ~n464 ;
  assign n466 = ~n406 & n454 ;
  assign n467 = ~n396 & n464 ;
  assign n468 = ( x107 & ~n454 ) | ( x107 & n467 ) | ( ~n454 & n467 ) ;
  assign n469 = ( ~n465 & n466 ) | ( ~n465 & n468 ) | ( n466 & n468 ) ;
  assign n470 = n396 & ~n454 ;
  assign n471 = ( x108 & n466 ) | ( x108 & n470 ) | ( n466 & n470 ) ;
  assign n472 = ( ~x108 & n466 ) | ( ~x108 & n470 ) | ( n466 & n470 ) ;
  assign n473 = ( x108 & ~n471 ) | ( x108 & n472 ) | ( ~n471 & n472 ) ;
  assign n474 = ( ~n344 & n469 ) | ( ~n344 & n473 ) | ( n469 & n473 ) ;
  assign n475 = ~n344 & n396 ;
  assign n476 = ( n412 & n454 ) | ( n412 & n475 ) | ( n454 & n475 ) ;
  assign n477 = ( ~x109 & n472 ) | ( ~x109 & n476 ) | ( n472 & n476 ) ;
  assign n478 = ( x109 & n472 ) | ( x109 & n476 ) | ( n472 & n476 ) ;
  assign n479 = ( x109 & n477 ) | ( x109 & ~n478 ) | ( n477 & ~n478 ) ;
  assign n480 = ( ~n298 & n474 ) | ( ~n298 & n479 ) | ( n474 & n479 ) ;
  assign n481 = ( n298 & ~n411 ) | ( n298 & n454 ) | ( ~n411 & n454 ) ;
  assign n482 = n298 & ~n411 ;
  assign n483 = ( ~n415 & n481 ) | ( ~n415 & n482 ) | ( n481 & n482 ) ;
  assign n484 = ( n415 & n481 ) | ( n415 & n482 ) | ( n481 & n482 ) ;
  assign n485 = ( n415 & n483 ) | ( n415 & ~n484 ) | ( n483 & ~n484 ) ;
  assign n486 = ( ~n258 & n480 ) | ( ~n258 & n485 ) | ( n480 & n485 ) ;
  assign n487 = ( n258 & ~n416 ) | ( n258 & n454 ) | ( ~n416 & n454 ) ;
  assign n488 = n258 & ~n416 ;
  assign n489 = ( n421 & n487 ) | ( n421 & n488 ) | ( n487 & n488 ) ;
  assign n490 = ( ~n421 & n487 ) | ( ~n421 & n488 ) | ( n487 & n488 ) ;
  assign n491 = ( n421 & ~n489 ) | ( n421 & n490 ) | ( ~n489 & n490 ) ;
  assign n492 = ( ~n225 & n486 ) | ( ~n225 & n491 ) | ( n486 & n491 ) ;
  assign n493 = ~n225 & n422 ;
  assign n494 = ( ~n225 & n422 ) | ( ~n225 & n454 ) | ( n422 & n454 ) ;
  assign n495 = ( ~n427 & n493 ) | ( ~n427 & n494 ) | ( n493 & n494 ) ;
  assign n496 = ( n427 & n493 ) | ( n427 & n494 ) | ( n493 & n494 ) ;
  assign n497 = ( n427 & n495 ) | ( n427 & ~n496 ) | ( n495 & ~n496 ) ;
  assign n498 = ( ~n197 & n492 ) | ( ~n197 & n497 ) | ( n492 & n497 ) ;
  assign n499 = ( n197 & ~n428 ) | ( n197 & n454 ) | ( ~n428 & n454 ) ;
  assign n500 = n197 & ~n428 ;
  assign n501 = ( n433 & n499 ) | ( n433 & n500 ) | ( n499 & n500 ) ;
  assign n502 = ( ~n433 & n499 ) | ( ~n433 & n500 ) | ( n499 & n500 ) ;
  assign n503 = ( n433 & ~n501 ) | ( n433 & n502 ) | ( ~n501 & n502 ) ;
  assign n504 = ( ~n170 & n498 ) | ( ~n170 & n503 ) | ( n498 & n503 ) ;
  assign n505 = ~n170 & n434 ;
  assign n506 = ( ~n170 & n434 ) | ( ~n170 & n454 ) | ( n434 & n454 ) ;
  assign n507 = ( ~n439 & n505 ) | ( ~n439 & n506 ) | ( n505 & n506 ) ;
  assign n508 = ( n439 & n505 ) | ( n439 & n506 ) | ( n505 & n506 ) ;
  assign n509 = ( n439 & n507 ) | ( n439 & ~n508 ) | ( n507 & ~n508 ) ;
  assign n510 = ( ~n142 & n504 ) | ( ~n142 & n509 ) | ( n504 & n509 ) ;
  assign n511 = ~n142 & n440 ;
  assign n512 = ( ~n142 & n440 ) | ( ~n142 & n454 ) | ( n440 & n454 ) ;
  assign n513 = ( ~n445 & n511 ) | ( ~n445 & n512 ) | ( n511 & n512 ) ;
  assign n514 = ( n445 & n511 ) | ( n445 & n512 ) | ( n511 & n512 ) ;
  assign n515 = ( n445 & n513 ) | ( n445 & ~n514 ) | ( n513 & ~n514 ) ;
  assign n516 = ( ~n132 & n510 ) | ( ~n132 & n515 ) | ( n510 & n515 ) ;
  assign n517 = ( ~n131 & n462 ) | ( ~n131 & n516 ) | ( n462 & n516 ) ;
  assign n518 = n457 | n517 ;
  assign n519 = n462 & ~n517 ;
  assign n520 = n457 & n516 ;
  assign n521 = n519 | n520 ;
  assign n522 = ( n132 & ~n510 ) | ( n132 & n518 ) | ( ~n510 & n518 ) ;
  assign n523 = n132 & ~n510 ;
  assign n524 = ( n515 & ~n522 ) | ( n515 & n523 ) | ( ~n522 & n523 ) ;
  assign n525 = ( n515 & n522 ) | ( n515 & n523 ) | ( n522 & n523 ) ;
  assign n526 = ( n522 & n524 ) | ( n522 & ~n525 ) | ( n524 & ~n525 ) ;
  assign n527 = ~n463 & n518 ;
  assign n528 = x102 | x103 ;
  assign n529 = x104 | n528 ;
  assign n530 = n454 & ~n529 ;
  assign n531 = ~n454 & n529 ;
  assign n532 = ( x105 & ~n518 ) | ( x105 & n531 ) | ( ~n518 & n531 ) ;
  assign n533 = ( n527 & ~n530 ) | ( n527 & n532 ) | ( ~n530 & n532 ) ;
  assign n534 = n454 & ~n518 ;
  assign n535 = ( x106 & n527 ) | ( x106 & n534 ) | ( n527 & n534 ) ;
  assign n536 = ( ~x106 & n527 ) | ( ~x106 & n534 ) | ( n527 & n534 ) ;
  assign n537 = ( x106 & ~n535 ) | ( x106 & n536 ) | ( ~n535 & n536 ) ;
  assign n538 = ( ~n396 & n533 ) | ( ~n396 & n537 ) | ( n533 & n537 ) ;
  assign n539 = ~n396 & n454 ;
  assign n540 = ( n470 & n518 ) | ( n470 & n539 ) | ( n518 & n539 ) ;
  assign n541 = ( x107 & n536 ) | ( x107 & n540 ) | ( n536 & n540 ) ;
  assign n542 = ( ~x107 & n536 ) | ( ~x107 & n540 ) | ( n536 & n540 ) ;
  assign n543 = ( x107 & ~n541 ) | ( x107 & n542 ) | ( ~n541 & n542 ) ;
  assign n544 = ( ~n344 & n538 ) | ( ~n344 & n543 ) | ( n538 & n543 ) ;
  assign n545 = ( n344 & ~n469 ) | ( n344 & n518 ) | ( ~n469 & n518 ) ;
  assign n546 = n344 & ~n469 ;
  assign n547 = ( n473 & n545 ) | ( n473 & n546 ) | ( n545 & n546 ) ;
  assign n548 = ( ~n473 & n545 ) | ( ~n473 & n546 ) | ( n545 & n546 ) ;
  assign n549 = ( n473 & ~n547 ) | ( n473 & n548 ) | ( ~n547 & n548 ) ;
  assign n550 = ( ~n298 & n544 ) | ( ~n298 & n549 ) | ( n544 & n549 ) ;
  assign n551 = ( n298 & ~n474 ) | ( n298 & n518 ) | ( ~n474 & n518 ) ;
  assign n552 = n298 & ~n474 ;
  assign n553 = ( n479 & n551 ) | ( n479 & n552 ) | ( n551 & n552 ) ;
  assign n554 = ( ~n479 & n551 ) | ( ~n479 & n552 ) | ( n551 & n552 ) ;
  assign n555 = ( n479 & ~n553 ) | ( n479 & n554 ) | ( ~n553 & n554 ) ;
  assign n556 = ( ~n258 & n550 ) | ( ~n258 & n555 ) | ( n550 & n555 ) ;
  assign n557 = ( n258 & ~n480 ) | ( n258 & n518 ) | ( ~n480 & n518 ) ;
  assign n558 = n258 & ~n480 ;
  assign n559 = ( n485 & n557 ) | ( n485 & n558 ) | ( n557 & n558 ) ;
  assign n560 = ( ~n485 & n557 ) | ( ~n485 & n558 ) | ( n557 & n558 ) ;
  assign n561 = ( n485 & ~n559 ) | ( n485 & n560 ) | ( ~n559 & n560 ) ;
  assign n562 = ( ~n225 & n556 ) | ( ~n225 & n561 ) | ( n556 & n561 ) ;
  assign n563 = n225 & ~n486 ;
  assign n564 = ( n225 & ~n486 ) | ( n225 & n518 ) | ( ~n486 & n518 ) ;
  assign n565 = ( n491 & n563 ) | ( n491 & n564 ) | ( n563 & n564 ) ;
  assign n566 = ( ~n491 & n563 ) | ( ~n491 & n564 ) | ( n563 & n564 ) ;
  assign n567 = ( n491 & ~n565 ) | ( n491 & n566 ) | ( ~n565 & n566 ) ;
  assign n568 = ( ~n197 & n562 ) | ( ~n197 & n567 ) | ( n562 & n567 ) ;
  assign n569 = ( n197 & ~n492 ) | ( n197 & n518 ) | ( ~n492 & n518 ) ;
  assign n570 = n197 & ~n492 ;
  assign n571 = ( n497 & n569 ) | ( n497 & n570 ) | ( n569 & n570 ) ;
  assign n572 = ( ~n497 & n569 ) | ( ~n497 & n570 ) | ( n569 & n570 ) ;
  assign n573 = ( n497 & ~n571 ) | ( n497 & n572 ) | ( ~n571 & n572 ) ;
  assign n574 = ( ~n170 & n568 ) | ( ~n170 & n573 ) | ( n568 & n573 ) ;
  assign n575 = ( n170 & ~n498 ) | ( n170 & n518 ) | ( ~n498 & n518 ) ;
  assign n576 = n170 & ~n498 ;
  assign n577 = ( n503 & n575 ) | ( n503 & n576 ) | ( n575 & n576 ) ;
  assign n578 = ( ~n503 & n575 ) | ( ~n503 & n576 ) | ( n575 & n576 ) ;
  assign n579 = ( n503 & ~n577 ) | ( n503 & n578 ) | ( ~n577 & n578 ) ;
  assign n580 = ( ~n142 & n574 ) | ( ~n142 & n579 ) | ( n574 & n579 ) ;
  assign n581 = ~n142 & n504 ;
  assign n582 = ( ~n142 & n504 ) | ( ~n142 & n518 ) | ( n504 & n518 ) ;
  assign n583 = ( ~n509 & n581 ) | ( ~n509 & n582 ) | ( n581 & n582 ) ;
  assign n584 = ( n509 & n581 ) | ( n509 & n582 ) | ( n581 & n582 ) ;
  assign n585 = ( n509 & n583 ) | ( n509 & ~n584 ) | ( n583 & ~n584 ) ;
  assign n586 = ( ~n132 & n580 ) | ( ~n132 & n585 ) | ( n580 & n585 ) ;
  assign n587 = ( ~n131 & n526 ) | ( ~n131 & n586 ) | ( n526 & n586 ) ;
  assign n588 = n521 | n587 ;
  assign n589 = n526 & ~n587 ;
  assign n590 = n521 & n586 ;
  assign n591 = n589 | n590 ;
  assign n592 = ( n132 & ~n580 ) | ( n132 & n588 ) | ( ~n580 & n588 ) ;
  assign n593 = n132 & ~n580 ;
  assign n594 = ( n585 & ~n592 ) | ( n585 & n593 ) | ( ~n592 & n593 ) ;
  assign n595 = ( n585 & n592 ) | ( n585 & n593 ) | ( n592 & n593 ) ;
  assign n596 = ( n592 & n594 ) | ( n592 & ~n595 ) | ( n594 & ~n595 ) ;
  assign n597 = x100 | x101 ;
  assign n598 = x102 | n597 ;
  assign n599 = ~n518 & n598 ;
  assign n600 = ( x103 & ~n588 ) | ( x103 & n599 ) | ( ~n588 & n599 ) ;
  assign n601 = ~n528 & n588 ;
  assign n602 = n518 & ~n598 ;
  assign n603 = ( n600 & n601 ) | ( n600 & ~n602 ) | ( n601 & ~n602 ) ;
  assign n604 = n518 & ~n588 ;
  assign n605 = ( x104 & n601 ) | ( x104 & n604 ) | ( n601 & n604 ) ;
  assign n606 = ( ~x104 & n601 ) | ( ~x104 & n604 ) | ( n601 & n604 ) ;
  assign n607 = ( x104 & ~n605 ) | ( x104 & n606 ) | ( ~n605 & n606 ) ;
  assign n608 = ( ~n454 & n603 ) | ( ~n454 & n607 ) | ( n603 & n607 ) ;
  assign n609 = ~n454 & n518 ;
  assign n610 = ( n534 & n588 ) | ( n534 & n609 ) | ( n588 & n609 ) ;
  assign n611 = ( x105 & n606 ) | ( x105 & n610 ) | ( n606 & n610 ) ;
  assign n612 = ( ~x105 & n606 ) | ( ~x105 & n610 ) | ( n606 & n610 ) ;
  assign n613 = ( x105 & ~n611 ) | ( x105 & n612 ) | ( ~n611 & n612 ) ;
  assign n614 = ( ~n396 & n608 ) | ( ~n396 & n613 ) | ( n608 & n613 ) ;
  assign n615 = ( n396 & ~n533 ) | ( n396 & n588 ) | ( ~n533 & n588 ) ;
  assign n616 = n396 & ~n533 ;
  assign n617 = ( n537 & n615 ) | ( n537 & n616 ) | ( n615 & n616 ) ;
  assign n618 = ( ~n537 & n615 ) | ( ~n537 & n616 ) | ( n615 & n616 ) ;
  assign n619 = ( n537 & ~n617 ) | ( n537 & n618 ) | ( ~n617 & n618 ) ;
  assign n620 = ( ~n344 & n614 ) | ( ~n344 & n619 ) | ( n614 & n619 ) ;
  assign n621 = ( n344 & ~n538 ) | ( n344 & n588 ) | ( ~n538 & n588 ) ;
  assign n622 = n344 & ~n538 ;
  assign n623 = ( n543 & n621 ) | ( n543 & n622 ) | ( n621 & n622 ) ;
  assign n624 = ( ~n543 & n621 ) | ( ~n543 & n622 ) | ( n621 & n622 ) ;
  assign n625 = ( n543 & ~n623 ) | ( n543 & n624 ) | ( ~n623 & n624 ) ;
  assign n626 = ( ~n298 & n620 ) | ( ~n298 & n625 ) | ( n620 & n625 ) ;
  assign n627 = ~n298 & n544 ;
  assign n628 = ( ~n298 & n544 ) | ( ~n298 & n588 ) | ( n544 & n588 ) ;
  assign n629 = ( ~n549 & n627 ) | ( ~n549 & n628 ) | ( n627 & n628 ) ;
  assign n630 = ( n549 & n627 ) | ( n549 & n628 ) | ( n627 & n628 ) ;
  assign n631 = ( n549 & n629 ) | ( n549 & ~n630 ) | ( n629 & ~n630 ) ;
  assign n632 = ( ~n258 & n626 ) | ( ~n258 & n631 ) | ( n626 & n631 ) ;
  assign n633 = ~n258 & n550 ;
  assign n634 = ( ~n258 & n550 ) | ( ~n258 & n588 ) | ( n550 & n588 ) ;
  assign n635 = ( ~n555 & n633 ) | ( ~n555 & n634 ) | ( n633 & n634 ) ;
  assign n636 = ( n555 & n633 ) | ( n555 & n634 ) | ( n633 & n634 ) ;
  assign n637 = ( n555 & n635 ) | ( n555 & ~n636 ) | ( n635 & ~n636 ) ;
  assign n638 = ( ~n225 & n632 ) | ( ~n225 & n637 ) | ( n632 & n637 ) ;
  assign n639 = ( n225 & ~n556 ) | ( n225 & n588 ) | ( ~n556 & n588 ) ;
  assign n640 = n225 & ~n556 ;
  assign n641 = ( n561 & n639 ) | ( n561 & n640 ) | ( n639 & n640 ) ;
  assign n642 = ( ~n561 & n639 ) | ( ~n561 & n640 ) | ( n639 & n640 ) ;
  assign n643 = ( n561 & ~n641 ) | ( n561 & n642 ) | ( ~n641 & n642 ) ;
  assign n644 = ( ~n197 & n638 ) | ( ~n197 & n643 ) | ( n638 & n643 ) ;
  assign n645 = ~n197 & n562 ;
  assign n646 = ( ~n197 & n562 ) | ( ~n197 & n588 ) | ( n562 & n588 ) ;
  assign n647 = ( n567 & n645 ) | ( n567 & n646 ) | ( n645 & n646 ) ;
  assign n648 = ( ~n567 & n645 ) | ( ~n567 & n646 ) | ( n645 & n646 ) ;
  assign n649 = ( n567 & ~n647 ) | ( n567 & n648 ) | ( ~n647 & n648 ) ;
  assign n650 = ( ~n170 & n644 ) | ( ~n170 & n649 ) | ( n644 & n649 ) ;
  assign n651 = ~n170 & n568 ;
  assign n652 = ( ~n170 & n568 ) | ( ~n170 & n588 ) | ( n568 & n588 ) ;
  assign n653 = ( ~n573 & n651 ) | ( ~n573 & n652 ) | ( n651 & n652 ) ;
  assign n654 = ( n573 & n651 ) | ( n573 & n652 ) | ( n651 & n652 ) ;
  assign n655 = ( n573 & n653 ) | ( n573 & ~n654 ) | ( n653 & ~n654 ) ;
  assign n656 = ( ~n142 & n650 ) | ( ~n142 & n655 ) | ( n650 & n655 ) ;
  assign n657 = ~n142 & n574 ;
  assign n658 = ( ~n142 & n574 ) | ( ~n142 & n588 ) | ( n574 & n588 ) ;
  assign n659 = ( n579 & n657 ) | ( n579 & n658 ) | ( n657 & n658 ) ;
  assign n660 = ( ~n579 & n657 ) | ( ~n579 & n658 ) | ( n657 & n658 ) ;
  assign n661 = ( n579 & ~n659 ) | ( n579 & n660 ) | ( ~n659 & n660 ) ;
  assign n662 = ( ~n132 & n656 ) | ( ~n132 & n661 ) | ( n656 & n661 ) ;
  assign n663 = ( ~n131 & n596 ) | ( ~n131 & n662 ) | ( n596 & n662 ) ;
  assign n664 = n591 | n663 ;
  assign n665 = ( n132 & ~n656 ) | ( n132 & n664 ) | ( ~n656 & n664 ) ;
  assign n666 = n132 & ~n656 ;
  assign n667 = ( n661 & ~n665 ) | ( n661 & n666 ) | ( ~n665 & n666 ) ;
  assign n668 = ( n661 & n665 ) | ( n661 & n666 ) | ( n665 & n666 ) ;
  assign n669 = ( n665 & n667 ) | ( n665 & ~n668 ) | ( n667 & ~n668 ) ;
  assign n670 = ~n597 & n664 ;
  assign n671 = x98 | x99 ;
  assign n672 = x100 | n671 ;
  assign n673 = n588 & ~n672 ;
  assign n674 = ~n588 & n672 ;
  assign n675 = ( x101 & ~n664 ) | ( x101 & n674 ) | ( ~n664 & n674 ) ;
  assign n676 = ( n670 & ~n673 ) | ( n670 & n675 ) | ( ~n673 & n675 ) ;
  assign n677 = n588 & ~n664 ;
  assign n678 = ( x102 & n670 ) | ( x102 & n677 ) | ( n670 & n677 ) ;
  assign n679 = ( ~x102 & n670 ) | ( ~x102 & n677 ) | ( n670 & n677 ) ;
  assign n680 = ( x102 & ~n678 ) | ( x102 & n679 ) | ( ~n678 & n679 ) ;
  assign n681 = ( ~n518 & n676 ) | ( ~n518 & n680 ) | ( n676 & n680 ) ;
  assign n682 = ~n518 & n588 ;
  assign n683 = ( n604 & n664 ) | ( n604 & n682 ) | ( n664 & n682 ) ;
  assign n684 = ( ~x103 & n679 ) | ( ~x103 & n683 ) | ( n679 & n683 ) ;
  assign n685 = ( x103 & n679 ) | ( x103 & n683 ) | ( n679 & n683 ) ;
  assign n686 = ( x103 & n684 ) | ( x103 & ~n685 ) | ( n684 & ~n685 ) ;
  assign n687 = ( ~n454 & n681 ) | ( ~n454 & n686 ) | ( n681 & n686 ) ;
  assign n688 = ( n454 & ~n603 ) | ( n454 & n664 ) | ( ~n603 & n664 ) ;
  assign n689 = n454 & ~n603 ;
  assign n690 = ( n607 & n688 ) | ( n607 & n689 ) | ( n688 & n689 ) ;
  assign n691 = ( ~n607 & n688 ) | ( ~n607 & n689 ) | ( n688 & n689 ) ;
  assign n692 = ( n607 & ~n690 ) | ( n607 & n691 ) | ( ~n690 & n691 ) ;
  assign n693 = ( ~n396 & n687 ) | ( ~n396 & n692 ) | ( n687 & n692 ) ;
  assign n694 = ( n396 & ~n608 ) | ( n396 & n664 ) | ( ~n608 & n664 ) ;
  assign n695 = n396 & ~n608 ;
  assign n696 = ( n613 & n694 ) | ( n613 & n695 ) | ( n694 & n695 ) ;
  assign n697 = ( ~n613 & n694 ) | ( ~n613 & n695 ) | ( n694 & n695 ) ;
  assign n698 = ( n613 & ~n696 ) | ( n613 & n697 ) | ( ~n696 & n697 ) ;
  assign n699 = ( ~n344 & n693 ) | ( ~n344 & n698 ) | ( n693 & n698 ) ;
  assign n700 = ( n344 & ~n614 ) | ( n344 & n664 ) | ( ~n614 & n664 ) ;
  assign n701 = n344 & ~n614 ;
  assign n702 = ( n619 & n700 ) | ( n619 & n701 ) | ( n700 & n701 ) ;
  assign n703 = ( ~n619 & n700 ) | ( ~n619 & n701 ) | ( n700 & n701 ) ;
  assign n704 = ( n619 & ~n702 ) | ( n619 & n703 ) | ( ~n702 & n703 ) ;
  assign n705 = ( ~n298 & n699 ) | ( ~n298 & n704 ) | ( n699 & n704 ) ;
  assign n706 = ( n298 & ~n620 ) | ( n298 & n664 ) | ( ~n620 & n664 ) ;
  assign n707 = n298 & ~n620 ;
  assign n708 = ( n625 & n706 ) | ( n625 & n707 ) | ( n706 & n707 ) ;
  assign n709 = ( ~n625 & n706 ) | ( ~n625 & n707 ) | ( n706 & n707 ) ;
  assign n710 = ( n625 & ~n708 ) | ( n625 & n709 ) | ( ~n708 & n709 ) ;
  assign n711 = ( ~n258 & n705 ) | ( ~n258 & n710 ) | ( n705 & n710 ) ;
  assign n712 = ~n258 & n626 ;
  assign n713 = ( ~n258 & n626 ) | ( ~n258 & n664 ) | ( n626 & n664 ) ;
  assign n714 = ( n631 & n712 ) | ( n631 & n713 ) | ( n712 & n713 ) ;
  assign n715 = ( ~n631 & n712 ) | ( ~n631 & n713 ) | ( n712 & n713 ) ;
  assign n716 = ( n631 & ~n714 ) | ( n631 & n715 ) | ( ~n714 & n715 ) ;
  assign n717 = ( ~n225 & n711 ) | ( ~n225 & n716 ) | ( n711 & n716 ) ;
  assign n718 = n225 & ~n632 ;
  assign n719 = ( n225 & ~n632 ) | ( n225 & n664 ) | ( ~n632 & n664 ) ;
  assign n720 = ( n637 & n718 ) | ( n637 & n719 ) | ( n718 & n719 ) ;
  assign n721 = ( ~n637 & n718 ) | ( ~n637 & n719 ) | ( n718 & n719 ) ;
  assign n722 = ( n637 & ~n720 ) | ( n637 & n721 ) | ( ~n720 & n721 ) ;
  assign n723 = ( ~n197 & n717 ) | ( ~n197 & n722 ) | ( n717 & n722 ) ;
  assign n724 = ( n197 & ~n638 ) | ( n197 & n664 ) | ( ~n638 & n664 ) ;
  assign n725 = n197 & ~n638 ;
  assign n726 = ( n643 & n724 ) | ( n643 & n725 ) | ( n724 & n725 ) ;
  assign n727 = ( ~n643 & n724 ) | ( ~n643 & n725 ) | ( n724 & n725 ) ;
  assign n728 = ( n643 & ~n726 ) | ( n643 & n727 ) | ( ~n726 & n727 ) ;
  assign n729 = ( ~n170 & n723 ) | ( ~n170 & n728 ) | ( n723 & n728 ) ;
  assign n730 = ~n170 & n644 ;
  assign n731 = ( ~n170 & n644 ) | ( ~n170 & n664 ) | ( n644 & n664 ) ;
  assign n732 = ( n649 & n730 ) | ( n649 & n731 ) | ( n730 & n731 ) ;
  assign n733 = ( ~n649 & n730 ) | ( ~n649 & n731 ) | ( n730 & n731 ) ;
  assign n734 = ( n649 & ~n732 ) | ( n649 & n733 ) | ( ~n732 & n733 ) ;
  assign n735 = ( ~n142 & n729 ) | ( ~n142 & n734 ) | ( n729 & n734 ) ;
  assign n736 = ~n142 & n650 ;
  assign n737 = ( ~n142 & n650 ) | ( ~n142 & n664 ) | ( n650 & n664 ) ;
  assign n738 = ( ~n655 & n736 ) | ( ~n655 & n737 ) | ( n736 & n737 ) ;
  assign n739 = ( n655 & n736 ) | ( n655 & n737 ) | ( n736 & n737 ) ;
  assign n740 = ( n655 & n738 ) | ( n655 & ~n739 ) | ( n738 & ~n739 ) ;
  assign n741 = ( ~n132 & n735 ) | ( ~n132 & n740 ) | ( n735 & n740 ) ;
  assign n742 = ( ~n131 & n669 ) | ( ~n131 & n741 ) | ( n669 & n741 ) ;
  assign n743 = n591 | n596 ;
  assign n744 = ( n596 & n662 ) | ( n596 & n743 ) | ( n662 & n743 ) ;
  assign n745 = ~n663 & n744 ;
  assign n746 = n742 | n745 ;
  assign n747 = x96 | x97 ;
  assign n748 = ~x98 & n747 ;
  assign n749 = x98 | n747 ;
  assign n750 = ( ~n746 & n748 ) | ( ~n746 & n749 ) | ( n748 & n749 ) ;
  assign n751 = ( ~x98 & n742 ) | ( ~x98 & n745 ) | ( n742 & n745 ) ;
  assign n752 = ~x99 & n751 ;
  assign n753 = x99 & ~n751 ;
  assign n754 = n752 | n753 ;
  assign n755 = ( ~n664 & n750 ) | ( ~n664 & n754 ) | ( n750 & n754 ) ;
  assign n756 = n664 & ~n746 ;
  assign n757 = ( ~x100 & n752 ) | ( ~x100 & n756 ) | ( n752 & n756 ) ;
  assign n758 = ( x100 & n752 ) | ( x100 & n756 ) | ( n752 & n756 ) ;
  assign n759 = ( x100 & n757 ) | ( x100 & ~n758 ) | ( n757 & ~n758 ) ;
  assign n760 = ( ~n588 & n755 ) | ( ~n588 & n759 ) | ( n755 & n759 ) ;
  assign n761 = ~x100 & n756 ;
  assign n762 = n673 | n674 ;
  assign n763 = n664 & n762 ;
  assign n764 = n664 | n762 ;
  assign n765 = ( n746 & n763 ) | ( n746 & ~n764 ) | ( n763 & ~n764 ) ;
  assign n766 = ( ~x101 & n761 ) | ( ~x101 & n765 ) | ( n761 & n765 ) ;
  assign n767 = ( x101 & n761 ) | ( x101 & n765 ) | ( n761 & n765 ) ;
  assign n768 = ( x101 & n766 ) | ( x101 & ~n767 ) | ( n766 & ~n767 ) ;
  assign n769 = ( ~n518 & n760 ) | ( ~n518 & n768 ) | ( n760 & n768 ) ;
  assign n770 = n518 & ~n676 ;
  assign n771 = ( n518 & ~n676 ) | ( n518 & n746 ) | ( ~n676 & n746 ) ;
  assign n772 = ( n680 & n770 ) | ( n680 & n771 ) | ( n770 & n771 ) ;
  assign n773 = ( ~n680 & n770 ) | ( ~n680 & n771 ) | ( n770 & n771 ) ;
  assign n774 = ( n680 & ~n772 ) | ( n680 & n773 ) | ( ~n772 & n773 ) ;
  assign n775 = ( ~n454 & n769 ) | ( ~n454 & n774 ) | ( n769 & n774 ) ;
  assign n776 = ( n454 & ~n681 ) | ( n454 & n746 ) | ( ~n681 & n746 ) ;
  assign n777 = n454 & ~n681 ;
  assign n778 = ( n686 & n776 ) | ( n686 & n777 ) | ( n776 & n777 ) ;
  assign n779 = ( ~n686 & n776 ) | ( ~n686 & n777 ) | ( n776 & n777 ) ;
  assign n780 = ( n686 & ~n778 ) | ( n686 & n779 ) | ( ~n778 & n779 ) ;
  assign n781 = ( ~n396 & n775 ) | ( ~n396 & n780 ) | ( n775 & n780 ) ;
  assign n782 = ( n396 & ~n687 ) | ( n396 & n746 ) | ( ~n687 & n746 ) ;
  assign n783 = n396 & ~n687 ;
  assign n784 = ( n692 & n782 ) | ( n692 & n783 ) | ( n782 & n783 ) ;
  assign n785 = ( ~n692 & n782 ) | ( ~n692 & n783 ) | ( n782 & n783 ) ;
  assign n786 = ( n692 & ~n784 ) | ( n692 & n785 ) | ( ~n784 & n785 ) ;
  assign n787 = ( ~n344 & n781 ) | ( ~n344 & n786 ) | ( n781 & n786 ) ;
  assign n788 = ~n344 & n693 ;
  assign n789 = ( ~n344 & n693 ) | ( ~n344 & n746 ) | ( n693 & n746 ) ;
  assign n790 = ( ~n698 & n788 ) | ( ~n698 & n789 ) | ( n788 & n789 ) ;
  assign n791 = ( n698 & n788 ) | ( n698 & n789 ) | ( n788 & n789 ) ;
  assign n792 = ( n698 & n790 ) | ( n698 & ~n791 ) | ( n790 & ~n791 ) ;
  assign n793 = ( ~n298 & n787 ) | ( ~n298 & n792 ) | ( n787 & n792 ) ;
  assign n794 = ~n298 & n699 ;
  assign n795 = ( ~n298 & n699 ) | ( ~n298 & n746 ) | ( n699 & n746 ) ;
  assign n796 = ( ~n704 & n794 ) | ( ~n704 & n795 ) | ( n794 & n795 ) ;
  assign n797 = ( n704 & n794 ) | ( n704 & n795 ) | ( n794 & n795 ) ;
  assign n798 = ( n704 & n796 ) | ( n704 & ~n797 ) | ( n796 & ~n797 ) ;
  assign n799 = ( ~n258 & n793 ) | ( ~n258 & n798 ) | ( n793 & n798 ) ;
  assign n800 = ( n258 & ~n705 ) | ( n258 & n746 ) | ( ~n705 & n746 ) ;
  assign n801 = n258 & ~n705 ;
  assign n802 = ( n710 & n800 ) | ( n710 & n801 ) | ( n800 & n801 ) ;
  assign n803 = ( ~n710 & n800 ) | ( ~n710 & n801 ) | ( n800 & n801 ) ;
  assign n804 = ( n710 & ~n802 ) | ( n710 & n803 ) | ( ~n802 & n803 ) ;
  assign n805 = ( ~n225 & n799 ) | ( ~n225 & n804 ) | ( n799 & n804 ) ;
  assign n806 = ( n225 & ~n711 ) | ( n225 & n746 ) | ( ~n711 & n746 ) ;
  assign n807 = n225 & ~n711 ;
  assign n808 = ( n716 & n806 ) | ( n716 & n807 ) | ( n806 & n807 ) ;
  assign n809 = ( ~n716 & n806 ) | ( ~n716 & n807 ) | ( n806 & n807 ) ;
  assign n810 = ( n716 & ~n808 ) | ( n716 & n809 ) | ( ~n808 & n809 ) ;
  assign n811 = ( ~n197 & n805 ) | ( ~n197 & n810 ) | ( n805 & n810 ) ;
  assign n812 = ( n197 & ~n717 ) | ( n197 & n746 ) | ( ~n717 & n746 ) ;
  assign n813 = n197 & ~n717 ;
  assign n814 = ( n722 & n812 ) | ( n722 & n813 ) | ( n812 & n813 ) ;
  assign n815 = ( ~n722 & n812 ) | ( ~n722 & n813 ) | ( n812 & n813 ) ;
  assign n816 = ( n722 & ~n814 ) | ( n722 & n815 ) | ( ~n814 & n815 ) ;
  assign n817 = ( ~n170 & n811 ) | ( ~n170 & n816 ) | ( n811 & n816 ) ;
  assign n818 = ( n170 & ~n723 ) | ( n170 & n746 ) | ( ~n723 & n746 ) ;
  assign n819 = n170 & ~n723 ;
  assign n820 = ( n728 & n818 ) | ( n728 & n819 ) | ( n818 & n819 ) ;
  assign n821 = ( ~n728 & n818 ) | ( ~n728 & n819 ) | ( n818 & n819 ) ;
  assign n822 = ( n728 & ~n820 ) | ( n728 & n821 ) | ( ~n820 & n821 ) ;
  assign n823 = ( ~n142 & n817 ) | ( ~n142 & n822 ) | ( n817 & n822 ) ;
  assign n824 = ( n142 & ~n729 ) | ( n142 & n746 ) | ( ~n729 & n746 ) ;
  assign n825 = n142 & ~n729 ;
  assign n826 = ( n734 & n824 ) | ( n734 & n825 ) | ( n824 & n825 ) ;
  assign n827 = ( ~n734 & n824 ) | ( ~n734 & n825 ) | ( n824 & n825 ) ;
  assign n828 = ( n734 & ~n826 ) | ( n734 & n827 ) | ( ~n826 & n827 ) ;
  assign n829 = ( ~n132 & n823 ) | ( ~n132 & n828 ) | ( n823 & n828 ) ;
  assign n830 = ( n132 & ~n735 ) | ( n132 & n746 ) | ( ~n735 & n746 ) ;
  assign n831 = n132 & ~n735 ;
  assign n832 = ( n740 & n830 ) | ( n740 & n831 ) | ( n830 & n831 ) ;
  assign n833 = ( ~n740 & n830 ) | ( ~n740 & n831 ) | ( n830 & n831 ) ;
  assign n834 = ( n740 & ~n832 ) | ( n740 & n833 ) | ( ~n832 & n833 ) ;
  assign n835 = ( ~n131 & n829 ) | ( ~n131 & n834 ) | ( n829 & n834 ) ;
  assign n836 = n669 | n745 ;
  assign n837 = ( n669 & n741 ) | ( n669 & n836 ) | ( n741 & n836 ) ;
  assign n838 = ~n742 & n837 ;
  assign n839 = n835 | n838 ;
  assign n840 = ( n829 & n835 ) | ( n829 & ~n838 ) | ( n835 & ~n838 ) ;
  assign n841 = ( n131 & n829 ) | ( n131 & n834 ) | ( n829 & n834 ) ;
  assign n842 = ~n840 & n841 ;
  assign n843 = x94 | x95 ;
  assign n844 = x96 | n843 ;
  assign n845 = n746 & ~n844 ;
  assign n846 = ~n747 & n839 ;
  assign n847 = ~n746 & n844 ;
  assign n848 = ( x97 & ~n839 ) | ( x97 & n847 ) | ( ~n839 & n847 ) ;
  assign n849 = ( ~n845 & n846 ) | ( ~n845 & n848 ) | ( n846 & n848 ) ;
  assign n850 = n746 & ~n839 ;
  assign n851 = ( x98 & n846 ) | ( x98 & n850 ) | ( n846 & n850 ) ;
  assign n852 = ( ~x98 & n846 ) | ( ~x98 & n850 ) | ( n846 & n850 ) ;
  assign n853 = ( x98 & ~n851 ) | ( x98 & n852 ) | ( ~n851 & n852 ) ;
  assign n854 = ( ~n664 & n849 ) | ( ~n664 & n853 ) | ( n849 & n853 ) ;
  assign n855 = ( n664 & ~n750 ) | ( n664 & n839 ) | ( ~n750 & n839 ) ;
  assign n856 = n664 & ~n750 ;
  assign n857 = ( n754 & n855 ) | ( n754 & n856 ) | ( n855 & n856 ) ;
  assign n858 = ( ~n754 & n855 ) | ( ~n754 & n856 ) | ( n855 & n856 ) ;
  assign n859 = ( n754 & ~n857 ) | ( n754 & n858 ) | ( ~n857 & n858 ) ;
  assign n860 = ( ~n588 & n854 ) | ( ~n588 & n859 ) | ( n854 & n859 ) ;
  assign n861 = ( n588 & ~n755 ) | ( n588 & n839 ) | ( ~n755 & n839 ) ;
  assign n862 = n588 & ~n755 ;
  assign n863 = ( n759 & n861 ) | ( n759 & n862 ) | ( n861 & n862 ) ;
  assign n864 = ( ~n759 & n861 ) | ( ~n759 & n862 ) | ( n861 & n862 ) ;
  assign n865 = ( n759 & ~n863 ) | ( n759 & n864 ) | ( ~n863 & n864 ) ;
  assign n866 = ( ~n518 & n860 ) | ( ~n518 & n865 ) | ( n860 & n865 ) ;
  assign n867 = ( n518 & ~n760 ) | ( n518 & n839 ) | ( ~n760 & n839 ) ;
  assign n868 = n518 & ~n760 ;
  assign n869 = ( n768 & n867 ) | ( n768 & n868 ) | ( n867 & n868 ) ;
  assign n870 = ( ~n768 & n867 ) | ( ~n768 & n868 ) | ( n867 & n868 ) ;
  assign n871 = ( n768 & ~n869 ) | ( n768 & n870 ) | ( ~n869 & n870 ) ;
  assign n872 = ( ~n454 & n866 ) | ( ~n454 & n871 ) | ( n866 & n871 ) ;
  assign n873 = ( n454 & ~n769 ) | ( n454 & n839 ) | ( ~n769 & n839 ) ;
  assign n874 = n454 & ~n769 ;
  assign n875 = ( n774 & n873 ) | ( n774 & n874 ) | ( n873 & n874 ) ;
  assign n876 = ( ~n774 & n873 ) | ( ~n774 & n874 ) | ( n873 & n874 ) ;
  assign n877 = ( n774 & ~n875 ) | ( n774 & n876 ) | ( ~n875 & n876 ) ;
  assign n878 = ( ~n396 & n872 ) | ( ~n396 & n877 ) | ( n872 & n877 ) ;
  assign n879 = ( n396 & ~n775 ) | ( n396 & n839 ) | ( ~n775 & n839 ) ;
  assign n880 = n396 & ~n775 ;
  assign n881 = ( n780 & n879 ) | ( n780 & n880 ) | ( n879 & n880 ) ;
  assign n882 = ( ~n780 & n879 ) | ( ~n780 & n880 ) | ( n879 & n880 ) ;
  assign n883 = ( n780 & ~n881 ) | ( n780 & n882 ) | ( ~n881 & n882 ) ;
  assign n884 = ( ~n344 & n878 ) | ( ~n344 & n883 ) | ( n878 & n883 ) ;
  assign n885 = ~n344 & n781 ;
  assign n886 = ( ~n344 & n781 ) | ( ~n344 & n839 ) | ( n781 & n839 ) ;
  assign n887 = ( ~n786 & n885 ) | ( ~n786 & n886 ) | ( n885 & n886 ) ;
  assign n888 = ( n786 & n885 ) | ( n786 & n886 ) | ( n885 & n886 ) ;
  assign n889 = ( n786 & n887 ) | ( n786 & ~n888 ) | ( n887 & ~n888 ) ;
  assign n890 = ( ~n298 & n884 ) | ( ~n298 & n889 ) | ( n884 & n889 ) ;
  assign n891 = n298 & ~n787 ;
  assign n892 = ( n298 & ~n787 ) | ( n298 & n839 ) | ( ~n787 & n839 ) ;
  assign n893 = ( n792 & n891 ) | ( n792 & n892 ) | ( n891 & n892 ) ;
  assign n894 = ( ~n792 & n891 ) | ( ~n792 & n892 ) | ( n891 & n892 ) ;
  assign n895 = ( n792 & ~n893 ) | ( n792 & n894 ) | ( ~n893 & n894 ) ;
  assign n896 = ( ~n258 & n890 ) | ( ~n258 & n895 ) | ( n890 & n895 ) ;
  assign n897 = ( n258 & ~n793 ) | ( n258 & n839 ) | ( ~n793 & n839 ) ;
  assign n898 = n258 & ~n793 ;
  assign n899 = ( n798 & n897 ) | ( n798 & n898 ) | ( n897 & n898 ) ;
  assign n900 = ( ~n798 & n897 ) | ( ~n798 & n898 ) | ( n897 & n898 ) ;
  assign n901 = ( n798 & ~n899 ) | ( n798 & n900 ) | ( ~n899 & n900 ) ;
  assign n902 = ( ~n225 & n896 ) | ( ~n225 & n901 ) | ( n896 & n901 ) ;
  assign n903 = ~n225 & n799 ;
  assign n904 = ( ~n225 & n799 ) | ( ~n225 & n839 ) | ( n799 & n839 ) ;
  assign n905 = ( ~n804 & n903 ) | ( ~n804 & n904 ) | ( n903 & n904 ) ;
  assign n906 = ( n804 & n903 ) | ( n804 & n904 ) | ( n903 & n904 ) ;
  assign n907 = ( n804 & n905 ) | ( n804 & ~n906 ) | ( n905 & ~n906 ) ;
  assign n908 = ( ~n197 & n902 ) | ( ~n197 & n907 ) | ( n902 & n907 ) ;
  assign n909 = ( n197 & ~n805 ) | ( n197 & n839 ) | ( ~n805 & n839 ) ;
  assign n910 = n197 & ~n805 ;
  assign n911 = ( n810 & n909 ) | ( n810 & n910 ) | ( n909 & n910 ) ;
  assign n912 = ( ~n810 & n909 ) | ( ~n810 & n910 ) | ( n909 & n910 ) ;
  assign n913 = ( n810 & ~n911 ) | ( n810 & n912 ) | ( ~n911 & n912 ) ;
  assign n914 = ( ~n170 & n908 ) | ( ~n170 & n913 ) | ( n908 & n913 ) ;
  assign n915 = n170 & ~n811 ;
  assign n916 = ( n170 & ~n811 ) | ( n170 & n839 ) | ( ~n811 & n839 ) ;
  assign n917 = ( n816 & n915 ) | ( n816 & n916 ) | ( n915 & n916 ) ;
  assign n918 = ( ~n816 & n915 ) | ( ~n816 & n916 ) | ( n915 & n916 ) ;
  assign n919 = ( n816 & ~n917 ) | ( n816 & n918 ) | ( ~n917 & n918 ) ;
  assign n920 = ( ~n142 & n914 ) | ( ~n142 & n919 ) | ( n914 & n919 ) ;
  assign n921 = ( n142 & ~n817 ) | ( n142 & n839 ) | ( ~n817 & n839 ) ;
  assign n922 = n142 & ~n817 ;
  assign n923 = ( n822 & n921 ) | ( n822 & n922 ) | ( n921 & n922 ) ;
  assign n924 = ( ~n822 & n921 ) | ( ~n822 & n922 ) | ( n921 & n922 ) ;
  assign n925 = ( n822 & ~n923 ) | ( n822 & n924 ) | ( ~n923 & n924 ) ;
  assign n926 = ( ~n132 & n920 ) | ( ~n132 & n925 ) | ( n920 & n925 ) ;
  assign n927 = ( n132 & ~n823 ) | ( n132 & n839 ) | ( ~n823 & n839 ) ;
  assign n928 = n132 & ~n823 ;
  assign n929 = ( n828 & n927 ) | ( n828 & n928 ) | ( n927 & n928 ) ;
  assign n930 = ( ~n828 & n927 ) | ( ~n828 & n928 ) | ( n927 & n928 ) ;
  assign n931 = ( n828 & ~n929 ) | ( n828 & n930 ) | ( ~n929 & n930 ) ;
  assign n932 = ( ~n131 & n926 ) | ( ~n131 & n931 ) | ( n926 & n931 ) ;
  assign n933 = n842 | n932 ;
  assign n934 = ~n843 & n933 ;
  assign n935 = ( ~x95 & n839 ) | ( ~x95 & n933 ) | ( n839 & n933 ) ;
  assign n936 = x95 & n933 ;
  assign n937 = ( x95 & ~n839 ) | ( x95 & n933 ) | ( ~n839 & n933 ) ;
  assign n938 = x92 | x93 ;
  assign n939 = x94 | n938 ;
  assign n940 = ( ~n936 & n937 ) | ( ~n936 & n939 ) | ( n937 & n939 ) ;
  assign n941 = ( n934 & ~n935 ) | ( n934 & n940 ) | ( ~n935 & n940 ) ;
  assign n942 = n839 & ~n933 ;
  assign n943 = ( x96 & n934 ) | ( x96 & n942 ) | ( n934 & n942 ) ;
  assign n944 = ( ~x96 & n934 ) | ( ~x96 & n942 ) | ( n934 & n942 ) ;
  assign n945 = ( x96 & ~n943 ) | ( x96 & n944 ) | ( ~n943 & n944 ) ;
  assign n946 = ( ~n746 & n941 ) | ( ~n746 & n945 ) | ( n941 & n945 ) ;
  assign n947 = ~n746 & n839 ;
  assign n948 = ( n850 & n933 ) | ( n850 & n947 ) | ( n933 & n947 ) ;
  assign n949 = ( x97 & n944 ) | ( x97 & n948 ) | ( n944 & n948 ) ;
  assign n950 = ( ~x97 & n944 ) | ( ~x97 & n948 ) | ( n944 & n948 ) ;
  assign n951 = ( x97 & ~n949 ) | ( x97 & n950 ) | ( ~n949 & n950 ) ;
  assign n952 = ( ~n664 & n946 ) | ( ~n664 & n951 ) | ( n946 & n951 ) ;
  assign n953 = ( n664 & ~n849 ) | ( n664 & n933 ) | ( ~n849 & n933 ) ;
  assign n954 = n664 & ~n849 ;
  assign n955 = ( n853 & n953 ) | ( n853 & n954 ) | ( n953 & n954 ) ;
  assign n956 = ( ~n853 & n953 ) | ( ~n853 & n954 ) | ( n953 & n954 ) ;
  assign n957 = ( n853 & ~n955 ) | ( n853 & n956 ) | ( ~n955 & n956 ) ;
  assign n958 = ( ~n588 & n952 ) | ( ~n588 & n957 ) | ( n952 & n957 ) ;
  assign n959 = ( n588 & ~n854 ) | ( n588 & n933 ) | ( ~n854 & n933 ) ;
  assign n960 = n588 & ~n854 ;
  assign n961 = ( n859 & n959 ) | ( n859 & n960 ) | ( n959 & n960 ) ;
  assign n962 = ( ~n859 & n959 ) | ( ~n859 & n960 ) | ( n959 & n960 ) ;
  assign n963 = ( n859 & ~n961 ) | ( n859 & n962 ) | ( ~n961 & n962 ) ;
  assign n964 = ( ~n518 & n958 ) | ( ~n518 & n963 ) | ( n958 & n963 ) ;
  assign n965 = ( n518 & ~n860 ) | ( n518 & n933 ) | ( ~n860 & n933 ) ;
  assign n966 = n518 & ~n860 ;
  assign n967 = ( n865 & n965 ) | ( n865 & n966 ) | ( n965 & n966 ) ;
  assign n968 = ( ~n865 & n965 ) | ( ~n865 & n966 ) | ( n965 & n966 ) ;
  assign n969 = ( n865 & ~n967 ) | ( n865 & n968 ) | ( ~n967 & n968 ) ;
  assign n970 = ( ~n454 & n964 ) | ( ~n454 & n969 ) | ( n964 & n969 ) ;
  assign n971 = ( n454 & ~n866 ) | ( n454 & n933 ) | ( ~n866 & n933 ) ;
  assign n972 = n454 & ~n866 ;
  assign n973 = ( n871 & n971 ) | ( n871 & n972 ) | ( n971 & n972 ) ;
  assign n974 = ( ~n871 & n971 ) | ( ~n871 & n972 ) | ( n971 & n972 ) ;
  assign n975 = ( n871 & ~n973 ) | ( n871 & n974 ) | ( ~n973 & n974 ) ;
  assign n976 = ( ~n396 & n970 ) | ( ~n396 & n975 ) | ( n970 & n975 ) ;
  assign n977 = ( n396 & ~n872 ) | ( n396 & n933 ) | ( ~n872 & n933 ) ;
  assign n978 = n396 & ~n872 ;
  assign n979 = ( n877 & n977 ) | ( n877 & n978 ) | ( n977 & n978 ) ;
  assign n980 = ( ~n877 & n977 ) | ( ~n877 & n978 ) | ( n977 & n978 ) ;
  assign n981 = ( n877 & ~n979 ) | ( n877 & n980 ) | ( ~n979 & n980 ) ;
  assign n982 = ( ~n344 & n976 ) | ( ~n344 & n981 ) | ( n976 & n981 ) ;
  assign n983 = ( n344 & ~n878 ) | ( n344 & n933 ) | ( ~n878 & n933 ) ;
  assign n984 = n344 & ~n878 ;
  assign n985 = ( n883 & n983 ) | ( n883 & n984 ) | ( n983 & n984 ) ;
  assign n986 = ( ~n883 & n983 ) | ( ~n883 & n984 ) | ( n983 & n984 ) ;
  assign n987 = ( n883 & ~n985 ) | ( n883 & n986 ) | ( ~n985 & n986 ) ;
  assign n988 = ( ~n298 & n982 ) | ( ~n298 & n987 ) | ( n982 & n987 ) ;
  assign n989 = n298 & ~n884 ;
  assign n990 = ( n298 & ~n884 ) | ( n298 & n933 ) | ( ~n884 & n933 ) ;
  assign n991 = ( n889 & n989 ) | ( n889 & n990 ) | ( n989 & n990 ) ;
  assign n992 = ( ~n889 & n989 ) | ( ~n889 & n990 ) | ( n989 & n990 ) ;
  assign n993 = ( n889 & ~n991 ) | ( n889 & n992 ) | ( ~n991 & n992 ) ;
  assign n994 = ( ~n258 & n988 ) | ( ~n258 & n993 ) | ( n988 & n993 ) ;
  assign n995 = ~n258 & n890 ;
  assign n996 = ( ~n258 & n890 ) | ( ~n258 & n933 ) | ( n890 & n933 ) ;
  assign n997 = ( ~n895 & n995 ) | ( ~n895 & n996 ) | ( n995 & n996 ) ;
  assign n998 = ( n895 & n995 ) | ( n895 & n996 ) | ( n995 & n996 ) ;
  assign n999 = ( n895 & n997 ) | ( n895 & ~n998 ) | ( n997 & ~n998 ) ;
  assign n1000 = ( ~n225 & n994 ) | ( ~n225 & n999 ) | ( n994 & n999 ) ;
  assign n1001 = ( n225 & ~n896 ) | ( n225 & n933 ) | ( ~n896 & n933 ) ;
  assign n1002 = n225 & ~n896 ;
  assign n1003 = ( n901 & n1001 ) | ( n901 & n1002 ) | ( n1001 & n1002 ) ;
  assign n1004 = ( ~n901 & n1001 ) | ( ~n901 & n1002 ) | ( n1001 & n1002 ) ;
  assign n1005 = ( n901 & ~n1003 ) | ( n901 & n1004 ) | ( ~n1003 & n1004 ) ;
  assign n1006 = ( ~n197 & n1000 ) | ( ~n197 & n1005 ) | ( n1000 & n1005 ) ;
  assign n1007 = ~n197 & n902 ;
  assign n1008 = ( ~n197 & n902 ) | ( ~n197 & n933 ) | ( n902 & n933 ) ;
  assign n1009 = ( n907 & n1007 ) | ( n907 & n1008 ) | ( n1007 & n1008 ) ;
  assign n1010 = ( ~n907 & n1007 ) | ( ~n907 & n1008 ) | ( n1007 & n1008 ) ;
  assign n1011 = ( n907 & ~n1009 ) | ( n907 & n1010 ) | ( ~n1009 & n1010 ) ;
  assign n1012 = ( ~n170 & n1006 ) | ( ~n170 & n1011 ) | ( n1006 & n1011 ) ;
  assign n1013 = ~n170 & n908 ;
  assign n1014 = ( ~n170 & n908 ) | ( ~n170 & n933 ) | ( n908 & n933 ) ;
  assign n1015 = ( ~n913 & n1013 ) | ( ~n913 & n1014 ) | ( n1013 & n1014 ) ;
  assign n1016 = ( n913 & n1013 ) | ( n913 & n1014 ) | ( n1013 & n1014 ) ;
  assign n1017 = ( n913 & n1015 ) | ( n913 & ~n1016 ) | ( n1015 & ~n1016 ) ;
  assign n1018 = ( ~n142 & n1012 ) | ( ~n142 & n1017 ) | ( n1012 & n1017 ) ;
  assign n1019 = ( n142 & ~n914 ) | ( n142 & n933 ) | ( ~n914 & n933 ) ;
  assign n1020 = n142 & ~n914 ;
  assign n1021 = ( n919 & n1019 ) | ( n919 & n1020 ) | ( n1019 & n1020 ) ;
  assign n1022 = ( ~n919 & n1019 ) | ( ~n919 & n1020 ) | ( n1019 & n1020 ) ;
  assign n1023 = ( n919 & ~n1021 ) | ( n919 & n1022 ) | ( ~n1021 & n1022 ) ;
  assign n1024 = ( ~n132 & n1018 ) | ( ~n132 & n1023 ) | ( n1018 & n1023 ) ;
  assign n1025 = n926 & n931 ;
  assign n1026 = n131 | n1025 ;
  assign n1027 = n1024 | n1026 ;
  assign n1028 = ( n132 & ~n920 ) | ( n132 & n933 ) | ( ~n920 & n933 ) ;
  assign n1029 = n132 & ~n920 ;
  assign n1030 = ( n925 & ~n1028 ) | ( n925 & n1029 ) | ( ~n1028 & n1029 ) ;
  assign n1031 = ( n925 & n1028 ) | ( n925 & n1029 ) | ( n1028 & n1029 ) ;
  assign n1032 = ( n1028 & n1030 ) | ( n1028 & ~n1031 ) | ( n1030 & ~n1031 ) ;
  assign n1033 = n1024 & n1032 ;
  assign n1034 = ( ~n131 & n1032 ) | ( ~n131 & n1033 ) | ( n1032 & n1033 ) ;
  assign n1035 = n842 | n931 ;
  assign n1036 = ( n926 & n931 ) | ( n926 & n1035 ) | ( n931 & n1035 ) ;
  assign n1037 = ( n131 & n1025 ) | ( n131 & ~n1036 ) | ( n1025 & ~n1036 ) ;
  assign n1038 = ( n1027 & n1034 ) | ( n1027 & ~n1037 ) | ( n1034 & ~n1037 ) ;
  assign n1039 = ~n1032 & n1037 ;
  assign n1040 = ( n1024 & n1032 ) | ( n1024 & ~n1039 ) | ( n1032 & ~n1039 ) ;
  assign n1041 = ( n131 & n1033 ) | ( n131 & ~n1040 ) | ( n1033 & ~n1040 ) ;
  assign n1042 = x90 | x91 ;
  assign n1043 = x92 | n1042 ;
  assign n1044 = n933 & ~n1043 ;
  assign n1045 = ~n938 & n1038 ;
  assign n1046 = ~n933 & n1043 ;
  assign n1047 = ( x93 & ~n1038 ) | ( x93 & n1046 ) | ( ~n1038 & n1046 ) ;
  assign n1048 = ( ~n1044 & n1045 ) | ( ~n1044 & n1047 ) | ( n1045 & n1047 ) ;
  assign n1049 = n933 & ~n1038 ;
  assign n1050 = ( ~x94 & n1045 ) | ( ~x94 & n1049 ) | ( n1045 & n1049 ) ;
  assign n1051 = ( x94 & n1045 ) | ( x94 & n1049 ) | ( n1045 & n1049 ) ;
  assign n1052 = ( x94 & n1050 ) | ( x94 & ~n1051 ) | ( n1050 & ~n1051 ) ;
  assign n1053 = ( ~n839 & n1048 ) | ( ~n839 & n1052 ) | ( n1048 & n1052 ) ;
  assign n1054 = ~n839 & n933 ;
  assign n1055 = ( n942 & n1038 ) | ( n942 & n1054 ) | ( n1038 & n1054 ) ;
  assign n1056 = ( x95 & n1050 ) | ( x95 & n1055 ) | ( n1050 & n1055 ) ;
  assign n1057 = ( ~x95 & n1050 ) | ( ~x95 & n1055 ) | ( n1050 & n1055 ) ;
  assign n1058 = ( x95 & ~n1056 ) | ( x95 & n1057 ) | ( ~n1056 & n1057 ) ;
  assign n1059 = ( ~n746 & n1053 ) | ( ~n746 & n1058 ) | ( n1053 & n1058 ) ;
  assign n1060 = ( n746 & ~n941 ) | ( n746 & n1038 ) | ( ~n941 & n1038 ) ;
  assign n1061 = n746 & ~n941 ;
  assign n1062 = ( n945 & n1060 ) | ( n945 & n1061 ) | ( n1060 & n1061 ) ;
  assign n1063 = ( ~n945 & n1060 ) | ( ~n945 & n1061 ) | ( n1060 & n1061 ) ;
  assign n1064 = ( n945 & ~n1062 ) | ( n945 & n1063 ) | ( ~n1062 & n1063 ) ;
  assign n1065 = ( ~n664 & n1059 ) | ( ~n664 & n1064 ) | ( n1059 & n1064 ) ;
  assign n1066 = ~n664 & n946 ;
  assign n1067 = ( ~n664 & n946 ) | ( ~n664 & n1038 ) | ( n946 & n1038 ) ;
  assign n1068 = ( ~n951 & n1066 ) | ( ~n951 & n1067 ) | ( n1066 & n1067 ) ;
  assign n1069 = ( n951 & n1066 ) | ( n951 & n1067 ) | ( n1066 & n1067 ) ;
  assign n1070 = ( n951 & n1068 ) | ( n951 & ~n1069 ) | ( n1068 & ~n1069 ) ;
  assign n1071 = ( ~n588 & n1065 ) | ( ~n588 & n1070 ) | ( n1065 & n1070 ) ;
  assign n1072 = ( n588 & ~n952 ) | ( n588 & n1038 ) | ( ~n952 & n1038 ) ;
  assign n1073 = n588 & ~n952 ;
  assign n1074 = ( n957 & n1072 ) | ( n957 & n1073 ) | ( n1072 & n1073 ) ;
  assign n1075 = ( ~n957 & n1072 ) | ( ~n957 & n1073 ) | ( n1072 & n1073 ) ;
  assign n1076 = ( n957 & ~n1074 ) | ( n957 & n1075 ) | ( ~n1074 & n1075 ) ;
  assign n1077 = ( ~n518 & n1071 ) | ( ~n518 & n1076 ) | ( n1071 & n1076 ) ;
  assign n1078 = ~n518 & n958 ;
  assign n1079 = ( ~n518 & n958 ) | ( ~n518 & n1038 ) | ( n958 & n1038 ) ;
  assign n1080 = ( n963 & n1078 ) | ( n963 & n1079 ) | ( n1078 & n1079 ) ;
  assign n1081 = ( ~n963 & n1078 ) | ( ~n963 & n1079 ) | ( n1078 & n1079 ) ;
  assign n1082 = ( n963 & ~n1080 ) | ( n963 & n1081 ) | ( ~n1080 & n1081 ) ;
  assign n1083 = ( ~n454 & n1077 ) | ( ~n454 & n1082 ) | ( n1077 & n1082 ) ;
  assign n1084 = ( n454 & ~n964 ) | ( n454 & n1038 ) | ( ~n964 & n1038 ) ;
  assign n1085 = n454 & ~n964 ;
  assign n1086 = ( n969 & n1084 ) | ( n969 & n1085 ) | ( n1084 & n1085 ) ;
  assign n1087 = ( ~n969 & n1084 ) | ( ~n969 & n1085 ) | ( n1084 & n1085 ) ;
  assign n1088 = ( n969 & ~n1086 ) | ( n969 & n1087 ) | ( ~n1086 & n1087 ) ;
  assign n1089 = ( ~n396 & n1083 ) | ( ~n396 & n1088 ) | ( n1083 & n1088 ) ;
  assign n1090 = ( n396 & ~n970 ) | ( n396 & n1038 ) | ( ~n970 & n1038 ) ;
  assign n1091 = n396 & ~n970 ;
  assign n1092 = ( n975 & n1090 ) | ( n975 & n1091 ) | ( n1090 & n1091 ) ;
  assign n1093 = ( ~n975 & n1090 ) | ( ~n975 & n1091 ) | ( n1090 & n1091 ) ;
  assign n1094 = ( n975 & ~n1092 ) | ( n975 & n1093 ) | ( ~n1092 & n1093 ) ;
  assign n1095 = ( ~n344 & n1089 ) | ( ~n344 & n1094 ) | ( n1089 & n1094 ) ;
  assign n1096 = ~n344 & n976 ;
  assign n1097 = ( ~n344 & n976 ) | ( ~n344 & n1038 ) | ( n976 & n1038 ) ;
  assign n1098 = ( n981 & n1096 ) | ( n981 & n1097 ) | ( n1096 & n1097 ) ;
  assign n1099 = ( ~n981 & n1096 ) | ( ~n981 & n1097 ) | ( n1096 & n1097 ) ;
  assign n1100 = ( n981 & ~n1098 ) | ( n981 & n1099 ) | ( ~n1098 & n1099 ) ;
  assign n1101 = ( ~n298 & n1095 ) | ( ~n298 & n1100 ) | ( n1095 & n1100 ) ;
  assign n1102 = ~n298 & n982 ;
  assign n1103 = ( ~n298 & n982 ) | ( ~n298 & n1038 ) | ( n982 & n1038 ) ;
  assign n1104 = ( ~n987 & n1102 ) | ( ~n987 & n1103 ) | ( n1102 & n1103 ) ;
  assign n1105 = ( n987 & n1102 ) | ( n987 & n1103 ) | ( n1102 & n1103 ) ;
  assign n1106 = ( n987 & n1104 ) | ( n987 & ~n1105 ) | ( n1104 & ~n1105 ) ;
  assign n1107 = ( ~n258 & n1101 ) | ( ~n258 & n1106 ) | ( n1101 & n1106 ) ;
  assign n1108 = ( n258 & ~n988 ) | ( n258 & n1038 ) | ( ~n988 & n1038 ) ;
  assign n1109 = n258 & ~n988 ;
  assign n1110 = ( n993 & n1108 ) | ( n993 & n1109 ) | ( n1108 & n1109 ) ;
  assign n1111 = ( ~n993 & n1108 ) | ( ~n993 & n1109 ) | ( n1108 & n1109 ) ;
  assign n1112 = ( n993 & ~n1110 ) | ( n993 & n1111 ) | ( ~n1110 & n1111 ) ;
  assign n1113 = ( ~n225 & n1107 ) | ( ~n225 & n1112 ) | ( n1107 & n1112 ) ;
  assign n1114 = ( n225 & ~n994 ) | ( n225 & n1038 ) | ( ~n994 & n1038 ) ;
  assign n1115 = n225 & ~n994 ;
  assign n1116 = ( n999 & n1114 ) | ( n999 & n1115 ) | ( n1114 & n1115 ) ;
  assign n1117 = ( ~n999 & n1114 ) | ( ~n999 & n1115 ) | ( n1114 & n1115 ) ;
  assign n1118 = ( n999 & ~n1116 ) | ( n999 & n1117 ) | ( ~n1116 & n1117 ) ;
  assign n1119 = ( ~n197 & n1113 ) | ( ~n197 & n1118 ) | ( n1113 & n1118 ) ;
  assign n1120 = ~n197 & n1000 ;
  assign n1121 = ( ~n197 & n1000 ) | ( ~n197 & n1038 ) | ( n1000 & n1038 ) ;
  assign n1122 = ( ~n1005 & n1120 ) | ( ~n1005 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1123 = ( n1005 & n1120 ) | ( n1005 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1124 = ( n1005 & n1122 ) | ( n1005 & ~n1123 ) | ( n1122 & ~n1123 ) ;
  assign n1125 = ( ~n170 & n1119 ) | ( ~n170 & n1124 ) | ( n1119 & n1124 ) ;
  assign n1126 = ( n170 & ~n1006 ) | ( n170 & n1038 ) | ( ~n1006 & n1038 ) ;
  assign n1127 = n170 & ~n1006 ;
  assign n1128 = ( n1011 & n1126 ) | ( n1011 & n1127 ) | ( n1126 & n1127 ) ;
  assign n1129 = ( ~n1011 & n1126 ) | ( ~n1011 & n1127 ) | ( n1126 & n1127 ) ;
  assign n1130 = ( n1011 & ~n1128 ) | ( n1011 & n1129 ) | ( ~n1128 & n1129 ) ;
  assign n1131 = ( ~n142 & n1125 ) | ( ~n142 & n1130 ) | ( n1125 & n1130 ) ;
  assign n1132 = ~n142 & n1012 ;
  assign n1133 = ( ~n142 & n1012 ) | ( ~n142 & n1038 ) | ( n1012 & n1038 ) ;
  assign n1134 = ( n1017 & n1132 ) | ( n1017 & n1133 ) | ( n1132 & n1133 ) ;
  assign n1135 = ( ~n1017 & n1132 ) | ( ~n1017 & n1133 ) | ( n1132 & n1133 ) ;
  assign n1136 = ( n1017 & ~n1134 ) | ( n1017 & n1135 ) | ( ~n1134 & n1135 ) ;
  assign n1137 = ( ~n132 & n1131 ) | ( ~n132 & n1136 ) | ( n1131 & n1136 ) ;
  assign n1138 = ~n926 & n931 ;
  assign n1139 = ( ~n926 & n931 ) | ( ~n926 & n1035 ) | ( n931 & n1035 ) ;
  assign n1140 = ( n1032 & ~n1138 ) | ( n1032 & n1139 ) | ( ~n1138 & n1139 ) ;
  assign n1141 = ( ~n1024 & n1032 ) | ( ~n1024 & n1140 ) | ( n1032 & n1140 ) ;
  assign n1142 = ~n1024 & n1032 ;
  assign n1143 = ( n131 & n1141 ) | ( n131 & ~n1142 ) | ( n1141 & ~n1142 ) ;
  assign n1144 = ~n132 & n1018 ;
  assign n1145 = ( ~n132 & n1018 ) | ( ~n132 & n1038 ) | ( n1018 & n1038 ) ;
  assign n1146 = ( n1023 & n1144 ) | ( n1023 & n1145 ) | ( n1144 & n1145 ) ;
  assign n1147 = ( ~n1023 & n1144 ) | ( ~n1023 & n1145 ) | ( n1144 & n1145 ) ;
  assign n1148 = ( n1023 & ~n1146 ) | ( n1023 & n1147 ) | ( ~n1146 & n1147 ) ;
  assign n1149 = ( ~n1041 & n1143 ) | ( ~n1041 & n1148 ) | ( n1143 & n1148 ) ;
  assign n1150 = ( ~n1041 & n1137 ) | ( ~n1041 & n1149 ) | ( n1137 & n1149 ) ;
  assign n1151 = n1137 & n1148 ;
  assign n1152 = n1137 | n1148 ;
  assign n1153 = ( n1041 & n1137 ) | ( n1041 & n1151 ) | ( n1137 & n1151 ) ;
  assign n1154 = ( n131 & ~n1152 ) | ( n131 & n1153 ) | ( ~n1152 & n1153 ) ;
  assign n1155 = n1143 & ~n1148 ;
  assign n1156 = ( n131 & ~n1137 ) | ( n131 & n1155 ) | ( ~n1137 & n1155 ) ;
  assign n1157 = ( n1151 & ~n1154 ) | ( n1151 & n1156 ) | ( ~n1154 & n1156 ) ;
  assign n1158 = x88 | x89 ;
  assign n1159 = x90 | n1158 ;
  assign n1160 = n1038 & ~n1159 ;
  assign n1161 = ~n1042 & n1150 ;
  assign n1162 = ~n1038 & n1159 ;
  assign n1163 = ( x91 & ~n1150 ) | ( x91 & n1162 ) | ( ~n1150 & n1162 ) ;
  assign n1164 = ( ~n1160 & n1161 ) | ( ~n1160 & n1163 ) | ( n1161 & n1163 ) ;
  assign n1165 = n1038 & ~n1150 ;
  assign n1166 = ( x92 & n1161 ) | ( x92 & n1165 ) | ( n1161 & n1165 ) ;
  assign n1167 = ( ~x92 & n1161 ) | ( ~x92 & n1165 ) | ( n1161 & n1165 ) ;
  assign n1168 = ( x92 & ~n1166 ) | ( x92 & n1167 ) | ( ~n1166 & n1167 ) ;
  assign n1169 = ( ~n933 & n1164 ) | ( ~n933 & n1168 ) | ( n1164 & n1168 ) ;
  assign n1170 = ~n933 & n1038 ;
  assign n1171 = ( n1049 & n1150 ) | ( n1049 & n1170 ) | ( n1150 & n1170 ) ;
  assign n1172 = ( x93 & n1167 ) | ( x93 & n1171 ) | ( n1167 & n1171 ) ;
  assign n1173 = ( ~x93 & n1167 ) | ( ~x93 & n1171 ) | ( n1167 & n1171 ) ;
  assign n1174 = ( x93 & ~n1172 ) | ( x93 & n1173 ) | ( ~n1172 & n1173 ) ;
  assign n1175 = ( ~n839 & n1169 ) | ( ~n839 & n1174 ) | ( n1169 & n1174 ) ;
  assign n1176 = ( n839 & ~n1048 ) | ( n839 & n1150 ) | ( ~n1048 & n1150 ) ;
  assign n1177 = n839 & ~n1048 ;
  assign n1178 = ( n1052 & n1176 ) | ( n1052 & n1177 ) | ( n1176 & n1177 ) ;
  assign n1179 = ( ~n1052 & n1176 ) | ( ~n1052 & n1177 ) | ( n1176 & n1177 ) ;
  assign n1180 = ( n1052 & ~n1178 ) | ( n1052 & n1179 ) | ( ~n1178 & n1179 ) ;
  assign n1181 = ( ~n746 & n1175 ) | ( ~n746 & n1180 ) | ( n1175 & n1180 ) ;
  assign n1182 = n746 & ~n1053 ;
  assign n1183 = ( n746 & ~n1053 ) | ( n746 & n1150 ) | ( ~n1053 & n1150 ) ;
  assign n1184 = ( n1058 & n1182 ) | ( n1058 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1185 = ( ~n1058 & n1182 ) | ( ~n1058 & n1183 ) | ( n1182 & n1183 ) ;
  assign n1186 = ( n1058 & ~n1184 ) | ( n1058 & n1185 ) | ( ~n1184 & n1185 ) ;
  assign n1187 = ( ~n664 & n1181 ) | ( ~n664 & n1186 ) | ( n1181 & n1186 ) ;
  assign n1188 = n664 & ~n1059 ;
  assign n1189 = ( n664 & ~n1059 ) | ( n664 & n1150 ) | ( ~n1059 & n1150 ) ;
  assign n1190 = ( n1064 & n1188 ) | ( n1064 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1191 = ( ~n1064 & n1188 ) | ( ~n1064 & n1189 ) | ( n1188 & n1189 ) ;
  assign n1192 = ( n1064 & ~n1190 ) | ( n1064 & n1191 ) | ( ~n1190 & n1191 ) ;
  assign n1193 = ( ~n588 & n1187 ) | ( ~n588 & n1192 ) | ( n1187 & n1192 ) ;
  assign n1194 = ~n588 & n1065 ;
  assign n1195 = ( ~n588 & n1065 ) | ( ~n588 & n1150 ) | ( n1065 & n1150 ) ;
  assign n1196 = ( n1070 & n1194 ) | ( n1070 & n1195 ) | ( n1194 & n1195 ) ;
  assign n1197 = ( ~n1070 & n1194 ) | ( ~n1070 & n1195 ) | ( n1194 & n1195 ) ;
  assign n1198 = ( n1070 & ~n1196 ) | ( n1070 & n1197 ) | ( ~n1196 & n1197 ) ;
  assign n1199 = ( ~n518 & n1193 ) | ( ~n518 & n1198 ) | ( n1193 & n1198 ) ;
  assign n1200 = ~n518 & n1071 ;
  assign n1201 = ( ~n518 & n1071 ) | ( ~n518 & n1150 ) | ( n1071 & n1150 ) ;
  assign n1202 = ( ~n1076 & n1200 ) | ( ~n1076 & n1201 ) | ( n1200 & n1201 ) ;
  assign n1203 = ( n1076 & n1200 ) | ( n1076 & n1201 ) | ( n1200 & n1201 ) ;
  assign n1204 = ( n1076 & n1202 ) | ( n1076 & ~n1203 ) | ( n1202 & ~n1203 ) ;
  assign n1205 = ( ~n454 & n1199 ) | ( ~n454 & n1204 ) | ( n1199 & n1204 ) ;
  assign n1206 = ~n454 & n1077 ;
  assign n1207 = ( ~n454 & n1077 ) | ( ~n454 & n1150 ) | ( n1077 & n1150 ) ;
  assign n1208 = ( n1082 & n1206 ) | ( n1082 & n1207 ) | ( n1206 & n1207 ) ;
  assign n1209 = ( ~n1082 & n1206 ) | ( ~n1082 & n1207 ) | ( n1206 & n1207 ) ;
  assign n1210 = ( n1082 & ~n1208 ) | ( n1082 & n1209 ) | ( ~n1208 & n1209 ) ;
  assign n1211 = ( ~n396 & n1205 ) | ( ~n396 & n1210 ) | ( n1205 & n1210 ) ;
  assign n1212 = ( n396 & ~n1083 ) | ( n396 & n1150 ) | ( ~n1083 & n1150 ) ;
  assign n1213 = n396 & ~n1083 ;
  assign n1214 = ( n1088 & n1212 ) | ( n1088 & n1213 ) | ( n1212 & n1213 ) ;
  assign n1215 = ( ~n1088 & n1212 ) | ( ~n1088 & n1213 ) | ( n1212 & n1213 ) ;
  assign n1216 = ( n1088 & ~n1214 ) | ( n1088 & n1215 ) | ( ~n1214 & n1215 ) ;
  assign n1217 = ( ~n344 & n1211 ) | ( ~n344 & n1216 ) | ( n1211 & n1216 ) ;
  assign n1218 = ( n344 & ~n1089 ) | ( n344 & n1150 ) | ( ~n1089 & n1150 ) ;
  assign n1219 = n344 & ~n1089 ;
  assign n1220 = ( n1094 & n1218 ) | ( n1094 & n1219 ) | ( n1218 & n1219 ) ;
  assign n1221 = ( ~n1094 & n1218 ) | ( ~n1094 & n1219 ) | ( n1218 & n1219 ) ;
  assign n1222 = ( n1094 & ~n1220 ) | ( n1094 & n1221 ) | ( ~n1220 & n1221 ) ;
  assign n1223 = ( ~n298 & n1217 ) | ( ~n298 & n1222 ) | ( n1217 & n1222 ) ;
  assign n1224 = ( n298 & ~n1095 ) | ( n298 & n1150 ) | ( ~n1095 & n1150 ) ;
  assign n1225 = n298 & ~n1095 ;
  assign n1226 = ( n1100 & n1224 ) | ( n1100 & n1225 ) | ( n1224 & n1225 ) ;
  assign n1227 = ( ~n1100 & n1224 ) | ( ~n1100 & n1225 ) | ( n1224 & n1225 ) ;
  assign n1228 = ( n1100 & ~n1226 ) | ( n1100 & n1227 ) | ( ~n1226 & n1227 ) ;
  assign n1229 = ( ~n258 & n1223 ) | ( ~n258 & n1228 ) | ( n1223 & n1228 ) ;
  assign n1230 = ( n258 & ~n1101 ) | ( n258 & n1150 ) | ( ~n1101 & n1150 ) ;
  assign n1231 = n258 & ~n1101 ;
  assign n1232 = ( n1106 & n1230 ) | ( n1106 & n1231 ) | ( n1230 & n1231 ) ;
  assign n1233 = ( ~n1106 & n1230 ) | ( ~n1106 & n1231 ) | ( n1230 & n1231 ) ;
  assign n1234 = ( n1106 & ~n1232 ) | ( n1106 & n1233 ) | ( ~n1232 & n1233 ) ;
  assign n1235 = ( ~n225 & n1229 ) | ( ~n225 & n1234 ) | ( n1229 & n1234 ) ;
  assign n1236 = ( n225 & ~n1107 ) | ( n225 & n1150 ) | ( ~n1107 & n1150 ) ;
  assign n1237 = n225 & ~n1107 ;
  assign n1238 = ( n1112 & n1236 ) | ( n1112 & n1237 ) | ( n1236 & n1237 ) ;
  assign n1239 = ( ~n1112 & n1236 ) | ( ~n1112 & n1237 ) | ( n1236 & n1237 ) ;
  assign n1240 = ( n1112 & ~n1238 ) | ( n1112 & n1239 ) | ( ~n1238 & n1239 ) ;
  assign n1241 = ( ~n197 & n1235 ) | ( ~n197 & n1240 ) | ( n1235 & n1240 ) ;
  assign n1242 = n197 & ~n1113 ;
  assign n1243 = ( n197 & ~n1113 ) | ( n197 & n1150 ) | ( ~n1113 & n1150 ) ;
  assign n1244 = ( n1118 & n1242 ) | ( n1118 & n1243 ) | ( n1242 & n1243 ) ;
  assign n1245 = ( ~n1118 & n1242 ) | ( ~n1118 & n1243 ) | ( n1242 & n1243 ) ;
  assign n1246 = ( n1118 & ~n1244 ) | ( n1118 & n1245 ) | ( ~n1244 & n1245 ) ;
  assign n1247 = ( ~n170 & n1241 ) | ( ~n170 & n1246 ) | ( n1241 & n1246 ) ;
  assign n1248 = ( n170 & ~n1119 ) | ( n170 & n1150 ) | ( ~n1119 & n1150 ) ;
  assign n1249 = n170 & ~n1119 ;
  assign n1250 = ( n1124 & n1248 ) | ( n1124 & n1249 ) | ( n1248 & n1249 ) ;
  assign n1251 = ( ~n1124 & n1248 ) | ( ~n1124 & n1249 ) | ( n1248 & n1249 ) ;
  assign n1252 = ( n1124 & ~n1250 ) | ( n1124 & n1251 ) | ( ~n1250 & n1251 ) ;
  assign n1253 = ( ~n142 & n1247 ) | ( ~n142 & n1252 ) | ( n1247 & n1252 ) ;
  assign n1254 = ~n142 & n1125 ;
  assign n1255 = ( ~n142 & n1125 ) | ( ~n142 & n1150 ) | ( n1125 & n1150 ) ;
  assign n1256 = ( n1130 & n1254 ) | ( n1130 & n1255 ) | ( n1254 & n1255 ) ;
  assign n1257 = ( ~n1130 & n1254 ) | ( ~n1130 & n1255 ) | ( n1254 & n1255 ) ;
  assign n1258 = ( n1130 & ~n1256 ) | ( n1130 & n1257 ) | ( ~n1256 & n1257 ) ;
  assign n1259 = ( ~n132 & n1253 ) | ( ~n132 & n1258 ) | ( n1253 & n1258 ) ;
  assign n1260 = ( n132 & ~n1131 ) | ( n132 & n1150 ) | ( ~n1131 & n1150 ) ;
  assign n1261 = n132 & ~n1131 ;
  assign n1262 = ( n1136 & n1260 ) | ( n1136 & n1261 ) | ( n1260 & n1261 ) ;
  assign n1263 = ( ~n1136 & n1260 ) | ( ~n1136 & n1261 ) | ( n1260 & n1261 ) ;
  assign n1264 = ( n1136 & ~n1262 ) | ( n1136 & n1263 ) | ( ~n1262 & n1263 ) ;
  assign n1265 = ( ~n131 & n1259 ) | ( ~n131 & n1264 ) | ( n1259 & n1264 ) ;
  assign n1266 = n1157 | n1265 ;
  assign n1267 = ~n1259 & n1264 ;
  assign n1268 = ( n132 & ~n1253 ) | ( n132 & n1266 ) | ( ~n1253 & n1266 ) ;
  assign n1269 = n132 & ~n1253 ;
  assign n1270 = ( n1258 & ~n1268 ) | ( n1258 & n1269 ) | ( ~n1268 & n1269 ) ;
  assign n1271 = ( n1258 & n1268 ) | ( n1258 & n1269 ) | ( n1268 & n1269 ) ;
  assign n1272 = ( n1268 & n1270 ) | ( n1268 & ~n1271 ) | ( n1270 & ~n1271 ) ;
  assign n1273 = ( ~n1259 & n1264 ) | ( ~n1259 & n1266 ) | ( n1264 & n1266 ) ;
  assign n1274 = ( ~n1267 & n1272 ) | ( ~n1267 & n1273 ) | ( n1272 & n1273 ) ;
  assign n1275 = ~n131 & n1274 ;
  assign n1276 = x89 & n1266 ;
  assign n1277 = x86 | x87 ;
  assign n1278 = x88 | n1277 ;
  assign n1279 = ( x89 & n1266 ) | ( x89 & n1278 ) | ( n1266 & n1278 ) ;
  assign n1280 = ( n1150 & n1276 ) | ( n1150 & ~n1279 ) | ( n1276 & ~n1279 ) ;
  assign n1281 = ( ~n1266 & n1276 ) | ( ~n1266 & n1278 ) | ( n1276 & n1278 ) ;
  assign n1282 = ( ~x88 & x89 ) | ( ~x88 & n1266 ) | ( x89 & n1266 ) ;
  assign n1283 = ( ~n1276 & n1281 ) | ( ~n1276 & n1282 ) | ( n1281 & n1282 ) ;
  assign n1284 = ~n1280 & n1283 ;
  assign n1285 = n1150 & ~n1266 ;
  assign n1286 = ~n1158 & n1266 ;
  assign n1287 = ( x90 & n1285 ) | ( x90 & n1286 ) | ( n1285 & n1286 ) ;
  assign n1288 = ( ~x90 & n1285 ) | ( ~x90 & n1286 ) | ( n1285 & n1286 ) ;
  assign n1289 = ( x90 & ~n1287 ) | ( x90 & n1288 ) | ( ~n1287 & n1288 ) ;
  assign n1290 = ( ~n1038 & n1284 ) | ( ~n1038 & n1289 ) | ( n1284 & n1289 ) ;
  assign n1291 = ~n1038 & n1150 ;
  assign n1292 = ( n1165 & n1266 ) | ( n1165 & n1291 ) | ( n1266 & n1291 ) ;
  assign n1293 = ( ~x91 & n1288 ) | ( ~x91 & n1292 ) | ( n1288 & n1292 ) ;
  assign n1294 = ( x91 & n1288 ) | ( x91 & n1292 ) | ( n1288 & n1292 ) ;
  assign n1295 = ( x91 & n1293 ) | ( x91 & ~n1294 ) | ( n1293 & ~n1294 ) ;
  assign n1296 = ( ~n933 & n1290 ) | ( ~n933 & n1295 ) | ( n1290 & n1295 ) ;
  assign n1297 = n933 & ~n1164 ;
  assign n1298 = ( n933 & ~n1164 ) | ( n933 & n1266 ) | ( ~n1164 & n1266 ) ;
  assign n1299 = ( n1168 & n1297 ) | ( n1168 & n1298 ) | ( n1297 & n1298 ) ;
  assign n1300 = ( ~n1168 & n1297 ) | ( ~n1168 & n1298 ) | ( n1297 & n1298 ) ;
  assign n1301 = ( n1168 & ~n1299 ) | ( n1168 & n1300 ) | ( ~n1299 & n1300 ) ;
  assign n1302 = ( ~n839 & n1296 ) | ( ~n839 & n1301 ) | ( n1296 & n1301 ) ;
  assign n1303 = ( n839 & ~n1169 ) | ( n839 & n1266 ) | ( ~n1169 & n1266 ) ;
  assign n1304 = n839 & ~n1169 ;
  assign n1305 = ( n1174 & n1303 ) | ( n1174 & n1304 ) | ( n1303 & n1304 ) ;
  assign n1306 = ( ~n1174 & n1303 ) | ( ~n1174 & n1304 ) | ( n1303 & n1304 ) ;
  assign n1307 = ( n1174 & ~n1305 ) | ( n1174 & n1306 ) | ( ~n1305 & n1306 ) ;
  assign n1308 = ( ~n746 & n1302 ) | ( ~n746 & n1307 ) | ( n1302 & n1307 ) ;
  assign n1309 = ( n746 & ~n1175 ) | ( n746 & n1266 ) | ( ~n1175 & n1266 ) ;
  assign n1310 = n746 & ~n1175 ;
  assign n1311 = ( n1180 & n1309 ) | ( n1180 & n1310 ) | ( n1309 & n1310 ) ;
  assign n1312 = ( ~n1180 & n1309 ) | ( ~n1180 & n1310 ) | ( n1309 & n1310 ) ;
  assign n1313 = ( n1180 & ~n1311 ) | ( n1180 & n1312 ) | ( ~n1311 & n1312 ) ;
  assign n1314 = ( ~n664 & n1308 ) | ( ~n664 & n1313 ) | ( n1308 & n1313 ) ;
  assign n1315 = ~n664 & n1181 ;
  assign n1316 = ( ~n664 & n1181 ) | ( ~n664 & n1266 ) | ( n1181 & n1266 ) ;
  assign n1317 = ( ~n1186 & n1315 ) | ( ~n1186 & n1316 ) | ( n1315 & n1316 ) ;
  assign n1318 = ( n1186 & n1315 ) | ( n1186 & n1316 ) | ( n1315 & n1316 ) ;
  assign n1319 = ( n1186 & n1317 ) | ( n1186 & ~n1318 ) | ( n1317 & ~n1318 ) ;
  assign n1320 = ( ~n588 & n1314 ) | ( ~n588 & n1319 ) | ( n1314 & n1319 ) ;
  assign n1321 = n588 & ~n1187 ;
  assign n1322 = ( n588 & ~n1187 ) | ( n588 & n1266 ) | ( ~n1187 & n1266 ) ;
  assign n1323 = ( ~n1192 & n1321 ) | ( ~n1192 & n1322 ) | ( n1321 & n1322 ) ;
  assign n1324 = ( n1192 & n1321 ) | ( n1192 & n1322 ) | ( n1321 & n1322 ) ;
  assign n1325 = ( n1192 & n1323 ) | ( n1192 & ~n1324 ) | ( n1323 & ~n1324 ) ;
  assign n1326 = ( ~n518 & n1320 ) | ( ~n518 & n1325 ) | ( n1320 & n1325 ) ;
  assign n1327 = ~n518 & n1193 ;
  assign n1328 = ( ~n518 & n1193 ) | ( ~n518 & n1266 ) | ( n1193 & n1266 ) ;
  assign n1329 = ( ~n1198 & n1327 ) | ( ~n1198 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1330 = ( n1198 & n1327 ) | ( n1198 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1331 = ( n1198 & n1329 ) | ( n1198 & ~n1330 ) | ( n1329 & ~n1330 ) ;
  assign n1332 = ( ~n454 & n1326 ) | ( ~n454 & n1331 ) | ( n1326 & n1331 ) ;
  assign n1333 = ( n454 & ~n1199 ) | ( n454 & n1266 ) | ( ~n1199 & n1266 ) ;
  assign n1334 = n454 & ~n1199 ;
  assign n1335 = ( n1204 & n1333 ) | ( n1204 & n1334 ) | ( n1333 & n1334 ) ;
  assign n1336 = ( ~n1204 & n1333 ) | ( ~n1204 & n1334 ) | ( n1333 & n1334 ) ;
  assign n1337 = ( n1204 & ~n1335 ) | ( n1204 & n1336 ) | ( ~n1335 & n1336 ) ;
  assign n1338 = ( ~n396 & n1332 ) | ( ~n396 & n1337 ) | ( n1332 & n1337 ) ;
  assign n1339 = ( n396 & ~n1205 ) | ( n396 & n1266 ) | ( ~n1205 & n1266 ) ;
  assign n1340 = n396 & ~n1205 ;
  assign n1341 = ( n1210 & n1339 ) | ( n1210 & n1340 ) | ( n1339 & n1340 ) ;
  assign n1342 = ( ~n1210 & n1339 ) | ( ~n1210 & n1340 ) | ( n1339 & n1340 ) ;
  assign n1343 = ( n1210 & ~n1341 ) | ( n1210 & n1342 ) | ( ~n1341 & n1342 ) ;
  assign n1344 = ( ~n344 & n1338 ) | ( ~n344 & n1343 ) | ( n1338 & n1343 ) ;
  assign n1345 = n344 & ~n1211 ;
  assign n1346 = ( n344 & ~n1211 ) | ( n344 & n1266 ) | ( ~n1211 & n1266 ) ;
  assign n1347 = ( ~n1216 & n1345 ) | ( ~n1216 & n1346 ) | ( n1345 & n1346 ) ;
  assign n1348 = ( n1216 & n1345 ) | ( n1216 & n1346 ) | ( n1345 & n1346 ) ;
  assign n1349 = ( n1216 & n1347 ) | ( n1216 & ~n1348 ) | ( n1347 & ~n1348 ) ;
  assign n1350 = ( ~n298 & n1344 ) | ( ~n298 & n1349 ) | ( n1344 & n1349 ) ;
  assign n1351 = ( n298 & ~n1217 ) | ( n298 & n1266 ) | ( ~n1217 & n1266 ) ;
  assign n1352 = n298 & ~n1217 ;
  assign n1353 = ( n1222 & n1351 ) | ( n1222 & n1352 ) | ( n1351 & n1352 ) ;
  assign n1354 = ( ~n1222 & n1351 ) | ( ~n1222 & n1352 ) | ( n1351 & n1352 ) ;
  assign n1355 = ( n1222 & ~n1353 ) | ( n1222 & n1354 ) | ( ~n1353 & n1354 ) ;
  assign n1356 = ( ~n258 & n1350 ) | ( ~n258 & n1355 ) | ( n1350 & n1355 ) ;
  assign n1357 = ( n258 & ~n1223 ) | ( n258 & n1266 ) | ( ~n1223 & n1266 ) ;
  assign n1358 = n258 & ~n1223 ;
  assign n1359 = ( n1228 & n1357 ) | ( n1228 & n1358 ) | ( n1357 & n1358 ) ;
  assign n1360 = ( ~n1228 & n1357 ) | ( ~n1228 & n1358 ) | ( n1357 & n1358 ) ;
  assign n1361 = ( n1228 & ~n1359 ) | ( n1228 & n1360 ) | ( ~n1359 & n1360 ) ;
  assign n1362 = ( ~n225 & n1356 ) | ( ~n225 & n1361 ) | ( n1356 & n1361 ) ;
  assign n1363 = ~n225 & n1229 ;
  assign n1364 = ( ~n225 & n1229 ) | ( ~n225 & n1266 ) | ( n1229 & n1266 ) ;
  assign n1365 = ( n1234 & n1363 ) | ( n1234 & n1364 ) | ( n1363 & n1364 ) ;
  assign n1366 = ( ~n1234 & n1363 ) | ( ~n1234 & n1364 ) | ( n1363 & n1364 ) ;
  assign n1367 = ( n1234 & ~n1365 ) | ( n1234 & n1366 ) | ( ~n1365 & n1366 ) ;
  assign n1368 = ( ~n197 & n1362 ) | ( ~n197 & n1367 ) | ( n1362 & n1367 ) ;
  assign n1369 = ( n197 & ~n1235 ) | ( n197 & n1266 ) | ( ~n1235 & n1266 ) ;
  assign n1370 = n197 & ~n1235 ;
  assign n1371 = ( n1240 & n1369 ) | ( n1240 & n1370 ) | ( n1369 & n1370 ) ;
  assign n1372 = ( ~n1240 & n1369 ) | ( ~n1240 & n1370 ) | ( n1369 & n1370 ) ;
  assign n1373 = ( n1240 & ~n1371 ) | ( n1240 & n1372 ) | ( ~n1371 & n1372 ) ;
  assign n1374 = ( ~n170 & n1368 ) | ( ~n170 & n1373 ) | ( n1368 & n1373 ) ;
  assign n1375 = ( n170 & ~n1241 ) | ( n170 & n1266 ) | ( ~n1241 & n1266 ) ;
  assign n1376 = n170 & ~n1241 ;
  assign n1377 = ( n1246 & n1375 ) | ( n1246 & n1376 ) | ( n1375 & n1376 ) ;
  assign n1378 = ( ~n1246 & n1375 ) | ( ~n1246 & n1376 ) | ( n1375 & n1376 ) ;
  assign n1379 = ( n1246 & ~n1377 ) | ( n1246 & n1378 ) | ( ~n1377 & n1378 ) ;
  assign n1380 = ( ~n142 & n1374 ) | ( ~n142 & n1379 ) | ( n1374 & n1379 ) ;
  assign n1381 = ~n142 & n1247 ;
  assign n1382 = ( ~n142 & n1247 ) | ( ~n142 & n1266 ) | ( n1247 & n1266 ) ;
  assign n1383 = ( n1252 & n1381 ) | ( n1252 & n1382 ) | ( n1381 & n1382 ) ;
  assign n1384 = ( ~n1252 & n1381 ) | ( ~n1252 & n1382 ) | ( n1381 & n1382 ) ;
  assign n1385 = ( n1252 & ~n1383 ) | ( n1252 & n1384 ) | ( ~n1383 & n1384 ) ;
  assign n1386 = ( ~n132 & n1380 ) | ( ~n132 & n1385 ) | ( n1380 & n1385 ) ;
  assign n1387 = ( ~n131 & n1275 ) | ( ~n131 & n1386 ) | ( n1275 & n1386 ) ;
  assign n1388 = n1152 & ~n1153 ;
  assign n1389 = n1259 & n1388 ;
  assign n1390 = ( ~n1265 & n1267 ) | ( ~n1265 & n1389 ) | ( n1267 & n1389 ) ;
  assign n1391 = n1272 & n1386 ;
  assign n1392 = ( ~n1387 & n1390 ) | ( ~n1387 & n1391 ) | ( n1390 & n1391 ) ;
  assign n1393 = n1387 | n1392 ;
  assign n1394 = ( n131 & n1272 ) | ( n131 & n1390 ) | ( n1272 & n1390 ) ;
  assign n1395 = ( n1272 & n1386 ) | ( n1272 & n1394 ) | ( n1386 & n1394 ) ;
  assign n1396 = ~n1391 & n1395 ;
  assign n1397 = x87 & ~n1393 ;
  assign n1398 = ( ~x87 & n1387 ) | ( ~x87 & n1392 ) | ( n1387 & n1392 ) ;
  assign n1399 = x84 | x85 ;
  assign n1400 = x86 | n1399 ;
  assign n1401 = ~n1266 & n1400 ;
  assign n1402 = n1398 | n1401 ;
  assign n1403 = n1266 & ~n1400 ;
  assign n1404 = ~x86 & n1398 ;
  assign n1405 = ( n1398 & n1403 ) | ( n1398 & ~n1404 ) | ( n1403 & ~n1404 ) ;
  assign n1406 = ( n1397 & n1402 ) | ( n1397 & ~n1405 ) | ( n1402 & ~n1405 ) ;
  assign n1407 = n1266 & ~n1393 ;
  assign n1408 = ( x88 & n1404 ) | ( x88 & n1407 ) | ( n1404 & n1407 ) ;
  assign n1409 = ( ~x88 & n1404 ) | ( ~x88 & n1407 ) | ( n1404 & n1407 ) ;
  assign n1410 = ( x88 & ~n1408 ) | ( x88 & n1409 ) | ( ~n1408 & n1409 ) ;
  assign n1411 = ( ~n1150 & n1406 ) | ( ~n1150 & n1410 ) | ( n1406 & n1410 ) ;
  assign n1412 = ~n1150 & n1266 ;
  assign n1413 = ( n1285 & n1393 ) | ( n1285 & n1412 ) | ( n1393 & n1412 ) ;
  assign n1414 = ( x89 & n1409 ) | ( x89 & n1413 ) | ( n1409 & n1413 ) ;
  assign n1415 = ( ~x89 & n1409 ) | ( ~x89 & n1413 ) | ( n1409 & n1413 ) ;
  assign n1416 = ( x89 & ~n1414 ) | ( x89 & n1415 ) | ( ~n1414 & n1415 ) ;
  assign n1417 = ( ~n1038 & n1411 ) | ( ~n1038 & n1416 ) | ( n1411 & n1416 ) ;
  assign n1418 = ( n1038 & ~n1284 ) | ( n1038 & n1393 ) | ( ~n1284 & n1393 ) ;
  assign n1419 = n1038 & ~n1284 ;
  assign n1420 = ( n1289 & n1418 ) | ( n1289 & n1419 ) | ( n1418 & n1419 ) ;
  assign n1421 = ( ~n1289 & n1418 ) | ( ~n1289 & n1419 ) | ( n1418 & n1419 ) ;
  assign n1422 = ( n1289 & ~n1420 ) | ( n1289 & n1421 ) | ( ~n1420 & n1421 ) ;
  assign n1423 = ( ~n933 & n1417 ) | ( ~n933 & n1422 ) | ( n1417 & n1422 ) ;
  assign n1424 = ( n933 & ~n1290 ) | ( n933 & n1393 ) | ( ~n1290 & n1393 ) ;
  assign n1425 = n933 & ~n1290 ;
  assign n1426 = ( n1295 & n1424 ) | ( n1295 & n1425 ) | ( n1424 & n1425 ) ;
  assign n1427 = ( ~n1295 & n1424 ) | ( ~n1295 & n1425 ) | ( n1424 & n1425 ) ;
  assign n1428 = ( n1295 & ~n1426 ) | ( n1295 & n1427 ) | ( ~n1426 & n1427 ) ;
  assign n1429 = ( ~n839 & n1423 ) | ( ~n839 & n1428 ) | ( n1423 & n1428 ) ;
  assign n1430 = ( n839 & ~n1296 ) | ( n839 & n1393 ) | ( ~n1296 & n1393 ) ;
  assign n1431 = n839 & ~n1296 ;
  assign n1432 = ( n1301 & n1430 ) | ( n1301 & n1431 ) | ( n1430 & n1431 ) ;
  assign n1433 = ( ~n1301 & n1430 ) | ( ~n1301 & n1431 ) | ( n1430 & n1431 ) ;
  assign n1434 = ( n1301 & ~n1432 ) | ( n1301 & n1433 ) | ( ~n1432 & n1433 ) ;
  assign n1435 = ( ~n746 & n1429 ) | ( ~n746 & n1434 ) | ( n1429 & n1434 ) ;
  assign n1436 = ( n746 & ~n1302 ) | ( n746 & n1393 ) | ( ~n1302 & n1393 ) ;
  assign n1437 = n746 & ~n1302 ;
  assign n1438 = ( n1307 & n1436 ) | ( n1307 & n1437 ) | ( n1436 & n1437 ) ;
  assign n1439 = ( ~n1307 & n1436 ) | ( ~n1307 & n1437 ) | ( n1436 & n1437 ) ;
  assign n1440 = ( n1307 & ~n1438 ) | ( n1307 & n1439 ) | ( ~n1438 & n1439 ) ;
  assign n1441 = ( ~n664 & n1435 ) | ( ~n664 & n1440 ) | ( n1435 & n1440 ) ;
  assign n1442 = n664 & ~n1308 ;
  assign n1443 = ( n664 & ~n1308 ) | ( n664 & n1393 ) | ( ~n1308 & n1393 ) ;
  assign n1444 = ( n1313 & n1442 ) | ( n1313 & n1443 ) | ( n1442 & n1443 ) ;
  assign n1445 = ( ~n1313 & n1442 ) | ( ~n1313 & n1443 ) | ( n1442 & n1443 ) ;
  assign n1446 = ( n1313 & ~n1444 ) | ( n1313 & n1445 ) | ( ~n1444 & n1445 ) ;
  assign n1447 = ( ~n588 & n1441 ) | ( ~n588 & n1446 ) | ( n1441 & n1446 ) ;
  assign n1448 = ( n588 & ~n1314 ) | ( n588 & n1393 ) | ( ~n1314 & n1393 ) ;
  assign n1449 = n588 & ~n1314 ;
  assign n1450 = ( n1319 & n1448 ) | ( n1319 & n1449 ) | ( n1448 & n1449 ) ;
  assign n1451 = ( ~n1319 & n1448 ) | ( ~n1319 & n1449 ) | ( n1448 & n1449 ) ;
  assign n1452 = ( n1319 & ~n1450 ) | ( n1319 & n1451 ) | ( ~n1450 & n1451 ) ;
  assign n1453 = ( ~n518 & n1447 ) | ( ~n518 & n1452 ) | ( n1447 & n1452 ) ;
  assign n1454 = ( n518 & ~n1320 ) | ( n518 & n1393 ) | ( ~n1320 & n1393 ) ;
  assign n1455 = n518 & ~n1320 ;
  assign n1456 = ( n1325 & n1454 ) | ( n1325 & n1455 ) | ( n1454 & n1455 ) ;
  assign n1457 = ( ~n1325 & n1454 ) | ( ~n1325 & n1455 ) | ( n1454 & n1455 ) ;
  assign n1458 = ( n1325 & ~n1456 ) | ( n1325 & n1457 ) | ( ~n1456 & n1457 ) ;
  assign n1459 = ( ~n454 & n1453 ) | ( ~n454 & n1458 ) | ( n1453 & n1458 ) ;
  assign n1460 = n454 & ~n1326 ;
  assign n1461 = ( n454 & ~n1326 ) | ( n454 & n1393 ) | ( ~n1326 & n1393 ) ;
  assign n1462 = ( ~n1331 & n1460 ) | ( ~n1331 & n1461 ) | ( n1460 & n1461 ) ;
  assign n1463 = ( n1331 & n1460 ) | ( n1331 & n1461 ) | ( n1460 & n1461 ) ;
  assign n1464 = ( n1331 & n1462 ) | ( n1331 & ~n1463 ) | ( n1462 & ~n1463 ) ;
  assign n1465 = ( ~n396 & n1459 ) | ( ~n396 & n1464 ) | ( n1459 & n1464 ) ;
  assign n1466 = ~n396 & n1332 ;
  assign n1467 = ( ~n396 & n1332 ) | ( ~n396 & n1393 ) | ( n1332 & n1393 ) ;
  assign n1468 = ( ~n1337 & n1466 ) | ( ~n1337 & n1467 ) | ( n1466 & n1467 ) ;
  assign n1469 = ( n1337 & n1466 ) | ( n1337 & n1467 ) | ( n1466 & n1467 ) ;
  assign n1470 = ( n1337 & n1468 ) | ( n1337 & ~n1469 ) | ( n1468 & ~n1469 ) ;
  assign n1471 = ( ~n344 & n1465 ) | ( ~n344 & n1470 ) | ( n1465 & n1470 ) ;
  assign n1472 = ( n344 & ~n1338 ) | ( n344 & n1393 ) | ( ~n1338 & n1393 ) ;
  assign n1473 = n344 & ~n1338 ;
  assign n1474 = ( n1343 & n1472 ) | ( n1343 & n1473 ) | ( n1472 & n1473 ) ;
  assign n1475 = ( ~n1343 & n1472 ) | ( ~n1343 & n1473 ) | ( n1472 & n1473 ) ;
  assign n1476 = ( n1343 & ~n1474 ) | ( n1343 & n1475 ) | ( ~n1474 & n1475 ) ;
  assign n1477 = ( ~n298 & n1471 ) | ( ~n298 & n1476 ) | ( n1471 & n1476 ) ;
  assign n1478 = ( n298 & ~n1344 ) | ( n298 & n1393 ) | ( ~n1344 & n1393 ) ;
  assign n1479 = n298 & ~n1344 ;
  assign n1480 = ( n1349 & n1478 ) | ( n1349 & n1479 ) | ( n1478 & n1479 ) ;
  assign n1481 = ( ~n1349 & n1478 ) | ( ~n1349 & n1479 ) | ( n1478 & n1479 ) ;
  assign n1482 = ( n1349 & ~n1480 ) | ( n1349 & n1481 ) | ( ~n1480 & n1481 ) ;
  assign n1483 = ( ~n258 & n1477 ) | ( ~n258 & n1482 ) | ( n1477 & n1482 ) ;
  assign n1484 = ( n258 & ~n1350 ) | ( n258 & n1393 ) | ( ~n1350 & n1393 ) ;
  assign n1485 = n258 & ~n1350 ;
  assign n1486 = ( n1355 & n1484 ) | ( n1355 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1487 = ( ~n1355 & n1484 ) | ( ~n1355 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1488 = ( n1355 & ~n1486 ) | ( n1355 & n1487 ) | ( ~n1486 & n1487 ) ;
  assign n1489 = ( ~n225 & n1483 ) | ( ~n225 & n1488 ) | ( n1483 & n1488 ) ;
  assign n1490 = ~n225 & n1356 ;
  assign n1491 = ( ~n225 & n1356 ) | ( ~n225 & n1393 ) | ( n1356 & n1393 ) ;
  assign n1492 = ( n1361 & n1490 ) | ( n1361 & n1491 ) | ( n1490 & n1491 ) ;
  assign n1493 = ( ~n1361 & n1490 ) | ( ~n1361 & n1491 ) | ( n1490 & n1491 ) ;
  assign n1494 = ( n1361 & ~n1492 ) | ( n1361 & n1493 ) | ( ~n1492 & n1493 ) ;
  assign n1495 = ( ~n197 & n1489 ) | ( ~n197 & n1494 ) | ( n1489 & n1494 ) ;
  assign n1496 = ~n197 & n1362 ;
  assign n1497 = ( ~n197 & n1362 ) | ( ~n197 & n1393 ) | ( n1362 & n1393 ) ;
  assign n1498 = ( n1367 & n1496 ) | ( n1367 & n1497 ) | ( n1496 & n1497 ) ;
  assign n1499 = ( ~n1367 & n1496 ) | ( ~n1367 & n1497 ) | ( n1496 & n1497 ) ;
  assign n1500 = ( n1367 & ~n1498 ) | ( n1367 & n1499 ) | ( ~n1498 & n1499 ) ;
  assign n1501 = ( ~n170 & n1495 ) | ( ~n170 & n1500 ) | ( n1495 & n1500 ) ;
  assign n1502 = ( n170 & ~n1368 ) | ( n170 & n1393 ) | ( ~n1368 & n1393 ) ;
  assign n1503 = n170 & ~n1368 ;
  assign n1504 = ( n1373 & n1502 ) | ( n1373 & n1503 ) | ( n1502 & n1503 ) ;
  assign n1505 = ( ~n1373 & n1502 ) | ( ~n1373 & n1503 ) | ( n1502 & n1503 ) ;
  assign n1506 = ( n1373 & ~n1504 ) | ( n1373 & n1505 ) | ( ~n1504 & n1505 ) ;
  assign n1507 = ( ~n142 & n1501 ) | ( ~n142 & n1506 ) | ( n1501 & n1506 ) ;
  assign n1508 = n142 & ~n1374 ;
  assign n1509 = ( n142 & ~n1374 ) | ( n142 & n1393 ) | ( ~n1374 & n1393 ) ;
  assign n1510 = ( n1379 & n1508 ) | ( n1379 & n1509 ) | ( n1508 & n1509 ) ;
  assign n1511 = ( ~n1379 & n1508 ) | ( ~n1379 & n1509 ) | ( n1508 & n1509 ) ;
  assign n1512 = ( n1379 & ~n1510 ) | ( n1379 & n1511 ) | ( ~n1510 & n1511 ) ;
  assign n1513 = ( ~n132 & n1507 ) | ( ~n132 & n1512 ) | ( n1507 & n1512 ) ;
  assign n1514 = ( n132 & ~n1380 ) | ( n132 & n1393 ) | ( ~n1380 & n1393 ) ;
  assign n1515 = n132 & ~n1380 ;
  assign n1516 = ( n1385 & n1514 ) | ( n1385 & n1515 ) | ( n1514 & n1515 ) ;
  assign n1517 = ( ~n1385 & n1514 ) | ( ~n1385 & n1515 ) | ( n1514 & n1515 ) ;
  assign n1518 = ( n1385 & ~n1516 ) | ( n1385 & n1517 ) | ( ~n1516 & n1517 ) ;
  assign n1519 = ( ~n131 & n1513 ) | ( ~n131 & n1518 ) | ( n1513 & n1518 ) ;
  assign n1520 = n1396 | n1519 ;
  assign n1521 = n1272 | n1386 ;
  assign n1522 = ( n1387 & n1391 ) | ( n1387 & ~n1521 ) | ( n1391 & ~n1521 ) ;
  assign n1523 = n1520 | n1522 ;
  assign n1524 = ~n1513 & n1518 ;
  assign n1525 = ( n1396 & n1513 ) | ( n1396 & n1518 ) | ( n1513 & n1518 ) ;
  assign n1526 = ( ~n1519 & n1524 ) | ( ~n1519 & n1525 ) | ( n1524 & n1525 ) ;
  assign n1527 = ( n132 & ~n1507 ) | ( n132 & n1523 ) | ( ~n1507 & n1523 ) ;
  assign n1528 = n132 & ~n1507 ;
  assign n1529 = ( n1512 & ~n1527 ) | ( n1512 & n1528 ) | ( ~n1527 & n1528 ) ;
  assign n1530 = ( n1512 & n1527 ) | ( n1512 & n1528 ) | ( n1527 & n1528 ) ;
  assign n1531 = ( n1527 & n1529 ) | ( n1527 & ~n1530 ) | ( n1529 & ~n1530 ) ;
  assign n1532 = n131 & ~n1531 ;
  assign n1533 = x82 | x83 ;
  assign n1534 = x84 | n1533 ;
  assign n1535 = ~n1393 & n1534 ;
  assign n1536 = n1399 & n1523 ;
  assign n1537 = ( x85 & n1523 ) | ( x85 & ~n1535 ) | ( n1523 & ~n1535 ) ;
  assign n1538 = n1393 & ~n1534 ;
  assign n1539 = n1537 & ~n1538 ;
  assign n1540 = ( n1535 & ~n1536 ) | ( n1535 & n1539 ) | ( ~n1536 & n1539 ) ;
  assign n1541 = n1393 | n1520 ;
  assign n1542 = ( x86 & n1536 ) | ( x86 & n1541 ) | ( n1536 & n1541 ) ;
  assign n1543 = ( ~x86 & n1536 ) | ( ~x86 & n1541 ) | ( n1536 & n1541 ) ;
  assign n1544 = ( x86 & ~n1542 ) | ( x86 & n1543 ) | ( ~n1542 & n1543 ) ;
  assign n1545 = ( ~n1266 & n1540 ) | ( ~n1266 & n1544 ) | ( n1540 & n1544 ) ;
  assign n1546 = n1541 & ~n1542 ;
  assign n1547 = ( ~n1266 & n1387 ) | ( ~n1266 & n1392 ) | ( n1387 & n1392 ) ;
  assign n1548 = ( n1407 & n1523 ) | ( n1407 & n1547 ) | ( n1523 & n1547 ) ;
  assign n1549 = ( x87 & n1546 ) | ( x87 & n1548 ) | ( n1546 & n1548 ) ;
  assign n1550 = ( ~x87 & n1546 ) | ( ~x87 & n1548 ) | ( n1546 & n1548 ) ;
  assign n1551 = ( x87 & ~n1549 ) | ( x87 & n1550 ) | ( ~n1549 & n1550 ) ;
  assign n1552 = ( ~n1150 & n1545 ) | ( ~n1150 & n1551 ) | ( n1545 & n1551 ) ;
  assign n1553 = ( n1150 & ~n1406 ) | ( n1150 & n1523 ) | ( ~n1406 & n1523 ) ;
  assign n1554 = n1150 & ~n1406 ;
  assign n1555 = ( n1410 & n1553 ) | ( n1410 & n1554 ) | ( n1553 & n1554 ) ;
  assign n1556 = ( ~n1410 & n1553 ) | ( ~n1410 & n1554 ) | ( n1553 & n1554 ) ;
  assign n1557 = ( n1410 & ~n1555 ) | ( n1410 & n1556 ) | ( ~n1555 & n1556 ) ;
  assign n1558 = ( ~n1038 & n1552 ) | ( ~n1038 & n1557 ) | ( n1552 & n1557 ) ;
  assign n1559 = ~n1038 & n1411 ;
  assign n1560 = ( ~n1038 & n1411 ) | ( ~n1038 & n1523 ) | ( n1411 & n1523 ) ;
  assign n1561 = ( ~n1416 & n1559 ) | ( ~n1416 & n1560 ) | ( n1559 & n1560 ) ;
  assign n1562 = ( n1416 & n1559 ) | ( n1416 & n1560 ) | ( n1559 & n1560 ) ;
  assign n1563 = ( n1416 & n1561 ) | ( n1416 & ~n1562 ) | ( n1561 & ~n1562 ) ;
  assign n1564 = ( ~n933 & n1558 ) | ( ~n933 & n1563 ) | ( n1558 & n1563 ) ;
  assign n1565 = ( n933 & ~n1417 ) | ( n933 & n1523 ) | ( ~n1417 & n1523 ) ;
  assign n1566 = n933 & ~n1417 ;
  assign n1567 = ( n1422 & n1565 ) | ( n1422 & n1566 ) | ( n1565 & n1566 ) ;
  assign n1568 = ( ~n1422 & n1565 ) | ( ~n1422 & n1566 ) | ( n1565 & n1566 ) ;
  assign n1569 = ( n1422 & ~n1567 ) | ( n1422 & n1568 ) | ( ~n1567 & n1568 ) ;
  assign n1570 = ( ~n839 & n1564 ) | ( ~n839 & n1569 ) | ( n1564 & n1569 ) ;
  assign n1571 = n839 & ~n1423 ;
  assign n1572 = ( n839 & ~n1423 ) | ( n839 & n1523 ) | ( ~n1423 & n1523 ) ;
  assign n1573 = ( n1428 & n1571 ) | ( n1428 & n1572 ) | ( n1571 & n1572 ) ;
  assign n1574 = ( ~n1428 & n1571 ) | ( ~n1428 & n1572 ) | ( n1571 & n1572 ) ;
  assign n1575 = ( n1428 & ~n1573 ) | ( n1428 & n1574 ) | ( ~n1573 & n1574 ) ;
  assign n1576 = ( ~n746 & n1570 ) | ( ~n746 & n1575 ) | ( n1570 & n1575 ) ;
  assign n1577 = ~n746 & n1429 ;
  assign n1578 = ( ~n746 & n1429 ) | ( ~n746 & n1523 ) | ( n1429 & n1523 ) ;
  assign n1579 = ( ~n1434 & n1577 ) | ( ~n1434 & n1578 ) | ( n1577 & n1578 ) ;
  assign n1580 = ( n1434 & n1577 ) | ( n1434 & n1578 ) | ( n1577 & n1578 ) ;
  assign n1581 = ( n1434 & n1579 ) | ( n1434 & ~n1580 ) | ( n1579 & ~n1580 ) ;
  assign n1582 = ( ~n664 & n1576 ) | ( ~n664 & n1581 ) | ( n1576 & n1581 ) ;
  assign n1583 = ~n664 & n1435 ;
  assign n1584 = ( ~n664 & n1435 ) | ( ~n664 & n1523 ) | ( n1435 & n1523 ) ;
  assign n1585 = ( ~n1440 & n1583 ) | ( ~n1440 & n1584 ) | ( n1583 & n1584 ) ;
  assign n1586 = ( n1440 & n1583 ) | ( n1440 & n1584 ) | ( n1583 & n1584 ) ;
  assign n1587 = ( n1440 & n1585 ) | ( n1440 & ~n1586 ) | ( n1585 & ~n1586 ) ;
  assign n1588 = ( ~n588 & n1582 ) | ( ~n588 & n1587 ) | ( n1582 & n1587 ) ;
  assign n1589 = ( n588 & ~n1441 ) | ( n588 & n1523 ) | ( ~n1441 & n1523 ) ;
  assign n1590 = n588 & ~n1441 ;
  assign n1591 = ( n1446 & n1589 ) | ( n1446 & n1590 ) | ( n1589 & n1590 ) ;
  assign n1592 = ( ~n1446 & n1589 ) | ( ~n1446 & n1590 ) | ( n1589 & n1590 ) ;
  assign n1593 = ( n1446 & ~n1591 ) | ( n1446 & n1592 ) | ( ~n1591 & n1592 ) ;
  assign n1594 = ( ~n518 & n1588 ) | ( ~n518 & n1593 ) | ( n1588 & n1593 ) ;
  assign n1595 = ~n518 & n1447 ;
  assign n1596 = ( ~n518 & n1447 ) | ( ~n518 & n1523 ) | ( n1447 & n1523 ) ;
  assign n1597 = ( ~n1452 & n1595 ) | ( ~n1452 & n1596 ) | ( n1595 & n1596 ) ;
  assign n1598 = ( n1452 & n1595 ) | ( n1452 & n1596 ) | ( n1595 & n1596 ) ;
  assign n1599 = ( n1452 & n1597 ) | ( n1452 & ~n1598 ) | ( n1597 & ~n1598 ) ;
  assign n1600 = ( ~n454 & n1594 ) | ( ~n454 & n1599 ) | ( n1594 & n1599 ) ;
  assign n1601 = ( n454 & ~n1453 ) | ( n454 & n1523 ) | ( ~n1453 & n1523 ) ;
  assign n1602 = n454 & ~n1453 ;
  assign n1603 = ( n1458 & n1601 ) | ( n1458 & n1602 ) | ( n1601 & n1602 ) ;
  assign n1604 = ( ~n1458 & n1601 ) | ( ~n1458 & n1602 ) | ( n1601 & n1602 ) ;
  assign n1605 = ( n1458 & ~n1603 ) | ( n1458 & n1604 ) | ( ~n1603 & n1604 ) ;
  assign n1606 = ( ~n396 & n1600 ) | ( ~n396 & n1605 ) | ( n1600 & n1605 ) ;
  assign n1607 = ( n396 & ~n1459 ) | ( n396 & n1523 ) | ( ~n1459 & n1523 ) ;
  assign n1608 = n396 & ~n1459 ;
  assign n1609 = ( n1464 & n1607 ) | ( n1464 & n1608 ) | ( n1607 & n1608 ) ;
  assign n1610 = ( ~n1464 & n1607 ) | ( ~n1464 & n1608 ) | ( n1607 & n1608 ) ;
  assign n1611 = ( n1464 & ~n1609 ) | ( n1464 & n1610 ) | ( ~n1609 & n1610 ) ;
  assign n1612 = ( ~n344 & n1606 ) | ( ~n344 & n1611 ) | ( n1606 & n1611 ) ;
  assign n1613 = ~n344 & n1465 ;
  assign n1614 = ( ~n344 & n1465 ) | ( ~n344 & n1523 ) | ( n1465 & n1523 ) ;
  assign n1615 = ( ~n1470 & n1613 ) | ( ~n1470 & n1614 ) | ( n1613 & n1614 ) ;
  assign n1616 = ( n1470 & n1613 ) | ( n1470 & n1614 ) | ( n1613 & n1614 ) ;
  assign n1617 = ( n1470 & n1615 ) | ( n1470 & ~n1616 ) | ( n1615 & ~n1616 ) ;
  assign n1618 = ( ~n298 & n1612 ) | ( ~n298 & n1617 ) | ( n1612 & n1617 ) ;
  assign n1619 = n298 & ~n1471 ;
  assign n1620 = ( n298 & ~n1471 ) | ( n298 & n1523 ) | ( ~n1471 & n1523 ) ;
  assign n1621 = ( ~n1476 & n1619 ) | ( ~n1476 & n1620 ) | ( n1619 & n1620 ) ;
  assign n1622 = ( n1476 & n1619 ) | ( n1476 & n1620 ) | ( n1619 & n1620 ) ;
  assign n1623 = ( n1476 & n1621 ) | ( n1476 & ~n1622 ) | ( n1621 & ~n1622 ) ;
  assign n1624 = ( ~n258 & n1618 ) | ( ~n258 & n1623 ) | ( n1618 & n1623 ) ;
  assign n1625 = ~n258 & n1477 ;
  assign n1626 = ( ~n258 & n1477 ) | ( ~n258 & n1523 ) | ( n1477 & n1523 ) ;
  assign n1627 = ( n1482 & n1625 ) | ( n1482 & n1626 ) | ( n1625 & n1626 ) ;
  assign n1628 = ( ~n1482 & n1625 ) | ( ~n1482 & n1626 ) | ( n1625 & n1626 ) ;
  assign n1629 = ( n1482 & ~n1627 ) | ( n1482 & n1628 ) | ( ~n1627 & n1628 ) ;
  assign n1630 = ( ~n225 & n1624 ) | ( ~n225 & n1629 ) | ( n1624 & n1629 ) ;
  assign n1631 = ( n225 & ~n1483 ) | ( n225 & n1523 ) | ( ~n1483 & n1523 ) ;
  assign n1632 = n225 & ~n1483 ;
  assign n1633 = ( n1488 & n1631 ) | ( n1488 & n1632 ) | ( n1631 & n1632 ) ;
  assign n1634 = ( ~n1488 & n1631 ) | ( ~n1488 & n1632 ) | ( n1631 & n1632 ) ;
  assign n1635 = ( n1488 & ~n1633 ) | ( n1488 & n1634 ) | ( ~n1633 & n1634 ) ;
  assign n1636 = ( ~n197 & n1630 ) | ( ~n197 & n1635 ) | ( n1630 & n1635 ) ;
  assign n1637 = ~n197 & n1489 ;
  assign n1638 = ( ~n197 & n1489 ) | ( ~n197 & n1523 ) | ( n1489 & n1523 ) ;
  assign n1639 = ( ~n1494 & n1637 ) | ( ~n1494 & n1638 ) | ( n1637 & n1638 ) ;
  assign n1640 = ( n1494 & n1637 ) | ( n1494 & n1638 ) | ( n1637 & n1638 ) ;
  assign n1641 = ( n1494 & n1639 ) | ( n1494 & ~n1640 ) | ( n1639 & ~n1640 ) ;
  assign n1642 = ( ~n170 & n1636 ) | ( ~n170 & n1641 ) | ( n1636 & n1641 ) ;
  assign n1643 = n170 & ~n1495 ;
  assign n1644 = ( n170 & ~n1495 ) | ( n170 & n1523 ) | ( ~n1495 & n1523 ) ;
  assign n1645 = ( n1500 & n1643 ) | ( n1500 & n1644 ) | ( n1643 & n1644 ) ;
  assign n1646 = ( ~n1500 & n1643 ) | ( ~n1500 & n1644 ) | ( n1643 & n1644 ) ;
  assign n1647 = ( n1500 & ~n1645 ) | ( n1500 & n1646 ) | ( ~n1645 & n1646 ) ;
  assign n1648 = ( ~n142 & n1642 ) | ( ~n142 & n1647 ) | ( n1642 & n1647 ) ;
  assign n1649 = ( n142 & ~n1501 ) | ( n142 & n1523 ) | ( ~n1501 & n1523 ) ;
  assign n1650 = n142 & ~n1501 ;
  assign n1651 = ( n1506 & n1649 ) | ( n1506 & n1650 ) | ( n1649 & n1650 ) ;
  assign n1652 = ( ~n1506 & n1649 ) | ( ~n1506 & n1650 ) | ( n1649 & n1650 ) ;
  assign n1653 = ( n1506 & ~n1651 ) | ( n1506 & n1652 ) | ( ~n1651 & n1652 ) ;
  assign n1654 = ( ~n132 & n1648 ) | ( ~n132 & n1653 ) | ( n1648 & n1653 ) ;
  assign n1655 = n1513 | n1518 ;
  assign n1656 = n1522 & ~n1655 ;
  assign n1657 = ( n1396 & n1518 ) | ( n1396 & ~n1524 ) | ( n1518 & ~n1524 ) ;
  assign n1658 = ( ~n131 & n1656 ) | ( ~n131 & n1657 ) | ( n1656 & n1657 ) ;
  assign n1659 = ( ~n131 & n1531 ) | ( ~n131 & n1658 ) | ( n1531 & n1658 ) ;
  assign n1660 = ( ~n1532 & n1654 ) | ( ~n1532 & n1659 ) | ( n1654 & n1659 ) ;
  assign n1661 = n1526 | n1660 ;
  assign n1662 = n1531 | n1654 ;
  assign n1663 = n1526 & ~n1531 ;
  assign n1664 = n1654 & ~n1663 ;
  assign n1665 = ( n131 & ~n1662 ) | ( n131 & n1664 ) | ( ~n1662 & n1664 ) ;
  assign n1666 = ( n132 & ~n1648 ) | ( n132 & n1661 ) | ( ~n1648 & n1661 ) ;
  assign n1667 = n132 & ~n1648 ;
  assign n1668 = ( n1653 & ~n1666 ) | ( n1653 & n1667 ) | ( ~n1666 & n1667 ) ;
  assign n1669 = ( n1653 & n1666 ) | ( n1653 & n1667 ) | ( n1666 & n1667 ) ;
  assign n1670 = ( n1666 & n1668 ) | ( n1666 & ~n1669 ) | ( n1668 & ~n1669 ) ;
  assign n1671 = n1665 & ~n1670 ;
  assign n1672 = x80 | x81 ;
  assign n1673 = x82 | n1672 ;
  assign n1674 = ~n1523 & n1673 ;
  assign n1675 = ( x83 & ~n1661 ) | ( x83 & n1674 ) | ( ~n1661 & n1674 ) ;
  assign n1676 = ~n1533 & n1661 ;
  assign n1677 = n1523 & ~n1673 ;
  assign n1678 = ( n1675 & n1676 ) | ( n1675 & ~n1677 ) | ( n1676 & ~n1677 ) ;
  assign n1679 = n1523 & ~n1661 ;
  assign n1680 = ( ~x84 & n1676 ) | ( ~x84 & n1679 ) | ( n1676 & n1679 ) ;
  assign n1681 = ( x84 & n1676 ) | ( x84 & n1679 ) | ( n1676 & n1679 ) ;
  assign n1682 = ( x84 & n1680 ) | ( x84 & ~n1681 ) | ( n1680 & ~n1681 ) ;
  assign n1683 = ( ~n1393 & n1678 ) | ( ~n1393 & n1682 ) | ( n1678 & n1682 ) ;
  assign n1684 = ( n1393 & n1523 ) | ( n1393 & ~n1661 ) | ( n1523 & ~n1661 ) ;
  assign n1685 = n1541 & ~n1684 ;
  assign n1686 = ( ~x85 & n1680 ) | ( ~x85 & n1685 ) | ( n1680 & n1685 ) ;
  assign n1687 = ( x85 & n1680 ) | ( x85 & n1685 ) | ( n1680 & n1685 ) ;
  assign n1688 = ( x85 & n1686 ) | ( x85 & ~n1687 ) | ( n1686 & ~n1687 ) ;
  assign n1689 = ( ~n1266 & n1683 ) | ( ~n1266 & n1688 ) | ( n1683 & n1688 ) ;
  assign n1690 = n1266 & ~n1540 ;
  assign n1691 = ( n1266 & ~n1540 ) | ( n1266 & n1661 ) | ( ~n1540 & n1661 ) ;
  assign n1692 = ( ~n1544 & n1690 ) | ( ~n1544 & n1691 ) | ( n1690 & n1691 ) ;
  assign n1693 = ( n1544 & n1690 ) | ( n1544 & n1691 ) | ( n1690 & n1691 ) ;
  assign n1694 = ( n1544 & n1692 ) | ( n1544 & ~n1693 ) | ( n1692 & ~n1693 ) ;
  assign n1695 = ( ~n1150 & n1689 ) | ( ~n1150 & n1694 ) | ( n1689 & n1694 ) ;
  assign n1696 = ( n1150 & ~n1545 ) | ( n1150 & n1661 ) | ( ~n1545 & n1661 ) ;
  assign n1697 = n1150 & ~n1545 ;
  assign n1698 = ( n1551 & n1696 ) | ( n1551 & n1697 ) | ( n1696 & n1697 ) ;
  assign n1699 = ( ~n1551 & n1696 ) | ( ~n1551 & n1697 ) | ( n1696 & n1697 ) ;
  assign n1700 = ( n1551 & ~n1698 ) | ( n1551 & n1699 ) | ( ~n1698 & n1699 ) ;
  assign n1701 = ( ~n1038 & n1695 ) | ( ~n1038 & n1700 ) | ( n1695 & n1700 ) ;
  assign n1702 = ~n1038 & n1552 ;
  assign n1703 = ( ~n1038 & n1552 ) | ( ~n1038 & n1661 ) | ( n1552 & n1661 ) ;
  assign n1704 = ( ~n1557 & n1702 ) | ( ~n1557 & n1703 ) | ( n1702 & n1703 ) ;
  assign n1705 = ( n1557 & n1702 ) | ( n1557 & n1703 ) | ( n1702 & n1703 ) ;
  assign n1706 = ( n1557 & n1704 ) | ( n1557 & ~n1705 ) | ( n1704 & ~n1705 ) ;
  assign n1707 = ( ~n933 & n1701 ) | ( ~n933 & n1706 ) | ( n1701 & n1706 ) ;
  assign n1708 = ~n933 & n1558 ;
  assign n1709 = ( ~n933 & n1558 ) | ( ~n933 & n1661 ) | ( n1558 & n1661 ) ;
  assign n1710 = ( ~n1563 & n1708 ) | ( ~n1563 & n1709 ) | ( n1708 & n1709 ) ;
  assign n1711 = ( n1563 & n1708 ) | ( n1563 & n1709 ) | ( n1708 & n1709 ) ;
  assign n1712 = ( n1563 & n1710 ) | ( n1563 & ~n1711 ) | ( n1710 & ~n1711 ) ;
  assign n1713 = ( ~n839 & n1707 ) | ( ~n839 & n1712 ) | ( n1707 & n1712 ) ;
  assign n1714 = ( n839 & ~n1564 ) | ( n839 & n1661 ) | ( ~n1564 & n1661 ) ;
  assign n1715 = n839 & ~n1564 ;
  assign n1716 = ( n1569 & n1714 ) | ( n1569 & n1715 ) | ( n1714 & n1715 ) ;
  assign n1717 = ( ~n1569 & n1714 ) | ( ~n1569 & n1715 ) | ( n1714 & n1715 ) ;
  assign n1718 = ( n1569 & ~n1716 ) | ( n1569 & n1717 ) | ( ~n1716 & n1717 ) ;
  assign n1719 = ( ~n746 & n1713 ) | ( ~n746 & n1718 ) | ( n1713 & n1718 ) ;
  assign n1720 = ( n746 & ~n1570 ) | ( n746 & n1661 ) | ( ~n1570 & n1661 ) ;
  assign n1721 = n746 & ~n1570 ;
  assign n1722 = ( n1575 & n1720 ) | ( n1575 & n1721 ) | ( n1720 & n1721 ) ;
  assign n1723 = ( ~n1575 & n1720 ) | ( ~n1575 & n1721 ) | ( n1720 & n1721 ) ;
  assign n1724 = ( n1575 & ~n1722 ) | ( n1575 & n1723 ) | ( ~n1722 & n1723 ) ;
  assign n1725 = ( ~n664 & n1719 ) | ( ~n664 & n1724 ) | ( n1719 & n1724 ) ;
  assign n1726 = ( n664 & ~n1576 ) | ( n664 & n1661 ) | ( ~n1576 & n1661 ) ;
  assign n1727 = n664 & ~n1576 ;
  assign n1728 = ( n1581 & n1726 ) | ( n1581 & n1727 ) | ( n1726 & n1727 ) ;
  assign n1729 = ( ~n1581 & n1726 ) | ( ~n1581 & n1727 ) | ( n1726 & n1727 ) ;
  assign n1730 = ( n1581 & ~n1728 ) | ( n1581 & n1729 ) | ( ~n1728 & n1729 ) ;
  assign n1731 = ( ~n588 & n1725 ) | ( ~n588 & n1730 ) | ( n1725 & n1730 ) ;
  assign n1732 = ( n588 & ~n1582 ) | ( n588 & n1661 ) | ( ~n1582 & n1661 ) ;
  assign n1733 = n588 & ~n1582 ;
  assign n1734 = ( n1587 & n1732 ) | ( n1587 & n1733 ) | ( n1732 & n1733 ) ;
  assign n1735 = ( ~n1587 & n1732 ) | ( ~n1587 & n1733 ) | ( n1732 & n1733 ) ;
  assign n1736 = ( n1587 & ~n1734 ) | ( n1587 & n1735 ) | ( ~n1734 & n1735 ) ;
  assign n1737 = ( ~n518 & n1731 ) | ( ~n518 & n1736 ) | ( n1731 & n1736 ) ;
  assign n1738 = ( n518 & ~n1588 ) | ( n518 & n1661 ) | ( ~n1588 & n1661 ) ;
  assign n1739 = n518 & ~n1588 ;
  assign n1740 = ( n1593 & n1738 ) | ( n1593 & n1739 ) | ( n1738 & n1739 ) ;
  assign n1741 = ( ~n1593 & n1738 ) | ( ~n1593 & n1739 ) | ( n1738 & n1739 ) ;
  assign n1742 = ( n1593 & ~n1740 ) | ( n1593 & n1741 ) | ( ~n1740 & n1741 ) ;
  assign n1743 = ( ~n454 & n1737 ) | ( ~n454 & n1742 ) | ( n1737 & n1742 ) ;
  assign n1744 = ~n454 & n1594 ;
  assign n1745 = ( ~n454 & n1594 ) | ( ~n454 & n1661 ) | ( n1594 & n1661 ) ;
  assign n1746 = ( ~n1599 & n1744 ) | ( ~n1599 & n1745 ) | ( n1744 & n1745 ) ;
  assign n1747 = ( n1599 & n1744 ) | ( n1599 & n1745 ) | ( n1744 & n1745 ) ;
  assign n1748 = ( n1599 & n1746 ) | ( n1599 & ~n1747 ) | ( n1746 & ~n1747 ) ;
  assign n1749 = ( ~n396 & n1743 ) | ( ~n396 & n1748 ) | ( n1743 & n1748 ) ;
  assign n1750 = ( n396 & ~n1600 ) | ( n396 & n1661 ) | ( ~n1600 & n1661 ) ;
  assign n1751 = n396 & ~n1600 ;
  assign n1752 = ( n1605 & n1750 ) | ( n1605 & n1751 ) | ( n1750 & n1751 ) ;
  assign n1753 = ( ~n1605 & n1750 ) | ( ~n1605 & n1751 ) | ( n1750 & n1751 ) ;
  assign n1754 = ( n1605 & ~n1752 ) | ( n1605 & n1753 ) | ( ~n1752 & n1753 ) ;
  assign n1755 = ( ~n344 & n1749 ) | ( ~n344 & n1754 ) | ( n1749 & n1754 ) ;
  assign n1756 = n344 & ~n1606 ;
  assign n1757 = ( n344 & ~n1606 ) | ( n344 & n1661 ) | ( ~n1606 & n1661 ) ;
  assign n1758 = ( n1611 & n1756 ) | ( n1611 & n1757 ) | ( n1756 & n1757 ) ;
  assign n1759 = ( ~n1611 & n1756 ) | ( ~n1611 & n1757 ) | ( n1756 & n1757 ) ;
  assign n1760 = ( n1611 & ~n1758 ) | ( n1611 & n1759 ) | ( ~n1758 & n1759 ) ;
  assign n1761 = ( ~n298 & n1755 ) | ( ~n298 & n1760 ) | ( n1755 & n1760 ) ;
  assign n1762 = ( n298 & ~n1612 ) | ( n298 & n1661 ) | ( ~n1612 & n1661 ) ;
  assign n1763 = n298 & ~n1612 ;
  assign n1764 = ( n1617 & n1762 ) | ( n1617 & n1763 ) | ( n1762 & n1763 ) ;
  assign n1765 = ( ~n1617 & n1762 ) | ( ~n1617 & n1763 ) | ( n1762 & n1763 ) ;
  assign n1766 = ( n1617 & ~n1764 ) | ( n1617 & n1765 ) | ( ~n1764 & n1765 ) ;
  assign n1767 = ( ~n258 & n1761 ) | ( ~n258 & n1766 ) | ( n1761 & n1766 ) ;
  assign n1768 = ( n258 & ~n1618 ) | ( n258 & n1661 ) | ( ~n1618 & n1661 ) ;
  assign n1769 = n258 & ~n1618 ;
  assign n1770 = ( n1623 & n1768 ) | ( n1623 & n1769 ) | ( n1768 & n1769 ) ;
  assign n1771 = ( ~n1623 & n1768 ) | ( ~n1623 & n1769 ) | ( n1768 & n1769 ) ;
  assign n1772 = ( n1623 & ~n1770 ) | ( n1623 & n1771 ) | ( ~n1770 & n1771 ) ;
  assign n1773 = ( ~n225 & n1767 ) | ( ~n225 & n1772 ) | ( n1767 & n1772 ) ;
  assign n1774 = ~n225 & n1624 ;
  assign n1775 = ( ~n225 & n1624 ) | ( ~n225 & n1661 ) | ( n1624 & n1661 ) ;
  assign n1776 = ( n1629 & n1774 ) | ( n1629 & n1775 ) | ( n1774 & n1775 ) ;
  assign n1777 = ( ~n1629 & n1774 ) | ( ~n1629 & n1775 ) | ( n1774 & n1775 ) ;
  assign n1778 = ( n1629 & ~n1776 ) | ( n1629 & n1777 ) | ( ~n1776 & n1777 ) ;
  assign n1779 = ( ~n197 & n1773 ) | ( ~n197 & n1778 ) | ( n1773 & n1778 ) ;
  assign n1780 = ( n197 & ~n1630 ) | ( n197 & n1661 ) | ( ~n1630 & n1661 ) ;
  assign n1781 = n197 & ~n1630 ;
  assign n1782 = ( n1635 & n1780 ) | ( n1635 & n1781 ) | ( n1780 & n1781 ) ;
  assign n1783 = ( ~n1635 & n1780 ) | ( ~n1635 & n1781 ) | ( n1780 & n1781 ) ;
  assign n1784 = ( n1635 & ~n1782 ) | ( n1635 & n1783 ) | ( ~n1782 & n1783 ) ;
  assign n1785 = ( ~n170 & n1779 ) | ( ~n170 & n1784 ) | ( n1779 & n1784 ) ;
  assign n1786 = ~n170 & n1636 ;
  assign n1787 = ( ~n170 & n1636 ) | ( ~n170 & n1661 ) | ( n1636 & n1661 ) ;
  assign n1788 = ( ~n1641 & n1786 ) | ( ~n1641 & n1787 ) | ( n1786 & n1787 ) ;
  assign n1789 = ( n1641 & n1786 ) | ( n1641 & n1787 ) | ( n1786 & n1787 ) ;
  assign n1790 = ( n1641 & n1788 ) | ( n1641 & ~n1789 ) | ( n1788 & ~n1789 ) ;
  assign n1791 = ( ~n142 & n1785 ) | ( ~n142 & n1790 ) | ( n1785 & n1790 ) ;
  assign n1792 = ( n142 & ~n1642 ) | ( n142 & n1661 ) | ( ~n1642 & n1661 ) ;
  assign n1793 = n142 & ~n1642 ;
  assign n1794 = ( n1647 & n1792 ) | ( n1647 & n1793 ) | ( n1792 & n1793 ) ;
  assign n1795 = ( ~n1647 & n1792 ) | ( ~n1647 & n1793 ) | ( n1792 & n1793 ) ;
  assign n1796 = ( n1647 & ~n1794 ) | ( n1647 & n1795 ) | ( ~n1794 & n1795 ) ;
  assign n1797 = ( ~n132 & n1791 ) | ( ~n132 & n1796 ) | ( n1791 & n1796 ) ;
  assign n1798 = n131 | n1670 ;
  assign n1799 = ( ~n1531 & n1654 ) | ( ~n1531 & n1659 ) | ( n1654 & n1659 ) ;
  assign n1800 = ( n1531 & ~n1662 ) | ( n1531 & n1799 ) | ( ~n1662 & n1799 ) ;
  assign n1801 = ( ~n1665 & n1798 ) | ( ~n1665 & n1800 ) | ( n1798 & n1800 ) ;
  assign n1802 = ( ~n1671 & n1797 ) | ( ~n1671 & n1801 ) | ( n1797 & n1801 ) ;
  assign n1803 = ~n1670 & n1797 ;
  assign n1804 = n1670 & ~n1797 ;
  assign n1805 = ( n1662 & ~n1664 ) | ( n1662 & n1670 ) | ( ~n1664 & n1670 ) ;
  assign n1806 = ( n1803 & n1804 ) | ( n1803 & n1805 ) | ( n1804 & n1805 ) ;
  assign n1807 = n131 & ~n1806 ;
  assign n1808 = ~n1672 & n1802 ;
  assign n1809 = x78 | x79 ;
  assign n1810 = x80 | n1809 ;
  assign n1811 = n1661 & ~n1810 ;
  assign n1812 = ~n1661 & n1810 ;
  assign n1813 = ( x81 & ~n1802 ) | ( x81 & n1812 ) | ( ~n1802 & n1812 ) ;
  assign n1814 = ( n1808 & ~n1811 ) | ( n1808 & n1813 ) | ( ~n1811 & n1813 ) ;
  assign n1815 = n1661 & ~n1802 ;
  assign n1816 = ( x82 & n1808 ) | ( x82 & n1815 ) | ( n1808 & n1815 ) ;
  assign n1817 = ( ~x82 & n1808 ) | ( ~x82 & n1815 ) | ( n1808 & n1815 ) ;
  assign n1818 = ( x82 & ~n1816 ) | ( x82 & n1817 ) | ( ~n1816 & n1817 ) ;
  assign n1819 = ( ~n1523 & n1814 ) | ( ~n1523 & n1818 ) | ( n1814 & n1818 ) ;
  assign n1820 = ~n1523 & n1661 ;
  assign n1821 = ( n1679 & n1802 ) | ( n1679 & n1820 ) | ( n1802 & n1820 ) ;
  assign n1822 = ( ~x83 & n1817 ) | ( ~x83 & n1821 ) | ( n1817 & n1821 ) ;
  assign n1823 = ( x83 & n1817 ) | ( x83 & n1821 ) | ( n1817 & n1821 ) ;
  assign n1824 = ( x83 & n1822 ) | ( x83 & ~n1823 ) | ( n1822 & ~n1823 ) ;
  assign n1825 = ( ~n1393 & n1819 ) | ( ~n1393 & n1824 ) | ( n1819 & n1824 ) ;
  assign n1826 = ( n1393 & ~n1678 ) | ( n1393 & n1802 ) | ( ~n1678 & n1802 ) ;
  assign n1827 = n1393 & ~n1678 ;
  assign n1828 = ( n1682 & n1826 ) | ( n1682 & n1827 ) | ( n1826 & n1827 ) ;
  assign n1829 = ( ~n1682 & n1826 ) | ( ~n1682 & n1827 ) | ( n1826 & n1827 ) ;
  assign n1830 = ( n1682 & ~n1828 ) | ( n1682 & n1829 ) | ( ~n1828 & n1829 ) ;
  assign n1831 = ( ~n1266 & n1825 ) | ( ~n1266 & n1830 ) | ( n1825 & n1830 ) ;
  assign n1832 = n1266 & ~n1683 ;
  assign n1833 = ( n1266 & ~n1683 ) | ( n1266 & n1802 ) | ( ~n1683 & n1802 ) ;
  assign n1834 = ( ~n1688 & n1832 ) | ( ~n1688 & n1833 ) | ( n1832 & n1833 ) ;
  assign n1835 = ( n1688 & n1832 ) | ( n1688 & n1833 ) | ( n1832 & n1833 ) ;
  assign n1836 = ( n1688 & n1834 ) | ( n1688 & ~n1835 ) | ( n1834 & ~n1835 ) ;
  assign n1837 = ( ~n1150 & n1831 ) | ( ~n1150 & n1836 ) | ( n1831 & n1836 ) ;
  assign n1838 = ( n1150 & ~n1689 ) | ( n1150 & n1802 ) | ( ~n1689 & n1802 ) ;
  assign n1839 = n1150 & ~n1689 ;
  assign n1840 = ( n1694 & n1838 ) | ( n1694 & n1839 ) | ( n1838 & n1839 ) ;
  assign n1841 = ( ~n1694 & n1838 ) | ( ~n1694 & n1839 ) | ( n1838 & n1839 ) ;
  assign n1842 = ( n1694 & ~n1840 ) | ( n1694 & n1841 ) | ( ~n1840 & n1841 ) ;
  assign n1843 = ( ~n1038 & n1837 ) | ( ~n1038 & n1842 ) | ( n1837 & n1842 ) ;
  assign n1844 = n1038 & ~n1695 ;
  assign n1845 = ( n1038 & ~n1695 ) | ( n1038 & n1802 ) | ( ~n1695 & n1802 ) ;
  assign n1846 = ( n1700 & n1844 ) | ( n1700 & n1845 ) | ( n1844 & n1845 ) ;
  assign n1847 = ( ~n1700 & n1844 ) | ( ~n1700 & n1845 ) | ( n1844 & n1845 ) ;
  assign n1848 = ( n1700 & ~n1846 ) | ( n1700 & n1847 ) | ( ~n1846 & n1847 ) ;
  assign n1849 = ( ~n933 & n1843 ) | ( ~n933 & n1848 ) | ( n1843 & n1848 ) ;
  assign n1850 = n933 & ~n1701 ;
  assign n1851 = ( n933 & ~n1701 ) | ( n933 & n1802 ) | ( ~n1701 & n1802 ) ;
  assign n1852 = ( n1706 & n1850 ) | ( n1706 & n1851 ) | ( n1850 & n1851 ) ;
  assign n1853 = ( ~n1706 & n1850 ) | ( ~n1706 & n1851 ) | ( n1850 & n1851 ) ;
  assign n1854 = ( n1706 & ~n1852 ) | ( n1706 & n1853 ) | ( ~n1852 & n1853 ) ;
  assign n1855 = ( ~n839 & n1849 ) | ( ~n839 & n1854 ) | ( n1849 & n1854 ) ;
  assign n1856 = ~n839 & n1707 ;
  assign n1857 = ( ~n839 & n1707 ) | ( ~n839 & n1802 ) | ( n1707 & n1802 ) ;
  assign n1858 = ( ~n1712 & n1856 ) | ( ~n1712 & n1857 ) | ( n1856 & n1857 ) ;
  assign n1859 = ( n1712 & n1856 ) | ( n1712 & n1857 ) | ( n1856 & n1857 ) ;
  assign n1860 = ( n1712 & n1858 ) | ( n1712 & ~n1859 ) | ( n1858 & ~n1859 ) ;
  assign n1861 = ( ~n746 & n1855 ) | ( ~n746 & n1860 ) | ( n1855 & n1860 ) ;
  assign n1862 = ~n746 & n1713 ;
  assign n1863 = ( ~n746 & n1713 ) | ( ~n746 & n1802 ) | ( n1713 & n1802 ) ;
  assign n1864 = ( ~n1718 & n1862 ) | ( ~n1718 & n1863 ) | ( n1862 & n1863 ) ;
  assign n1865 = ( n1718 & n1862 ) | ( n1718 & n1863 ) | ( n1862 & n1863 ) ;
  assign n1866 = ( n1718 & n1864 ) | ( n1718 & ~n1865 ) | ( n1864 & ~n1865 ) ;
  assign n1867 = ( ~n664 & n1861 ) | ( ~n664 & n1866 ) | ( n1861 & n1866 ) ;
  assign n1868 = ~n664 & n1719 ;
  assign n1869 = ( ~n664 & n1719 ) | ( ~n664 & n1802 ) | ( n1719 & n1802 ) ;
  assign n1870 = ( ~n1724 & n1868 ) | ( ~n1724 & n1869 ) | ( n1868 & n1869 ) ;
  assign n1871 = ( n1724 & n1868 ) | ( n1724 & n1869 ) | ( n1868 & n1869 ) ;
  assign n1872 = ( n1724 & n1870 ) | ( n1724 & ~n1871 ) | ( n1870 & ~n1871 ) ;
  assign n1873 = ( ~n588 & n1867 ) | ( ~n588 & n1872 ) | ( n1867 & n1872 ) ;
  assign n1874 = ~n588 & n1725 ;
  assign n1875 = ( ~n588 & n1725 ) | ( ~n588 & n1802 ) | ( n1725 & n1802 ) ;
  assign n1876 = ( ~n1730 & n1874 ) | ( ~n1730 & n1875 ) | ( n1874 & n1875 ) ;
  assign n1877 = ( n1730 & n1874 ) | ( n1730 & n1875 ) | ( n1874 & n1875 ) ;
  assign n1878 = ( n1730 & n1876 ) | ( n1730 & ~n1877 ) | ( n1876 & ~n1877 ) ;
  assign n1879 = ( ~n518 & n1873 ) | ( ~n518 & n1878 ) | ( n1873 & n1878 ) ;
  assign n1880 = ~n518 & n1731 ;
  assign n1881 = ( ~n518 & n1731 ) | ( ~n518 & n1802 ) | ( n1731 & n1802 ) ;
  assign n1882 = ( ~n1736 & n1880 ) | ( ~n1736 & n1881 ) | ( n1880 & n1881 ) ;
  assign n1883 = ( n1736 & n1880 ) | ( n1736 & n1881 ) | ( n1880 & n1881 ) ;
  assign n1884 = ( n1736 & n1882 ) | ( n1736 & ~n1883 ) | ( n1882 & ~n1883 ) ;
  assign n1885 = ( ~n454 & n1879 ) | ( ~n454 & n1884 ) | ( n1879 & n1884 ) ;
  assign n1886 = ( n454 & ~n1737 ) | ( n454 & n1802 ) | ( ~n1737 & n1802 ) ;
  assign n1887 = n454 & ~n1737 ;
  assign n1888 = ( n1742 & n1886 ) | ( n1742 & n1887 ) | ( n1886 & n1887 ) ;
  assign n1889 = ( ~n1742 & n1886 ) | ( ~n1742 & n1887 ) | ( n1886 & n1887 ) ;
  assign n1890 = ( n1742 & ~n1888 ) | ( n1742 & n1889 ) | ( ~n1888 & n1889 ) ;
  assign n1891 = ( ~n396 & n1885 ) | ( ~n396 & n1890 ) | ( n1885 & n1890 ) ;
  assign n1892 = ( n396 & ~n1743 ) | ( n396 & n1802 ) | ( ~n1743 & n1802 ) ;
  assign n1893 = n396 & ~n1743 ;
  assign n1894 = ( n1748 & n1892 ) | ( n1748 & n1893 ) | ( n1892 & n1893 ) ;
  assign n1895 = ( ~n1748 & n1892 ) | ( ~n1748 & n1893 ) | ( n1892 & n1893 ) ;
  assign n1896 = ( n1748 & ~n1894 ) | ( n1748 & n1895 ) | ( ~n1894 & n1895 ) ;
  assign n1897 = ( ~n344 & n1891 ) | ( ~n344 & n1896 ) | ( n1891 & n1896 ) ;
  assign n1898 = n344 & ~n1749 ;
  assign n1899 = ( n344 & ~n1749 ) | ( n344 & n1802 ) | ( ~n1749 & n1802 ) ;
  assign n1900 = ( n1754 & n1898 ) | ( n1754 & n1899 ) | ( n1898 & n1899 ) ;
  assign n1901 = ( ~n1754 & n1898 ) | ( ~n1754 & n1899 ) | ( n1898 & n1899 ) ;
  assign n1902 = ( n1754 & ~n1900 ) | ( n1754 & n1901 ) | ( ~n1900 & n1901 ) ;
  assign n1903 = ( ~n298 & n1897 ) | ( ~n298 & n1902 ) | ( n1897 & n1902 ) ;
  assign n1904 = ~n298 & n1755 ;
  assign n1905 = ( ~n298 & n1755 ) | ( ~n298 & n1802 ) | ( n1755 & n1802 ) ;
  assign n1906 = ( ~n1760 & n1904 ) | ( ~n1760 & n1905 ) | ( n1904 & n1905 ) ;
  assign n1907 = ( n1760 & n1904 ) | ( n1760 & n1905 ) | ( n1904 & n1905 ) ;
  assign n1908 = ( n1760 & n1906 ) | ( n1760 & ~n1907 ) | ( n1906 & ~n1907 ) ;
  assign n1909 = ( ~n258 & n1903 ) | ( ~n258 & n1908 ) | ( n1903 & n1908 ) ;
  assign n1910 = ( n258 & ~n1761 ) | ( n258 & n1802 ) | ( ~n1761 & n1802 ) ;
  assign n1911 = n258 & ~n1761 ;
  assign n1912 = ( n1766 & n1910 ) | ( n1766 & n1911 ) | ( n1910 & n1911 ) ;
  assign n1913 = ( ~n1766 & n1910 ) | ( ~n1766 & n1911 ) | ( n1910 & n1911 ) ;
  assign n1914 = ( n1766 & ~n1912 ) | ( n1766 & n1913 ) | ( ~n1912 & n1913 ) ;
  assign n1915 = ( ~n225 & n1909 ) | ( ~n225 & n1914 ) | ( n1909 & n1914 ) ;
  assign n1916 = ~n225 & n1767 ;
  assign n1917 = ( ~n225 & n1767 ) | ( ~n225 & n1802 ) | ( n1767 & n1802 ) ;
  assign n1918 = ( ~n1772 & n1916 ) | ( ~n1772 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1919 = ( n1772 & n1916 ) | ( n1772 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1920 = ( n1772 & n1918 ) | ( n1772 & ~n1919 ) | ( n1918 & ~n1919 ) ;
  assign n1921 = ( ~n197 & n1915 ) | ( ~n197 & n1920 ) | ( n1915 & n1920 ) ;
  assign n1922 = ~n197 & n1773 ;
  assign n1923 = ( ~n197 & n1773 ) | ( ~n197 & n1802 ) | ( n1773 & n1802 ) ;
  assign n1924 = ( n1778 & n1922 ) | ( n1778 & n1923 ) | ( n1922 & n1923 ) ;
  assign n1925 = ( ~n1778 & n1922 ) | ( ~n1778 & n1923 ) | ( n1922 & n1923 ) ;
  assign n1926 = ( n1778 & ~n1924 ) | ( n1778 & n1925 ) | ( ~n1924 & n1925 ) ;
  assign n1927 = ( ~n170 & n1921 ) | ( ~n170 & n1926 ) | ( n1921 & n1926 ) ;
  assign n1928 = ~n170 & n1779 ;
  assign n1929 = ( ~n170 & n1779 ) | ( ~n170 & n1802 ) | ( n1779 & n1802 ) ;
  assign n1930 = ( ~n1784 & n1928 ) | ( ~n1784 & n1929 ) | ( n1928 & n1929 ) ;
  assign n1931 = ( n1784 & n1928 ) | ( n1784 & n1929 ) | ( n1928 & n1929 ) ;
  assign n1932 = ( n1784 & n1930 ) | ( n1784 & ~n1931 ) | ( n1930 & ~n1931 ) ;
  assign n1933 = ( ~n142 & n1927 ) | ( ~n142 & n1932 ) | ( n1927 & n1932 ) ;
  assign n1934 = ( n142 & ~n1785 ) | ( n142 & n1802 ) | ( ~n1785 & n1802 ) ;
  assign n1935 = n142 & ~n1785 ;
  assign n1936 = ( n1790 & n1934 ) | ( n1790 & n1935 ) | ( n1934 & n1935 ) ;
  assign n1937 = ( ~n1790 & n1934 ) | ( ~n1790 & n1935 ) | ( n1934 & n1935 ) ;
  assign n1938 = ( n1790 & ~n1936 ) | ( n1790 & n1937 ) | ( ~n1936 & n1937 ) ;
  assign n1939 = ( ~n132 & n1933 ) | ( ~n132 & n1938 ) | ( n1933 & n1938 ) ;
  assign n1940 = ~n132 & n1791 ;
  assign n1941 = ( ~n132 & n1791 ) | ( ~n132 & n1802 ) | ( n1791 & n1802 ) ;
  assign n1942 = ( n1796 & n1940 ) | ( n1796 & n1941 ) | ( n1940 & n1941 ) ;
  assign n1943 = ( ~n1796 & n1940 ) | ( ~n1796 & n1941 ) | ( n1940 & n1941 ) ;
  assign n1944 = ( n1796 & ~n1942 ) | ( n1796 & n1943 ) | ( ~n1942 & n1943 ) ;
  assign n1945 = ( n1797 & n1800 ) | ( n1797 & ~n1804 ) | ( n1800 & ~n1804 ) ;
  assign n1946 = ( ~n1803 & n1944 ) | ( ~n1803 & n1945 ) | ( n1944 & n1945 ) ;
  assign n1947 = n131 | n1946 ;
  assign n1948 = ( ~n1807 & n1944 ) | ( ~n1807 & n1947 ) | ( n1944 & n1947 ) ;
  assign n1949 = ( ~n1807 & n1939 ) | ( ~n1807 & n1948 ) | ( n1939 & n1948 ) ;
  assign n1950 = ( n142 & ~n1927 ) | ( n142 & n1949 ) | ( ~n1927 & n1949 ) ;
  assign n1951 = n142 & ~n1927 ;
  assign n1952 = ( n1932 & ~n1950 ) | ( n1932 & n1951 ) | ( ~n1950 & n1951 ) ;
  assign n1953 = ( n1932 & n1950 ) | ( n1932 & n1951 ) | ( n1950 & n1951 ) ;
  assign n1954 = ( n1950 & n1952 ) | ( n1950 & ~n1953 ) | ( n1952 & ~n1953 ) ;
  assign n1955 = n1802 | n1949 ;
  assign n1956 = ~x80 & n1955 ;
  assign n1957 = ~n1661 & n1802 ;
  assign n1958 = ( n1810 & n1815 ) | ( n1810 & n1957 ) | ( n1815 & n1957 ) ;
  assign n1959 = n1949 & ~n1958 ;
  assign n1960 = ( ~n1661 & n1802 ) | ( ~n1661 & n1809 ) | ( n1802 & n1809 ) ;
  assign n1961 = n1815 | n1960 ;
  assign n1962 = ( n1949 & n1958 ) | ( n1949 & ~n1961 ) | ( n1958 & ~n1961 ) ;
  assign n1963 = ( n1956 & ~n1959 ) | ( n1956 & n1962 ) | ( ~n1959 & n1962 ) ;
  assign n1964 = x81 & ~n1963 ;
  assign n1965 = ~x81 & n1963 ;
  assign n1966 = n1964 | n1965 ;
  assign n1967 = n1809 & n1949 ;
  assign n1968 = ~x79 & n1967 ;
  assign n1969 = x76 | x77 ;
  assign n1970 = x78 | n1969 ;
  assign n1971 = x79 & n1949 ;
  assign n1972 = x79 | n1949 ;
  assign n1973 = ~n1802 & n1970 ;
  assign n1974 = ( ~n1971 & n1972 ) | ( ~n1971 & n1973 ) | ( n1972 & n1973 ) ;
  assign n1975 = ( ~n1802 & n1970 ) | ( ~n1802 & n1974 ) | ( n1970 & n1974 ) ;
  assign n1976 = ~n1968 & n1975 ;
  assign n1977 = ( ~x80 & n1955 ) | ( ~x80 & n1967 ) | ( n1955 & n1967 ) ;
  assign n1978 = ( x80 & n1955 ) | ( x80 & n1967 ) | ( n1955 & n1967 ) ;
  assign n1979 = ( x80 & n1977 ) | ( x80 & ~n1978 ) | ( n1977 & ~n1978 ) ;
  assign n1980 = ( ~n1661 & n1976 ) | ( ~n1661 & n1979 ) | ( n1976 & n1979 ) ;
  assign n1981 = ( ~n1523 & n1966 ) | ( ~n1523 & n1980 ) | ( n1966 & n1980 ) ;
  assign n1982 = n1523 & ~n1814 ;
  assign n1983 = ( n1523 & ~n1814 ) | ( n1523 & n1949 ) | ( ~n1814 & n1949 ) ;
  assign n1984 = ( n1818 & n1982 ) | ( n1818 & n1983 ) | ( n1982 & n1983 ) ;
  assign n1985 = ( ~n1818 & n1982 ) | ( ~n1818 & n1983 ) | ( n1982 & n1983 ) ;
  assign n1986 = ( n1818 & ~n1984 ) | ( n1818 & n1985 ) | ( ~n1984 & n1985 ) ;
  assign n1987 = ( ~n1393 & n1981 ) | ( ~n1393 & n1986 ) | ( n1981 & n1986 ) ;
  assign n1988 = n1393 & ~n1819 ;
  assign n1989 = ( n1393 & ~n1819 ) | ( n1393 & n1949 ) | ( ~n1819 & n1949 ) ;
  assign n1990 = ( ~n1824 & n1988 ) | ( ~n1824 & n1989 ) | ( n1988 & n1989 ) ;
  assign n1991 = ( n1824 & n1988 ) | ( n1824 & n1989 ) | ( n1988 & n1989 ) ;
  assign n1992 = ( n1824 & n1990 ) | ( n1824 & ~n1991 ) | ( n1990 & ~n1991 ) ;
  assign n1993 = ( ~n1266 & n1987 ) | ( ~n1266 & n1992 ) | ( n1987 & n1992 ) ;
  assign n1994 = ( n1266 & ~n1825 ) | ( n1266 & n1949 ) | ( ~n1825 & n1949 ) ;
  assign n1995 = n1266 & ~n1825 ;
  assign n1996 = ( n1830 & n1994 ) | ( n1830 & n1995 ) | ( n1994 & n1995 ) ;
  assign n1997 = ( ~n1830 & n1994 ) | ( ~n1830 & n1995 ) | ( n1994 & n1995 ) ;
  assign n1998 = ( n1830 & ~n1996 ) | ( n1830 & n1997 ) | ( ~n1996 & n1997 ) ;
  assign n1999 = ( ~n1150 & n1993 ) | ( ~n1150 & n1998 ) | ( n1993 & n1998 ) ;
  assign n2000 = ~n1150 & n1831 ;
  assign n2001 = ( ~n1150 & n1831 ) | ( ~n1150 & n1949 ) | ( n1831 & n1949 ) ;
  assign n2002 = ( ~n1836 & n2000 ) | ( ~n1836 & n2001 ) | ( n2000 & n2001 ) ;
  assign n2003 = ( n1836 & n2000 ) | ( n1836 & n2001 ) | ( n2000 & n2001 ) ;
  assign n2004 = ( n1836 & n2002 ) | ( n1836 & ~n2003 ) | ( n2002 & ~n2003 ) ;
  assign n2005 = ( ~n1038 & n1999 ) | ( ~n1038 & n2004 ) | ( n1999 & n2004 ) ;
  assign n2006 = ~n1038 & n1837 ;
  assign n2007 = ( ~n1038 & n1837 ) | ( ~n1038 & n1949 ) | ( n1837 & n1949 ) ;
  assign n2008 = ( n1842 & n2006 ) | ( n1842 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2009 = ( ~n1842 & n2006 ) | ( ~n1842 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2010 = ( n1842 & ~n2008 ) | ( n1842 & n2009 ) | ( ~n2008 & n2009 ) ;
  assign n2011 = ( ~n933 & n2005 ) | ( ~n933 & n2010 ) | ( n2005 & n2010 ) ;
  assign n2012 = ( n933 & ~n1843 ) | ( n933 & n1949 ) | ( ~n1843 & n1949 ) ;
  assign n2013 = n933 & ~n1843 ;
  assign n2014 = ( n1848 & n2012 ) | ( n1848 & n2013 ) | ( n2012 & n2013 ) ;
  assign n2015 = ( ~n1848 & n2012 ) | ( ~n1848 & n2013 ) | ( n2012 & n2013 ) ;
  assign n2016 = ( n1848 & ~n2014 ) | ( n1848 & n2015 ) | ( ~n2014 & n2015 ) ;
  assign n2017 = ( ~n839 & n2011 ) | ( ~n839 & n2016 ) | ( n2011 & n2016 ) ;
  assign n2018 = ( n839 & ~n1849 ) | ( n839 & n1949 ) | ( ~n1849 & n1949 ) ;
  assign n2019 = n839 & ~n1849 ;
  assign n2020 = ( n1854 & n2018 ) | ( n1854 & n2019 ) | ( n2018 & n2019 ) ;
  assign n2021 = ( ~n1854 & n2018 ) | ( ~n1854 & n2019 ) | ( n2018 & n2019 ) ;
  assign n2022 = ( n1854 & ~n2020 ) | ( n1854 & n2021 ) | ( ~n2020 & n2021 ) ;
  assign n2023 = ( ~n746 & n2017 ) | ( ~n746 & n2022 ) | ( n2017 & n2022 ) ;
  assign n2024 = ( n746 & ~n1855 ) | ( n746 & n1949 ) | ( ~n1855 & n1949 ) ;
  assign n2025 = n746 & ~n1855 ;
  assign n2026 = ( n1860 & n2024 ) | ( n1860 & n2025 ) | ( n2024 & n2025 ) ;
  assign n2027 = ( ~n1860 & n2024 ) | ( ~n1860 & n2025 ) | ( n2024 & n2025 ) ;
  assign n2028 = ( n1860 & ~n2026 ) | ( n1860 & n2027 ) | ( ~n2026 & n2027 ) ;
  assign n2029 = ( ~n664 & n2023 ) | ( ~n664 & n2028 ) | ( n2023 & n2028 ) ;
  assign n2030 = n664 & ~n1861 ;
  assign n2031 = ( n664 & ~n1861 ) | ( n664 & n1949 ) | ( ~n1861 & n1949 ) ;
  assign n2032 = ( n1866 & n2030 ) | ( n1866 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2033 = ( ~n1866 & n2030 ) | ( ~n1866 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2034 = ( n1866 & ~n2032 ) | ( n1866 & n2033 ) | ( ~n2032 & n2033 ) ;
  assign n2035 = ( ~n588 & n2029 ) | ( ~n588 & n2034 ) | ( n2029 & n2034 ) ;
  assign n2036 = ( n588 & ~n1867 ) | ( n588 & n1949 ) | ( ~n1867 & n1949 ) ;
  assign n2037 = n588 & ~n1867 ;
  assign n2038 = ( n1872 & n2036 ) | ( n1872 & n2037 ) | ( n2036 & n2037 ) ;
  assign n2039 = ( ~n1872 & n2036 ) | ( ~n1872 & n2037 ) | ( n2036 & n2037 ) ;
  assign n2040 = ( n1872 & ~n2038 ) | ( n1872 & n2039 ) | ( ~n2038 & n2039 ) ;
  assign n2041 = ( ~n518 & n2035 ) | ( ~n518 & n2040 ) | ( n2035 & n2040 ) ;
  assign n2042 = ( n518 & ~n1873 ) | ( n518 & n1949 ) | ( ~n1873 & n1949 ) ;
  assign n2043 = n518 & ~n1873 ;
  assign n2044 = ( n1878 & n2042 ) | ( n1878 & n2043 ) | ( n2042 & n2043 ) ;
  assign n2045 = ( ~n1878 & n2042 ) | ( ~n1878 & n2043 ) | ( n2042 & n2043 ) ;
  assign n2046 = ( n1878 & ~n2044 ) | ( n1878 & n2045 ) | ( ~n2044 & n2045 ) ;
  assign n2047 = ( ~n454 & n2041 ) | ( ~n454 & n2046 ) | ( n2041 & n2046 ) ;
  assign n2048 = ~n454 & n1879 ;
  assign n2049 = ( ~n454 & n1879 ) | ( ~n454 & n1949 ) | ( n1879 & n1949 ) ;
  assign n2050 = ( n1884 & n2048 ) | ( n1884 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2051 = ( ~n1884 & n2048 ) | ( ~n1884 & n2049 ) | ( n2048 & n2049 ) ;
  assign n2052 = ( n1884 & ~n2050 ) | ( n1884 & n2051 ) | ( ~n2050 & n2051 ) ;
  assign n2053 = ( ~n396 & n2047 ) | ( ~n396 & n2052 ) | ( n2047 & n2052 ) ;
  assign n2054 = n396 & ~n1885 ;
  assign n2055 = ( n396 & ~n1885 ) | ( n396 & n1949 ) | ( ~n1885 & n1949 ) ;
  assign n2056 = ( n1890 & n2054 ) | ( n1890 & n2055 ) | ( n2054 & n2055 ) ;
  assign n2057 = ( ~n1890 & n2054 ) | ( ~n1890 & n2055 ) | ( n2054 & n2055 ) ;
  assign n2058 = ( n1890 & ~n2056 ) | ( n1890 & n2057 ) | ( ~n2056 & n2057 ) ;
  assign n2059 = ( ~n344 & n2053 ) | ( ~n344 & n2058 ) | ( n2053 & n2058 ) ;
  assign n2060 = ( n344 & ~n1891 ) | ( n344 & n1949 ) | ( ~n1891 & n1949 ) ;
  assign n2061 = n344 & ~n1891 ;
  assign n2062 = ( n1896 & n2060 ) | ( n1896 & n2061 ) | ( n2060 & n2061 ) ;
  assign n2063 = ( ~n1896 & n2060 ) | ( ~n1896 & n2061 ) | ( n2060 & n2061 ) ;
  assign n2064 = ( n1896 & ~n2062 ) | ( n1896 & n2063 ) | ( ~n2062 & n2063 ) ;
  assign n2065 = ( ~n298 & n2059 ) | ( ~n298 & n2064 ) | ( n2059 & n2064 ) ;
  assign n2066 = ( n298 & ~n1897 ) | ( n298 & n1949 ) | ( ~n1897 & n1949 ) ;
  assign n2067 = n298 & ~n1897 ;
  assign n2068 = ( n1902 & n2066 ) | ( n1902 & n2067 ) | ( n2066 & n2067 ) ;
  assign n2069 = ( ~n1902 & n2066 ) | ( ~n1902 & n2067 ) | ( n2066 & n2067 ) ;
  assign n2070 = ( n1902 & ~n2068 ) | ( n1902 & n2069 ) | ( ~n2068 & n2069 ) ;
  assign n2071 = ( ~n258 & n2065 ) | ( ~n258 & n2070 ) | ( n2065 & n2070 ) ;
  assign n2072 = ( n258 & ~n1903 ) | ( n258 & n1949 ) | ( ~n1903 & n1949 ) ;
  assign n2073 = n258 & ~n1903 ;
  assign n2074 = ( n1908 & n2072 ) | ( n1908 & n2073 ) | ( n2072 & n2073 ) ;
  assign n2075 = ( ~n1908 & n2072 ) | ( ~n1908 & n2073 ) | ( n2072 & n2073 ) ;
  assign n2076 = ( n1908 & ~n2074 ) | ( n1908 & n2075 ) | ( ~n2074 & n2075 ) ;
  assign n2077 = ( ~n225 & n2071 ) | ( ~n225 & n2076 ) | ( n2071 & n2076 ) ;
  assign n2078 = n225 & ~n1909 ;
  assign n2079 = ( n225 & ~n1909 ) | ( n225 & n1949 ) | ( ~n1909 & n1949 ) ;
  assign n2080 = ( ~n1914 & n2078 ) | ( ~n1914 & n2079 ) | ( n2078 & n2079 ) ;
  assign n2081 = ( n1914 & n2078 ) | ( n1914 & n2079 ) | ( n2078 & n2079 ) ;
  assign n2082 = ( n1914 & n2080 ) | ( n1914 & ~n2081 ) | ( n2080 & ~n2081 ) ;
  assign n2083 = ( ~n197 & n2077 ) | ( ~n197 & n2082 ) | ( n2077 & n2082 ) ;
  assign n2084 = ~n197 & n1915 ;
  assign n2085 = ( ~n197 & n1915 ) | ( ~n197 & n1949 ) | ( n1915 & n1949 ) ;
  assign n2086 = ( n1920 & n2084 ) | ( n1920 & n2085 ) | ( n2084 & n2085 ) ;
  assign n2087 = ( ~n1920 & n2084 ) | ( ~n1920 & n2085 ) | ( n2084 & n2085 ) ;
  assign n2088 = ( n1920 & ~n2086 ) | ( n1920 & n2087 ) | ( ~n2086 & n2087 ) ;
  assign n2089 = ( ~n170 & n2083 ) | ( ~n170 & n2088 ) | ( n2083 & n2088 ) ;
  assign n2090 = ( n170 & ~n1921 ) | ( n170 & n1949 ) | ( ~n1921 & n1949 ) ;
  assign n2091 = n170 & ~n1921 ;
  assign n2092 = ( n1926 & n2090 ) | ( n1926 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2093 = ( ~n1926 & n2090 ) | ( ~n1926 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2094 = ( n1926 & ~n2092 ) | ( n1926 & n2093 ) | ( ~n2092 & n2093 ) ;
  assign n2095 = ( ~n142 & n2089 ) | ( ~n142 & n2094 ) | ( n2089 & n2094 ) ;
  assign n2096 = ( ~n132 & n1954 ) | ( ~n132 & n2095 ) | ( n1954 & n2095 ) ;
  assign n2097 = ( n131 & n1939 ) | ( n131 & ~n1944 ) | ( n1939 & ~n1944 ) ;
  assign n2098 = n1806 & ~n1944 ;
  assign n2099 = n1939 & n2098 ;
  assign n2100 = ( n131 & ~n2097 ) | ( n131 & n2099 ) | ( ~n2097 & n2099 ) ;
  assign n2101 = ~n132 & n1933 ;
  assign n2102 = ( ~n132 & n1933 ) | ( ~n132 & n1949 ) | ( n1933 & n1949 ) ;
  assign n2103 = ( ~n1938 & n2101 ) | ( ~n1938 & n2102 ) | ( n2101 & n2102 ) ;
  assign n2104 = ( n1938 & n2101 ) | ( n1938 & n2102 ) | ( n2101 & n2102 ) ;
  assign n2105 = ( n1938 & n2103 ) | ( n1938 & ~n2104 ) | ( n2103 & ~n2104 ) ;
  assign n2106 = ( n1939 & ~n1944 ) | ( n1939 & n1946 ) | ( ~n1944 & n1946 ) ;
  assign n2107 = ~n2097 & n2106 ;
  assign n2108 = ( n2100 & ~n2105 ) | ( n2100 & n2107 ) | ( ~n2105 & n2107 ) ;
  assign n2109 = ( ~n2096 & n2100 ) | ( ~n2096 & n2108 ) | ( n2100 & n2108 ) ;
  assign n2110 = ( ~n131 & n2096 ) | ( ~n131 & n2105 ) | ( n2096 & n2105 ) ;
  assign n2111 = n2109 | n2110 ;
  assign n2112 = ( ~n132 & n2095 ) | ( ~n132 & n2111 ) | ( n2095 & n2111 ) ;
  assign n2113 = ~n132 & n2095 ;
  assign n2114 = ( n1954 & n2112 ) | ( n1954 & ~n2113 ) | ( n2112 & ~n2113 ) ;
  assign n2115 = ( ~n1954 & n2112 ) | ( ~n1954 & n2113 ) | ( n2112 & n2113 ) ;
  assign n2116 = ( ~n2112 & n2114 ) | ( ~n2112 & n2115 ) | ( n2114 & n2115 ) ;
  assign n2117 = x77 | n2111 ;
  assign n2118 = x74 | x75 ;
  assign n2119 = x76 | n2118 ;
  assign n2120 = n1949 & ~n2119 ;
  assign n2121 = n2117 & ~n2120 ;
  assign n2122 = n1969 & n2111 ;
  assign n2123 = x77 & n2111 ;
  assign n2124 = ~n1949 & n2119 ;
  assign n2125 = ( ~n2117 & n2123 ) | ( ~n2117 & n2124 ) | ( n2123 & n2124 ) ;
  assign n2126 = ( n2121 & ~n2122 ) | ( n2121 & n2125 ) | ( ~n2122 & n2125 ) ;
  assign n2127 = n1949 | n2111 ;
  assign n2128 = ( ~x78 & n2122 ) | ( ~x78 & n2127 ) | ( n2122 & n2127 ) ;
  assign n2129 = ( x78 & n2122 ) | ( x78 & n2127 ) | ( n2122 & n2127 ) ;
  assign n2130 = ( x78 & n2128 ) | ( x78 & ~n2129 ) | ( n2128 & ~n2129 ) ;
  assign n2131 = ( ~n1802 & n2126 ) | ( ~n1802 & n2130 ) | ( n2126 & n2130 ) ;
  assign n2132 = ( x79 & n1949 ) | ( x79 & ~n1967 ) | ( n1949 & ~n1967 ) ;
  assign n2133 = ( ~x79 & n1809 ) | ( ~x79 & n1969 ) | ( n1809 & n1969 ) ;
  assign n2134 = ( n1968 & ~n1975 ) | ( n1968 & n2133 ) | ( ~n1975 & n2133 ) ;
  assign n2135 = ( n1802 & n1974 ) | ( n1802 & ~n2134 ) | ( n1974 & ~n2134 ) ;
  assign n2136 = n2111 & ~n2135 ;
  assign n2137 = ~n1971 & n1973 ;
  assign n2138 = ~x78 & n1971 ;
  assign n2139 = ( n1972 & n1976 ) | ( n1972 & n2138 ) | ( n1976 & n2138 ) ;
  assign n2140 = ( n2111 & n2138 ) | ( n2111 & n2139 ) | ( n2138 & n2139 ) ;
  assign n2141 = ~n2137 & n2140 ;
  assign n2142 = ( n2132 & n2136 ) | ( n2132 & ~n2141 ) | ( n2136 & ~n2141 ) ;
  assign n2143 = ( ~n1661 & n2131 ) | ( ~n1661 & n2142 ) | ( n2131 & n2142 ) ;
  assign n2144 = n1661 & ~n1976 ;
  assign n2145 = ( n1661 & ~n1976 ) | ( n1661 & n2111 ) | ( ~n1976 & n2111 ) ;
  assign n2146 = ( n1979 & n2144 ) | ( n1979 & n2145 ) | ( n2144 & n2145 ) ;
  assign n2147 = ( ~n1979 & n2144 ) | ( ~n1979 & n2145 ) | ( n2144 & n2145 ) ;
  assign n2148 = ( n1979 & ~n2146 ) | ( n1979 & n2147 ) | ( ~n2146 & n2147 ) ;
  assign n2149 = ( ~n1523 & n2143 ) | ( ~n1523 & n2148 ) | ( n2143 & n2148 ) ;
  assign n2150 = n1523 & ~n1980 ;
  assign n2151 = ( n1523 & ~n1980 ) | ( n1523 & n2111 ) | ( ~n1980 & n2111 ) ;
  assign n2152 = ( ~n1966 & n2150 ) | ( ~n1966 & n2151 ) | ( n2150 & n2151 ) ;
  assign n2153 = ( n1966 & n2150 ) | ( n1966 & n2151 ) | ( n2150 & n2151 ) ;
  assign n2154 = ( n1966 & n2152 ) | ( n1966 & ~n2153 ) | ( n2152 & ~n2153 ) ;
  assign n2155 = ( ~n1393 & n2149 ) | ( ~n1393 & n2154 ) | ( n2149 & n2154 ) ;
  assign n2156 = ( n1393 & ~n1981 ) | ( n1393 & n2111 ) | ( ~n1981 & n2111 ) ;
  assign n2157 = n1393 & ~n1981 ;
  assign n2158 = ( n1986 & n2156 ) | ( n1986 & n2157 ) | ( n2156 & n2157 ) ;
  assign n2159 = ( ~n1986 & n2156 ) | ( ~n1986 & n2157 ) | ( n2156 & n2157 ) ;
  assign n2160 = ( n1986 & ~n2158 ) | ( n1986 & n2159 ) | ( ~n2158 & n2159 ) ;
  assign n2161 = ( ~n1266 & n2155 ) | ( ~n1266 & n2160 ) | ( n2155 & n2160 ) ;
  assign n2162 = ( n1266 & ~n1987 ) | ( n1266 & n2111 ) | ( ~n1987 & n2111 ) ;
  assign n2163 = n1266 & ~n1987 ;
  assign n2164 = ( n1992 & n2162 ) | ( n1992 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2165 = ( ~n1992 & n2162 ) | ( ~n1992 & n2163 ) | ( n2162 & n2163 ) ;
  assign n2166 = ( n1992 & ~n2164 ) | ( n1992 & n2165 ) | ( ~n2164 & n2165 ) ;
  assign n2167 = ( ~n1150 & n2161 ) | ( ~n1150 & n2166 ) | ( n2161 & n2166 ) ;
  assign n2168 = ( n1150 & ~n1993 ) | ( n1150 & n2111 ) | ( ~n1993 & n2111 ) ;
  assign n2169 = n1150 & ~n1993 ;
  assign n2170 = ( n1998 & n2168 ) | ( n1998 & n2169 ) | ( n2168 & n2169 ) ;
  assign n2171 = ( ~n1998 & n2168 ) | ( ~n1998 & n2169 ) | ( n2168 & n2169 ) ;
  assign n2172 = ( n1998 & ~n2170 ) | ( n1998 & n2171 ) | ( ~n2170 & n2171 ) ;
  assign n2173 = ( ~n1038 & n2167 ) | ( ~n1038 & n2172 ) | ( n2167 & n2172 ) ;
  assign n2174 = n1038 & ~n1999 ;
  assign n2175 = ( n1038 & ~n1999 ) | ( n1038 & n2111 ) | ( ~n1999 & n2111 ) ;
  assign n2176 = ( n2004 & n2174 ) | ( n2004 & n2175 ) | ( n2174 & n2175 ) ;
  assign n2177 = ( ~n2004 & n2174 ) | ( ~n2004 & n2175 ) | ( n2174 & n2175 ) ;
  assign n2178 = ( n2004 & ~n2176 ) | ( n2004 & n2177 ) | ( ~n2176 & n2177 ) ;
  assign n2179 = ( ~n933 & n2173 ) | ( ~n933 & n2178 ) | ( n2173 & n2178 ) ;
  assign n2180 = ( n933 & ~n2005 ) | ( n933 & n2111 ) | ( ~n2005 & n2111 ) ;
  assign n2181 = n933 & ~n2005 ;
  assign n2182 = ( n2010 & n2180 ) | ( n2010 & n2181 ) | ( n2180 & n2181 ) ;
  assign n2183 = ( ~n2010 & n2180 ) | ( ~n2010 & n2181 ) | ( n2180 & n2181 ) ;
  assign n2184 = ( n2010 & ~n2182 ) | ( n2010 & n2183 ) | ( ~n2182 & n2183 ) ;
  assign n2185 = ( ~n839 & n2179 ) | ( ~n839 & n2184 ) | ( n2179 & n2184 ) ;
  assign n2186 = n839 & ~n2011 ;
  assign n2187 = ( n839 & ~n2011 ) | ( n839 & n2111 ) | ( ~n2011 & n2111 ) ;
  assign n2188 = ( n2016 & n2186 ) | ( n2016 & n2187 ) | ( n2186 & n2187 ) ;
  assign n2189 = ( ~n2016 & n2186 ) | ( ~n2016 & n2187 ) | ( n2186 & n2187 ) ;
  assign n2190 = ( n2016 & ~n2188 ) | ( n2016 & n2189 ) | ( ~n2188 & n2189 ) ;
  assign n2191 = ( ~n746 & n2185 ) | ( ~n746 & n2190 ) | ( n2185 & n2190 ) ;
  assign n2192 = ( n746 & ~n2017 ) | ( n746 & n2111 ) | ( ~n2017 & n2111 ) ;
  assign n2193 = n746 & ~n2017 ;
  assign n2194 = ( n2022 & n2192 ) | ( n2022 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2195 = ( ~n2022 & n2192 ) | ( ~n2022 & n2193 ) | ( n2192 & n2193 ) ;
  assign n2196 = ( n2022 & ~n2194 ) | ( n2022 & n2195 ) | ( ~n2194 & n2195 ) ;
  assign n2197 = ( ~n664 & n2191 ) | ( ~n664 & n2196 ) | ( n2191 & n2196 ) ;
  assign n2198 = ( n664 & ~n2023 ) | ( n664 & n2111 ) | ( ~n2023 & n2111 ) ;
  assign n2199 = n664 & ~n2023 ;
  assign n2200 = ( n2028 & n2198 ) | ( n2028 & n2199 ) | ( n2198 & n2199 ) ;
  assign n2201 = ( ~n2028 & n2198 ) | ( ~n2028 & n2199 ) | ( n2198 & n2199 ) ;
  assign n2202 = ( n2028 & ~n2200 ) | ( n2028 & n2201 ) | ( ~n2200 & n2201 ) ;
  assign n2203 = ( ~n588 & n2197 ) | ( ~n588 & n2202 ) | ( n2197 & n2202 ) ;
  assign n2204 = ( n588 & ~n2029 ) | ( n588 & n2111 ) | ( ~n2029 & n2111 ) ;
  assign n2205 = n588 & ~n2029 ;
  assign n2206 = ( n2034 & n2204 ) | ( n2034 & n2205 ) | ( n2204 & n2205 ) ;
  assign n2207 = ( ~n2034 & n2204 ) | ( ~n2034 & n2205 ) | ( n2204 & n2205 ) ;
  assign n2208 = ( n2034 & ~n2206 ) | ( n2034 & n2207 ) | ( ~n2206 & n2207 ) ;
  assign n2209 = ( ~n518 & n2203 ) | ( ~n518 & n2208 ) | ( n2203 & n2208 ) ;
  assign n2210 = ~n518 & n2035 ;
  assign n2211 = ( ~n518 & n2035 ) | ( ~n518 & n2111 ) | ( n2035 & n2111 ) ;
  assign n2212 = ( ~n2040 & n2210 ) | ( ~n2040 & n2211 ) | ( n2210 & n2211 ) ;
  assign n2213 = ( n2040 & n2210 ) | ( n2040 & n2211 ) | ( n2210 & n2211 ) ;
  assign n2214 = ( n2040 & n2212 ) | ( n2040 & ~n2213 ) | ( n2212 & ~n2213 ) ;
  assign n2215 = ( ~n454 & n2209 ) | ( ~n454 & n2214 ) | ( n2209 & n2214 ) ;
  assign n2216 = ( n454 & ~n2041 ) | ( n454 & n2111 ) | ( ~n2041 & n2111 ) ;
  assign n2217 = n454 & ~n2041 ;
  assign n2218 = ( n2046 & n2216 ) | ( n2046 & n2217 ) | ( n2216 & n2217 ) ;
  assign n2219 = ( ~n2046 & n2216 ) | ( ~n2046 & n2217 ) | ( n2216 & n2217 ) ;
  assign n2220 = ( n2046 & ~n2218 ) | ( n2046 & n2219 ) | ( ~n2218 & n2219 ) ;
  assign n2221 = ( ~n396 & n2215 ) | ( ~n396 & n2220 ) | ( n2215 & n2220 ) ;
  assign n2222 = ~n396 & n2047 ;
  assign n2223 = ( ~n396 & n2047 ) | ( ~n396 & n2111 ) | ( n2047 & n2111 ) ;
  assign n2224 = ( n2052 & n2222 ) | ( n2052 & n2223 ) | ( n2222 & n2223 ) ;
  assign n2225 = ( ~n2052 & n2222 ) | ( ~n2052 & n2223 ) | ( n2222 & n2223 ) ;
  assign n2226 = ( n2052 & ~n2224 ) | ( n2052 & n2225 ) | ( ~n2224 & n2225 ) ;
  assign n2227 = ( ~n344 & n2221 ) | ( ~n344 & n2226 ) | ( n2221 & n2226 ) ;
  assign n2228 = ~n344 & n2053 ;
  assign n2229 = ( ~n344 & n2053 ) | ( ~n344 & n2111 ) | ( n2053 & n2111 ) ;
  assign n2230 = ( n2058 & n2228 ) | ( n2058 & n2229 ) | ( n2228 & n2229 ) ;
  assign n2231 = ( ~n2058 & n2228 ) | ( ~n2058 & n2229 ) | ( n2228 & n2229 ) ;
  assign n2232 = ( n2058 & ~n2230 ) | ( n2058 & n2231 ) | ( ~n2230 & n2231 ) ;
  assign n2233 = ( ~n298 & n2227 ) | ( ~n298 & n2232 ) | ( n2227 & n2232 ) ;
  assign n2234 = ( n298 & ~n2059 ) | ( n298 & n2111 ) | ( ~n2059 & n2111 ) ;
  assign n2235 = n298 & ~n2059 ;
  assign n2236 = ( n2064 & n2234 ) | ( n2064 & n2235 ) | ( n2234 & n2235 ) ;
  assign n2237 = ( ~n2064 & n2234 ) | ( ~n2064 & n2235 ) | ( n2234 & n2235 ) ;
  assign n2238 = ( n2064 & ~n2236 ) | ( n2064 & n2237 ) | ( ~n2236 & n2237 ) ;
  assign n2239 = ( ~n258 & n2233 ) | ( ~n258 & n2238 ) | ( n2233 & n2238 ) ;
  assign n2240 = ~n258 & n2065 ;
  assign n2241 = ( ~n258 & n2065 ) | ( ~n258 & n2111 ) | ( n2065 & n2111 ) ;
  assign n2242 = ( n2070 & n2240 ) | ( n2070 & n2241 ) | ( n2240 & n2241 ) ;
  assign n2243 = ( ~n2070 & n2240 ) | ( ~n2070 & n2241 ) | ( n2240 & n2241 ) ;
  assign n2244 = ( n2070 & ~n2242 ) | ( n2070 & n2243 ) | ( ~n2242 & n2243 ) ;
  assign n2245 = ( ~n225 & n2239 ) | ( ~n225 & n2244 ) | ( n2239 & n2244 ) ;
  assign n2246 = n225 & ~n2071 ;
  assign n2247 = ( n225 & ~n2071 ) | ( n225 & n2111 ) | ( ~n2071 & n2111 ) ;
  assign n2248 = ( n2076 & n2246 ) | ( n2076 & n2247 ) | ( n2246 & n2247 ) ;
  assign n2249 = ( ~n2076 & n2246 ) | ( ~n2076 & n2247 ) | ( n2246 & n2247 ) ;
  assign n2250 = ( n2076 & ~n2248 ) | ( n2076 & n2249 ) | ( ~n2248 & n2249 ) ;
  assign n2251 = ( ~n197 & n2245 ) | ( ~n197 & n2250 ) | ( n2245 & n2250 ) ;
  assign n2252 = ~n197 & n2077 ;
  assign n2253 = ( ~n197 & n2077 ) | ( ~n197 & n2111 ) | ( n2077 & n2111 ) ;
  assign n2254 = ( ~n2082 & n2252 ) | ( ~n2082 & n2253 ) | ( n2252 & n2253 ) ;
  assign n2255 = ( n2082 & n2252 ) | ( n2082 & n2253 ) | ( n2252 & n2253 ) ;
  assign n2256 = ( n2082 & n2254 ) | ( n2082 & ~n2255 ) | ( n2254 & ~n2255 ) ;
  assign n2257 = ( ~n170 & n2251 ) | ( ~n170 & n2256 ) | ( n2251 & n2256 ) ;
  assign n2258 = ~n170 & n2083 ;
  assign n2259 = ( ~n170 & n2083 ) | ( ~n170 & n2111 ) | ( n2083 & n2111 ) ;
  assign n2260 = ( n2088 & n2258 ) | ( n2088 & n2259 ) | ( n2258 & n2259 ) ;
  assign n2261 = ( ~n2088 & n2258 ) | ( ~n2088 & n2259 ) | ( n2258 & n2259 ) ;
  assign n2262 = ( n2088 & ~n2260 ) | ( n2088 & n2261 ) | ( ~n2260 & n2261 ) ;
  assign n2263 = ( ~n142 & n2257 ) | ( ~n142 & n2262 ) | ( n2257 & n2262 ) ;
  assign n2264 = ( n142 & ~n2089 ) | ( n142 & n2111 ) | ( ~n2089 & n2111 ) ;
  assign n2265 = n142 & ~n2089 ;
  assign n2266 = ( n2094 & n2264 ) | ( n2094 & n2265 ) | ( n2264 & n2265 ) ;
  assign n2267 = ( ~n2094 & n2264 ) | ( ~n2094 & n2265 ) | ( n2264 & n2265 ) ;
  assign n2268 = ( n2094 & ~n2266 ) | ( n2094 & n2267 ) | ( ~n2266 & n2267 ) ;
  assign n2269 = ( ~n132 & n2263 ) | ( ~n132 & n2268 ) | ( n2263 & n2268 ) ;
  assign n2270 = ( n2096 & n2100 ) | ( n2096 & n2105 ) | ( n2100 & n2105 ) ;
  assign n2271 = n2109 | n2270 ;
  assign n2272 = n2116 & ~n2269 ;
  assign n2273 = ( n2269 & n2271 ) | ( n2269 & ~n2272 ) | ( n2271 & ~n2272 ) ;
  assign n2274 = ( ~n131 & n2116 ) | ( ~n131 & n2273 ) | ( n2116 & n2273 ) ;
  assign n2275 = n2105 & ~n2110 ;
  assign n2276 = ( ~n2110 & n2270 ) | ( ~n2110 & n2275 ) | ( n2270 & n2275 ) ;
  assign n2277 = n2274 | n2276 ;
  assign n2278 = ( n131 & ~n2116 ) | ( n131 & n2269 ) | ( ~n2116 & n2269 ) ;
  assign n2279 = n2273 & ~n2278 ;
  assign n2280 = ( n131 & n2116 ) | ( n131 & ~n2276 ) | ( n2116 & ~n2276 ) ;
  assign n2281 = n2269 & ~n2280 ;
  assign n2282 = ( n131 & n2272 ) | ( n131 & n2281 ) | ( n2272 & n2281 ) ;
  assign n2283 = n2279 | n2282 ;
  assign n2284 = ~x75 & n2277 ;
  assign n2285 = x74 & n2284 ;
  assign n2286 = x75 & ~n2277 ;
  assign n2287 = n2284 | n2286 ;
  assign n2288 = x72 | x73 ;
  assign n2289 = x74 | n2288 ;
  assign n2290 = ( ~n2111 & n2287 ) | ( ~n2111 & n2289 ) | ( n2287 & n2289 ) ;
  assign n2291 = ~n2285 & n2290 ;
  assign n2292 = n2118 & n2277 ;
  assign n2293 = n2111 | n2277 ;
  assign n2294 = ( x76 & n2292 ) | ( x76 & n2293 ) | ( n2292 & n2293 ) ;
  assign n2295 = ( x76 & ~n2292 ) | ( x76 & n2293 ) | ( ~n2292 & n2293 ) ;
  assign n2296 = ( n2292 & ~n2294 ) | ( n2292 & n2295 ) | ( ~n2294 & n2295 ) ;
  assign n2297 = ( ~n1949 & n2291 ) | ( ~n1949 & n2296 ) | ( n2291 & n2296 ) ;
  assign n2298 = ~n2124 & n2277 ;
  assign n2299 = ( n2120 & n2124 ) | ( n2120 & n2277 ) | ( n2124 & n2277 ) ;
  assign n2300 = ( n2294 & n2298 ) | ( n2294 & ~n2299 ) | ( n2298 & ~n2299 ) ;
  assign n2301 = ( x77 & n2111 ) | ( x77 & n2300 ) | ( n2111 & n2300 ) ;
  assign n2302 = ( ~x77 & n2111 ) | ( ~x77 & n2300 ) | ( n2111 & n2300 ) ;
  assign n2303 = ( x77 & ~n2301 ) | ( x77 & n2302 ) | ( ~n2301 & n2302 ) ;
  assign n2304 = ( ~n1802 & n2297 ) | ( ~n1802 & n2303 ) | ( n2297 & n2303 ) ;
  assign n2305 = ~n1802 & n2126 ;
  assign n2306 = ( ~n1802 & n2126 ) | ( ~n1802 & n2277 ) | ( n2126 & n2277 ) ;
  assign n2307 = ( n2130 & n2305 ) | ( n2130 & n2306 ) | ( n2305 & n2306 ) ;
  assign n2308 = ( ~n2130 & n2305 ) | ( ~n2130 & n2306 ) | ( n2305 & n2306 ) ;
  assign n2309 = ( n2130 & ~n2307 ) | ( n2130 & n2308 ) | ( ~n2307 & n2308 ) ;
  assign n2310 = ( ~n1661 & n2304 ) | ( ~n1661 & n2309 ) | ( n2304 & n2309 ) ;
  assign n2311 = ( n1661 & ~n2131 ) | ( n1661 & n2277 ) | ( ~n2131 & n2277 ) ;
  assign n2312 = n1661 & ~n2131 ;
  assign n2313 = ( n2142 & n2311 ) | ( n2142 & n2312 ) | ( n2311 & n2312 ) ;
  assign n2314 = ( ~n2142 & n2311 ) | ( ~n2142 & n2312 ) | ( n2311 & n2312 ) ;
  assign n2315 = ( n2142 & ~n2313 ) | ( n2142 & n2314 ) | ( ~n2313 & n2314 ) ;
  assign n2316 = ( ~n1523 & n2310 ) | ( ~n1523 & n2315 ) | ( n2310 & n2315 ) ;
  assign n2317 = ( n1523 & ~n2143 ) | ( n1523 & n2277 ) | ( ~n2143 & n2277 ) ;
  assign n2318 = n1523 & ~n2143 ;
  assign n2319 = ( n2148 & n2317 ) | ( n2148 & n2318 ) | ( n2317 & n2318 ) ;
  assign n2320 = ( ~n2148 & n2317 ) | ( ~n2148 & n2318 ) | ( n2317 & n2318 ) ;
  assign n2321 = ( n2148 & ~n2319 ) | ( n2148 & n2320 ) | ( ~n2319 & n2320 ) ;
  assign n2322 = ( ~n1393 & n2316 ) | ( ~n1393 & n2321 ) | ( n2316 & n2321 ) ;
  assign n2323 = ~n1393 & n2149 ;
  assign n2324 = ( ~n1393 & n2149 ) | ( ~n1393 & n2277 ) | ( n2149 & n2277 ) ;
  assign n2325 = ( ~n2154 & n2323 ) | ( ~n2154 & n2324 ) | ( n2323 & n2324 ) ;
  assign n2326 = ( n2154 & n2323 ) | ( n2154 & n2324 ) | ( n2323 & n2324 ) ;
  assign n2327 = ( n2154 & n2325 ) | ( n2154 & ~n2326 ) | ( n2325 & ~n2326 ) ;
  assign n2328 = ( ~n1266 & n2322 ) | ( ~n1266 & n2327 ) | ( n2322 & n2327 ) ;
  assign n2329 = ~n1266 & n2155 ;
  assign n2330 = ( ~n1266 & n2155 ) | ( ~n1266 & n2277 ) | ( n2155 & n2277 ) ;
  assign n2331 = ( ~n2160 & n2329 ) | ( ~n2160 & n2330 ) | ( n2329 & n2330 ) ;
  assign n2332 = ( n2160 & n2329 ) | ( n2160 & n2330 ) | ( n2329 & n2330 ) ;
  assign n2333 = ( n2160 & n2331 ) | ( n2160 & ~n2332 ) | ( n2331 & ~n2332 ) ;
  assign n2334 = ( ~n1150 & n2328 ) | ( ~n1150 & n2333 ) | ( n2328 & n2333 ) ;
  assign n2335 = ( n1150 & ~n2161 ) | ( n1150 & n2277 ) | ( ~n2161 & n2277 ) ;
  assign n2336 = n1150 & ~n2161 ;
  assign n2337 = ( n2166 & n2335 ) | ( n2166 & n2336 ) | ( n2335 & n2336 ) ;
  assign n2338 = ( ~n2166 & n2335 ) | ( ~n2166 & n2336 ) | ( n2335 & n2336 ) ;
  assign n2339 = ( n2166 & ~n2337 ) | ( n2166 & n2338 ) | ( ~n2337 & n2338 ) ;
  assign n2340 = ( ~n1038 & n2334 ) | ( ~n1038 & n2339 ) | ( n2334 & n2339 ) ;
  assign n2341 = ~n1038 & n2167 ;
  assign n2342 = ( ~n1038 & n2167 ) | ( ~n1038 & n2277 ) | ( n2167 & n2277 ) ;
  assign n2343 = ( ~n2172 & n2341 ) | ( ~n2172 & n2342 ) | ( n2341 & n2342 ) ;
  assign n2344 = ( n2172 & n2341 ) | ( n2172 & n2342 ) | ( n2341 & n2342 ) ;
  assign n2345 = ( n2172 & n2343 ) | ( n2172 & ~n2344 ) | ( n2343 & ~n2344 ) ;
  assign n2346 = ( ~n933 & n2340 ) | ( ~n933 & n2345 ) | ( n2340 & n2345 ) ;
  assign n2347 = ~n933 & n2173 ;
  assign n2348 = ( ~n933 & n2173 ) | ( ~n933 & n2277 ) | ( n2173 & n2277 ) ;
  assign n2349 = ( ~n2178 & n2347 ) | ( ~n2178 & n2348 ) | ( n2347 & n2348 ) ;
  assign n2350 = ( n2178 & n2347 ) | ( n2178 & n2348 ) | ( n2347 & n2348 ) ;
  assign n2351 = ( n2178 & n2349 ) | ( n2178 & ~n2350 ) | ( n2349 & ~n2350 ) ;
  assign n2352 = ( ~n839 & n2346 ) | ( ~n839 & n2351 ) | ( n2346 & n2351 ) ;
  assign n2353 = ~n839 & n2179 ;
  assign n2354 = ( ~n839 & n2179 ) | ( ~n839 & n2277 ) | ( n2179 & n2277 ) ;
  assign n2355 = ( ~n2184 & n2353 ) | ( ~n2184 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2356 = ( n2184 & n2353 ) | ( n2184 & n2354 ) | ( n2353 & n2354 ) ;
  assign n2357 = ( n2184 & n2355 ) | ( n2184 & ~n2356 ) | ( n2355 & ~n2356 ) ;
  assign n2358 = ( ~n746 & n2352 ) | ( ~n746 & n2357 ) | ( n2352 & n2357 ) ;
  assign n2359 = ( n746 & ~n2185 ) | ( n746 & n2277 ) | ( ~n2185 & n2277 ) ;
  assign n2360 = n746 & ~n2185 ;
  assign n2361 = ( n2190 & n2359 ) | ( n2190 & n2360 ) | ( n2359 & n2360 ) ;
  assign n2362 = ( ~n2190 & n2359 ) | ( ~n2190 & n2360 ) | ( n2359 & n2360 ) ;
  assign n2363 = ( n2190 & ~n2361 ) | ( n2190 & n2362 ) | ( ~n2361 & n2362 ) ;
  assign n2364 = ( ~n664 & n2358 ) | ( ~n664 & n2363 ) | ( n2358 & n2363 ) ;
  assign n2365 = ( n664 & ~n2191 ) | ( n664 & n2277 ) | ( ~n2191 & n2277 ) ;
  assign n2366 = n664 & ~n2191 ;
  assign n2367 = ( n2196 & n2365 ) | ( n2196 & n2366 ) | ( n2365 & n2366 ) ;
  assign n2368 = ( ~n2196 & n2365 ) | ( ~n2196 & n2366 ) | ( n2365 & n2366 ) ;
  assign n2369 = ( n2196 & ~n2367 ) | ( n2196 & n2368 ) | ( ~n2367 & n2368 ) ;
  assign n2370 = ( ~n588 & n2364 ) | ( ~n588 & n2369 ) | ( n2364 & n2369 ) ;
  assign n2371 = n588 & ~n2197 ;
  assign n2372 = ( n588 & ~n2197 ) | ( n588 & n2277 ) | ( ~n2197 & n2277 ) ;
  assign n2373 = ( n2202 & n2371 ) | ( n2202 & n2372 ) | ( n2371 & n2372 ) ;
  assign n2374 = ( ~n2202 & n2371 ) | ( ~n2202 & n2372 ) | ( n2371 & n2372 ) ;
  assign n2375 = ( n2202 & ~n2373 ) | ( n2202 & n2374 ) | ( ~n2373 & n2374 ) ;
  assign n2376 = ( ~n518 & n2370 ) | ( ~n518 & n2375 ) | ( n2370 & n2375 ) ;
  assign n2377 = ( n518 & ~n2203 ) | ( n518 & n2277 ) | ( ~n2203 & n2277 ) ;
  assign n2378 = n518 & ~n2203 ;
  assign n2379 = ( n2208 & n2377 ) | ( n2208 & n2378 ) | ( n2377 & n2378 ) ;
  assign n2380 = ( ~n2208 & n2377 ) | ( ~n2208 & n2378 ) | ( n2377 & n2378 ) ;
  assign n2381 = ( n2208 & ~n2379 ) | ( n2208 & n2380 ) | ( ~n2379 & n2380 ) ;
  assign n2382 = ( ~n454 & n2376 ) | ( ~n454 & n2381 ) | ( n2376 & n2381 ) ;
  assign n2383 = ~n454 & n2209 ;
  assign n2384 = ( ~n454 & n2209 ) | ( ~n454 & n2277 ) | ( n2209 & n2277 ) ;
  assign n2385 = ( ~n2214 & n2383 ) | ( ~n2214 & n2384 ) | ( n2383 & n2384 ) ;
  assign n2386 = ( n2214 & n2383 ) | ( n2214 & n2384 ) | ( n2383 & n2384 ) ;
  assign n2387 = ( n2214 & n2385 ) | ( n2214 & ~n2386 ) | ( n2385 & ~n2386 ) ;
  assign n2388 = ( ~n396 & n2382 ) | ( ~n396 & n2387 ) | ( n2382 & n2387 ) ;
  assign n2389 = ~n396 & n2215 ;
  assign n2390 = ( ~n396 & n2215 ) | ( ~n396 & n2277 ) | ( n2215 & n2277 ) ;
  assign n2391 = ( n2220 & n2389 ) | ( n2220 & n2390 ) | ( n2389 & n2390 ) ;
  assign n2392 = ( ~n2220 & n2389 ) | ( ~n2220 & n2390 ) | ( n2389 & n2390 ) ;
  assign n2393 = ( n2220 & ~n2391 ) | ( n2220 & n2392 ) | ( ~n2391 & n2392 ) ;
  assign n2394 = ( ~n344 & n2388 ) | ( ~n344 & n2393 ) | ( n2388 & n2393 ) ;
  assign n2395 = ( n344 & ~n2221 ) | ( n344 & n2277 ) | ( ~n2221 & n2277 ) ;
  assign n2396 = n344 & ~n2221 ;
  assign n2397 = ( n2226 & n2395 ) | ( n2226 & n2396 ) | ( n2395 & n2396 ) ;
  assign n2398 = ( ~n2226 & n2395 ) | ( ~n2226 & n2396 ) | ( n2395 & n2396 ) ;
  assign n2399 = ( n2226 & ~n2397 ) | ( n2226 & n2398 ) | ( ~n2397 & n2398 ) ;
  assign n2400 = ( ~n298 & n2394 ) | ( ~n298 & n2399 ) | ( n2394 & n2399 ) ;
  assign n2401 = ~n298 & n2227 ;
  assign n2402 = ( ~n298 & n2227 ) | ( ~n298 & n2277 ) | ( n2227 & n2277 ) ;
  assign n2403 = ( n2232 & n2401 ) | ( n2232 & n2402 ) | ( n2401 & n2402 ) ;
  assign n2404 = ( ~n2232 & n2401 ) | ( ~n2232 & n2402 ) | ( n2401 & n2402 ) ;
  assign n2405 = ( n2232 & ~n2403 ) | ( n2232 & n2404 ) | ( ~n2403 & n2404 ) ;
  assign n2406 = ( ~n258 & n2400 ) | ( ~n258 & n2405 ) | ( n2400 & n2405 ) ;
  assign n2407 = ( n258 & ~n2233 ) | ( n258 & n2277 ) | ( ~n2233 & n2277 ) ;
  assign n2408 = n258 & ~n2233 ;
  assign n2409 = ( n2238 & n2407 ) | ( n2238 & n2408 ) | ( n2407 & n2408 ) ;
  assign n2410 = ( ~n2238 & n2407 ) | ( ~n2238 & n2408 ) | ( n2407 & n2408 ) ;
  assign n2411 = ( n2238 & ~n2409 ) | ( n2238 & n2410 ) | ( ~n2409 & n2410 ) ;
  assign n2412 = ( ~n225 & n2406 ) | ( ~n225 & n2411 ) | ( n2406 & n2411 ) ;
  assign n2413 = ( n225 & ~n2239 ) | ( n225 & n2277 ) | ( ~n2239 & n2277 ) ;
  assign n2414 = n225 & ~n2239 ;
  assign n2415 = ( n2244 & n2413 ) | ( n2244 & n2414 ) | ( n2413 & n2414 ) ;
  assign n2416 = ( ~n2244 & n2413 ) | ( ~n2244 & n2414 ) | ( n2413 & n2414 ) ;
  assign n2417 = ( n2244 & ~n2415 ) | ( n2244 & n2416 ) | ( ~n2415 & n2416 ) ;
  assign n2418 = ( ~n197 & n2412 ) | ( ~n197 & n2417 ) | ( n2412 & n2417 ) ;
  assign n2419 = ( n197 & ~n2245 ) | ( n197 & n2277 ) | ( ~n2245 & n2277 ) ;
  assign n2420 = n197 & ~n2245 ;
  assign n2421 = ( n2250 & n2419 ) | ( n2250 & n2420 ) | ( n2419 & n2420 ) ;
  assign n2422 = ( ~n2250 & n2419 ) | ( ~n2250 & n2420 ) | ( n2419 & n2420 ) ;
  assign n2423 = ( n2250 & ~n2421 ) | ( n2250 & n2422 ) | ( ~n2421 & n2422 ) ;
  assign n2424 = ( ~n170 & n2418 ) | ( ~n170 & n2423 ) | ( n2418 & n2423 ) ;
  assign n2425 = ( n170 & ~n2251 ) | ( n170 & n2277 ) | ( ~n2251 & n2277 ) ;
  assign n2426 = n170 & ~n2251 ;
  assign n2427 = ( n2256 & n2425 ) | ( n2256 & n2426 ) | ( n2425 & n2426 ) ;
  assign n2428 = ( ~n2256 & n2425 ) | ( ~n2256 & n2426 ) | ( n2425 & n2426 ) ;
  assign n2429 = ( n2256 & ~n2427 ) | ( n2256 & n2428 ) | ( ~n2427 & n2428 ) ;
  assign n2430 = ( ~n142 & n2424 ) | ( ~n142 & n2429 ) | ( n2424 & n2429 ) ;
  assign n2431 = ( n142 & ~n2257 ) | ( n142 & n2277 ) | ( ~n2257 & n2277 ) ;
  assign n2432 = n142 & ~n2257 ;
  assign n2433 = ( n2262 & n2431 ) | ( n2262 & n2432 ) | ( n2431 & n2432 ) ;
  assign n2434 = ( ~n2262 & n2431 ) | ( ~n2262 & n2432 ) | ( n2431 & n2432 ) ;
  assign n2435 = ( n2262 & ~n2433 ) | ( n2262 & n2434 ) | ( ~n2433 & n2434 ) ;
  assign n2436 = ( ~n132 & n2430 ) | ( ~n132 & n2435 ) | ( n2430 & n2435 ) ;
  assign n2437 = ( n132 & ~n2263 ) | ( n132 & n2277 ) | ( ~n2263 & n2277 ) ;
  assign n2438 = n132 & ~n2263 ;
  assign n2439 = ( n2268 & n2437 ) | ( n2268 & n2438 ) | ( n2437 & n2438 ) ;
  assign n2440 = ( ~n2268 & n2437 ) | ( ~n2268 & n2438 ) | ( n2437 & n2438 ) ;
  assign n2441 = ( n2268 & ~n2439 ) | ( n2268 & n2440 ) | ( ~n2439 & n2440 ) ;
  assign n2442 = ( ~n131 & n2436 ) | ( ~n131 & n2441 ) | ( n2436 & n2441 ) ;
  assign n2443 = n2283 | n2442 ;
  assign n2444 = x70 | x71 ;
  assign n2445 = x72 | n2444 ;
  assign n2446 = x73 | n2443 ;
  assign n2447 = ( ~n2277 & n2445 ) | ( ~n2277 & n2446 ) | ( n2445 & n2446 ) ;
  assign n2448 = n2288 & n2443 ;
  assign n2449 = ( ~x73 & n2277 ) | ( ~x73 & n2445 ) | ( n2277 & n2445 ) ;
  assign n2450 = n2445 & ~n2449 ;
  assign n2451 = ( n2447 & ~n2448 ) | ( n2447 & n2450 ) | ( ~n2448 & n2450 ) ;
  assign n2452 = n2277 | n2443 ;
  assign n2453 = ( x74 & n2448 ) | ( x74 & n2452 ) | ( n2448 & n2452 ) ;
  assign n2454 = ( ~x74 & n2448 ) | ( ~x74 & n2452 ) | ( n2448 & n2452 ) ;
  assign n2455 = ( x74 & ~n2453 ) | ( x74 & n2454 ) | ( ~n2453 & n2454 ) ;
  assign n2456 = ( ~n2111 & n2451 ) | ( ~n2111 & n2455 ) | ( n2451 & n2455 ) ;
  assign n2457 = x74 & ~x75 ;
  assign n2458 = ( n2111 & n2287 ) | ( n2111 & n2289 ) | ( n2287 & n2289 ) ;
  assign n2459 = ( n2111 & n2290 ) | ( n2111 & ~n2458 ) | ( n2290 & ~n2458 ) ;
  assign n2460 = n2443 & ~n2459 ;
  assign n2461 = x74 | n2287 ;
  assign n2462 = ( ~n2443 & n2457 ) | ( ~n2443 & n2461 ) | ( n2457 & n2461 ) ;
  assign n2463 = ( ~n2457 & n2460 ) | ( ~n2457 & n2462 ) | ( n2460 & n2462 ) ;
  assign n2464 = ( ~n1949 & n2456 ) | ( ~n1949 & n2463 ) | ( n2456 & n2463 ) ;
  assign n2465 = n1949 & ~n2291 ;
  assign n2466 = ( n1949 & ~n2291 ) | ( n1949 & n2443 ) | ( ~n2291 & n2443 ) ;
  assign n2467 = ( ~n2296 & n2465 ) | ( ~n2296 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2468 = ( n2296 & n2465 ) | ( n2296 & n2466 ) | ( n2465 & n2466 ) ;
  assign n2469 = ( n2296 & n2467 ) | ( n2296 & ~n2468 ) | ( n2467 & ~n2468 ) ;
  assign n2470 = ( ~n1802 & n2464 ) | ( ~n1802 & n2469 ) | ( n2464 & n2469 ) ;
  assign n2471 = ( n1802 & ~n2297 ) | ( n1802 & n2443 ) | ( ~n2297 & n2443 ) ;
  assign n2472 = n1802 & ~n2297 ;
  assign n2473 = ( n2303 & n2471 ) | ( n2303 & n2472 ) | ( n2471 & n2472 ) ;
  assign n2474 = ( ~n2303 & n2471 ) | ( ~n2303 & n2472 ) | ( n2471 & n2472 ) ;
  assign n2475 = ( n2303 & ~n2473 ) | ( n2303 & n2474 ) | ( ~n2473 & n2474 ) ;
  assign n2476 = ( ~n1661 & n2470 ) | ( ~n1661 & n2475 ) | ( n2470 & n2475 ) ;
  assign n2477 = ( n1661 & ~n2304 ) | ( n1661 & n2443 ) | ( ~n2304 & n2443 ) ;
  assign n2478 = n1661 & ~n2304 ;
  assign n2479 = ( n2309 & n2477 ) | ( n2309 & n2478 ) | ( n2477 & n2478 ) ;
  assign n2480 = ( ~n2309 & n2477 ) | ( ~n2309 & n2478 ) | ( n2477 & n2478 ) ;
  assign n2481 = ( n2309 & ~n2479 ) | ( n2309 & n2480 ) | ( ~n2479 & n2480 ) ;
  assign n2482 = ( ~n1523 & n2476 ) | ( ~n1523 & n2481 ) | ( n2476 & n2481 ) ;
  assign n2483 = ( n1523 & ~n2310 ) | ( n1523 & n2443 ) | ( ~n2310 & n2443 ) ;
  assign n2484 = n1523 & ~n2310 ;
  assign n2485 = ( n2315 & n2483 ) | ( n2315 & n2484 ) | ( n2483 & n2484 ) ;
  assign n2486 = ( ~n2315 & n2483 ) | ( ~n2315 & n2484 ) | ( n2483 & n2484 ) ;
  assign n2487 = ( n2315 & ~n2485 ) | ( n2315 & n2486 ) | ( ~n2485 & n2486 ) ;
  assign n2488 = ( ~n1393 & n2482 ) | ( ~n1393 & n2487 ) | ( n2482 & n2487 ) ;
  assign n2489 = ~n1393 & n2316 ;
  assign n2490 = ( ~n1393 & n2316 ) | ( ~n1393 & n2443 ) | ( n2316 & n2443 ) ;
  assign n2491 = ( n2321 & n2489 ) | ( n2321 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2492 = ( ~n2321 & n2489 ) | ( ~n2321 & n2490 ) | ( n2489 & n2490 ) ;
  assign n2493 = ( n2321 & ~n2491 ) | ( n2321 & n2492 ) | ( ~n2491 & n2492 ) ;
  assign n2494 = ( ~n1266 & n2488 ) | ( ~n1266 & n2493 ) | ( n2488 & n2493 ) ;
  assign n2495 = ( n1266 & ~n2322 ) | ( n1266 & n2443 ) | ( ~n2322 & n2443 ) ;
  assign n2496 = n1266 & ~n2322 ;
  assign n2497 = ( n2327 & n2495 ) | ( n2327 & n2496 ) | ( n2495 & n2496 ) ;
  assign n2498 = ( ~n2327 & n2495 ) | ( ~n2327 & n2496 ) | ( n2495 & n2496 ) ;
  assign n2499 = ( n2327 & ~n2497 ) | ( n2327 & n2498 ) | ( ~n2497 & n2498 ) ;
  assign n2500 = ( ~n1150 & n2494 ) | ( ~n1150 & n2499 ) | ( n2494 & n2499 ) ;
  assign n2501 = ~n1150 & n2328 ;
  assign n2502 = ( ~n1150 & n2328 ) | ( ~n1150 & n2443 ) | ( n2328 & n2443 ) ;
  assign n2503 = ( ~n2333 & n2501 ) | ( ~n2333 & n2502 ) | ( n2501 & n2502 ) ;
  assign n2504 = ( n2333 & n2501 ) | ( n2333 & n2502 ) | ( n2501 & n2502 ) ;
  assign n2505 = ( n2333 & n2503 ) | ( n2333 & ~n2504 ) | ( n2503 & ~n2504 ) ;
  assign n2506 = ( ~n1038 & n2500 ) | ( ~n1038 & n2505 ) | ( n2500 & n2505 ) ;
  assign n2507 = ( n1038 & ~n2334 ) | ( n1038 & n2443 ) | ( ~n2334 & n2443 ) ;
  assign n2508 = n1038 & ~n2334 ;
  assign n2509 = ( n2339 & n2507 ) | ( n2339 & n2508 ) | ( n2507 & n2508 ) ;
  assign n2510 = ( ~n2339 & n2507 ) | ( ~n2339 & n2508 ) | ( n2507 & n2508 ) ;
  assign n2511 = ( n2339 & ~n2509 ) | ( n2339 & n2510 ) | ( ~n2509 & n2510 ) ;
  assign n2512 = ( ~n933 & n2506 ) | ( ~n933 & n2511 ) | ( n2506 & n2511 ) ;
  assign n2513 = ~n933 & n2340 ;
  assign n2514 = ( ~n933 & n2340 ) | ( ~n933 & n2443 ) | ( n2340 & n2443 ) ;
  assign n2515 = ( n2345 & n2513 ) | ( n2345 & n2514 ) | ( n2513 & n2514 ) ;
  assign n2516 = ( ~n2345 & n2513 ) | ( ~n2345 & n2514 ) | ( n2513 & n2514 ) ;
  assign n2517 = ( n2345 & ~n2515 ) | ( n2345 & n2516 ) | ( ~n2515 & n2516 ) ;
  assign n2518 = ( ~n839 & n2512 ) | ( ~n839 & n2517 ) | ( n2512 & n2517 ) ;
  assign n2519 = ~n839 & n2346 ;
  assign n2520 = ( ~n839 & n2346 ) | ( ~n839 & n2443 ) | ( n2346 & n2443 ) ;
  assign n2521 = ( n2351 & n2519 ) | ( n2351 & n2520 ) | ( n2519 & n2520 ) ;
  assign n2522 = ( ~n2351 & n2519 ) | ( ~n2351 & n2520 ) | ( n2519 & n2520 ) ;
  assign n2523 = ( n2351 & ~n2521 ) | ( n2351 & n2522 ) | ( ~n2521 & n2522 ) ;
  assign n2524 = ( ~n746 & n2518 ) | ( ~n746 & n2523 ) | ( n2518 & n2523 ) ;
  assign n2525 = ( n746 & ~n2352 ) | ( n746 & n2443 ) | ( ~n2352 & n2443 ) ;
  assign n2526 = n746 & ~n2352 ;
  assign n2527 = ( n2357 & n2525 ) | ( n2357 & n2526 ) | ( n2525 & n2526 ) ;
  assign n2528 = ( ~n2357 & n2525 ) | ( ~n2357 & n2526 ) | ( n2525 & n2526 ) ;
  assign n2529 = ( n2357 & ~n2527 ) | ( n2357 & n2528 ) | ( ~n2527 & n2528 ) ;
  assign n2530 = ( ~n664 & n2524 ) | ( ~n664 & n2529 ) | ( n2524 & n2529 ) ;
  assign n2531 = ( n664 & ~n2358 ) | ( n664 & n2443 ) | ( ~n2358 & n2443 ) ;
  assign n2532 = n664 & ~n2358 ;
  assign n2533 = ( n2363 & n2531 ) | ( n2363 & n2532 ) | ( n2531 & n2532 ) ;
  assign n2534 = ( ~n2363 & n2531 ) | ( ~n2363 & n2532 ) | ( n2531 & n2532 ) ;
  assign n2535 = ( n2363 & ~n2533 ) | ( n2363 & n2534 ) | ( ~n2533 & n2534 ) ;
  assign n2536 = ( ~n588 & n2530 ) | ( ~n588 & n2535 ) | ( n2530 & n2535 ) ;
  assign n2537 = ~n588 & n2364 ;
  assign n2538 = ( ~n588 & n2364 ) | ( ~n588 & n2443 ) | ( n2364 & n2443 ) ;
  assign n2539 = ( ~n2369 & n2537 ) | ( ~n2369 & n2538 ) | ( n2537 & n2538 ) ;
  assign n2540 = ( n2369 & n2537 ) | ( n2369 & n2538 ) | ( n2537 & n2538 ) ;
  assign n2541 = ( n2369 & n2539 ) | ( n2369 & ~n2540 ) | ( n2539 & ~n2540 ) ;
  assign n2542 = ( ~n518 & n2536 ) | ( ~n518 & n2541 ) | ( n2536 & n2541 ) ;
  assign n2543 = n518 & ~n2370 ;
  assign n2544 = ( n518 & ~n2370 ) | ( n518 & n2443 ) | ( ~n2370 & n2443 ) ;
  assign n2545 = ( n2375 & n2543 ) | ( n2375 & n2544 ) | ( n2543 & n2544 ) ;
  assign n2546 = ( ~n2375 & n2543 ) | ( ~n2375 & n2544 ) | ( n2543 & n2544 ) ;
  assign n2547 = ( n2375 & ~n2545 ) | ( n2375 & n2546 ) | ( ~n2545 & n2546 ) ;
  assign n2548 = ( ~n454 & n2542 ) | ( ~n454 & n2547 ) | ( n2542 & n2547 ) ;
  assign n2549 = ~n454 & n2376 ;
  assign n2550 = ( ~n454 & n2376 ) | ( ~n454 & n2443 ) | ( n2376 & n2443 ) ;
  assign n2551 = ( ~n2381 & n2549 ) | ( ~n2381 & n2550 ) | ( n2549 & n2550 ) ;
  assign n2552 = ( n2381 & n2549 ) | ( n2381 & n2550 ) | ( n2549 & n2550 ) ;
  assign n2553 = ( n2381 & n2551 ) | ( n2381 & ~n2552 ) | ( n2551 & ~n2552 ) ;
  assign n2554 = ( ~n396 & n2548 ) | ( ~n396 & n2553 ) | ( n2548 & n2553 ) ;
  assign n2555 = ( n396 & ~n2382 ) | ( n396 & n2443 ) | ( ~n2382 & n2443 ) ;
  assign n2556 = n396 & ~n2382 ;
  assign n2557 = ( n2387 & n2555 ) | ( n2387 & n2556 ) | ( n2555 & n2556 ) ;
  assign n2558 = ( ~n2387 & n2555 ) | ( ~n2387 & n2556 ) | ( n2555 & n2556 ) ;
  assign n2559 = ( n2387 & ~n2557 ) | ( n2387 & n2558 ) | ( ~n2557 & n2558 ) ;
  assign n2560 = ( ~n344 & n2554 ) | ( ~n344 & n2559 ) | ( n2554 & n2559 ) ;
  assign n2561 = ~n344 & n2388 ;
  assign n2562 = ( ~n344 & n2388 ) | ( ~n344 & n2443 ) | ( n2388 & n2443 ) ;
  assign n2563 = ( n2393 & n2561 ) | ( n2393 & n2562 ) | ( n2561 & n2562 ) ;
  assign n2564 = ( ~n2393 & n2561 ) | ( ~n2393 & n2562 ) | ( n2561 & n2562 ) ;
  assign n2565 = ( n2393 & ~n2563 ) | ( n2393 & n2564 ) | ( ~n2563 & n2564 ) ;
  assign n2566 = ( ~n298 & n2560 ) | ( ~n298 & n2565 ) | ( n2560 & n2565 ) ;
  assign n2567 = ~n298 & n2394 ;
  assign n2568 = ( ~n298 & n2394 ) | ( ~n298 & n2443 ) | ( n2394 & n2443 ) ;
  assign n2569 = ( ~n2399 & n2567 ) | ( ~n2399 & n2568 ) | ( n2567 & n2568 ) ;
  assign n2570 = ( n2399 & n2567 ) | ( n2399 & n2568 ) | ( n2567 & n2568 ) ;
  assign n2571 = ( n2399 & n2569 ) | ( n2399 & ~n2570 ) | ( n2569 & ~n2570 ) ;
  assign n2572 = ( ~n258 & n2566 ) | ( ~n258 & n2571 ) | ( n2566 & n2571 ) ;
  assign n2573 = ( n258 & ~n2400 ) | ( n258 & n2443 ) | ( ~n2400 & n2443 ) ;
  assign n2574 = n258 & ~n2400 ;
  assign n2575 = ( n2405 & n2573 ) | ( n2405 & n2574 ) | ( n2573 & n2574 ) ;
  assign n2576 = ( ~n2405 & n2573 ) | ( ~n2405 & n2574 ) | ( n2573 & n2574 ) ;
  assign n2577 = ( n2405 & ~n2575 ) | ( n2405 & n2576 ) | ( ~n2575 & n2576 ) ;
  assign n2578 = ( ~n225 & n2572 ) | ( ~n225 & n2577 ) | ( n2572 & n2577 ) ;
  assign n2579 = ( n225 & ~n2406 ) | ( n225 & n2443 ) | ( ~n2406 & n2443 ) ;
  assign n2580 = n225 & ~n2406 ;
  assign n2581 = ( n2411 & n2579 ) | ( n2411 & n2580 ) | ( n2579 & n2580 ) ;
  assign n2582 = ( ~n2411 & n2579 ) | ( ~n2411 & n2580 ) | ( n2579 & n2580 ) ;
  assign n2583 = ( n2411 & ~n2581 ) | ( n2411 & n2582 ) | ( ~n2581 & n2582 ) ;
  assign n2584 = ( ~n197 & n2578 ) | ( ~n197 & n2583 ) | ( n2578 & n2583 ) ;
  assign n2585 = ( n197 & ~n2412 ) | ( n197 & n2443 ) | ( ~n2412 & n2443 ) ;
  assign n2586 = n197 & ~n2412 ;
  assign n2587 = ( n2417 & n2585 ) | ( n2417 & n2586 ) | ( n2585 & n2586 ) ;
  assign n2588 = ( ~n2417 & n2585 ) | ( ~n2417 & n2586 ) | ( n2585 & n2586 ) ;
  assign n2589 = ( n2417 & ~n2587 ) | ( n2417 & n2588 ) | ( ~n2587 & n2588 ) ;
  assign n2590 = ( ~n170 & n2584 ) | ( ~n170 & n2589 ) | ( n2584 & n2589 ) ;
  assign n2591 = ~n170 & n2418 ;
  assign n2592 = ( ~n170 & n2418 ) | ( ~n170 & n2443 ) | ( n2418 & n2443 ) ;
  assign n2593 = ( n2423 & n2591 ) | ( n2423 & n2592 ) | ( n2591 & n2592 ) ;
  assign n2594 = ( ~n2423 & n2591 ) | ( ~n2423 & n2592 ) | ( n2591 & n2592 ) ;
  assign n2595 = ( n2423 & ~n2593 ) | ( n2423 & n2594 ) | ( ~n2593 & n2594 ) ;
  assign n2596 = ( ~n142 & n2590 ) | ( ~n142 & n2595 ) | ( n2590 & n2595 ) ;
  assign n2597 = ~n142 & n2424 ;
  assign n2598 = ( ~n142 & n2424 ) | ( ~n142 & n2443 ) | ( n2424 & n2443 ) ;
  assign n2599 = ( n2429 & n2597 ) | ( n2429 & n2598 ) | ( n2597 & n2598 ) ;
  assign n2600 = ( ~n2429 & n2597 ) | ( ~n2429 & n2598 ) | ( n2597 & n2598 ) ;
  assign n2601 = ( n2429 & ~n2599 ) | ( n2429 & n2600 ) | ( ~n2599 & n2600 ) ;
  assign n2602 = ( ~n132 & n2596 ) | ( ~n132 & n2601 ) | ( n2596 & n2601 ) ;
  assign n2603 = ( ~n132 & n2430 ) | ( ~n132 & n2443 ) | ( n2430 & n2443 ) ;
  assign n2604 = ~n132 & n2430 ;
  assign n2605 = ( ~n2435 & n2603 ) | ( ~n2435 & n2604 ) | ( n2603 & n2604 ) ;
  assign n2606 = ( n2435 & n2603 ) | ( n2435 & n2604 ) | ( n2603 & n2604 ) ;
  assign n2607 = ( n2435 & n2605 ) | ( n2435 & ~n2606 ) | ( n2605 & ~n2606 ) ;
  assign n2608 = ( ~n131 & n2602 ) | ( ~n131 & n2607 ) | ( n2602 & n2607 ) ;
  assign n2609 = n131 | n2436 ;
  assign n2610 = ( n131 & n2436 ) | ( n131 & ~n2441 ) | ( n2436 & ~n2441 ) ;
  assign n2611 = n2279 & ~n2436 ;
  assign n2612 = n2282 & n2436 ;
  assign n2613 = ( ~n2441 & n2611 ) | ( ~n2441 & n2612 ) | ( n2611 & n2612 ) ;
  assign n2614 = ( n2609 & ~n2610 ) | ( n2609 & n2613 ) | ( ~n2610 & n2613 ) ;
  assign n2615 = n2608 | n2614 ;
  assign n2616 = ~n2607 & n2614 ;
  assign n2617 = ( ~n131 & n2602 ) | ( ~n131 & n2616 ) | ( n2602 & n2616 ) ;
  assign n2618 = ( n2607 & ~n2608 ) | ( n2607 & n2617 ) | ( ~n2608 & n2617 ) ;
  assign n2619 = x68 | x69 ;
  assign n2620 = x70 | n2619 ;
  assign n2621 = ~n2443 & n2620 ;
  assign n2622 = ( x71 & ~n2615 ) | ( x71 & n2621 ) | ( ~n2615 & n2621 ) ;
  assign n2623 = ~n2444 & n2615 ;
  assign n2624 = n2443 & ~n2620 ;
  assign n2625 = ( n2622 & n2623 ) | ( n2622 & ~n2624 ) | ( n2623 & ~n2624 ) ;
  assign n2626 = n2443 & ~n2615 ;
  assign n2627 = ( x72 & n2623 ) | ( x72 & n2626 ) | ( n2623 & n2626 ) ;
  assign n2628 = ( ~x72 & n2623 ) | ( ~x72 & n2626 ) | ( n2623 & n2626 ) ;
  assign n2629 = ( x72 & ~n2627 ) | ( x72 & n2628 ) | ( ~n2627 & n2628 ) ;
  assign n2630 = ( ~n2277 & n2625 ) | ( ~n2277 & n2629 ) | ( n2625 & n2629 ) ;
  assign n2631 = ( n2277 & n2443 ) | ( n2277 & n2445 ) | ( n2443 & n2445 ) ;
  assign n2632 = ( n2277 & n2443 ) | ( n2277 & ~n2615 ) | ( n2443 & ~n2615 ) ;
  assign n2633 = n2631 & ~n2632 ;
  assign n2634 = ( n2443 & n2445 ) | ( n2443 & n2615 ) | ( n2445 & n2615 ) ;
  assign n2635 = n2277 | n2634 ;
  assign n2636 = ( n2628 & n2631 ) | ( n2628 & ~n2635 ) | ( n2631 & ~n2635 ) ;
  assign n2637 = ( x73 & n2633 ) | ( x73 & n2636 ) | ( n2633 & n2636 ) ;
  assign n2638 = ( ~x73 & n2633 ) | ( ~x73 & n2636 ) | ( n2633 & n2636 ) ;
  assign n2639 = ( x73 & ~n2637 ) | ( x73 & n2638 ) | ( ~n2637 & n2638 ) ;
  assign n2640 = ( ~n2111 & n2630 ) | ( ~n2111 & n2639 ) | ( n2630 & n2639 ) ;
  assign n2641 = n2111 & ~n2451 ;
  assign n2642 = ( n2111 & ~n2451 ) | ( n2111 & n2615 ) | ( ~n2451 & n2615 ) ;
  assign n2643 = ( n2455 & n2641 ) | ( n2455 & n2642 ) | ( n2641 & n2642 ) ;
  assign n2644 = ( ~n2455 & n2641 ) | ( ~n2455 & n2642 ) | ( n2641 & n2642 ) ;
  assign n2645 = ( n2455 & ~n2643 ) | ( n2455 & n2644 ) | ( ~n2643 & n2644 ) ;
  assign n2646 = ( ~n1949 & n2640 ) | ( ~n1949 & n2645 ) | ( n2640 & n2645 ) ;
  assign n2647 = ~n1949 & n2456 ;
  assign n2648 = ( ~n1949 & n2456 ) | ( ~n1949 & n2615 ) | ( n2456 & n2615 ) ;
  assign n2649 = ( ~n2463 & n2647 ) | ( ~n2463 & n2648 ) | ( n2647 & n2648 ) ;
  assign n2650 = ( n2463 & n2647 ) | ( n2463 & n2648 ) | ( n2647 & n2648 ) ;
  assign n2651 = ( n2463 & n2649 ) | ( n2463 & ~n2650 ) | ( n2649 & ~n2650 ) ;
  assign n2652 = ( ~n1802 & n2646 ) | ( ~n1802 & n2651 ) | ( n2646 & n2651 ) ;
  assign n2653 = ( n1802 & ~n2464 ) | ( n1802 & n2615 ) | ( ~n2464 & n2615 ) ;
  assign n2654 = n1802 & ~n2464 ;
  assign n2655 = ( n2469 & n2653 ) | ( n2469 & n2654 ) | ( n2653 & n2654 ) ;
  assign n2656 = ( ~n2469 & n2653 ) | ( ~n2469 & n2654 ) | ( n2653 & n2654 ) ;
  assign n2657 = ( n2469 & ~n2655 ) | ( n2469 & n2656 ) | ( ~n2655 & n2656 ) ;
  assign n2658 = ( ~n1661 & n2652 ) | ( ~n1661 & n2657 ) | ( n2652 & n2657 ) ;
  assign n2659 = ( n1661 & ~n2470 ) | ( n1661 & n2615 ) | ( ~n2470 & n2615 ) ;
  assign n2660 = n1661 & ~n2470 ;
  assign n2661 = ( n2475 & n2659 ) | ( n2475 & n2660 ) | ( n2659 & n2660 ) ;
  assign n2662 = ( ~n2475 & n2659 ) | ( ~n2475 & n2660 ) | ( n2659 & n2660 ) ;
  assign n2663 = ( n2475 & ~n2661 ) | ( n2475 & n2662 ) | ( ~n2661 & n2662 ) ;
  assign n2664 = ( ~n1523 & n2658 ) | ( ~n1523 & n2663 ) | ( n2658 & n2663 ) ;
  assign n2665 = ~n1523 & n2476 ;
  assign n2666 = ( ~n1523 & n2476 ) | ( ~n1523 & n2615 ) | ( n2476 & n2615 ) ;
  assign n2667 = ( ~n2481 & n2665 ) | ( ~n2481 & n2666 ) | ( n2665 & n2666 ) ;
  assign n2668 = ( n2481 & n2665 ) | ( n2481 & n2666 ) | ( n2665 & n2666 ) ;
  assign n2669 = ( n2481 & n2667 ) | ( n2481 & ~n2668 ) | ( n2667 & ~n2668 ) ;
  assign n2670 = ( ~n1393 & n2664 ) | ( ~n1393 & n2669 ) | ( n2664 & n2669 ) ;
  assign n2671 = ( n1393 & ~n2482 ) | ( n1393 & n2615 ) | ( ~n2482 & n2615 ) ;
  assign n2672 = n1393 & ~n2482 ;
  assign n2673 = ( n2487 & n2671 ) | ( n2487 & n2672 ) | ( n2671 & n2672 ) ;
  assign n2674 = ( ~n2487 & n2671 ) | ( ~n2487 & n2672 ) | ( n2671 & n2672 ) ;
  assign n2675 = ( n2487 & ~n2673 ) | ( n2487 & n2674 ) | ( ~n2673 & n2674 ) ;
  assign n2676 = ( ~n1266 & n2670 ) | ( ~n1266 & n2675 ) | ( n2670 & n2675 ) ;
  assign n2677 = ( n1266 & ~n2488 ) | ( n1266 & n2615 ) | ( ~n2488 & n2615 ) ;
  assign n2678 = n1266 & ~n2488 ;
  assign n2679 = ( n2493 & n2677 ) | ( n2493 & n2678 ) | ( n2677 & n2678 ) ;
  assign n2680 = ( ~n2493 & n2677 ) | ( ~n2493 & n2678 ) | ( n2677 & n2678 ) ;
  assign n2681 = ( n2493 & ~n2679 ) | ( n2493 & n2680 ) | ( ~n2679 & n2680 ) ;
  assign n2682 = ( ~n1150 & n2676 ) | ( ~n1150 & n2681 ) | ( n2676 & n2681 ) ;
  assign n2683 = ( n1150 & ~n2494 ) | ( n1150 & n2615 ) | ( ~n2494 & n2615 ) ;
  assign n2684 = n1150 & ~n2494 ;
  assign n2685 = ( n2499 & n2683 ) | ( n2499 & n2684 ) | ( n2683 & n2684 ) ;
  assign n2686 = ( ~n2499 & n2683 ) | ( ~n2499 & n2684 ) | ( n2683 & n2684 ) ;
  assign n2687 = ( n2499 & ~n2685 ) | ( n2499 & n2686 ) | ( ~n2685 & n2686 ) ;
  assign n2688 = ( ~n1038 & n2682 ) | ( ~n1038 & n2687 ) | ( n2682 & n2687 ) ;
  assign n2689 = ( n1038 & ~n2500 ) | ( n1038 & n2615 ) | ( ~n2500 & n2615 ) ;
  assign n2690 = n1038 & ~n2500 ;
  assign n2691 = ( n2505 & n2689 ) | ( n2505 & n2690 ) | ( n2689 & n2690 ) ;
  assign n2692 = ( ~n2505 & n2689 ) | ( ~n2505 & n2690 ) | ( n2689 & n2690 ) ;
  assign n2693 = ( n2505 & ~n2691 ) | ( n2505 & n2692 ) | ( ~n2691 & n2692 ) ;
  assign n2694 = ( ~n933 & n2688 ) | ( ~n933 & n2693 ) | ( n2688 & n2693 ) ;
  assign n2695 = ~n933 & n2506 ;
  assign n2696 = ( ~n933 & n2506 ) | ( ~n933 & n2615 ) | ( n2506 & n2615 ) ;
  assign n2697 = ( ~n2511 & n2695 ) | ( ~n2511 & n2696 ) | ( n2695 & n2696 ) ;
  assign n2698 = ( n2511 & n2695 ) | ( n2511 & n2696 ) | ( n2695 & n2696 ) ;
  assign n2699 = ( n2511 & n2697 ) | ( n2511 & ~n2698 ) | ( n2697 & ~n2698 ) ;
  assign n2700 = ( ~n839 & n2694 ) | ( ~n839 & n2699 ) | ( n2694 & n2699 ) ;
  assign n2701 = ~n839 & n2512 ;
  assign n2702 = ( ~n839 & n2512 ) | ( ~n839 & n2615 ) | ( n2512 & n2615 ) ;
  assign n2703 = ( ~n2517 & n2701 ) | ( ~n2517 & n2702 ) | ( n2701 & n2702 ) ;
  assign n2704 = ( n2517 & n2701 ) | ( n2517 & n2702 ) | ( n2701 & n2702 ) ;
  assign n2705 = ( n2517 & n2703 ) | ( n2517 & ~n2704 ) | ( n2703 & ~n2704 ) ;
  assign n2706 = ( ~n746 & n2700 ) | ( ~n746 & n2705 ) | ( n2700 & n2705 ) ;
  assign n2707 = ~n746 & n2518 ;
  assign n2708 = ( ~n746 & n2518 ) | ( ~n746 & n2615 ) | ( n2518 & n2615 ) ;
  assign n2709 = ( n2523 & n2707 ) | ( n2523 & n2708 ) | ( n2707 & n2708 ) ;
  assign n2710 = ( ~n2523 & n2707 ) | ( ~n2523 & n2708 ) | ( n2707 & n2708 ) ;
  assign n2711 = ( n2523 & ~n2709 ) | ( n2523 & n2710 ) | ( ~n2709 & n2710 ) ;
  assign n2712 = ( ~n664 & n2706 ) | ( ~n664 & n2711 ) | ( n2706 & n2711 ) ;
  assign n2713 = ~n664 & n2524 ;
  assign n2714 = ( ~n664 & n2524 ) | ( ~n664 & n2615 ) | ( n2524 & n2615 ) ;
  assign n2715 = ( ~n2529 & n2713 ) | ( ~n2529 & n2714 ) | ( n2713 & n2714 ) ;
  assign n2716 = ( n2529 & n2713 ) | ( n2529 & n2714 ) | ( n2713 & n2714 ) ;
  assign n2717 = ( n2529 & n2715 ) | ( n2529 & ~n2716 ) | ( n2715 & ~n2716 ) ;
  assign n2718 = ( ~n588 & n2712 ) | ( ~n588 & n2717 ) | ( n2712 & n2717 ) ;
  assign n2719 = ( n588 & ~n2530 ) | ( n588 & n2615 ) | ( ~n2530 & n2615 ) ;
  assign n2720 = n588 & ~n2530 ;
  assign n2721 = ( n2535 & n2719 ) | ( n2535 & n2720 ) | ( n2719 & n2720 ) ;
  assign n2722 = ( ~n2535 & n2719 ) | ( ~n2535 & n2720 ) | ( n2719 & n2720 ) ;
  assign n2723 = ( n2535 & ~n2721 ) | ( n2535 & n2722 ) | ( ~n2721 & n2722 ) ;
  assign n2724 = ( ~n518 & n2718 ) | ( ~n518 & n2723 ) | ( n2718 & n2723 ) ;
  assign n2725 = ~n518 & n2536 ;
  assign n2726 = ( ~n518 & n2536 ) | ( ~n518 & n2615 ) | ( n2536 & n2615 ) ;
  assign n2727 = ( n2541 & n2725 ) | ( n2541 & n2726 ) | ( n2725 & n2726 ) ;
  assign n2728 = ( ~n2541 & n2725 ) | ( ~n2541 & n2726 ) | ( n2725 & n2726 ) ;
  assign n2729 = ( n2541 & ~n2727 ) | ( n2541 & n2728 ) | ( ~n2727 & n2728 ) ;
  assign n2730 = ( ~n454 & n2724 ) | ( ~n454 & n2729 ) | ( n2724 & n2729 ) ;
  assign n2731 = ~n454 & n2542 ;
  assign n2732 = ( ~n454 & n2542 ) | ( ~n454 & n2615 ) | ( n2542 & n2615 ) ;
  assign n2733 = ( ~n2547 & n2731 ) | ( ~n2547 & n2732 ) | ( n2731 & n2732 ) ;
  assign n2734 = ( n2547 & n2731 ) | ( n2547 & n2732 ) | ( n2731 & n2732 ) ;
  assign n2735 = ( n2547 & n2733 ) | ( n2547 & ~n2734 ) | ( n2733 & ~n2734 ) ;
  assign n2736 = ( ~n396 & n2730 ) | ( ~n396 & n2735 ) | ( n2730 & n2735 ) ;
  assign n2737 = ( n396 & ~n2548 ) | ( n396 & n2615 ) | ( ~n2548 & n2615 ) ;
  assign n2738 = n396 & ~n2548 ;
  assign n2739 = ( n2553 & n2737 ) | ( n2553 & n2738 ) | ( n2737 & n2738 ) ;
  assign n2740 = ( ~n2553 & n2737 ) | ( ~n2553 & n2738 ) | ( n2737 & n2738 ) ;
  assign n2741 = ( n2553 & ~n2739 ) | ( n2553 & n2740 ) | ( ~n2739 & n2740 ) ;
  assign n2742 = ( ~n344 & n2736 ) | ( ~n344 & n2741 ) | ( n2736 & n2741 ) ;
  assign n2743 = ( n344 & ~n2554 ) | ( n344 & n2615 ) | ( ~n2554 & n2615 ) ;
  assign n2744 = n344 & ~n2554 ;
  assign n2745 = ( n2559 & n2743 ) | ( n2559 & n2744 ) | ( n2743 & n2744 ) ;
  assign n2746 = ( ~n2559 & n2743 ) | ( ~n2559 & n2744 ) | ( n2743 & n2744 ) ;
  assign n2747 = ( n2559 & ~n2745 ) | ( n2559 & n2746 ) | ( ~n2745 & n2746 ) ;
  assign n2748 = ( ~n298 & n2742 ) | ( ~n298 & n2747 ) | ( n2742 & n2747 ) ;
  assign n2749 = ( n298 & ~n2560 ) | ( n298 & n2615 ) | ( ~n2560 & n2615 ) ;
  assign n2750 = n298 & ~n2560 ;
  assign n2751 = ( n2565 & n2749 ) | ( n2565 & n2750 ) | ( n2749 & n2750 ) ;
  assign n2752 = ( ~n2565 & n2749 ) | ( ~n2565 & n2750 ) | ( n2749 & n2750 ) ;
  assign n2753 = ( n2565 & ~n2751 ) | ( n2565 & n2752 ) | ( ~n2751 & n2752 ) ;
  assign n2754 = ( ~n258 & n2748 ) | ( ~n258 & n2753 ) | ( n2748 & n2753 ) ;
  assign n2755 = ~n258 & n2566 ;
  assign n2756 = ( ~n258 & n2566 ) | ( ~n258 & n2615 ) | ( n2566 & n2615 ) ;
  assign n2757 = ( ~n2571 & n2755 ) | ( ~n2571 & n2756 ) | ( n2755 & n2756 ) ;
  assign n2758 = ( n2571 & n2755 ) | ( n2571 & n2756 ) | ( n2755 & n2756 ) ;
  assign n2759 = ( n2571 & n2757 ) | ( n2571 & ~n2758 ) | ( n2757 & ~n2758 ) ;
  assign n2760 = ( ~n225 & n2754 ) | ( ~n225 & n2759 ) | ( n2754 & n2759 ) ;
  assign n2761 = ( n225 & ~n2572 ) | ( n225 & n2615 ) | ( ~n2572 & n2615 ) ;
  assign n2762 = n225 & ~n2572 ;
  assign n2763 = ( n2577 & n2761 ) | ( n2577 & n2762 ) | ( n2761 & n2762 ) ;
  assign n2764 = ( ~n2577 & n2761 ) | ( ~n2577 & n2762 ) | ( n2761 & n2762 ) ;
  assign n2765 = ( n2577 & ~n2763 ) | ( n2577 & n2764 ) | ( ~n2763 & n2764 ) ;
  assign n2766 = ( ~n197 & n2760 ) | ( ~n197 & n2765 ) | ( n2760 & n2765 ) ;
  assign n2767 = ( n197 & ~n2578 ) | ( n197 & n2615 ) | ( ~n2578 & n2615 ) ;
  assign n2768 = n197 & ~n2578 ;
  assign n2769 = ( n2583 & n2767 ) | ( n2583 & n2768 ) | ( n2767 & n2768 ) ;
  assign n2770 = ( ~n2583 & n2767 ) | ( ~n2583 & n2768 ) | ( n2767 & n2768 ) ;
  assign n2771 = ( n2583 & ~n2769 ) | ( n2583 & n2770 ) | ( ~n2769 & n2770 ) ;
  assign n2772 = ( ~n170 & n2766 ) | ( ~n170 & n2771 ) | ( n2766 & n2771 ) ;
  assign n2773 = ~n170 & n2584 ;
  assign n2774 = ( ~n170 & n2584 ) | ( ~n170 & n2615 ) | ( n2584 & n2615 ) ;
  assign n2775 = ( ~n2589 & n2773 ) | ( ~n2589 & n2774 ) | ( n2773 & n2774 ) ;
  assign n2776 = ( n2589 & n2773 ) | ( n2589 & n2774 ) | ( n2773 & n2774 ) ;
  assign n2777 = ( n2589 & n2775 ) | ( n2589 & ~n2776 ) | ( n2775 & ~n2776 ) ;
  assign n2778 = ( ~n142 & n2772 ) | ( ~n142 & n2777 ) | ( n2772 & n2777 ) ;
  assign n2779 = ( n142 & ~n2590 ) | ( n142 & n2615 ) | ( ~n2590 & n2615 ) ;
  assign n2780 = n142 & ~n2590 ;
  assign n2781 = ( n2595 & n2779 ) | ( n2595 & n2780 ) | ( n2779 & n2780 ) ;
  assign n2782 = ( ~n2595 & n2779 ) | ( ~n2595 & n2780 ) | ( n2779 & n2780 ) ;
  assign n2783 = ( n2595 & ~n2781 ) | ( n2595 & n2782 ) | ( ~n2781 & n2782 ) ;
  assign n2784 = ( ~n132 & n2778 ) | ( ~n132 & n2783 ) | ( n2778 & n2783 ) ;
  assign n2785 = n132 & ~n2596 ;
  assign n2786 = ( n132 & ~n2596 ) | ( n132 & n2615 ) | ( ~n2596 & n2615 ) ;
  assign n2787 = ( n2601 & n2785 ) | ( n2601 & n2786 ) | ( n2785 & n2786 ) ;
  assign n2788 = ( ~n2601 & n2785 ) | ( ~n2601 & n2786 ) | ( n2785 & n2786 ) ;
  assign n2789 = ( n2601 & ~n2787 ) | ( n2601 & n2788 ) | ( ~n2787 & n2788 ) ;
  assign n2790 = ( ~n131 & n2784 ) | ( ~n131 & n2789 ) | ( n2784 & n2789 ) ;
  assign n2791 = n2618 | n2790 ;
  assign n2792 = n2618 | n2789 ;
  assign n2793 = ( n2784 & n2789 ) | ( n2784 & n2792 ) | ( n2789 & n2792 ) ;
  assign n2794 = n131 & ~n2784 ;
  assign n2795 = ~n131 & n2602 ;
  assign n2796 = n2607 & n2795 ;
  assign n2797 = ~n2602 & n2617 ;
  assign n2798 = ( ~n2789 & n2796 ) | ( ~n2789 & n2797 ) | ( n2796 & n2797 ) ;
  assign n2799 = ( n2789 & ~n2794 ) | ( n2789 & n2798 ) | ( ~n2794 & n2798 ) ;
  assign n2800 = n2793 & ~n2799 ;
  assign n2801 = n2784 & n2789 ;
  assign n2802 = ( n131 & ~n2784 ) | ( n131 & n2798 ) | ( ~n2784 & n2798 ) ;
  assign n2803 = ( ~n131 & n2801 ) | ( ~n131 & n2802 ) | ( n2801 & n2802 ) ;
  assign n2804 = n2800 | n2803 ;
  assign n2805 = ( n132 & ~n2778 ) | ( n132 & n2791 ) | ( ~n2778 & n2791 ) ;
  assign n2806 = n132 & ~n2778 ;
  assign n2807 = ( n2783 & ~n2805 ) | ( n2783 & n2806 ) | ( ~n2805 & n2806 ) ;
  assign n2808 = ( n2783 & n2805 ) | ( n2783 & n2806 ) | ( n2805 & n2806 ) ;
  assign n2809 = ( n2805 & n2807 ) | ( n2805 & ~n2808 ) | ( n2807 & ~n2808 ) ;
  assign n2810 = x66 | x67 ;
  assign n2811 = x68 | n2810 ;
  assign n2812 = n2615 & ~n2811 ;
  assign n2813 = ~n2619 & n2791 ;
  assign n2814 = ~n2615 & n2811 ;
  assign n2815 = ( x69 & ~n2791 ) | ( x69 & n2814 ) | ( ~n2791 & n2814 ) ;
  assign n2816 = ( ~n2812 & n2813 ) | ( ~n2812 & n2815 ) | ( n2813 & n2815 ) ;
  assign n2817 = n2615 & ~n2791 ;
  assign n2818 = ( x70 & n2813 ) | ( x70 & n2817 ) | ( n2813 & n2817 ) ;
  assign n2819 = ( ~x70 & n2813 ) | ( ~x70 & n2817 ) | ( n2813 & n2817 ) ;
  assign n2820 = ( x70 & ~n2818 ) | ( x70 & n2819 ) | ( ~n2818 & n2819 ) ;
  assign n2821 = ( ~n2443 & n2816 ) | ( ~n2443 & n2820 ) | ( n2816 & n2820 ) ;
  assign n2822 = ~n2443 & n2615 ;
  assign n2823 = ( n2626 & n2791 ) | ( n2626 & n2822 ) | ( n2791 & n2822 ) ;
  assign n2824 = ( ~x71 & n2819 ) | ( ~x71 & n2823 ) | ( n2819 & n2823 ) ;
  assign n2825 = ( x71 & n2819 ) | ( x71 & n2823 ) | ( n2819 & n2823 ) ;
  assign n2826 = ( x71 & n2824 ) | ( x71 & ~n2825 ) | ( n2824 & ~n2825 ) ;
  assign n2827 = ( ~n2277 & n2821 ) | ( ~n2277 & n2826 ) | ( n2821 & n2826 ) ;
  assign n2828 = n2277 & ~n2625 ;
  assign n2829 = ( n2277 & ~n2625 ) | ( n2277 & n2791 ) | ( ~n2625 & n2791 ) ;
  assign n2830 = ( ~n2629 & n2828 ) | ( ~n2629 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2831 = ( n2629 & n2828 ) | ( n2629 & n2829 ) | ( n2828 & n2829 ) ;
  assign n2832 = ( n2629 & n2830 ) | ( n2629 & ~n2831 ) | ( n2830 & ~n2831 ) ;
  assign n2833 = ( ~n2111 & n2827 ) | ( ~n2111 & n2832 ) | ( n2827 & n2832 ) ;
  assign n2834 = ( n2111 & ~n2630 ) | ( n2111 & n2791 ) | ( ~n2630 & n2791 ) ;
  assign n2835 = n2111 & ~n2630 ;
  assign n2836 = ( n2639 & n2834 ) | ( n2639 & n2835 ) | ( n2834 & n2835 ) ;
  assign n2837 = ( ~n2639 & n2834 ) | ( ~n2639 & n2835 ) | ( n2834 & n2835 ) ;
  assign n2838 = ( n2639 & ~n2836 ) | ( n2639 & n2837 ) | ( ~n2836 & n2837 ) ;
  assign n2839 = ( ~n1949 & n2833 ) | ( ~n1949 & n2838 ) | ( n2833 & n2838 ) ;
  assign n2840 = ( n1949 & ~n2640 ) | ( n1949 & n2791 ) | ( ~n2640 & n2791 ) ;
  assign n2841 = n1949 & ~n2640 ;
  assign n2842 = ( n2645 & n2840 ) | ( n2645 & n2841 ) | ( n2840 & n2841 ) ;
  assign n2843 = ( ~n2645 & n2840 ) | ( ~n2645 & n2841 ) | ( n2840 & n2841 ) ;
  assign n2844 = ( n2645 & ~n2842 ) | ( n2645 & n2843 ) | ( ~n2842 & n2843 ) ;
  assign n2845 = ( ~n1802 & n2839 ) | ( ~n1802 & n2844 ) | ( n2839 & n2844 ) ;
  assign n2846 = ~n1802 & n2646 ;
  assign n2847 = ( ~n1802 & n2646 ) | ( ~n1802 & n2791 ) | ( n2646 & n2791 ) ;
  assign n2848 = ( n2651 & n2846 ) | ( n2651 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2849 = ( ~n2651 & n2846 ) | ( ~n2651 & n2847 ) | ( n2846 & n2847 ) ;
  assign n2850 = ( n2651 & ~n2848 ) | ( n2651 & n2849 ) | ( ~n2848 & n2849 ) ;
  assign n2851 = ( ~n1661 & n2845 ) | ( ~n1661 & n2850 ) | ( n2845 & n2850 ) ;
  assign n2852 = ~n1661 & n2652 ;
  assign n2853 = ( ~n1661 & n2652 ) | ( ~n1661 & n2791 ) | ( n2652 & n2791 ) ;
  assign n2854 = ( n2657 & n2852 ) | ( n2657 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2855 = ( ~n2657 & n2852 ) | ( ~n2657 & n2853 ) | ( n2852 & n2853 ) ;
  assign n2856 = ( n2657 & ~n2854 ) | ( n2657 & n2855 ) | ( ~n2854 & n2855 ) ;
  assign n2857 = ( ~n1523 & n2851 ) | ( ~n1523 & n2856 ) | ( n2851 & n2856 ) ;
  assign n2858 = ( n1523 & ~n2658 ) | ( n1523 & n2791 ) | ( ~n2658 & n2791 ) ;
  assign n2859 = n1523 & ~n2658 ;
  assign n2860 = ( n2663 & n2858 ) | ( n2663 & n2859 ) | ( n2858 & n2859 ) ;
  assign n2861 = ( ~n2663 & n2858 ) | ( ~n2663 & n2859 ) | ( n2858 & n2859 ) ;
  assign n2862 = ( n2663 & ~n2860 ) | ( n2663 & n2861 ) | ( ~n2860 & n2861 ) ;
  assign n2863 = ( ~n1393 & n2857 ) | ( ~n1393 & n2862 ) | ( n2857 & n2862 ) ;
  assign n2864 = ~n1393 & n2664 ;
  assign n2865 = ( ~n1393 & n2664 ) | ( ~n1393 & n2791 ) | ( n2664 & n2791 ) ;
  assign n2866 = ( n2669 & n2864 ) | ( n2669 & n2865 ) | ( n2864 & n2865 ) ;
  assign n2867 = ( ~n2669 & n2864 ) | ( ~n2669 & n2865 ) | ( n2864 & n2865 ) ;
  assign n2868 = ( n2669 & ~n2866 ) | ( n2669 & n2867 ) | ( ~n2866 & n2867 ) ;
  assign n2869 = ( ~n1266 & n2863 ) | ( ~n1266 & n2868 ) | ( n2863 & n2868 ) ;
  assign n2870 = ( n1266 & ~n2670 ) | ( n1266 & n2791 ) | ( ~n2670 & n2791 ) ;
  assign n2871 = n1266 & ~n2670 ;
  assign n2872 = ( n2675 & n2870 ) | ( n2675 & n2871 ) | ( n2870 & n2871 ) ;
  assign n2873 = ( ~n2675 & n2870 ) | ( ~n2675 & n2871 ) | ( n2870 & n2871 ) ;
  assign n2874 = ( n2675 & ~n2872 ) | ( n2675 & n2873 ) | ( ~n2872 & n2873 ) ;
  assign n2875 = ( ~n1150 & n2869 ) | ( ~n1150 & n2874 ) | ( n2869 & n2874 ) ;
  assign n2876 = ( n1150 & ~n2676 ) | ( n1150 & n2791 ) | ( ~n2676 & n2791 ) ;
  assign n2877 = n1150 & ~n2676 ;
  assign n2878 = ( n2681 & n2876 ) | ( n2681 & n2877 ) | ( n2876 & n2877 ) ;
  assign n2879 = ( ~n2681 & n2876 ) | ( ~n2681 & n2877 ) | ( n2876 & n2877 ) ;
  assign n2880 = ( n2681 & ~n2878 ) | ( n2681 & n2879 ) | ( ~n2878 & n2879 ) ;
  assign n2881 = ( ~n1038 & n2875 ) | ( ~n1038 & n2880 ) | ( n2875 & n2880 ) ;
  assign n2882 = ~n1038 & n2682 ;
  assign n2883 = ( ~n1038 & n2682 ) | ( ~n1038 & n2791 ) | ( n2682 & n2791 ) ;
  assign n2884 = ( ~n2687 & n2882 ) | ( ~n2687 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2885 = ( n2687 & n2882 ) | ( n2687 & n2883 ) | ( n2882 & n2883 ) ;
  assign n2886 = ( n2687 & n2884 ) | ( n2687 & ~n2885 ) | ( n2884 & ~n2885 ) ;
  assign n2887 = ( ~n933 & n2881 ) | ( ~n933 & n2886 ) | ( n2881 & n2886 ) ;
  assign n2888 = ( n933 & ~n2688 ) | ( n933 & n2791 ) | ( ~n2688 & n2791 ) ;
  assign n2889 = n933 & ~n2688 ;
  assign n2890 = ( n2693 & n2888 ) | ( n2693 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2891 = ( ~n2693 & n2888 ) | ( ~n2693 & n2889 ) | ( n2888 & n2889 ) ;
  assign n2892 = ( n2693 & ~n2890 ) | ( n2693 & n2891 ) | ( ~n2890 & n2891 ) ;
  assign n2893 = ( ~n839 & n2887 ) | ( ~n839 & n2892 ) | ( n2887 & n2892 ) ;
  assign n2894 = ~n839 & n2694 ;
  assign n2895 = ( ~n839 & n2694 ) | ( ~n839 & n2791 ) | ( n2694 & n2791 ) ;
  assign n2896 = ( ~n2699 & n2894 ) | ( ~n2699 & n2895 ) | ( n2894 & n2895 ) ;
  assign n2897 = ( n2699 & n2894 ) | ( n2699 & n2895 ) | ( n2894 & n2895 ) ;
  assign n2898 = ( n2699 & n2896 ) | ( n2699 & ~n2897 ) | ( n2896 & ~n2897 ) ;
  assign n2899 = ( ~n746 & n2893 ) | ( ~n746 & n2898 ) | ( n2893 & n2898 ) ;
  assign n2900 = ~n746 & n2700 ;
  assign n2901 = ( ~n746 & n2700 ) | ( ~n746 & n2791 ) | ( n2700 & n2791 ) ;
  assign n2902 = ( n2705 & n2900 ) | ( n2705 & n2901 ) | ( n2900 & n2901 ) ;
  assign n2903 = ( ~n2705 & n2900 ) | ( ~n2705 & n2901 ) | ( n2900 & n2901 ) ;
  assign n2904 = ( n2705 & ~n2902 ) | ( n2705 & n2903 ) | ( ~n2902 & n2903 ) ;
  assign n2905 = ( ~n664 & n2899 ) | ( ~n664 & n2904 ) | ( n2899 & n2904 ) ;
  assign n2906 = ( n664 & ~n2706 ) | ( n664 & n2791 ) | ( ~n2706 & n2791 ) ;
  assign n2907 = n664 & ~n2706 ;
  assign n2908 = ( n2711 & n2906 ) | ( n2711 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2909 = ( ~n2711 & n2906 ) | ( ~n2711 & n2907 ) | ( n2906 & n2907 ) ;
  assign n2910 = ( n2711 & ~n2908 ) | ( n2711 & n2909 ) | ( ~n2908 & n2909 ) ;
  assign n2911 = ( ~n588 & n2905 ) | ( ~n588 & n2910 ) | ( n2905 & n2910 ) ;
  assign n2912 = ( n588 & ~n2712 ) | ( n588 & n2791 ) | ( ~n2712 & n2791 ) ;
  assign n2913 = n588 & ~n2712 ;
  assign n2914 = ( n2717 & n2912 ) | ( n2717 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2915 = ( ~n2717 & n2912 ) | ( ~n2717 & n2913 ) | ( n2912 & n2913 ) ;
  assign n2916 = ( n2717 & ~n2914 ) | ( n2717 & n2915 ) | ( ~n2914 & n2915 ) ;
  assign n2917 = ( ~n518 & n2911 ) | ( ~n518 & n2916 ) | ( n2911 & n2916 ) ;
  assign n2918 = n518 & ~n2718 ;
  assign n2919 = ( n518 & ~n2718 ) | ( n518 & n2791 ) | ( ~n2718 & n2791 ) ;
  assign n2920 = ( n2723 & n2918 ) | ( n2723 & n2919 ) | ( n2918 & n2919 ) ;
  assign n2921 = ( ~n2723 & n2918 ) | ( ~n2723 & n2919 ) | ( n2918 & n2919 ) ;
  assign n2922 = ( n2723 & ~n2920 ) | ( n2723 & n2921 ) | ( ~n2920 & n2921 ) ;
  assign n2923 = ( ~n454 & n2917 ) | ( ~n454 & n2922 ) | ( n2917 & n2922 ) ;
  assign n2924 = ( n454 & ~n2724 ) | ( n454 & n2791 ) | ( ~n2724 & n2791 ) ;
  assign n2925 = n454 & ~n2724 ;
  assign n2926 = ( n2729 & n2924 ) | ( n2729 & n2925 ) | ( n2924 & n2925 ) ;
  assign n2927 = ( ~n2729 & n2924 ) | ( ~n2729 & n2925 ) | ( n2924 & n2925 ) ;
  assign n2928 = ( n2729 & ~n2926 ) | ( n2729 & n2927 ) | ( ~n2926 & n2927 ) ;
  assign n2929 = ( ~n396 & n2923 ) | ( ~n396 & n2928 ) | ( n2923 & n2928 ) ;
  assign n2930 = ~n396 & n2730 ;
  assign n2931 = ( ~n396 & n2730 ) | ( ~n396 & n2791 ) | ( n2730 & n2791 ) ;
  assign n2932 = ( n2735 & n2930 ) | ( n2735 & n2931 ) | ( n2930 & n2931 ) ;
  assign n2933 = ( ~n2735 & n2930 ) | ( ~n2735 & n2931 ) | ( n2930 & n2931 ) ;
  assign n2934 = ( n2735 & ~n2932 ) | ( n2735 & n2933 ) | ( ~n2932 & n2933 ) ;
  assign n2935 = ( ~n344 & n2929 ) | ( ~n344 & n2934 ) | ( n2929 & n2934 ) ;
  assign n2936 = ( n344 & ~n2736 ) | ( n344 & n2791 ) | ( ~n2736 & n2791 ) ;
  assign n2937 = n344 & ~n2736 ;
  assign n2938 = ( n2741 & n2936 ) | ( n2741 & n2937 ) | ( n2936 & n2937 ) ;
  assign n2939 = ( ~n2741 & n2936 ) | ( ~n2741 & n2937 ) | ( n2936 & n2937 ) ;
  assign n2940 = ( n2741 & ~n2938 ) | ( n2741 & n2939 ) | ( ~n2938 & n2939 ) ;
  assign n2941 = ( ~n298 & n2935 ) | ( ~n298 & n2940 ) | ( n2935 & n2940 ) ;
  assign n2942 = ( n298 & ~n2742 ) | ( n298 & n2791 ) | ( ~n2742 & n2791 ) ;
  assign n2943 = n298 & ~n2742 ;
  assign n2944 = ( n2747 & n2942 ) | ( n2747 & n2943 ) | ( n2942 & n2943 ) ;
  assign n2945 = ( ~n2747 & n2942 ) | ( ~n2747 & n2943 ) | ( n2942 & n2943 ) ;
  assign n2946 = ( n2747 & ~n2944 ) | ( n2747 & n2945 ) | ( ~n2944 & n2945 ) ;
  assign n2947 = ( ~n258 & n2941 ) | ( ~n258 & n2946 ) | ( n2941 & n2946 ) ;
  assign n2948 = ( n258 & ~n2748 ) | ( n258 & n2791 ) | ( ~n2748 & n2791 ) ;
  assign n2949 = n258 & ~n2748 ;
  assign n2950 = ( n2753 & n2948 ) | ( n2753 & n2949 ) | ( n2948 & n2949 ) ;
  assign n2951 = ( ~n2753 & n2948 ) | ( ~n2753 & n2949 ) | ( n2948 & n2949 ) ;
  assign n2952 = ( n2753 & ~n2950 ) | ( n2753 & n2951 ) | ( ~n2950 & n2951 ) ;
  assign n2953 = ( ~n225 & n2947 ) | ( ~n225 & n2952 ) | ( n2947 & n2952 ) ;
  assign n2954 = ( n225 & ~n2754 ) | ( n225 & n2791 ) | ( ~n2754 & n2791 ) ;
  assign n2955 = n225 & ~n2754 ;
  assign n2956 = ( n2759 & n2954 ) | ( n2759 & n2955 ) | ( n2954 & n2955 ) ;
  assign n2957 = ( ~n2759 & n2954 ) | ( ~n2759 & n2955 ) | ( n2954 & n2955 ) ;
  assign n2958 = ( n2759 & ~n2956 ) | ( n2759 & n2957 ) | ( ~n2956 & n2957 ) ;
  assign n2959 = ( ~n197 & n2953 ) | ( ~n197 & n2958 ) | ( n2953 & n2958 ) ;
  assign n2960 = ( n197 & ~n2760 ) | ( n197 & n2791 ) | ( ~n2760 & n2791 ) ;
  assign n2961 = n197 & ~n2760 ;
  assign n2962 = ( n2765 & n2960 ) | ( n2765 & n2961 ) | ( n2960 & n2961 ) ;
  assign n2963 = ( ~n2765 & n2960 ) | ( ~n2765 & n2961 ) | ( n2960 & n2961 ) ;
  assign n2964 = ( n2765 & ~n2962 ) | ( n2765 & n2963 ) | ( ~n2962 & n2963 ) ;
  assign n2965 = ( ~n170 & n2959 ) | ( ~n170 & n2964 ) | ( n2959 & n2964 ) ;
  assign n2966 = ( n170 & ~n2766 ) | ( n170 & n2791 ) | ( ~n2766 & n2791 ) ;
  assign n2967 = n170 & ~n2766 ;
  assign n2968 = ( n2771 & n2966 ) | ( n2771 & n2967 ) | ( n2966 & n2967 ) ;
  assign n2969 = ( ~n2771 & n2966 ) | ( ~n2771 & n2967 ) | ( n2966 & n2967 ) ;
  assign n2970 = ( n2771 & ~n2968 ) | ( n2771 & n2969 ) | ( ~n2968 & n2969 ) ;
  assign n2971 = ( ~n142 & n2965 ) | ( ~n142 & n2970 ) | ( n2965 & n2970 ) ;
  assign n2972 = ( n142 & ~n2772 ) | ( n142 & n2791 ) | ( ~n2772 & n2791 ) ;
  assign n2973 = n142 & ~n2772 ;
  assign n2974 = ( n2777 & n2972 ) | ( n2777 & n2973 ) | ( n2972 & n2973 ) ;
  assign n2975 = ( ~n2777 & n2972 ) | ( ~n2777 & n2973 ) | ( n2972 & n2973 ) ;
  assign n2976 = ( n2777 & ~n2974 ) | ( n2777 & n2975 ) | ( ~n2974 & n2975 ) ;
  assign n2977 = ( ~n132 & n2971 ) | ( ~n132 & n2976 ) | ( n2971 & n2976 ) ;
  assign n2978 = ( ~n131 & n2809 ) | ( ~n131 & n2977 ) | ( n2809 & n2977 ) ;
  assign n2979 = n2804 | n2978 ;
  assign n2980 = ( n142 & ~n2965 ) | ( n142 & n2979 ) | ( ~n2965 & n2979 ) ;
  assign n2981 = n142 & ~n2965 ;
  assign n2982 = ( n2970 & ~n2980 ) | ( n2970 & n2981 ) | ( ~n2980 & n2981 ) ;
  assign n2983 = ( n2970 & n2980 ) | ( n2970 & n2981 ) | ( n2980 & n2981 ) ;
  assign n2984 = ( n2980 & n2982 ) | ( n2980 & ~n2983 ) | ( n2982 & ~n2983 ) ;
  assign n2985 = ~n2810 & n2979 ;
  assign n2986 = x64 | x65 ;
  assign n2987 = x66 | n2986 ;
  assign n2988 = n2791 & ~n2987 ;
  assign n2989 = ~n2791 & n2987 ;
  assign n2990 = ( x67 & ~n2979 ) | ( x67 & n2989 ) | ( ~n2979 & n2989 ) ;
  assign n2991 = ( n2985 & ~n2988 ) | ( n2985 & n2990 ) | ( ~n2988 & n2990 ) ;
  assign n2992 = n2791 & ~n2979 ;
  assign n2993 = ( x68 & n2985 ) | ( x68 & n2992 ) | ( n2985 & n2992 ) ;
  assign n2994 = ( ~x68 & n2985 ) | ( ~x68 & n2992 ) | ( n2985 & n2992 ) ;
  assign n2995 = ( x68 & ~n2993 ) | ( x68 & n2994 ) | ( ~n2993 & n2994 ) ;
  assign n2996 = ( ~n2615 & n2991 ) | ( ~n2615 & n2995 ) | ( n2991 & n2995 ) ;
  assign n2997 = ~n2615 & n2791 ;
  assign n2998 = ( n2817 & n2979 ) | ( n2817 & n2997 ) | ( n2979 & n2997 ) ;
  assign n2999 = ( ~x69 & n2994 ) | ( ~x69 & n2998 ) | ( n2994 & n2998 ) ;
  assign n3000 = ( x69 & n2994 ) | ( x69 & n2998 ) | ( n2994 & n2998 ) ;
  assign n3001 = ( x69 & n2999 ) | ( x69 & ~n3000 ) | ( n2999 & ~n3000 ) ;
  assign n3002 = ( ~n2443 & n2996 ) | ( ~n2443 & n3001 ) | ( n2996 & n3001 ) ;
  assign n3003 = ( n2443 & ~n2816 ) | ( n2443 & n2979 ) | ( ~n2816 & n2979 ) ;
  assign n3004 = n2443 & ~n2816 ;
  assign n3005 = ( n2820 & n3003 ) | ( n2820 & n3004 ) | ( n3003 & n3004 ) ;
  assign n3006 = ( ~n2820 & n3003 ) | ( ~n2820 & n3004 ) | ( n3003 & n3004 ) ;
  assign n3007 = ( n2820 & ~n3005 ) | ( n2820 & n3006 ) | ( ~n3005 & n3006 ) ;
  assign n3008 = ( ~n2277 & n3002 ) | ( ~n2277 & n3007 ) | ( n3002 & n3007 ) ;
  assign n3009 = ~n2277 & n2821 ;
  assign n3010 = ( ~n2277 & n2821 ) | ( ~n2277 & n2979 ) | ( n2821 & n2979 ) ;
  assign n3011 = ( ~n2826 & n3009 ) | ( ~n2826 & n3010 ) | ( n3009 & n3010 ) ;
  assign n3012 = ( n2826 & n3009 ) | ( n2826 & n3010 ) | ( n3009 & n3010 ) ;
  assign n3013 = ( n2826 & n3011 ) | ( n2826 & ~n3012 ) | ( n3011 & ~n3012 ) ;
  assign n3014 = ( ~n2111 & n3008 ) | ( ~n2111 & n3013 ) | ( n3008 & n3013 ) ;
  assign n3015 = n2111 & ~n2827 ;
  assign n3016 = ( n2111 & ~n2827 ) | ( n2111 & n2979 ) | ( ~n2827 & n2979 ) ;
  assign n3017 = ( n2832 & n3015 ) | ( n2832 & n3016 ) | ( n3015 & n3016 ) ;
  assign n3018 = ( ~n2832 & n3015 ) | ( ~n2832 & n3016 ) | ( n3015 & n3016 ) ;
  assign n3019 = ( n2832 & ~n3017 ) | ( n2832 & n3018 ) | ( ~n3017 & n3018 ) ;
  assign n3020 = ( ~n1949 & n3014 ) | ( ~n1949 & n3019 ) | ( n3014 & n3019 ) ;
  assign n3021 = ~n1949 & n2833 ;
  assign n3022 = ( ~n1949 & n2833 ) | ( ~n1949 & n2979 ) | ( n2833 & n2979 ) ;
  assign n3023 = ( n2838 & n3021 ) | ( n2838 & n3022 ) | ( n3021 & n3022 ) ;
  assign n3024 = ( ~n2838 & n3021 ) | ( ~n2838 & n3022 ) | ( n3021 & n3022 ) ;
  assign n3025 = ( n2838 & ~n3023 ) | ( n2838 & n3024 ) | ( ~n3023 & n3024 ) ;
  assign n3026 = ( ~n1802 & n3020 ) | ( ~n1802 & n3025 ) | ( n3020 & n3025 ) ;
  assign n3027 = ~n1802 & n2839 ;
  assign n3028 = ( ~n1802 & n2839 ) | ( ~n1802 & n2979 ) | ( n2839 & n2979 ) ;
  assign n3029 = ( ~n2844 & n3027 ) | ( ~n2844 & n3028 ) | ( n3027 & n3028 ) ;
  assign n3030 = ( n2844 & n3027 ) | ( n2844 & n3028 ) | ( n3027 & n3028 ) ;
  assign n3031 = ( n2844 & n3029 ) | ( n2844 & ~n3030 ) | ( n3029 & ~n3030 ) ;
  assign n3032 = ( ~n1661 & n3026 ) | ( ~n1661 & n3031 ) | ( n3026 & n3031 ) ;
  assign n3033 = ( n1661 & ~n2845 ) | ( n1661 & n2979 ) | ( ~n2845 & n2979 ) ;
  assign n3034 = n1661 & ~n2845 ;
  assign n3035 = ( n2850 & n3033 ) | ( n2850 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3036 = ( ~n2850 & n3033 ) | ( ~n2850 & n3034 ) | ( n3033 & n3034 ) ;
  assign n3037 = ( n2850 & ~n3035 ) | ( n2850 & n3036 ) | ( ~n3035 & n3036 ) ;
  assign n3038 = ( ~n1523 & n3032 ) | ( ~n1523 & n3037 ) | ( n3032 & n3037 ) ;
  assign n3039 = ( n1523 & ~n2851 ) | ( n1523 & n2979 ) | ( ~n2851 & n2979 ) ;
  assign n3040 = n1523 & ~n2851 ;
  assign n3041 = ( n2856 & n3039 ) | ( n2856 & n3040 ) | ( n3039 & n3040 ) ;
  assign n3042 = ( ~n2856 & n3039 ) | ( ~n2856 & n3040 ) | ( n3039 & n3040 ) ;
  assign n3043 = ( n2856 & ~n3041 ) | ( n2856 & n3042 ) | ( ~n3041 & n3042 ) ;
  assign n3044 = ( ~n1393 & n3038 ) | ( ~n1393 & n3043 ) | ( n3038 & n3043 ) ;
  assign n3045 = ( n1393 & ~n2857 ) | ( n1393 & n2979 ) | ( ~n2857 & n2979 ) ;
  assign n3046 = n1393 & ~n2857 ;
  assign n3047 = ( n2862 & n3045 ) | ( n2862 & n3046 ) | ( n3045 & n3046 ) ;
  assign n3048 = ( ~n2862 & n3045 ) | ( ~n2862 & n3046 ) | ( n3045 & n3046 ) ;
  assign n3049 = ( n2862 & ~n3047 ) | ( n2862 & n3048 ) | ( ~n3047 & n3048 ) ;
  assign n3050 = ( ~n1266 & n3044 ) | ( ~n1266 & n3049 ) | ( n3044 & n3049 ) ;
  assign n3051 = ( n1266 & ~n2863 ) | ( n1266 & n2979 ) | ( ~n2863 & n2979 ) ;
  assign n3052 = n1266 & ~n2863 ;
  assign n3053 = ( n2868 & n3051 ) | ( n2868 & n3052 ) | ( n3051 & n3052 ) ;
  assign n3054 = ( ~n2868 & n3051 ) | ( ~n2868 & n3052 ) | ( n3051 & n3052 ) ;
  assign n3055 = ( n2868 & ~n3053 ) | ( n2868 & n3054 ) | ( ~n3053 & n3054 ) ;
  assign n3056 = ( ~n1150 & n3050 ) | ( ~n1150 & n3055 ) | ( n3050 & n3055 ) ;
  assign n3057 = ( n1150 & ~n2869 ) | ( n1150 & n2979 ) | ( ~n2869 & n2979 ) ;
  assign n3058 = n1150 & ~n2869 ;
  assign n3059 = ( n2874 & n3057 ) | ( n2874 & n3058 ) | ( n3057 & n3058 ) ;
  assign n3060 = ( ~n2874 & n3057 ) | ( ~n2874 & n3058 ) | ( n3057 & n3058 ) ;
  assign n3061 = ( n2874 & ~n3059 ) | ( n2874 & n3060 ) | ( ~n3059 & n3060 ) ;
  assign n3062 = ( ~n1038 & n3056 ) | ( ~n1038 & n3061 ) | ( n3056 & n3061 ) ;
  assign n3063 = n1038 & ~n2875 ;
  assign n3064 = ( n1038 & ~n2875 ) | ( n1038 & n2979 ) | ( ~n2875 & n2979 ) ;
  assign n3065 = ( ~n2880 & n3063 ) | ( ~n2880 & n3064 ) | ( n3063 & n3064 ) ;
  assign n3066 = ( n2880 & n3063 ) | ( n2880 & n3064 ) | ( n3063 & n3064 ) ;
  assign n3067 = ( n2880 & n3065 ) | ( n2880 & ~n3066 ) | ( n3065 & ~n3066 ) ;
  assign n3068 = ( ~n933 & n3062 ) | ( ~n933 & n3067 ) | ( n3062 & n3067 ) ;
  assign n3069 = ( n933 & ~n2881 ) | ( n933 & n2979 ) | ( ~n2881 & n2979 ) ;
  assign n3070 = n933 & ~n2881 ;
  assign n3071 = ( n2886 & n3069 ) | ( n2886 & n3070 ) | ( n3069 & n3070 ) ;
  assign n3072 = ( ~n2886 & n3069 ) | ( ~n2886 & n3070 ) | ( n3069 & n3070 ) ;
  assign n3073 = ( n2886 & ~n3071 ) | ( n2886 & n3072 ) | ( ~n3071 & n3072 ) ;
  assign n3074 = ( ~n839 & n3068 ) | ( ~n839 & n3073 ) | ( n3068 & n3073 ) ;
  assign n3075 = ~n839 & n2887 ;
  assign n3076 = ( ~n839 & n2887 ) | ( ~n839 & n2979 ) | ( n2887 & n2979 ) ;
  assign n3077 = ( ~n2892 & n3075 ) | ( ~n2892 & n3076 ) | ( n3075 & n3076 ) ;
  assign n3078 = ( n2892 & n3075 ) | ( n2892 & n3076 ) | ( n3075 & n3076 ) ;
  assign n3079 = ( n2892 & n3077 ) | ( n2892 & ~n3078 ) | ( n3077 & ~n3078 ) ;
  assign n3080 = ( ~n746 & n3074 ) | ( ~n746 & n3079 ) | ( n3074 & n3079 ) ;
  assign n3081 = ( n746 & ~n2893 ) | ( n746 & n2979 ) | ( ~n2893 & n2979 ) ;
  assign n3082 = n746 & ~n2893 ;
  assign n3083 = ( n2898 & n3081 ) | ( n2898 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3084 = ( ~n2898 & n3081 ) | ( ~n2898 & n3082 ) | ( n3081 & n3082 ) ;
  assign n3085 = ( n2898 & ~n3083 ) | ( n2898 & n3084 ) | ( ~n3083 & n3084 ) ;
  assign n3086 = ( ~n664 & n3080 ) | ( ~n664 & n3085 ) | ( n3080 & n3085 ) ;
  assign n3087 = ( n664 & ~n2899 ) | ( n664 & n2979 ) | ( ~n2899 & n2979 ) ;
  assign n3088 = n664 & ~n2899 ;
  assign n3089 = ( n2904 & n3087 ) | ( n2904 & n3088 ) | ( n3087 & n3088 ) ;
  assign n3090 = ( ~n2904 & n3087 ) | ( ~n2904 & n3088 ) | ( n3087 & n3088 ) ;
  assign n3091 = ( n2904 & ~n3089 ) | ( n2904 & n3090 ) | ( ~n3089 & n3090 ) ;
  assign n3092 = ( ~n588 & n3086 ) | ( ~n588 & n3091 ) | ( n3086 & n3091 ) ;
  assign n3093 = ( n588 & ~n2905 ) | ( n588 & n2979 ) | ( ~n2905 & n2979 ) ;
  assign n3094 = n588 & ~n2905 ;
  assign n3095 = ( n2910 & n3093 ) | ( n2910 & n3094 ) | ( n3093 & n3094 ) ;
  assign n3096 = ( ~n2910 & n3093 ) | ( ~n2910 & n3094 ) | ( n3093 & n3094 ) ;
  assign n3097 = ( n2910 & ~n3095 ) | ( n2910 & n3096 ) | ( ~n3095 & n3096 ) ;
  assign n3098 = ( ~n518 & n3092 ) | ( ~n518 & n3097 ) | ( n3092 & n3097 ) ;
  assign n3099 = ~n518 & n2911 ;
  assign n3100 = ( ~n518 & n2911 ) | ( ~n518 & n2979 ) | ( n2911 & n2979 ) ;
  assign n3101 = ( n2916 & n3099 ) | ( n2916 & n3100 ) | ( n3099 & n3100 ) ;
  assign n3102 = ( ~n2916 & n3099 ) | ( ~n2916 & n3100 ) | ( n3099 & n3100 ) ;
  assign n3103 = ( n2916 & ~n3101 ) | ( n2916 & n3102 ) | ( ~n3101 & n3102 ) ;
  assign n3104 = ( ~n454 & n3098 ) | ( ~n454 & n3103 ) | ( n3098 & n3103 ) ;
  assign n3105 = ~n454 & n2917 ;
  assign n3106 = ( ~n454 & n2917 ) | ( ~n454 & n2979 ) | ( n2917 & n2979 ) ;
  assign n3107 = ( n2922 & n3105 ) | ( n2922 & n3106 ) | ( n3105 & n3106 ) ;
  assign n3108 = ( ~n2922 & n3105 ) | ( ~n2922 & n3106 ) | ( n3105 & n3106 ) ;
  assign n3109 = ( n2922 & ~n3107 ) | ( n2922 & n3108 ) | ( ~n3107 & n3108 ) ;
  assign n3110 = ( ~n396 & n3104 ) | ( ~n396 & n3109 ) | ( n3104 & n3109 ) ;
  assign n3111 = n396 & ~n2923 ;
  assign n3112 = ( n396 & ~n2923 ) | ( n396 & n2979 ) | ( ~n2923 & n2979 ) ;
  assign n3113 = ( n2928 & n3111 ) | ( n2928 & n3112 ) | ( n3111 & n3112 ) ;
  assign n3114 = ( ~n2928 & n3111 ) | ( ~n2928 & n3112 ) | ( n3111 & n3112 ) ;
  assign n3115 = ( n2928 & ~n3113 ) | ( n2928 & n3114 ) | ( ~n3113 & n3114 ) ;
  assign n3116 = ( ~n344 & n3110 ) | ( ~n344 & n3115 ) | ( n3110 & n3115 ) ;
  assign n3117 = n344 & ~n2929 ;
  assign n3118 = ( n344 & ~n2929 ) | ( n344 & n2979 ) | ( ~n2929 & n2979 ) ;
  assign n3119 = ( ~n2934 & n3117 ) | ( ~n2934 & n3118 ) | ( n3117 & n3118 ) ;
  assign n3120 = ( n2934 & n3117 ) | ( n2934 & n3118 ) | ( n3117 & n3118 ) ;
  assign n3121 = ( n2934 & n3119 ) | ( n2934 & ~n3120 ) | ( n3119 & ~n3120 ) ;
  assign n3122 = ( ~n298 & n3116 ) | ( ~n298 & n3121 ) | ( n3116 & n3121 ) ;
  assign n3123 = ( n298 & ~n2935 ) | ( n298 & n2979 ) | ( ~n2935 & n2979 ) ;
  assign n3124 = n298 & ~n2935 ;
  assign n3125 = ( n2940 & n3123 ) | ( n2940 & n3124 ) | ( n3123 & n3124 ) ;
  assign n3126 = ( ~n2940 & n3123 ) | ( ~n2940 & n3124 ) | ( n3123 & n3124 ) ;
  assign n3127 = ( n2940 & ~n3125 ) | ( n2940 & n3126 ) | ( ~n3125 & n3126 ) ;
  assign n3128 = ( ~n258 & n3122 ) | ( ~n258 & n3127 ) | ( n3122 & n3127 ) ;
  assign n3129 = ( n258 & ~n2941 ) | ( n258 & n2979 ) | ( ~n2941 & n2979 ) ;
  assign n3130 = n258 & ~n2941 ;
  assign n3131 = ( n2946 & n3129 ) | ( n2946 & n3130 ) | ( n3129 & n3130 ) ;
  assign n3132 = ( ~n2946 & n3129 ) | ( ~n2946 & n3130 ) | ( n3129 & n3130 ) ;
  assign n3133 = ( n2946 & ~n3131 ) | ( n2946 & n3132 ) | ( ~n3131 & n3132 ) ;
  assign n3134 = ( ~n225 & n3128 ) | ( ~n225 & n3133 ) | ( n3128 & n3133 ) ;
  assign n3135 = ( n225 & ~n2947 ) | ( n225 & n2979 ) | ( ~n2947 & n2979 ) ;
  assign n3136 = n225 & ~n2947 ;
  assign n3137 = ( n2952 & n3135 ) | ( n2952 & n3136 ) | ( n3135 & n3136 ) ;
  assign n3138 = ( ~n2952 & n3135 ) | ( ~n2952 & n3136 ) | ( n3135 & n3136 ) ;
  assign n3139 = ( n2952 & ~n3137 ) | ( n2952 & n3138 ) | ( ~n3137 & n3138 ) ;
  assign n3140 = ( ~n197 & n3134 ) | ( ~n197 & n3139 ) | ( n3134 & n3139 ) ;
  assign n3141 = ( n197 & ~n2953 ) | ( n197 & n2979 ) | ( ~n2953 & n2979 ) ;
  assign n3142 = n197 & ~n2953 ;
  assign n3143 = ( n2958 & n3141 ) | ( n2958 & n3142 ) | ( n3141 & n3142 ) ;
  assign n3144 = ( ~n2958 & n3141 ) | ( ~n2958 & n3142 ) | ( n3141 & n3142 ) ;
  assign n3145 = ( n2958 & ~n3143 ) | ( n2958 & n3144 ) | ( ~n3143 & n3144 ) ;
  assign n3146 = ( ~n170 & n3140 ) | ( ~n170 & n3145 ) | ( n3140 & n3145 ) ;
  assign n3147 = ( n170 & ~n2959 ) | ( n170 & n2979 ) | ( ~n2959 & n2979 ) ;
  assign n3148 = n170 & ~n2959 ;
  assign n3149 = ( n2964 & n3147 ) | ( n2964 & n3148 ) | ( n3147 & n3148 ) ;
  assign n3150 = ( ~n2964 & n3147 ) | ( ~n2964 & n3148 ) | ( n3147 & n3148 ) ;
  assign n3151 = ( n2964 & ~n3149 ) | ( n2964 & n3150 ) | ( ~n3149 & n3150 ) ;
  assign n3152 = ( ~n142 & n3146 ) | ( ~n142 & n3151 ) | ( n3146 & n3151 ) ;
  assign n3153 = ( ~n132 & n2984 ) | ( ~n132 & n3152 ) | ( n2984 & n3152 ) ;
  assign n3154 = n2809 & ~n2977 ;
  assign n3155 = n2804 | n2809 ;
  assign n3156 = ~n2809 & n2977 ;
  assign n3157 = ( n3154 & n3155 ) | ( n3154 & n3156 ) | ( n3155 & n3156 ) ;
  assign n3158 = n131 & ~n3157 ;
  assign n3159 = ( n132 & ~n2971 ) | ( n132 & n2979 ) | ( ~n2971 & n2979 ) ;
  assign n3160 = n132 & ~n2971 ;
  assign n3161 = ( n2976 & n3159 ) | ( n2976 & n3160 ) | ( n3159 & n3160 ) ;
  assign n3162 = ( ~n2976 & n3159 ) | ( ~n2976 & n3160 ) | ( n3159 & n3160 ) ;
  assign n3163 = ( n2976 & ~n3161 ) | ( n2976 & n3162 ) | ( ~n3161 & n3162 ) ;
  assign n3164 = ( n2809 & ~n2977 ) | ( n2809 & n3155 ) | ( ~n2977 & n3155 ) ;
  assign n3165 = ( ~n3154 & n3163 ) | ( ~n3154 & n3164 ) | ( n3163 & n3164 ) ;
  assign n3166 = n131 & n3157 ;
  assign n3167 = ( ~n3158 & n3165 ) | ( ~n3158 & n3166 ) | ( n3165 & n3166 ) ;
  assign n3168 = n3158 & ~n3163 ;
  assign n3169 = ( n3153 & n3167 ) | ( n3153 & ~n3168 ) | ( n3167 & ~n3168 ) ;
  assign n3170 = ( ~n131 & n3153 ) | ( ~n131 & n3163 ) | ( n3153 & n3163 ) ;
  assign n3171 = ( ~n131 & n3163 ) | ( ~n131 & n3165 ) | ( n3163 & n3165 ) ;
  assign n3172 = ( n131 & ~n3158 ) | ( n131 & n3163 ) | ( ~n3158 & n3163 ) ;
  assign n3173 = ( n131 & ~n3153 ) | ( n131 & n3163 ) | ( ~n3153 & n3163 ) ;
  assign n3174 = n3172 & ~n3173 ;
  assign n3175 = ( ~n3170 & n3171 ) | ( ~n3170 & n3174 ) | ( n3171 & n3174 ) ;
  assign n3176 = x62 | x63 ;
  assign n3177 = x64 | n3176 ;
  assign n3178 = ~n2979 & n3177 ;
  assign n3179 = ( x65 & ~n3169 ) | ( x65 & n3178 ) | ( ~n3169 & n3178 ) ;
  assign n3180 = ~n2986 & n3169 ;
  assign n3181 = n2979 & ~n3177 ;
  assign n3182 = ( n3179 & n3180 ) | ( n3179 & ~n3181 ) | ( n3180 & ~n3181 ) ;
  assign n3183 = n2979 & ~n3169 ;
  assign n3184 = ( x66 & n3180 ) | ( x66 & n3183 ) | ( n3180 & n3183 ) ;
  assign n3185 = ( ~x66 & n3180 ) | ( ~x66 & n3183 ) | ( n3180 & n3183 ) ;
  assign n3186 = ( x66 & ~n3184 ) | ( x66 & n3185 ) | ( ~n3184 & n3185 ) ;
  assign n3187 = ( ~n2791 & n3182 ) | ( ~n2791 & n3186 ) | ( n3182 & n3186 ) ;
  assign n3188 = ~n2791 & n2979 ;
  assign n3189 = ( n2992 & n3169 ) | ( n2992 & n3188 ) | ( n3169 & n3188 ) ;
  assign n3190 = ( ~x67 & n3185 ) | ( ~x67 & n3189 ) | ( n3185 & n3189 ) ;
  assign n3191 = ( x67 & n3185 ) | ( x67 & n3189 ) | ( n3185 & n3189 ) ;
  assign n3192 = ( x67 & n3190 ) | ( x67 & ~n3191 ) | ( n3190 & ~n3191 ) ;
  assign n3193 = ( ~n2615 & n3187 ) | ( ~n2615 & n3192 ) | ( n3187 & n3192 ) ;
  assign n3194 = ( n2615 & ~n2991 ) | ( n2615 & n3169 ) | ( ~n2991 & n3169 ) ;
  assign n3195 = n2615 & ~n2991 ;
  assign n3196 = ( n2995 & n3194 ) | ( n2995 & n3195 ) | ( n3194 & n3195 ) ;
  assign n3197 = ( ~n2995 & n3194 ) | ( ~n2995 & n3195 ) | ( n3194 & n3195 ) ;
  assign n3198 = ( n2995 & ~n3196 ) | ( n2995 & n3197 ) | ( ~n3196 & n3197 ) ;
  assign n3199 = ( ~n2443 & n3193 ) | ( ~n2443 & n3198 ) | ( n3193 & n3198 ) ;
  assign n3200 = n2443 & ~n2996 ;
  assign n3201 = ( n2443 & ~n2996 ) | ( n2443 & n3169 ) | ( ~n2996 & n3169 ) ;
  assign n3202 = ( n3001 & n3200 ) | ( n3001 & n3201 ) | ( n3200 & n3201 ) ;
  assign n3203 = ( ~n3001 & n3200 ) | ( ~n3001 & n3201 ) | ( n3200 & n3201 ) ;
  assign n3204 = ( n3001 & ~n3202 ) | ( n3001 & n3203 ) | ( ~n3202 & n3203 ) ;
  assign n3205 = ( ~n2277 & n3199 ) | ( ~n2277 & n3204 ) | ( n3199 & n3204 ) ;
  assign n3206 = ( n2277 & ~n3002 ) | ( n2277 & n3169 ) | ( ~n3002 & n3169 ) ;
  assign n3207 = n2277 & ~n3002 ;
  assign n3208 = ( n3007 & n3206 ) | ( n3007 & n3207 ) | ( n3206 & n3207 ) ;
  assign n3209 = ( ~n3007 & n3206 ) | ( ~n3007 & n3207 ) | ( n3206 & n3207 ) ;
  assign n3210 = ( n3007 & ~n3208 ) | ( n3007 & n3209 ) | ( ~n3208 & n3209 ) ;
  assign n3211 = ( ~n2111 & n3205 ) | ( ~n2111 & n3210 ) | ( n3205 & n3210 ) ;
  assign n3212 = ~n2111 & n3008 ;
  assign n3213 = ( ~n2111 & n3008 ) | ( ~n2111 & n3169 ) | ( n3008 & n3169 ) ;
  assign n3214 = ( n3013 & n3212 ) | ( n3013 & n3213 ) | ( n3212 & n3213 ) ;
  assign n3215 = ( ~n3013 & n3212 ) | ( ~n3013 & n3213 ) | ( n3212 & n3213 ) ;
  assign n3216 = ( n3013 & ~n3214 ) | ( n3013 & n3215 ) | ( ~n3214 & n3215 ) ;
  assign n3217 = ( ~n1949 & n3211 ) | ( ~n1949 & n3216 ) | ( n3211 & n3216 ) ;
  assign n3218 = n1949 & ~n3014 ;
  assign n3219 = ( n1949 & ~n3014 ) | ( n1949 & n3169 ) | ( ~n3014 & n3169 ) ;
  assign n3220 = ( n3019 & n3218 ) | ( n3019 & n3219 ) | ( n3218 & n3219 ) ;
  assign n3221 = ( ~n3019 & n3218 ) | ( ~n3019 & n3219 ) | ( n3218 & n3219 ) ;
  assign n3222 = ( n3019 & ~n3220 ) | ( n3019 & n3221 ) | ( ~n3220 & n3221 ) ;
  assign n3223 = ( ~n1802 & n3217 ) | ( ~n1802 & n3222 ) | ( n3217 & n3222 ) ;
  assign n3224 = ~n1802 & n3020 ;
  assign n3225 = ( ~n1802 & n3020 ) | ( ~n1802 & n3169 ) | ( n3020 & n3169 ) ;
  assign n3226 = ( n3025 & n3224 ) | ( n3025 & n3225 ) | ( n3224 & n3225 ) ;
  assign n3227 = ( ~n3025 & n3224 ) | ( ~n3025 & n3225 ) | ( n3224 & n3225 ) ;
  assign n3228 = ( n3025 & ~n3226 ) | ( n3025 & n3227 ) | ( ~n3226 & n3227 ) ;
  assign n3229 = ( ~n1661 & n3223 ) | ( ~n1661 & n3228 ) | ( n3223 & n3228 ) ;
  assign n3230 = ~n1661 & n3026 ;
  assign n3231 = ( ~n1661 & n3026 ) | ( ~n1661 & n3169 ) | ( n3026 & n3169 ) ;
  assign n3232 = ( ~n3031 & n3230 ) | ( ~n3031 & n3231 ) | ( n3230 & n3231 ) ;
  assign n3233 = ( n3031 & n3230 ) | ( n3031 & n3231 ) | ( n3230 & n3231 ) ;
  assign n3234 = ( n3031 & n3232 ) | ( n3031 & ~n3233 ) | ( n3232 & ~n3233 ) ;
  assign n3235 = ( ~n1523 & n3229 ) | ( ~n1523 & n3234 ) | ( n3229 & n3234 ) ;
  assign n3236 = ( n1523 & ~n3032 ) | ( n1523 & n3169 ) | ( ~n3032 & n3169 ) ;
  assign n3237 = n1523 & ~n3032 ;
  assign n3238 = ( n3037 & n3236 ) | ( n3037 & n3237 ) | ( n3236 & n3237 ) ;
  assign n3239 = ( ~n3037 & n3236 ) | ( ~n3037 & n3237 ) | ( n3236 & n3237 ) ;
  assign n3240 = ( n3037 & ~n3238 ) | ( n3037 & n3239 ) | ( ~n3238 & n3239 ) ;
  assign n3241 = ( ~n1393 & n3235 ) | ( ~n1393 & n3240 ) | ( n3235 & n3240 ) ;
  assign n3242 = ( n1393 & ~n3038 ) | ( n1393 & n3169 ) | ( ~n3038 & n3169 ) ;
  assign n3243 = n1393 & ~n3038 ;
  assign n3244 = ( n3043 & n3242 ) | ( n3043 & n3243 ) | ( n3242 & n3243 ) ;
  assign n3245 = ( ~n3043 & n3242 ) | ( ~n3043 & n3243 ) | ( n3242 & n3243 ) ;
  assign n3246 = ( n3043 & ~n3244 ) | ( n3043 & n3245 ) | ( ~n3244 & n3245 ) ;
  assign n3247 = ( ~n1266 & n3241 ) | ( ~n1266 & n3246 ) | ( n3241 & n3246 ) ;
  assign n3248 = ( n1266 & ~n3044 ) | ( n1266 & n3169 ) | ( ~n3044 & n3169 ) ;
  assign n3249 = n1266 & ~n3044 ;
  assign n3250 = ( n3049 & n3248 ) | ( n3049 & n3249 ) | ( n3248 & n3249 ) ;
  assign n3251 = ( ~n3049 & n3248 ) | ( ~n3049 & n3249 ) | ( n3248 & n3249 ) ;
  assign n3252 = ( n3049 & ~n3250 ) | ( n3049 & n3251 ) | ( ~n3250 & n3251 ) ;
  assign n3253 = ( ~n1150 & n3247 ) | ( ~n1150 & n3252 ) | ( n3247 & n3252 ) ;
  assign n3254 = ( n1150 & ~n3050 ) | ( n1150 & n3169 ) | ( ~n3050 & n3169 ) ;
  assign n3255 = n1150 & ~n3050 ;
  assign n3256 = ( n3055 & n3254 ) | ( n3055 & n3255 ) | ( n3254 & n3255 ) ;
  assign n3257 = ( ~n3055 & n3254 ) | ( ~n3055 & n3255 ) | ( n3254 & n3255 ) ;
  assign n3258 = ( n3055 & ~n3256 ) | ( n3055 & n3257 ) | ( ~n3256 & n3257 ) ;
  assign n3259 = ( ~n1038 & n3253 ) | ( ~n1038 & n3258 ) | ( n3253 & n3258 ) ;
  assign n3260 = ( ~n1038 & n3056 ) | ( ~n1038 & n3169 ) | ( n3056 & n3169 ) ;
  assign n3261 = ~n1038 & n3056 ;
  assign n3262 = ( ~n3061 & n3260 ) | ( ~n3061 & n3261 ) | ( n3260 & n3261 ) ;
  assign n3263 = ( n3061 & n3260 ) | ( n3061 & n3261 ) | ( n3260 & n3261 ) ;
  assign n3264 = ( n3061 & n3262 ) | ( n3061 & ~n3263 ) | ( n3262 & ~n3263 ) ;
  assign n3265 = ( ~n933 & n3259 ) | ( ~n933 & n3264 ) | ( n3259 & n3264 ) ;
  assign n3266 = ( n933 & ~n3062 ) | ( n933 & n3169 ) | ( ~n3062 & n3169 ) ;
  assign n3267 = n933 & ~n3062 ;
  assign n3268 = ( n3067 & n3266 ) | ( n3067 & n3267 ) | ( n3266 & n3267 ) ;
  assign n3269 = ( ~n3067 & n3266 ) | ( ~n3067 & n3267 ) | ( n3266 & n3267 ) ;
  assign n3270 = ( n3067 & ~n3268 ) | ( n3067 & n3269 ) | ( ~n3268 & n3269 ) ;
  assign n3271 = ( ~n839 & n3265 ) | ( ~n839 & n3270 ) | ( n3265 & n3270 ) ;
  assign n3272 = ( n839 & ~n3068 ) | ( n839 & n3169 ) | ( ~n3068 & n3169 ) ;
  assign n3273 = n839 & ~n3068 ;
  assign n3274 = ( n3073 & n3272 ) | ( n3073 & n3273 ) | ( n3272 & n3273 ) ;
  assign n3275 = ( ~n3073 & n3272 ) | ( ~n3073 & n3273 ) | ( n3272 & n3273 ) ;
  assign n3276 = ( n3073 & ~n3274 ) | ( n3073 & n3275 ) | ( ~n3274 & n3275 ) ;
  assign n3277 = ( ~n746 & n3271 ) | ( ~n746 & n3276 ) | ( n3271 & n3276 ) ;
  assign n3278 = ~n746 & n3074 ;
  assign n3279 = ( ~n746 & n3074 ) | ( ~n746 & n3169 ) | ( n3074 & n3169 ) ;
  assign n3280 = ( n3079 & n3278 ) | ( n3079 & n3279 ) | ( n3278 & n3279 ) ;
  assign n3281 = ( ~n3079 & n3278 ) | ( ~n3079 & n3279 ) | ( n3278 & n3279 ) ;
  assign n3282 = ( n3079 & ~n3280 ) | ( n3079 & n3281 ) | ( ~n3280 & n3281 ) ;
  assign n3283 = ( ~n664 & n3277 ) | ( ~n664 & n3282 ) | ( n3277 & n3282 ) ;
  assign n3284 = ( n664 & ~n3080 ) | ( n664 & n3169 ) | ( ~n3080 & n3169 ) ;
  assign n3285 = n664 & ~n3080 ;
  assign n3286 = ( n3085 & n3284 ) | ( n3085 & n3285 ) | ( n3284 & n3285 ) ;
  assign n3287 = ( ~n3085 & n3284 ) | ( ~n3085 & n3285 ) | ( n3284 & n3285 ) ;
  assign n3288 = ( n3085 & ~n3286 ) | ( n3085 & n3287 ) | ( ~n3286 & n3287 ) ;
  assign n3289 = ( ~n588 & n3283 ) | ( ~n588 & n3288 ) | ( n3283 & n3288 ) ;
  assign n3290 = ( n588 & ~n3086 ) | ( n588 & n3169 ) | ( ~n3086 & n3169 ) ;
  assign n3291 = n588 & ~n3086 ;
  assign n3292 = ( n3091 & n3290 ) | ( n3091 & n3291 ) | ( n3290 & n3291 ) ;
  assign n3293 = ( ~n3091 & n3290 ) | ( ~n3091 & n3291 ) | ( n3290 & n3291 ) ;
  assign n3294 = ( n3091 & ~n3292 ) | ( n3091 & n3293 ) | ( ~n3292 & n3293 ) ;
  assign n3295 = ( ~n518 & n3289 ) | ( ~n518 & n3294 ) | ( n3289 & n3294 ) ;
  assign n3296 = ~n518 & n3092 ;
  assign n3297 = ( ~n518 & n3092 ) | ( ~n518 & n3169 ) | ( n3092 & n3169 ) ;
  assign n3298 = ( n3097 & n3296 ) | ( n3097 & n3297 ) | ( n3296 & n3297 ) ;
  assign n3299 = ( ~n3097 & n3296 ) | ( ~n3097 & n3297 ) | ( n3296 & n3297 ) ;
  assign n3300 = ( n3097 & ~n3298 ) | ( n3097 & n3299 ) | ( ~n3298 & n3299 ) ;
  assign n3301 = ( ~n454 & n3295 ) | ( ~n454 & n3300 ) | ( n3295 & n3300 ) ;
  assign n3302 = ( n454 & ~n3098 ) | ( n454 & n3169 ) | ( ~n3098 & n3169 ) ;
  assign n3303 = n454 & ~n3098 ;
  assign n3304 = ( n3103 & n3302 ) | ( n3103 & n3303 ) | ( n3302 & n3303 ) ;
  assign n3305 = ( ~n3103 & n3302 ) | ( ~n3103 & n3303 ) | ( n3302 & n3303 ) ;
  assign n3306 = ( n3103 & ~n3304 ) | ( n3103 & n3305 ) | ( ~n3304 & n3305 ) ;
  assign n3307 = ( ~n396 & n3301 ) | ( ~n396 & n3306 ) | ( n3301 & n3306 ) ;
  assign n3308 = ( n396 & ~n3104 ) | ( n396 & n3169 ) | ( ~n3104 & n3169 ) ;
  assign n3309 = n396 & ~n3104 ;
  assign n3310 = ( n3109 & n3308 ) | ( n3109 & n3309 ) | ( n3308 & n3309 ) ;
  assign n3311 = ( ~n3109 & n3308 ) | ( ~n3109 & n3309 ) | ( n3308 & n3309 ) ;
  assign n3312 = ( n3109 & ~n3310 ) | ( n3109 & n3311 ) | ( ~n3310 & n3311 ) ;
  assign n3313 = ( ~n344 & n3307 ) | ( ~n344 & n3312 ) | ( n3307 & n3312 ) ;
  assign n3314 = ~n344 & n3110 ;
  assign n3315 = ( ~n344 & n3110 ) | ( ~n344 & n3169 ) | ( n3110 & n3169 ) ;
  assign n3316 = ( ~n3115 & n3314 ) | ( ~n3115 & n3315 ) | ( n3314 & n3315 ) ;
  assign n3317 = ( n3115 & n3314 ) | ( n3115 & n3315 ) | ( n3314 & n3315 ) ;
  assign n3318 = ( n3115 & n3316 ) | ( n3115 & ~n3317 ) | ( n3316 & ~n3317 ) ;
  assign n3319 = ( ~n298 & n3313 ) | ( ~n298 & n3318 ) | ( n3313 & n3318 ) ;
  assign n3320 = ( n298 & ~n3116 ) | ( n298 & n3169 ) | ( ~n3116 & n3169 ) ;
  assign n3321 = n298 & ~n3116 ;
  assign n3322 = ( n3121 & n3320 ) | ( n3121 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3323 = ( ~n3121 & n3320 ) | ( ~n3121 & n3321 ) | ( n3320 & n3321 ) ;
  assign n3324 = ( n3121 & ~n3322 ) | ( n3121 & n3323 ) | ( ~n3322 & n3323 ) ;
  assign n3325 = ( ~n258 & n3319 ) | ( ~n258 & n3324 ) | ( n3319 & n3324 ) ;
  assign n3326 = ~n258 & n3122 ;
  assign n3327 = ( ~n258 & n3122 ) | ( ~n258 & n3169 ) | ( n3122 & n3169 ) ;
  assign n3328 = ( ~n3127 & n3326 ) | ( ~n3127 & n3327 ) | ( n3326 & n3327 ) ;
  assign n3329 = ( n3127 & n3326 ) | ( n3127 & n3327 ) | ( n3326 & n3327 ) ;
  assign n3330 = ( n3127 & n3328 ) | ( n3127 & ~n3329 ) | ( n3328 & ~n3329 ) ;
  assign n3331 = ( ~n225 & n3325 ) | ( ~n225 & n3330 ) | ( n3325 & n3330 ) ;
  assign n3332 = ( n225 & ~n3128 ) | ( n225 & n3169 ) | ( ~n3128 & n3169 ) ;
  assign n3333 = n225 & ~n3128 ;
  assign n3334 = ( n3133 & n3332 ) | ( n3133 & n3333 ) | ( n3332 & n3333 ) ;
  assign n3335 = ( ~n3133 & n3332 ) | ( ~n3133 & n3333 ) | ( n3332 & n3333 ) ;
  assign n3336 = ( n3133 & ~n3334 ) | ( n3133 & n3335 ) | ( ~n3334 & n3335 ) ;
  assign n3337 = ( ~n197 & n3331 ) | ( ~n197 & n3336 ) | ( n3331 & n3336 ) ;
  assign n3338 = ( n197 & ~n3134 ) | ( n197 & n3169 ) | ( ~n3134 & n3169 ) ;
  assign n3339 = n197 & ~n3134 ;
  assign n3340 = ( n3139 & n3338 ) | ( n3139 & n3339 ) | ( n3338 & n3339 ) ;
  assign n3341 = ( ~n3139 & n3338 ) | ( ~n3139 & n3339 ) | ( n3338 & n3339 ) ;
  assign n3342 = ( n3139 & ~n3340 ) | ( n3139 & n3341 ) | ( ~n3340 & n3341 ) ;
  assign n3343 = ( ~n170 & n3337 ) | ( ~n170 & n3342 ) | ( n3337 & n3342 ) ;
  assign n3344 = ~n170 & n3140 ;
  assign n3345 = ( ~n170 & n3140 ) | ( ~n170 & n3169 ) | ( n3140 & n3169 ) ;
  assign n3346 = ( ~n3145 & n3344 ) | ( ~n3145 & n3345 ) | ( n3344 & n3345 ) ;
  assign n3347 = ( n3145 & n3344 ) | ( n3145 & n3345 ) | ( n3344 & n3345 ) ;
  assign n3348 = ( n3145 & n3346 ) | ( n3145 & ~n3347 ) | ( n3346 & ~n3347 ) ;
  assign n3349 = ( ~n142 & n3343 ) | ( ~n142 & n3348 ) | ( n3343 & n3348 ) ;
  assign n3350 = ~n142 & n3146 ;
  assign n3351 = ( ~n142 & n3146 ) | ( ~n142 & n3169 ) | ( n3146 & n3169 ) ;
  assign n3352 = ( ~n3151 & n3350 ) | ( ~n3151 & n3351 ) | ( n3350 & n3351 ) ;
  assign n3353 = ( n3151 & n3350 ) | ( n3151 & n3351 ) | ( n3350 & n3351 ) ;
  assign n3354 = ( n3151 & n3352 ) | ( n3151 & ~n3353 ) | ( n3352 & ~n3353 ) ;
  assign n3355 = ( ~n132 & n3349 ) | ( ~n132 & n3354 ) | ( n3349 & n3354 ) ;
  assign n3356 = ( ~n132 & n3152 ) | ( ~n132 & n3169 ) | ( n3152 & n3169 ) ;
  assign n3357 = ~n132 & n3152 ;
  assign n3358 = ( ~n2984 & n3356 ) | ( ~n2984 & n3357 ) | ( n3356 & n3357 ) ;
  assign n3359 = ( n2984 & n3356 ) | ( n2984 & n3357 ) | ( n3356 & n3357 ) ;
  assign n3360 = ( n2984 & n3358 ) | ( n2984 & ~n3359 ) | ( n3358 & ~n3359 ) ;
  assign n3361 = ( ~n131 & n3355 ) | ( ~n131 & n3360 ) | ( n3355 & n3360 ) ;
  assign n3362 = n3175 | n3361 ;
  assign n3363 = ~n3355 & n3360 ;
  assign n3364 = n3153 | n3163 ;
  assign n3365 = ( n3355 & n3360 ) | ( n3355 & ~n3364 ) | ( n3360 & ~n3364 ) ;
  assign n3366 = n3157 & ~n3163 ;
  assign n3367 = n3153 & ~n3366 ;
  assign n3368 = ( n3355 & n3360 ) | ( n3355 & ~n3367 ) | ( n3360 & ~n3367 ) ;
  assign n3369 = ( n3363 & ~n3365 ) | ( n3363 & n3368 ) | ( ~n3365 & n3368 ) ;
  assign n3370 = n131 & ~n3369 ;
  assign n3371 = x60 | x61 ;
  assign n3372 = x62 | n3371 ;
  assign n3373 = n3169 & ~n3372 ;
  assign n3374 = ~n3176 & n3362 ;
  assign n3375 = ~n3169 & n3372 ;
  assign n3376 = ( x63 & ~n3362 ) | ( x63 & n3375 ) | ( ~n3362 & n3375 ) ;
  assign n3377 = ( ~n3373 & n3374 ) | ( ~n3373 & n3376 ) | ( n3374 & n3376 ) ;
  assign n3378 = n3169 & ~n3362 ;
  assign n3379 = ( ~x64 & n3374 ) | ( ~x64 & n3378 ) | ( n3374 & n3378 ) ;
  assign n3380 = ( x64 & n3374 ) | ( x64 & n3378 ) | ( n3374 & n3378 ) ;
  assign n3381 = ( x64 & n3379 ) | ( x64 & ~n3380 ) | ( n3379 & ~n3380 ) ;
  assign n3382 = ( ~n2979 & n3377 ) | ( ~n2979 & n3381 ) | ( n3377 & n3381 ) ;
  assign n3383 = ~n2979 & n3169 ;
  assign n3384 = ( n3183 & n3362 ) | ( n3183 & n3383 ) | ( n3362 & n3383 ) ;
  assign n3385 = ( x65 & n3379 ) | ( x65 & n3384 ) | ( n3379 & n3384 ) ;
  assign n3386 = ( ~x65 & n3379 ) | ( ~x65 & n3384 ) | ( n3379 & n3384 ) ;
  assign n3387 = ( x65 & ~n3385 ) | ( x65 & n3386 ) | ( ~n3385 & n3386 ) ;
  assign n3388 = ( ~n2791 & n3382 ) | ( ~n2791 & n3387 ) | ( n3382 & n3387 ) ;
  assign n3389 = n2791 & ~n3182 ;
  assign n3390 = ( n2791 & ~n3182 ) | ( n2791 & n3362 ) | ( ~n3182 & n3362 ) ;
  assign n3391 = ( ~n3186 & n3389 ) | ( ~n3186 & n3390 ) | ( n3389 & n3390 ) ;
  assign n3392 = ( n3186 & n3389 ) | ( n3186 & n3390 ) | ( n3389 & n3390 ) ;
  assign n3393 = ( n3186 & n3391 ) | ( n3186 & ~n3392 ) | ( n3391 & ~n3392 ) ;
  assign n3394 = ( ~n2615 & n3388 ) | ( ~n2615 & n3393 ) | ( n3388 & n3393 ) ;
  assign n3395 = n2615 & ~n3187 ;
  assign n3396 = ( n2615 & ~n3187 ) | ( n2615 & n3362 ) | ( ~n3187 & n3362 ) ;
  assign n3397 = ( n3192 & n3395 ) | ( n3192 & n3396 ) | ( n3395 & n3396 ) ;
  assign n3398 = ( ~n3192 & n3395 ) | ( ~n3192 & n3396 ) | ( n3395 & n3396 ) ;
  assign n3399 = ( n3192 & ~n3397 ) | ( n3192 & n3398 ) | ( ~n3397 & n3398 ) ;
  assign n3400 = ( ~n2443 & n3394 ) | ( ~n2443 & n3399 ) | ( n3394 & n3399 ) ;
  assign n3401 = ( n2443 & ~n3193 ) | ( n2443 & n3362 ) | ( ~n3193 & n3362 ) ;
  assign n3402 = n2443 & ~n3193 ;
  assign n3403 = ( n3198 & n3401 ) | ( n3198 & n3402 ) | ( n3401 & n3402 ) ;
  assign n3404 = ( ~n3198 & n3401 ) | ( ~n3198 & n3402 ) | ( n3401 & n3402 ) ;
  assign n3405 = ( n3198 & ~n3403 ) | ( n3198 & n3404 ) | ( ~n3403 & n3404 ) ;
  assign n3406 = ( ~n2277 & n3400 ) | ( ~n2277 & n3405 ) | ( n3400 & n3405 ) ;
  assign n3407 = ~n2277 & n3199 ;
  assign n3408 = ( ~n2277 & n3199 ) | ( ~n2277 & n3362 ) | ( n3199 & n3362 ) ;
  assign n3409 = ( n3204 & n3407 ) | ( n3204 & n3408 ) | ( n3407 & n3408 ) ;
  assign n3410 = ( ~n3204 & n3407 ) | ( ~n3204 & n3408 ) | ( n3407 & n3408 ) ;
  assign n3411 = ( n3204 & ~n3409 ) | ( n3204 & n3410 ) | ( ~n3409 & n3410 ) ;
  assign n3412 = ( ~n2111 & n3406 ) | ( ~n2111 & n3411 ) | ( n3406 & n3411 ) ;
  assign n3413 = ( n2111 & ~n3205 ) | ( n2111 & n3362 ) | ( ~n3205 & n3362 ) ;
  assign n3414 = n2111 & ~n3205 ;
  assign n3415 = ( n3210 & n3413 ) | ( n3210 & n3414 ) | ( n3413 & n3414 ) ;
  assign n3416 = ( ~n3210 & n3413 ) | ( ~n3210 & n3414 ) | ( n3413 & n3414 ) ;
  assign n3417 = ( n3210 & ~n3415 ) | ( n3210 & n3416 ) | ( ~n3415 & n3416 ) ;
  assign n3418 = ( ~n1949 & n3412 ) | ( ~n1949 & n3417 ) | ( n3412 & n3417 ) ;
  assign n3419 = ~n1949 & n3211 ;
  assign n3420 = ( ~n1949 & n3211 ) | ( ~n1949 & n3362 ) | ( n3211 & n3362 ) ;
  assign n3421 = ( n3216 & n3419 ) | ( n3216 & n3420 ) | ( n3419 & n3420 ) ;
  assign n3422 = ( ~n3216 & n3419 ) | ( ~n3216 & n3420 ) | ( n3419 & n3420 ) ;
  assign n3423 = ( n3216 & ~n3421 ) | ( n3216 & n3422 ) | ( ~n3421 & n3422 ) ;
  assign n3424 = ( ~n1802 & n3418 ) | ( ~n1802 & n3423 ) | ( n3418 & n3423 ) ;
  assign n3425 = ( n1802 & ~n3217 ) | ( n1802 & n3362 ) | ( ~n3217 & n3362 ) ;
  assign n3426 = n1802 & ~n3217 ;
  assign n3427 = ( n3222 & n3425 ) | ( n3222 & n3426 ) | ( n3425 & n3426 ) ;
  assign n3428 = ( ~n3222 & n3425 ) | ( ~n3222 & n3426 ) | ( n3425 & n3426 ) ;
  assign n3429 = ( n3222 & ~n3427 ) | ( n3222 & n3428 ) | ( ~n3427 & n3428 ) ;
  assign n3430 = ( ~n1661 & n3424 ) | ( ~n1661 & n3429 ) | ( n3424 & n3429 ) ;
  assign n3431 = ~n1661 & n3223 ;
  assign n3432 = ( ~n1661 & n3223 ) | ( ~n1661 & n3362 ) | ( n3223 & n3362 ) ;
  assign n3433 = ( n3228 & n3431 ) | ( n3228 & n3432 ) | ( n3431 & n3432 ) ;
  assign n3434 = ( ~n3228 & n3431 ) | ( ~n3228 & n3432 ) | ( n3431 & n3432 ) ;
  assign n3435 = ( n3228 & ~n3433 ) | ( n3228 & n3434 ) | ( ~n3433 & n3434 ) ;
  assign n3436 = ( ~n1523 & n3430 ) | ( ~n1523 & n3435 ) | ( n3430 & n3435 ) ;
  assign n3437 = ~n1523 & n3229 ;
  assign n3438 = ( ~n1523 & n3229 ) | ( ~n1523 & n3362 ) | ( n3229 & n3362 ) ;
  assign n3439 = ( ~n3234 & n3437 ) | ( ~n3234 & n3438 ) | ( n3437 & n3438 ) ;
  assign n3440 = ( n3234 & n3437 ) | ( n3234 & n3438 ) | ( n3437 & n3438 ) ;
  assign n3441 = ( n3234 & n3439 ) | ( n3234 & ~n3440 ) | ( n3439 & ~n3440 ) ;
  assign n3442 = ( ~n1393 & n3436 ) | ( ~n1393 & n3441 ) | ( n3436 & n3441 ) ;
  assign n3443 = ~n1393 & n3235 ;
  assign n3444 = ( ~n1393 & n3235 ) | ( ~n1393 & n3362 ) | ( n3235 & n3362 ) ;
  assign n3445 = ( n3240 & n3443 ) | ( n3240 & n3444 ) | ( n3443 & n3444 ) ;
  assign n3446 = ( ~n3240 & n3443 ) | ( ~n3240 & n3444 ) | ( n3443 & n3444 ) ;
  assign n3447 = ( n3240 & ~n3445 ) | ( n3240 & n3446 ) | ( ~n3445 & n3446 ) ;
  assign n3448 = ( ~n1266 & n3442 ) | ( ~n1266 & n3447 ) | ( n3442 & n3447 ) ;
  assign n3449 = ~n1266 & n3241 ;
  assign n3450 = ( ~n1266 & n3241 ) | ( ~n1266 & n3362 ) | ( n3241 & n3362 ) ;
  assign n3451 = ( n3246 & n3449 ) | ( n3246 & n3450 ) | ( n3449 & n3450 ) ;
  assign n3452 = ( ~n3246 & n3449 ) | ( ~n3246 & n3450 ) | ( n3449 & n3450 ) ;
  assign n3453 = ( n3246 & ~n3451 ) | ( n3246 & n3452 ) | ( ~n3451 & n3452 ) ;
  assign n3454 = ( ~n1150 & n3448 ) | ( ~n1150 & n3453 ) | ( n3448 & n3453 ) ;
  assign n3455 = ( n1150 & ~n3247 ) | ( n1150 & n3362 ) | ( ~n3247 & n3362 ) ;
  assign n3456 = n1150 & ~n3247 ;
  assign n3457 = ( n3252 & n3455 ) | ( n3252 & n3456 ) | ( n3455 & n3456 ) ;
  assign n3458 = ( ~n3252 & n3455 ) | ( ~n3252 & n3456 ) | ( n3455 & n3456 ) ;
  assign n3459 = ( n3252 & ~n3457 ) | ( n3252 & n3458 ) | ( ~n3457 & n3458 ) ;
  assign n3460 = ( ~n1038 & n3454 ) | ( ~n1038 & n3459 ) | ( n3454 & n3459 ) ;
  assign n3461 = n1038 & ~n3253 ;
  assign n3462 = ( n1038 & ~n3253 ) | ( n1038 & n3362 ) | ( ~n3253 & n3362 ) ;
  assign n3463 = ( ~n3258 & n3461 ) | ( ~n3258 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3464 = ( n3258 & n3461 ) | ( n3258 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3465 = ( n3258 & n3463 ) | ( n3258 & ~n3464 ) | ( n3463 & ~n3464 ) ;
  assign n3466 = ( ~n933 & n3460 ) | ( ~n933 & n3465 ) | ( n3460 & n3465 ) ;
  assign n3467 = ~n933 & n3259 ;
  assign n3468 = ( ~n933 & n3259 ) | ( ~n933 & n3362 ) | ( n3259 & n3362 ) ;
  assign n3469 = ( ~n3264 & n3467 ) | ( ~n3264 & n3468 ) | ( n3467 & n3468 ) ;
  assign n3470 = ( n3264 & n3467 ) | ( n3264 & n3468 ) | ( n3467 & n3468 ) ;
  assign n3471 = ( n3264 & n3469 ) | ( n3264 & ~n3470 ) | ( n3469 & ~n3470 ) ;
  assign n3472 = ( ~n839 & n3466 ) | ( ~n839 & n3471 ) | ( n3466 & n3471 ) ;
  assign n3473 = ( n839 & ~n3265 ) | ( n839 & n3362 ) | ( ~n3265 & n3362 ) ;
  assign n3474 = n839 & ~n3265 ;
  assign n3475 = ( n3270 & n3473 ) | ( n3270 & n3474 ) | ( n3473 & n3474 ) ;
  assign n3476 = ( ~n3270 & n3473 ) | ( ~n3270 & n3474 ) | ( n3473 & n3474 ) ;
  assign n3477 = ( n3270 & ~n3475 ) | ( n3270 & n3476 ) | ( ~n3475 & n3476 ) ;
  assign n3478 = ( ~n746 & n3472 ) | ( ~n746 & n3477 ) | ( n3472 & n3477 ) ;
  assign n3479 = ( n746 & ~n3271 ) | ( n746 & n3362 ) | ( ~n3271 & n3362 ) ;
  assign n3480 = n746 & ~n3271 ;
  assign n3481 = ( n3276 & n3479 ) | ( n3276 & n3480 ) | ( n3479 & n3480 ) ;
  assign n3482 = ( ~n3276 & n3479 ) | ( ~n3276 & n3480 ) | ( n3479 & n3480 ) ;
  assign n3483 = ( n3276 & ~n3481 ) | ( n3276 & n3482 ) | ( ~n3481 & n3482 ) ;
  assign n3484 = ( ~n664 & n3478 ) | ( ~n664 & n3483 ) | ( n3478 & n3483 ) ;
  assign n3485 = ~n664 & n3277 ;
  assign n3486 = ( ~n664 & n3277 ) | ( ~n664 & n3362 ) | ( n3277 & n3362 ) ;
  assign n3487 = ( ~n3282 & n3485 ) | ( ~n3282 & n3486 ) | ( n3485 & n3486 ) ;
  assign n3488 = ( n3282 & n3485 ) | ( n3282 & n3486 ) | ( n3485 & n3486 ) ;
  assign n3489 = ( n3282 & n3487 ) | ( n3282 & ~n3488 ) | ( n3487 & ~n3488 ) ;
  assign n3490 = ( ~n588 & n3484 ) | ( ~n588 & n3489 ) | ( n3484 & n3489 ) ;
  assign n3491 = ( n588 & ~n3283 ) | ( n588 & n3362 ) | ( ~n3283 & n3362 ) ;
  assign n3492 = n588 & ~n3283 ;
  assign n3493 = ( n3288 & n3491 ) | ( n3288 & n3492 ) | ( n3491 & n3492 ) ;
  assign n3494 = ( ~n3288 & n3491 ) | ( ~n3288 & n3492 ) | ( n3491 & n3492 ) ;
  assign n3495 = ( n3288 & ~n3493 ) | ( n3288 & n3494 ) | ( ~n3493 & n3494 ) ;
  assign n3496 = ( ~n518 & n3490 ) | ( ~n518 & n3495 ) | ( n3490 & n3495 ) ;
  assign n3497 = ~n518 & n3289 ;
  assign n3498 = ( ~n518 & n3289 ) | ( ~n518 & n3362 ) | ( n3289 & n3362 ) ;
  assign n3499 = ( ~n3294 & n3497 ) | ( ~n3294 & n3498 ) | ( n3497 & n3498 ) ;
  assign n3500 = ( n3294 & n3497 ) | ( n3294 & n3498 ) | ( n3497 & n3498 ) ;
  assign n3501 = ( n3294 & n3499 ) | ( n3294 & ~n3500 ) | ( n3499 & ~n3500 ) ;
  assign n3502 = ( ~n454 & n3496 ) | ( ~n454 & n3501 ) | ( n3496 & n3501 ) ;
  assign n3503 = ~n454 & n3295 ;
  assign n3504 = ( ~n454 & n3295 ) | ( ~n454 & n3362 ) | ( n3295 & n3362 ) ;
  assign n3505 = ( n3300 & n3503 ) | ( n3300 & n3504 ) | ( n3503 & n3504 ) ;
  assign n3506 = ( ~n3300 & n3503 ) | ( ~n3300 & n3504 ) | ( n3503 & n3504 ) ;
  assign n3507 = ( n3300 & ~n3505 ) | ( n3300 & n3506 ) | ( ~n3505 & n3506 ) ;
  assign n3508 = ( ~n396 & n3502 ) | ( ~n396 & n3507 ) | ( n3502 & n3507 ) ;
  assign n3509 = n396 & ~n3301 ;
  assign n3510 = ( n396 & ~n3301 ) | ( n396 & n3362 ) | ( ~n3301 & n3362 ) ;
  assign n3511 = ( ~n3306 & n3509 ) | ( ~n3306 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3512 = ( n3306 & n3509 ) | ( n3306 & n3510 ) | ( n3509 & n3510 ) ;
  assign n3513 = ( n3306 & n3511 ) | ( n3306 & ~n3512 ) | ( n3511 & ~n3512 ) ;
  assign n3514 = ( ~n344 & n3508 ) | ( ~n344 & n3513 ) | ( n3508 & n3513 ) ;
  assign n3515 = n344 & ~n3307 ;
  assign n3516 = ( n344 & ~n3307 ) | ( n344 & n3362 ) | ( ~n3307 & n3362 ) ;
  assign n3517 = ( n3312 & n3515 ) | ( n3312 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3518 = ( ~n3312 & n3515 ) | ( ~n3312 & n3516 ) | ( n3515 & n3516 ) ;
  assign n3519 = ( n3312 & ~n3517 ) | ( n3312 & n3518 ) | ( ~n3517 & n3518 ) ;
  assign n3520 = ( ~n298 & n3514 ) | ( ~n298 & n3519 ) | ( n3514 & n3519 ) ;
  assign n3521 = ( n298 & ~n3313 ) | ( n298 & n3362 ) | ( ~n3313 & n3362 ) ;
  assign n3522 = n298 & ~n3313 ;
  assign n3523 = ( n3318 & n3521 ) | ( n3318 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3524 = ( ~n3318 & n3521 ) | ( ~n3318 & n3522 ) | ( n3521 & n3522 ) ;
  assign n3525 = ( n3318 & ~n3523 ) | ( n3318 & n3524 ) | ( ~n3523 & n3524 ) ;
  assign n3526 = ( ~n258 & n3520 ) | ( ~n258 & n3525 ) | ( n3520 & n3525 ) ;
  assign n3527 = ~n258 & n3319 ;
  assign n3528 = ( ~n258 & n3319 ) | ( ~n258 & n3362 ) | ( n3319 & n3362 ) ;
  assign n3529 = ( ~n3324 & n3527 ) | ( ~n3324 & n3528 ) | ( n3527 & n3528 ) ;
  assign n3530 = ( n3324 & n3527 ) | ( n3324 & n3528 ) | ( n3527 & n3528 ) ;
  assign n3531 = ( n3324 & n3529 ) | ( n3324 & ~n3530 ) | ( n3529 & ~n3530 ) ;
  assign n3532 = ( ~n225 & n3526 ) | ( ~n225 & n3531 ) | ( n3526 & n3531 ) ;
  assign n3533 = ( n225 & ~n3325 ) | ( n225 & n3362 ) | ( ~n3325 & n3362 ) ;
  assign n3534 = n225 & ~n3325 ;
  assign n3535 = ( n3330 & n3533 ) | ( n3330 & n3534 ) | ( n3533 & n3534 ) ;
  assign n3536 = ( ~n3330 & n3533 ) | ( ~n3330 & n3534 ) | ( n3533 & n3534 ) ;
  assign n3537 = ( n3330 & ~n3535 ) | ( n3330 & n3536 ) | ( ~n3535 & n3536 ) ;
  assign n3538 = ( ~n197 & n3532 ) | ( ~n197 & n3537 ) | ( n3532 & n3537 ) ;
  assign n3539 = ( n197 & ~n3331 ) | ( n197 & n3362 ) | ( ~n3331 & n3362 ) ;
  assign n3540 = n197 & ~n3331 ;
  assign n3541 = ( n3336 & n3539 ) | ( n3336 & n3540 ) | ( n3539 & n3540 ) ;
  assign n3542 = ( ~n3336 & n3539 ) | ( ~n3336 & n3540 ) | ( n3539 & n3540 ) ;
  assign n3543 = ( n3336 & ~n3541 ) | ( n3336 & n3542 ) | ( ~n3541 & n3542 ) ;
  assign n3544 = ( ~n170 & n3538 ) | ( ~n170 & n3543 ) | ( n3538 & n3543 ) ;
  assign n3545 = n170 & ~n3337 ;
  assign n3546 = ( n170 & ~n3337 ) | ( n170 & n3362 ) | ( ~n3337 & n3362 ) ;
  assign n3547 = ( n3342 & n3545 ) | ( n3342 & n3546 ) | ( n3545 & n3546 ) ;
  assign n3548 = ( ~n3342 & n3545 ) | ( ~n3342 & n3546 ) | ( n3545 & n3546 ) ;
  assign n3549 = ( n3342 & ~n3547 ) | ( n3342 & n3548 ) | ( ~n3547 & n3548 ) ;
  assign n3550 = ( ~n142 & n3544 ) | ( ~n142 & n3549 ) | ( n3544 & n3549 ) ;
  assign n3551 = ( n142 & ~n3343 ) | ( n142 & n3362 ) | ( ~n3343 & n3362 ) ;
  assign n3552 = n142 & ~n3343 ;
  assign n3553 = ( n3348 & n3551 ) | ( n3348 & n3552 ) | ( n3551 & n3552 ) ;
  assign n3554 = ( ~n3348 & n3551 ) | ( ~n3348 & n3552 ) | ( n3551 & n3552 ) ;
  assign n3555 = ( n3348 & ~n3553 ) | ( n3348 & n3554 ) | ( ~n3553 & n3554 ) ;
  assign n3556 = ( ~n132 & n3550 ) | ( ~n132 & n3555 ) | ( n3550 & n3555 ) ;
  assign n3557 = ( n132 & ~n3349 ) | ( n132 & n3362 ) | ( ~n3349 & n3362 ) ;
  assign n3558 = n132 & ~n3349 ;
  assign n3559 = ( n3354 & n3557 ) | ( n3354 & n3558 ) | ( n3557 & n3558 ) ;
  assign n3560 = ( ~n3354 & n3557 ) | ( ~n3354 & n3558 ) | ( n3557 & n3558 ) ;
  assign n3561 = ( n3354 & ~n3559 ) | ( n3354 & n3560 ) | ( ~n3559 & n3560 ) ;
  assign n3562 = n131 & n3369 ;
  assign n3563 = ( ~n3355 & n3360 ) | ( ~n3355 & n3362 ) | ( n3360 & n3362 ) ;
  assign n3564 = ( ~n3363 & n3562 ) | ( ~n3363 & n3563 ) | ( n3562 & n3563 ) ;
  assign n3565 = ~n3556 & n3564 ;
  assign n3566 = n3561 | n3565 ;
  assign n3567 = ( ~n3370 & n3556 ) | ( ~n3370 & n3566 ) | ( n3556 & n3566 ) ;
  assign n3568 = n3556 | n3561 ;
  assign n3569 = ~n3561 & n3562 ;
  assign n3570 = n3556 & ~n3569 ;
  assign n3571 = ( n131 & ~n3568 ) | ( n131 & n3570 ) | ( ~n3568 & n3570 ) ;
  assign n3572 = n3362 & ~n3567 ;
  assign n3573 = ~n3371 & n3567 ;
  assign n3574 = ( x62 & n3572 ) | ( x62 & n3573 ) | ( n3572 & n3573 ) ;
  assign n3575 = ( ~x62 & n3572 ) | ( ~x62 & n3573 ) | ( n3572 & n3573 ) ;
  assign n3576 = ( x62 & ~n3574 ) | ( x62 & n3575 ) | ( ~n3574 & n3575 ) ;
  assign n3577 = x58 | x59 ;
  assign n3578 = x60 | n3577 ;
  assign n3579 = n3362 & ~n3578 ;
  assign n3580 = ~n3362 & n3578 ;
  assign n3581 = ( x61 & ~n3567 ) | ( x61 & n3580 ) | ( ~n3567 & n3580 ) ;
  assign n3582 = ( n3573 & ~n3579 ) | ( n3573 & n3581 ) | ( ~n3579 & n3581 ) ;
  assign n3583 = ( ~n3169 & n3576 ) | ( ~n3169 & n3582 ) | ( n3576 & n3582 ) ;
  assign n3584 = ~n3169 & n3362 ;
  assign n3585 = ( n3378 & n3567 ) | ( n3378 & n3584 ) | ( n3567 & n3584 ) ;
  assign n3586 = ( x63 & n3575 ) | ( x63 & n3585 ) | ( n3575 & n3585 ) ;
  assign n3587 = ( ~x63 & n3575 ) | ( ~x63 & n3585 ) | ( n3575 & n3585 ) ;
  assign n3588 = ( x63 & ~n3586 ) | ( x63 & n3587 ) | ( ~n3586 & n3587 ) ;
  assign n3589 = ( ~n2979 & n3583 ) | ( ~n2979 & n3588 ) | ( n3583 & n3588 ) ;
  assign n3590 = n2979 & ~n3377 ;
  assign n3591 = ( n2979 & ~n3377 ) | ( n2979 & n3567 ) | ( ~n3377 & n3567 ) ;
  assign n3592 = ( ~n3381 & n3590 ) | ( ~n3381 & n3591 ) | ( n3590 & n3591 ) ;
  assign n3593 = ( n3381 & n3590 ) | ( n3381 & n3591 ) | ( n3590 & n3591 ) ;
  assign n3594 = ( n3381 & n3592 ) | ( n3381 & ~n3593 ) | ( n3592 & ~n3593 ) ;
  assign n3595 = ( ~n2791 & n3589 ) | ( ~n2791 & n3594 ) | ( n3589 & n3594 ) ;
  assign n3596 = n2791 & ~n3382 ;
  assign n3597 = ( n2791 & ~n3382 ) | ( n2791 & n3567 ) | ( ~n3382 & n3567 ) ;
  assign n3598 = ( n3387 & n3596 ) | ( n3387 & n3597 ) | ( n3596 & n3597 ) ;
  assign n3599 = ( ~n3387 & n3596 ) | ( ~n3387 & n3597 ) | ( n3596 & n3597 ) ;
  assign n3600 = ( n3387 & ~n3598 ) | ( n3387 & n3599 ) | ( ~n3598 & n3599 ) ;
  assign n3601 = ( ~n2615 & n3595 ) | ( ~n2615 & n3600 ) | ( n3595 & n3600 ) ;
  assign n3602 = n2615 & ~n3388 ;
  assign n3603 = ( n2615 & ~n3388 ) | ( n2615 & n3567 ) | ( ~n3388 & n3567 ) ;
  assign n3604 = ( n3393 & n3602 ) | ( n3393 & n3603 ) | ( n3602 & n3603 ) ;
  assign n3605 = ( ~n3393 & n3602 ) | ( ~n3393 & n3603 ) | ( n3602 & n3603 ) ;
  assign n3606 = ( n3393 & ~n3604 ) | ( n3393 & n3605 ) | ( ~n3604 & n3605 ) ;
  assign n3607 = ( ~n2443 & n3601 ) | ( ~n2443 & n3606 ) | ( n3601 & n3606 ) ;
  assign n3608 = ~n2443 & n3394 ;
  assign n3609 = ( ~n2443 & n3394 ) | ( ~n2443 & n3567 ) | ( n3394 & n3567 ) ;
  assign n3610 = ( ~n3399 & n3608 ) | ( ~n3399 & n3609 ) | ( n3608 & n3609 ) ;
  assign n3611 = ( n3399 & n3608 ) | ( n3399 & n3609 ) | ( n3608 & n3609 ) ;
  assign n3612 = ( n3399 & n3610 ) | ( n3399 & ~n3611 ) | ( n3610 & ~n3611 ) ;
  assign n3613 = ( ~n2277 & n3607 ) | ( ~n2277 & n3612 ) | ( n3607 & n3612 ) ;
  assign n3614 = n2277 & ~n3400 ;
  assign n3615 = ( n2277 & ~n3400 ) | ( n2277 & n3567 ) | ( ~n3400 & n3567 ) ;
  assign n3616 = ( n3405 & n3614 ) | ( n3405 & n3615 ) | ( n3614 & n3615 ) ;
  assign n3617 = ( ~n3405 & n3614 ) | ( ~n3405 & n3615 ) | ( n3614 & n3615 ) ;
  assign n3618 = ( n3405 & ~n3616 ) | ( n3405 & n3617 ) | ( ~n3616 & n3617 ) ;
  assign n3619 = ( ~n2111 & n3613 ) | ( ~n2111 & n3618 ) | ( n3613 & n3618 ) ;
  assign n3620 = ~n2111 & n3406 ;
  assign n3621 = ( ~n2111 & n3406 ) | ( ~n2111 & n3567 ) | ( n3406 & n3567 ) ;
  assign n3622 = ( n3411 & n3620 ) | ( n3411 & n3621 ) | ( n3620 & n3621 ) ;
  assign n3623 = ( ~n3411 & n3620 ) | ( ~n3411 & n3621 ) | ( n3620 & n3621 ) ;
  assign n3624 = ( n3411 & ~n3622 ) | ( n3411 & n3623 ) | ( ~n3622 & n3623 ) ;
  assign n3625 = ( ~n1949 & n3619 ) | ( ~n1949 & n3624 ) | ( n3619 & n3624 ) ;
  assign n3626 = ( n1949 & ~n3412 ) | ( n1949 & n3567 ) | ( ~n3412 & n3567 ) ;
  assign n3627 = n1949 & ~n3412 ;
  assign n3628 = ( n3417 & n3626 ) | ( n3417 & n3627 ) | ( n3626 & n3627 ) ;
  assign n3629 = ( ~n3417 & n3626 ) | ( ~n3417 & n3627 ) | ( n3626 & n3627 ) ;
  assign n3630 = ( n3417 & ~n3628 ) | ( n3417 & n3629 ) | ( ~n3628 & n3629 ) ;
  assign n3631 = ( ~n1802 & n3625 ) | ( ~n1802 & n3630 ) | ( n3625 & n3630 ) ;
  assign n3632 = ( n1802 & ~n3418 ) | ( n1802 & n3567 ) | ( ~n3418 & n3567 ) ;
  assign n3633 = n1802 & ~n3418 ;
  assign n3634 = ( n3423 & n3632 ) | ( n3423 & n3633 ) | ( n3632 & n3633 ) ;
  assign n3635 = ( ~n3423 & n3632 ) | ( ~n3423 & n3633 ) | ( n3632 & n3633 ) ;
  assign n3636 = ( n3423 & ~n3634 ) | ( n3423 & n3635 ) | ( ~n3634 & n3635 ) ;
  assign n3637 = ( ~n1661 & n3631 ) | ( ~n1661 & n3636 ) | ( n3631 & n3636 ) ;
  assign n3638 = ( n1661 & ~n3424 ) | ( n1661 & n3567 ) | ( ~n3424 & n3567 ) ;
  assign n3639 = n1661 & ~n3424 ;
  assign n3640 = ( n3429 & n3638 ) | ( n3429 & n3639 ) | ( n3638 & n3639 ) ;
  assign n3641 = ( ~n3429 & n3638 ) | ( ~n3429 & n3639 ) | ( n3638 & n3639 ) ;
  assign n3642 = ( n3429 & ~n3640 ) | ( n3429 & n3641 ) | ( ~n3640 & n3641 ) ;
  assign n3643 = ( ~n1523 & n3637 ) | ( ~n1523 & n3642 ) | ( n3637 & n3642 ) ;
  assign n3644 = n1523 & ~n3430 ;
  assign n3645 = ( n1523 & ~n3430 ) | ( n1523 & n3567 ) | ( ~n3430 & n3567 ) ;
  assign n3646 = ( n3435 & n3644 ) | ( n3435 & n3645 ) | ( n3644 & n3645 ) ;
  assign n3647 = ( ~n3435 & n3644 ) | ( ~n3435 & n3645 ) | ( n3644 & n3645 ) ;
  assign n3648 = ( n3435 & ~n3646 ) | ( n3435 & n3647 ) | ( ~n3646 & n3647 ) ;
  assign n3649 = ( ~n1393 & n3643 ) | ( ~n1393 & n3648 ) | ( n3643 & n3648 ) ;
  assign n3650 = ( n1393 & ~n3436 ) | ( n1393 & n3567 ) | ( ~n3436 & n3567 ) ;
  assign n3651 = n1393 & ~n3436 ;
  assign n3652 = ( n3441 & n3650 ) | ( n3441 & n3651 ) | ( n3650 & n3651 ) ;
  assign n3653 = ( ~n3441 & n3650 ) | ( ~n3441 & n3651 ) | ( n3650 & n3651 ) ;
  assign n3654 = ( n3441 & ~n3652 ) | ( n3441 & n3653 ) | ( ~n3652 & n3653 ) ;
  assign n3655 = ( ~n1266 & n3649 ) | ( ~n1266 & n3654 ) | ( n3649 & n3654 ) ;
  assign n3656 = ( n1266 & ~n3442 ) | ( n1266 & n3567 ) | ( ~n3442 & n3567 ) ;
  assign n3657 = n1266 & ~n3442 ;
  assign n3658 = ( n3447 & n3656 ) | ( n3447 & n3657 ) | ( n3656 & n3657 ) ;
  assign n3659 = ( ~n3447 & n3656 ) | ( ~n3447 & n3657 ) | ( n3656 & n3657 ) ;
  assign n3660 = ( n3447 & ~n3658 ) | ( n3447 & n3659 ) | ( ~n3658 & n3659 ) ;
  assign n3661 = ( ~n1150 & n3655 ) | ( ~n1150 & n3660 ) | ( n3655 & n3660 ) ;
  assign n3662 = ( n1150 & ~n3448 ) | ( n1150 & n3567 ) | ( ~n3448 & n3567 ) ;
  assign n3663 = n1150 & ~n3448 ;
  assign n3664 = ( n3453 & n3662 ) | ( n3453 & n3663 ) | ( n3662 & n3663 ) ;
  assign n3665 = ( ~n3453 & n3662 ) | ( ~n3453 & n3663 ) | ( n3662 & n3663 ) ;
  assign n3666 = ( n3453 & ~n3664 ) | ( n3453 & n3665 ) | ( ~n3664 & n3665 ) ;
  assign n3667 = ( ~n1038 & n3661 ) | ( ~n1038 & n3666 ) | ( n3661 & n3666 ) ;
  assign n3668 = ~n1038 & n3454 ;
  assign n3669 = ( ~n1038 & n3454 ) | ( ~n1038 & n3567 ) | ( n3454 & n3567 ) ;
  assign n3670 = ( ~n3459 & n3668 ) | ( ~n3459 & n3669 ) | ( n3668 & n3669 ) ;
  assign n3671 = ( n3459 & n3668 ) | ( n3459 & n3669 ) | ( n3668 & n3669 ) ;
  assign n3672 = ( n3459 & n3670 ) | ( n3459 & ~n3671 ) | ( n3670 & ~n3671 ) ;
  assign n3673 = ( ~n933 & n3667 ) | ( ~n933 & n3672 ) | ( n3667 & n3672 ) ;
  assign n3674 = n933 & ~n3460 ;
  assign n3675 = ( n933 & ~n3460 ) | ( n933 & n3567 ) | ( ~n3460 & n3567 ) ;
  assign n3676 = ( ~n3465 & n3674 ) | ( ~n3465 & n3675 ) | ( n3674 & n3675 ) ;
  assign n3677 = ( n3465 & n3674 ) | ( n3465 & n3675 ) | ( n3674 & n3675 ) ;
  assign n3678 = ( n3465 & n3676 ) | ( n3465 & ~n3677 ) | ( n3676 & ~n3677 ) ;
  assign n3679 = ( ~n839 & n3673 ) | ( ~n839 & n3678 ) | ( n3673 & n3678 ) ;
  assign n3680 = ( n839 & ~n3466 ) | ( n839 & n3567 ) | ( ~n3466 & n3567 ) ;
  assign n3681 = n839 & ~n3466 ;
  assign n3682 = ( n3471 & n3680 ) | ( n3471 & n3681 ) | ( n3680 & n3681 ) ;
  assign n3683 = ( ~n3471 & n3680 ) | ( ~n3471 & n3681 ) | ( n3680 & n3681 ) ;
  assign n3684 = ( n3471 & ~n3682 ) | ( n3471 & n3683 ) | ( ~n3682 & n3683 ) ;
  assign n3685 = ( ~n746 & n3679 ) | ( ~n746 & n3684 ) | ( n3679 & n3684 ) ;
  assign n3686 = ( n746 & ~n3472 ) | ( n746 & n3567 ) | ( ~n3472 & n3567 ) ;
  assign n3687 = n746 & ~n3472 ;
  assign n3688 = ( n3477 & n3686 ) | ( n3477 & n3687 ) | ( n3686 & n3687 ) ;
  assign n3689 = ( ~n3477 & n3686 ) | ( ~n3477 & n3687 ) | ( n3686 & n3687 ) ;
  assign n3690 = ( n3477 & ~n3688 ) | ( n3477 & n3689 ) | ( ~n3688 & n3689 ) ;
  assign n3691 = ( ~n664 & n3685 ) | ( ~n664 & n3690 ) | ( n3685 & n3690 ) ;
  assign n3692 = ( n664 & ~n3478 ) | ( n664 & n3567 ) | ( ~n3478 & n3567 ) ;
  assign n3693 = n664 & ~n3478 ;
  assign n3694 = ( n3483 & n3692 ) | ( n3483 & n3693 ) | ( n3692 & n3693 ) ;
  assign n3695 = ( ~n3483 & n3692 ) | ( ~n3483 & n3693 ) | ( n3692 & n3693 ) ;
  assign n3696 = ( n3483 & ~n3694 ) | ( n3483 & n3695 ) | ( ~n3694 & n3695 ) ;
  assign n3697 = ( ~n588 & n3691 ) | ( ~n588 & n3696 ) | ( n3691 & n3696 ) ;
  assign n3698 = ( n588 & ~n3484 ) | ( n588 & n3567 ) | ( ~n3484 & n3567 ) ;
  assign n3699 = n588 & ~n3484 ;
  assign n3700 = ( n3489 & n3698 ) | ( n3489 & n3699 ) | ( n3698 & n3699 ) ;
  assign n3701 = ( ~n3489 & n3698 ) | ( ~n3489 & n3699 ) | ( n3698 & n3699 ) ;
  assign n3702 = ( n3489 & ~n3700 ) | ( n3489 & n3701 ) | ( ~n3700 & n3701 ) ;
  assign n3703 = ( ~n518 & n3697 ) | ( ~n518 & n3702 ) | ( n3697 & n3702 ) ;
  assign n3704 = ( n518 & ~n3490 ) | ( n518 & n3567 ) | ( ~n3490 & n3567 ) ;
  assign n3705 = n518 & ~n3490 ;
  assign n3706 = ( n3495 & n3704 ) | ( n3495 & n3705 ) | ( n3704 & n3705 ) ;
  assign n3707 = ( ~n3495 & n3704 ) | ( ~n3495 & n3705 ) | ( n3704 & n3705 ) ;
  assign n3708 = ( n3495 & ~n3706 ) | ( n3495 & n3707 ) | ( ~n3706 & n3707 ) ;
  assign n3709 = ( ~n454 & n3703 ) | ( ~n454 & n3708 ) | ( n3703 & n3708 ) ;
  assign n3710 = n454 & ~n3496 ;
  assign n3711 = ( n454 & ~n3496 ) | ( n454 & n3567 ) | ( ~n3496 & n3567 ) ;
  assign n3712 = ( ~n3501 & n3710 ) | ( ~n3501 & n3711 ) | ( n3710 & n3711 ) ;
  assign n3713 = ( n3501 & n3710 ) | ( n3501 & n3711 ) | ( n3710 & n3711 ) ;
  assign n3714 = ( n3501 & n3712 ) | ( n3501 & ~n3713 ) | ( n3712 & ~n3713 ) ;
  assign n3715 = ( ~n396 & n3709 ) | ( ~n396 & n3714 ) | ( n3709 & n3714 ) ;
  assign n3716 = ( n396 & ~n3502 ) | ( n396 & n3567 ) | ( ~n3502 & n3567 ) ;
  assign n3717 = n396 & ~n3502 ;
  assign n3718 = ( n3507 & n3716 ) | ( n3507 & n3717 ) | ( n3716 & n3717 ) ;
  assign n3719 = ( ~n3507 & n3716 ) | ( ~n3507 & n3717 ) | ( n3716 & n3717 ) ;
  assign n3720 = ( n3507 & ~n3718 ) | ( n3507 & n3719 ) | ( ~n3718 & n3719 ) ;
  assign n3721 = ( ~n344 & n3715 ) | ( ~n344 & n3720 ) | ( n3715 & n3720 ) ;
  assign n3722 = ~n344 & n3508 ;
  assign n3723 = ( ~n344 & n3508 ) | ( ~n344 & n3567 ) | ( n3508 & n3567 ) ;
  assign n3724 = ( ~n3513 & n3722 ) | ( ~n3513 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3725 = ( n3513 & n3722 ) | ( n3513 & n3723 ) | ( n3722 & n3723 ) ;
  assign n3726 = ( n3513 & n3724 ) | ( n3513 & ~n3725 ) | ( n3724 & ~n3725 ) ;
  assign n3727 = ( ~n298 & n3721 ) | ( ~n298 & n3726 ) | ( n3721 & n3726 ) ;
  assign n3728 = ~n298 & n3514 ;
  assign n3729 = ( ~n298 & n3514 ) | ( ~n298 & n3567 ) | ( n3514 & n3567 ) ;
  assign n3730 = ( ~n3519 & n3728 ) | ( ~n3519 & n3729 ) | ( n3728 & n3729 ) ;
  assign n3731 = ( n3519 & n3728 ) | ( n3519 & n3729 ) | ( n3728 & n3729 ) ;
  assign n3732 = ( n3519 & n3730 ) | ( n3519 & ~n3731 ) | ( n3730 & ~n3731 ) ;
  assign n3733 = ( ~n258 & n3727 ) | ( ~n258 & n3732 ) | ( n3727 & n3732 ) ;
  assign n3734 = ~n258 & n3520 ;
  assign n3735 = ( ~n258 & n3520 ) | ( ~n258 & n3567 ) | ( n3520 & n3567 ) ;
  assign n3736 = ( ~n3525 & n3734 ) | ( ~n3525 & n3735 ) | ( n3734 & n3735 ) ;
  assign n3737 = ( n3525 & n3734 ) | ( n3525 & n3735 ) | ( n3734 & n3735 ) ;
  assign n3738 = ( n3525 & n3736 ) | ( n3525 & ~n3737 ) | ( n3736 & ~n3737 ) ;
  assign n3739 = ( ~n225 & n3733 ) | ( ~n225 & n3738 ) | ( n3733 & n3738 ) ;
  assign n3740 = ~n225 & n3526 ;
  assign n3741 = ( ~n225 & n3526 ) | ( ~n225 & n3567 ) | ( n3526 & n3567 ) ;
  assign n3742 = ( n3531 & n3740 ) | ( n3531 & n3741 ) | ( n3740 & n3741 ) ;
  assign n3743 = ( ~n3531 & n3740 ) | ( ~n3531 & n3741 ) | ( n3740 & n3741 ) ;
  assign n3744 = ( n3531 & ~n3742 ) | ( n3531 & n3743 ) | ( ~n3742 & n3743 ) ;
  assign n3745 = ( ~n197 & n3739 ) | ( ~n197 & n3744 ) | ( n3739 & n3744 ) ;
  assign n3746 = n197 & ~n3532 ;
  assign n3747 = ( n197 & ~n3532 ) | ( n197 & n3567 ) | ( ~n3532 & n3567 ) ;
  assign n3748 = ( n3537 & n3746 ) | ( n3537 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3749 = ( ~n3537 & n3746 ) | ( ~n3537 & n3747 ) | ( n3746 & n3747 ) ;
  assign n3750 = ( n3537 & ~n3748 ) | ( n3537 & n3749 ) | ( ~n3748 & n3749 ) ;
  assign n3751 = ( ~n170 & n3745 ) | ( ~n170 & n3750 ) | ( n3745 & n3750 ) ;
  assign n3752 = n170 & ~n3538 ;
  assign n3753 = ( n170 & ~n3538 ) | ( n170 & n3567 ) | ( ~n3538 & n3567 ) ;
  assign n3754 = ( n3543 & n3752 ) | ( n3543 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3755 = ( ~n3543 & n3752 ) | ( ~n3543 & n3753 ) | ( n3752 & n3753 ) ;
  assign n3756 = ( n3543 & ~n3754 ) | ( n3543 & n3755 ) | ( ~n3754 & n3755 ) ;
  assign n3757 = ( ~n142 & n3751 ) | ( ~n142 & n3756 ) | ( n3751 & n3756 ) ;
  assign n3758 = ~n142 & n3544 ;
  assign n3759 = ( ~n142 & n3544 ) | ( ~n142 & n3567 ) | ( n3544 & n3567 ) ;
  assign n3760 = ( n3549 & n3758 ) | ( n3549 & n3759 ) | ( n3758 & n3759 ) ;
  assign n3761 = ( ~n3549 & n3758 ) | ( ~n3549 & n3759 ) | ( n3758 & n3759 ) ;
  assign n3762 = ( n3549 & ~n3760 ) | ( n3549 & n3761 ) | ( ~n3760 & n3761 ) ;
  assign n3763 = ( ~n132 & n3757 ) | ( ~n132 & n3762 ) | ( n3757 & n3762 ) ;
  assign n3764 = ( n132 & ~n3550 ) | ( n132 & n3567 ) | ( ~n3550 & n3567 ) ;
  assign n3765 = n132 & ~n3550 ;
  assign n3766 = ( n3555 & n3764 ) | ( n3555 & n3765 ) | ( n3764 & n3765 ) ;
  assign n3767 = ( ~n3555 & n3764 ) | ( ~n3555 & n3765 ) | ( n3764 & n3765 ) ;
  assign n3768 = ( n3555 & ~n3766 ) | ( n3555 & n3767 ) | ( ~n3766 & n3767 ) ;
  assign n3769 = ~n3556 & n3561 ;
  assign n3770 = ( n131 & n3566 ) | ( n131 & ~n3769 ) | ( n3566 & ~n3769 ) ;
  assign n3771 = ( ~n3571 & n3768 ) | ( ~n3571 & n3770 ) | ( n3768 & n3770 ) ;
  assign n3772 = ( ~n3571 & n3763 ) | ( ~n3571 & n3771 ) | ( n3763 & n3771 ) ;
  assign n3773 = ~n3763 & n3768 ;
  assign n3774 = n3763 & ~n3768 ;
  assign n3775 = ( n3568 & n3570 ) | ( n3568 & n3774 ) | ( n3570 & n3774 ) ;
  assign n3776 = ( ~n3570 & n3773 ) | ( ~n3570 & n3775 ) | ( n3773 & n3775 ) ;
  assign n3777 = n131 & ~n3776 ;
  assign n3778 = x56 | x57 ;
  assign n3779 = x58 | n3778 ;
  assign n3780 = ~n3567 & n3779 ;
  assign n3781 = ( x59 & ~n3772 ) | ( x59 & n3780 ) | ( ~n3772 & n3780 ) ;
  assign n3782 = n3567 & ~n3779 ;
  assign n3783 = ~n3577 & n3772 ;
  assign n3784 = ( n3781 & ~n3782 ) | ( n3781 & n3783 ) | ( ~n3782 & n3783 ) ;
  assign n3785 = n3567 & ~n3772 ;
  assign n3786 = ( x60 & n3783 ) | ( x60 & n3785 ) | ( n3783 & n3785 ) ;
  assign n3787 = ( ~x60 & n3783 ) | ( ~x60 & n3785 ) | ( n3783 & n3785 ) ;
  assign n3788 = ( x60 & ~n3786 ) | ( x60 & n3787 ) | ( ~n3786 & n3787 ) ;
  assign n3789 = ( ~n3362 & n3784 ) | ( ~n3362 & n3788 ) | ( n3784 & n3788 ) ;
  assign n3790 = ~n3362 & n3567 ;
  assign n3791 = ( n3572 & n3772 ) | ( n3572 & n3790 ) | ( n3772 & n3790 ) ;
  assign n3792 = ( ~x61 & n3787 ) | ( ~x61 & n3791 ) | ( n3787 & n3791 ) ;
  assign n3793 = ( x61 & n3787 ) | ( x61 & n3791 ) | ( n3787 & n3791 ) ;
  assign n3794 = ( x61 & n3792 ) | ( x61 & ~n3793 ) | ( n3792 & ~n3793 ) ;
  assign n3795 = ( ~n3169 & n3789 ) | ( ~n3169 & n3794 ) | ( n3789 & n3794 ) ;
  assign n3796 = n3169 & ~n3582 ;
  assign n3797 = ( n3169 & ~n3582 ) | ( n3169 & n3772 ) | ( ~n3582 & n3772 ) ;
  assign n3798 = ( ~n3576 & n3796 ) | ( ~n3576 & n3797 ) | ( n3796 & n3797 ) ;
  assign n3799 = ( n3576 & n3796 ) | ( n3576 & n3797 ) | ( n3796 & n3797 ) ;
  assign n3800 = ( n3576 & n3798 ) | ( n3576 & ~n3799 ) | ( n3798 & ~n3799 ) ;
  assign n3801 = ( ~n2979 & n3795 ) | ( ~n2979 & n3800 ) | ( n3795 & n3800 ) ;
  assign n3802 = ( n2979 & ~n3583 ) | ( n2979 & n3772 ) | ( ~n3583 & n3772 ) ;
  assign n3803 = n2979 & ~n3583 ;
  assign n3804 = ( n3588 & n3802 ) | ( n3588 & n3803 ) | ( n3802 & n3803 ) ;
  assign n3805 = ( ~n3588 & n3802 ) | ( ~n3588 & n3803 ) | ( n3802 & n3803 ) ;
  assign n3806 = ( n3588 & ~n3804 ) | ( n3588 & n3805 ) | ( ~n3804 & n3805 ) ;
  assign n3807 = ( ~n2791 & n3801 ) | ( ~n2791 & n3806 ) | ( n3801 & n3806 ) ;
  assign n3808 = ~n2791 & n3589 ;
  assign n3809 = ( ~n2791 & n3589 ) | ( ~n2791 & n3772 ) | ( n3589 & n3772 ) ;
  assign n3810 = ( ~n3594 & n3808 ) | ( ~n3594 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3811 = ( n3594 & n3808 ) | ( n3594 & n3809 ) | ( n3808 & n3809 ) ;
  assign n3812 = ( n3594 & n3810 ) | ( n3594 & ~n3811 ) | ( n3810 & ~n3811 ) ;
  assign n3813 = ( ~n2615 & n3807 ) | ( ~n2615 & n3812 ) | ( n3807 & n3812 ) ;
  assign n3814 = ~n2615 & n3595 ;
  assign n3815 = ( ~n2615 & n3595 ) | ( ~n2615 & n3772 ) | ( n3595 & n3772 ) ;
  assign n3816 = ( n3600 & n3814 ) | ( n3600 & n3815 ) | ( n3814 & n3815 ) ;
  assign n3817 = ( ~n3600 & n3814 ) | ( ~n3600 & n3815 ) | ( n3814 & n3815 ) ;
  assign n3818 = ( n3600 & ~n3816 ) | ( n3600 & n3817 ) | ( ~n3816 & n3817 ) ;
  assign n3819 = ( ~n2443 & n3813 ) | ( ~n2443 & n3818 ) | ( n3813 & n3818 ) ;
  assign n3820 = ( n2443 & ~n3601 ) | ( n2443 & n3772 ) | ( ~n3601 & n3772 ) ;
  assign n3821 = n2443 & ~n3601 ;
  assign n3822 = ( n3606 & n3820 ) | ( n3606 & n3821 ) | ( n3820 & n3821 ) ;
  assign n3823 = ( ~n3606 & n3820 ) | ( ~n3606 & n3821 ) | ( n3820 & n3821 ) ;
  assign n3824 = ( n3606 & ~n3822 ) | ( n3606 & n3823 ) | ( ~n3822 & n3823 ) ;
  assign n3825 = ( ~n2277 & n3819 ) | ( ~n2277 & n3824 ) | ( n3819 & n3824 ) ;
  assign n3826 = ~n2277 & n3607 ;
  assign n3827 = ( ~n2277 & n3607 ) | ( ~n2277 & n3772 ) | ( n3607 & n3772 ) ;
  assign n3828 = ( ~n3612 & n3826 ) | ( ~n3612 & n3827 ) | ( n3826 & n3827 ) ;
  assign n3829 = ( n3612 & n3826 ) | ( n3612 & n3827 ) | ( n3826 & n3827 ) ;
  assign n3830 = ( n3612 & n3828 ) | ( n3612 & ~n3829 ) | ( n3828 & ~n3829 ) ;
  assign n3831 = ( ~n2111 & n3825 ) | ( ~n2111 & n3830 ) | ( n3825 & n3830 ) ;
  assign n3832 = ~n2111 & n3613 ;
  assign n3833 = ( ~n2111 & n3613 ) | ( ~n2111 & n3772 ) | ( n3613 & n3772 ) ;
  assign n3834 = ( ~n3618 & n3832 ) | ( ~n3618 & n3833 ) | ( n3832 & n3833 ) ;
  assign n3835 = ( n3618 & n3832 ) | ( n3618 & n3833 ) | ( n3832 & n3833 ) ;
  assign n3836 = ( n3618 & n3834 ) | ( n3618 & ~n3835 ) | ( n3834 & ~n3835 ) ;
  assign n3837 = ( ~n1949 & n3831 ) | ( ~n1949 & n3836 ) | ( n3831 & n3836 ) ;
  assign n3838 = ( n1949 & ~n3619 ) | ( n1949 & n3772 ) | ( ~n3619 & n3772 ) ;
  assign n3839 = n1949 & ~n3619 ;
  assign n3840 = ( n3624 & n3838 ) | ( n3624 & n3839 ) | ( n3838 & n3839 ) ;
  assign n3841 = ( ~n3624 & n3838 ) | ( ~n3624 & n3839 ) | ( n3838 & n3839 ) ;
  assign n3842 = ( n3624 & ~n3840 ) | ( n3624 & n3841 ) | ( ~n3840 & n3841 ) ;
  assign n3843 = ( ~n1802 & n3837 ) | ( ~n1802 & n3842 ) | ( n3837 & n3842 ) ;
  assign n3844 = ~n1802 & n3625 ;
  assign n3845 = ( ~n1802 & n3625 ) | ( ~n1802 & n3772 ) | ( n3625 & n3772 ) ;
  assign n3846 = ( n3630 & n3844 ) | ( n3630 & n3845 ) | ( n3844 & n3845 ) ;
  assign n3847 = ( ~n3630 & n3844 ) | ( ~n3630 & n3845 ) | ( n3844 & n3845 ) ;
  assign n3848 = ( n3630 & ~n3846 ) | ( n3630 & n3847 ) | ( ~n3846 & n3847 ) ;
  assign n3849 = ( ~n1661 & n3843 ) | ( ~n1661 & n3848 ) | ( n3843 & n3848 ) ;
  assign n3850 = ~n1661 & n3631 ;
  assign n3851 = ( ~n1661 & n3631 ) | ( ~n1661 & n3772 ) | ( n3631 & n3772 ) ;
  assign n3852 = ( ~n3636 & n3850 ) | ( ~n3636 & n3851 ) | ( n3850 & n3851 ) ;
  assign n3853 = ( n3636 & n3850 ) | ( n3636 & n3851 ) | ( n3850 & n3851 ) ;
  assign n3854 = ( n3636 & n3852 ) | ( n3636 & ~n3853 ) | ( n3852 & ~n3853 ) ;
  assign n3855 = ( ~n1523 & n3849 ) | ( ~n1523 & n3854 ) | ( n3849 & n3854 ) ;
  assign n3856 = ~n1523 & n3637 ;
  assign n3857 = ( ~n1523 & n3637 ) | ( ~n1523 & n3772 ) | ( n3637 & n3772 ) ;
  assign n3858 = ( ~n3642 & n3856 ) | ( ~n3642 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3859 = ( n3642 & n3856 ) | ( n3642 & n3857 ) | ( n3856 & n3857 ) ;
  assign n3860 = ( n3642 & n3858 ) | ( n3642 & ~n3859 ) | ( n3858 & ~n3859 ) ;
  assign n3861 = ( ~n1393 & n3855 ) | ( ~n1393 & n3860 ) | ( n3855 & n3860 ) ;
  assign n3862 = ( n1393 & ~n3643 ) | ( n1393 & n3772 ) | ( ~n3643 & n3772 ) ;
  assign n3863 = n1393 & ~n3643 ;
  assign n3864 = ( n3648 & n3862 ) | ( n3648 & n3863 ) | ( n3862 & n3863 ) ;
  assign n3865 = ( ~n3648 & n3862 ) | ( ~n3648 & n3863 ) | ( n3862 & n3863 ) ;
  assign n3866 = ( n3648 & ~n3864 ) | ( n3648 & n3865 ) | ( ~n3864 & n3865 ) ;
  assign n3867 = ( ~n1266 & n3861 ) | ( ~n1266 & n3866 ) | ( n3861 & n3866 ) ;
  assign n3868 = ~n1266 & n3649 ;
  assign n3869 = ( ~n1266 & n3649 ) | ( ~n1266 & n3772 ) | ( n3649 & n3772 ) ;
  assign n3870 = ( ~n3654 & n3868 ) | ( ~n3654 & n3869 ) | ( n3868 & n3869 ) ;
  assign n3871 = ( n3654 & n3868 ) | ( n3654 & n3869 ) | ( n3868 & n3869 ) ;
  assign n3872 = ( n3654 & n3870 ) | ( n3654 & ~n3871 ) | ( n3870 & ~n3871 ) ;
  assign n3873 = ( ~n1150 & n3867 ) | ( ~n1150 & n3872 ) | ( n3867 & n3872 ) ;
  assign n3874 = ~n1150 & n3655 ;
  assign n3875 = ( ~n1150 & n3655 ) | ( ~n1150 & n3772 ) | ( n3655 & n3772 ) ;
  assign n3876 = ( ~n3660 & n3874 ) | ( ~n3660 & n3875 ) | ( n3874 & n3875 ) ;
  assign n3877 = ( n3660 & n3874 ) | ( n3660 & n3875 ) | ( n3874 & n3875 ) ;
  assign n3878 = ( n3660 & n3876 ) | ( n3660 & ~n3877 ) | ( n3876 & ~n3877 ) ;
  assign n3879 = ( ~n1038 & n3873 ) | ( ~n1038 & n3878 ) | ( n3873 & n3878 ) ;
  assign n3880 = ( n1038 & ~n3661 ) | ( n1038 & n3772 ) | ( ~n3661 & n3772 ) ;
  assign n3881 = n1038 & ~n3661 ;
  assign n3882 = ( n3666 & n3880 ) | ( n3666 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3883 = ( ~n3666 & n3880 ) | ( ~n3666 & n3881 ) | ( n3880 & n3881 ) ;
  assign n3884 = ( n3666 & ~n3882 ) | ( n3666 & n3883 ) | ( ~n3882 & n3883 ) ;
  assign n3885 = ( ~n933 & n3879 ) | ( ~n933 & n3884 ) | ( n3879 & n3884 ) ;
  assign n3886 = ( n933 & ~n3667 ) | ( n933 & n3772 ) | ( ~n3667 & n3772 ) ;
  assign n3887 = n933 & ~n3667 ;
  assign n3888 = ( n3672 & n3886 ) | ( n3672 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3889 = ( ~n3672 & n3886 ) | ( ~n3672 & n3887 ) | ( n3886 & n3887 ) ;
  assign n3890 = ( n3672 & ~n3888 ) | ( n3672 & n3889 ) | ( ~n3888 & n3889 ) ;
  assign n3891 = ( ~n839 & n3885 ) | ( ~n839 & n3890 ) | ( n3885 & n3890 ) ;
  assign n3892 = ( n839 & ~n3673 ) | ( n839 & n3772 ) | ( ~n3673 & n3772 ) ;
  assign n3893 = n839 & ~n3673 ;
  assign n3894 = ( n3678 & n3892 ) | ( n3678 & n3893 ) | ( n3892 & n3893 ) ;
  assign n3895 = ( ~n3678 & n3892 ) | ( ~n3678 & n3893 ) | ( n3892 & n3893 ) ;
  assign n3896 = ( n3678 & ~n3894 ) | ( n3678 & n3895 ) | ( ~n3894 & n3895 ) ;
  assign n3897 = ( ~n746 & n3891 ) | ( ~n746 & n3896 ) | ( n3891 & n3896 ) ;
  assign n3898 = ( n746 & ~n3679 ) | ( n746 & n3772 ) | ( ~n3679 & n3772 ) ;
  assign n3899 = n746 & ~n3679 ;
  assign n3900 = ( n3684 & n3898 ) | ( n3684 & n3899 ) | ( n3898 & n3899 ) ;
  assign n3901 = ( ~n3684 & n3898 ) | ( ~n3684 & n3899 ) | ( n3898 & n3899 ) ;
  assign n3902 = ( n3684 & ~n3900 ) | ( n3684 & n3901 ) | ( ~n3900 & n3901 ) ;
  assign n3903 = ( ~n664 & n3897 ) | ( ~n664 & n3902 ) | ( n3897 & n3902 ) ;
  assign n3904 = ( n664 & ~n3685 ) | ( n664 & n3772 ) | ( ~n3685 & n3772 ) ;
  assign n3905 = n664 & ~n3685 ;
  assign n3906 = ( n3690 & n3904 ) | ( n3690 & n3905 ) | ( n3904 & n3905 ) ;
  assign n3907 = ( ~n3690 & n3904 ) | ( ~n3690 & n3905 ) | ( n3904 & n3905 ) ;
  assign n3908 = ( n3690 & ~n3906 ) | ( n3690 & n3907 ) | ( ~n3906 & n3907 ) ;
  assign n3909 = ( ~n588 & n3903 ) | ( ~n588 & n3908 ) | ( n3903 & n3908 ) ;
  assign n3910 = ~n588 & n3691 ;
  assign n3911 = ( ~n588 & n3691 ) | ( ~n588 & n3772 ) | ( n3691 & n3772 ) ;
  assign n3912 = ( ~n3696 & n3910 ) | ( ~n3696 & n3911 ) | ( n3910 & n3911 ) ;
  assign n3913 = ( n3696 & n3910 ) | ( n3696 & n3911 ) | ( n3910 & n3911 ) ;
  assign n3914 = ( n3696 & n3912 ) | ( n3696 & ~n3913 ) | ( n3912 & ~n3913 ) ;
  assign n3915 = ( ~n518 & n3909 ) | ( ~n518 & n3914 ) | ( n3909 & n3914 ) ;
  assign n3916 = ~n518 & n3697 ;
  assign n3917 = ( ~n518 & n3697 ) | ( ~n518 & n3772 ) | ( n3697 & n3772 ) ;
  assign n3918 = ( ~n3702 & n3916 ) | ( ~n3702 & n3917 ) | ( n3916 & n3917 ) ;
  assign n3919 = ( n3702 & n3916 ) | ( n3702 & n3917 ) | ( n3916 & n3917 ) ;
  assign n3920 = ( n3702 & n3918 ) | ( n3702 & ~n3919 ) | ( n3918 & ~n3919 ) ;
  assign n3921 = ( ~n454 & n3915 ) | ( ~n454 & n3920 ) | ( n3915 & n3920 ) ;
  assign n3922 = ~n454 & n3703 ;
  assign n3923 = ( ~n454 & n3703 ) | ( ~n454 & n3772 ) | ( n3703 & n3772 ) ;
  assign n3924 = ( n3708 & n3922 ) | ( n3708 & n3923 ) | ( n3922 & n3923 ) ;
  assign n3925 = ( ~n3708 & n3922 ) | ( ~n3708 & n3923 ) | ( n3922 & n3923 ) ;
  assign n3926 = ( n3708 & ~n3924 ) | ( n3708 & n3925 ) | ( ~n3924 & n3925 ) ;
  assign n3927 = ( ~n396 & n3921 ) | ( ~n396 & n3926 ) | ( n3921 & n3926 ) ;
  assign n3928 = ( n396 & ~n3709 ) | ( n396 & n3772 ) | ( ~n3709 & n3772 ) ;
  assign n3929 = n396 & ~n3709 ;
  assign n3930 = ( n3714 & n3928 ) | ( n3714 & n3929 ) | ( n3928 & n3929 ) ;
  assign n3931 = ( ~n3714 & n3928 ) | ( ~n3714 & n3929 ) | ( n3928 & n3929 ) ;
  assign n3932 = ( n3714 & ~n3930 ) | ( n3714 & n3931 ) | ( ~n3930 & n3931 ) ;
  assign n3933 = ( ~n344 & n3927 ) | ( ~n344 & n3932 ) | ( n3927 & n3932 ) ;
  assign n3934 = ( n344 & ~n3715 ) | ( n344 & n3772 ) | ( ~n3715 & n3772 ) ;
  assign n3935 = n344 & ~n3715 ;
  assign n3936 = ( n3720 & n3934 ) | ( n3720 & n3935 ) | ( n3934 & n3935 ) ;
  assign n3937 = ( ~n3720 & n3934 ) | ( ~n3720 & n3935 ) | ( n3934 & n3935 ) ;
  assign n3938 = ( n3720 & ~n3936 ) | ( n3720 & n3937 ) | ( ~n3936 & n3937 ) ;
  assign n3939 = ( ~n298 & n3933 ) | ( ~n298 & n3938 ) | ( n3933 & n3938 ) ;
  assign n3940 = ( n298 & ~n3721 ) | ( n298 & n3772 ) | ( ~n3721 & n3772 ) ;
  assign n3941 = n298 & ~n3721 ;
  assign n3942 = ( n3726 & n3940 ) | ( n3726 & n3941 ) | ( n3940 & n3941 ) ;
  assign n3943 = ( ~n3726 & n3940 ) | ( ~n3726 & n3941 ) | ( n3940 & n3941 ) ;
  assign n3944 = ( n3726 & ~n3942 ) | ( n3726 & n3943 ) | ( ~n3942 & n3943 ) ;
  assign n3945 = ( ~n258 & n3939 ) | ( ~n258 & n3944 ) | ( n3939 & n3944 ) ;
  assign n3946 = ( n258 & ~n3727 ) | ( n258 & n3772 ) | ( ~n3727 & n3772 ) ;
  assign n3947 = n258 & ~n3727 ;
  assign n3948 = ( n3732 & n3946 ) | ( n3732 & n3947 ) | ( n3946 & n3947 ) ;
  assign n3949 = ( ~n3732 & n3946 ) | ( ~n3732 & n3947 ) | ( n3946 & n3947 ) ;
  assign n3950 = ( n3732 & ~n3948 ) | ( n3732 & n3949 ) | ( ~n3948 & n3949 ) ;
  assign n3951 = ( ~n225 & n3945 ) | ( ~n225 & n3950 ) | ( n3945 & n3950 ) ;
  assign n3952 = ( n225 & ~n3733 ) | ( n225 & n3772 ) | ( ~n3733 & n3772 ) ;
  assign n3953 = n225 & ~n3733 ;
  assign n3954 = ( n3738 & n3952 ) | ( n3738 & n3953 ) | ( n3952 & n3953 ) ;
  assign n3955 = ( ~n3738 & n3952 ) | ( ~n3738 & n3953 ) | ( n3952 & n3953 ) ;
  assign n3956 = ( n3738 & ~n3954 ) | ( n3738 & n3955 ) | ( ~n3954 & n3955 ) ;
  assign n3957 = ( ~n197 & n3951 ) | ( ~n197 & n3956 ) | ( n3951 & n3956 ) ;
  assign n3958 = ( n197 & ~n3739 ) | ( n197 & n3772 ) | ( ~n3739 & n3772 ) ;
  assign n3959 = n197 & ~n3739 ;
  assign n3960 = ( n3744 & n3958 ) | ( n3744 & n3959 ) | ( n3958 & n3959 ) ;
  assign n3961 = ( ~n3744 & n3958 ) | ( ~n3744 & n3959 ) | ( n3958 & n3959 ) ;
  assign n3962 = ( n3744 & ~n3960 ) | ( n3744 & n3961 ) | ( ~n3960 & n3961 ) ;
  assign n3963 = ( ~n170 & n3957 ) | ( ~n170 & n3962 ) | ( n3957 & n3962 ) ;
  assign n3964 = ~n170 & n3745 ;
  assign n3965 = ( ~n170 & n3745 ) | ( ~n170 & n3772 ) | ( n3745 & n3772 ) ;
  assign n3966 = ( ~n3750 & n3964 ) | ( ~n3750 & n3965 ) | ( n3964 & n3965 ) ;
  assign n3967 = ( n3750 & n3964 ) | ( n3750 & n3965 ) | ( n3964 & n3965 ) ;
  assign n3968 = ( n3750 & n3966 ) | ( n3750 & ~n3967 ) | ( n3966 & ~n3967 ) ;
  assign n3969 = ( ~n142 & n3963 ) | ( ~n142 & n3968 ) | ( n3963 & n3968 ) ;
  assign n3970 = ( n142 & ~n3751 ) | ( n142 & n3772 ) | ( ~n3751 & n3772 ) ;
  assign n3971 = n142 & ~n3751 ;
  assign n3972 = ( n3756 & n3970 ) | ( n3756 & n3971 ) | ( n3970 & n3971 ) ;
  assign n3973 = ( ~n3756 & n3970 ) | ( ~n3756 & n3971 ) | ( n3970 & n3971 ) ;
  assign n3974 = ( n3756 & ~n3972 ) | ( n3756 & n3973 ) | ( ~n3972 & n3973 ) ;
  assign n3975 = ( ~n132 & n3969 ) | ( ~n132 & n3974 ) | ( n3969 & n3974 ) ;
  assign n3976 = ( n3763 & ~n3768 ) | ( n3763 & n3771 ) | ( ~n3768 & n3771 ) ;
  assign n3977 = ~n3774 & n3976 ;
  assign n3978 = n131 | n3977 ;
  assign n3979 = ( n132 & ~n3757 ) | ( n132 & n3772 ) | ( ~n3757 & n3772 ) ;
  assign n3980 = n132 & ~n3757 ;
  assign n3981 = ( n3762 & n3979 ) | ( n3762 & n3980 ) | ( n3979 & n3980 ) ;
  assign n3982 = ( ~n3762 & n3979 ) | ( ~n3762 & n3980 ) | ( n3979 & n3980 ) ;
  assign n3983 = ( n3762 & ~n3981 ) | ( n3762 & n3982 ) | ( ~n3981 & n3982 ) ;
  assign n3984 = ( ~n3777 & n3978 ) | ( ~n3777 & n3983 ) | ( n3978 & n3983 ) ;
  assign n3985 = ( ~n3777 & n3975 ) | ( ~n3777 & n3984 ) | ( n3975 & n3984 ) ;
  assign n3986 = ~n3975 & n3977 ;
  assign n3987 = ( ~n131 & n3983 ) | ( ~n131 & n3986 ) | ( n3983 & n3986 ) ;
  assign n3988 = ~n3975 & n3983 ;
  assign n3989 = x54 | x55 ;
  assign n3990 = x56 | n3989 ;
  assign n3991 = n3772 & ~n3990 ;
  assign n3992 = ~n3778 & n3985 ;
  assign n3993 = ~n3772 & n3990 ;
  assign n3994 = ( x57 & ~n3985 ) | ( x57 & n3993 ) | ( ~n3985 & n3993 ) ;
  assign n3995 = ( ~n3991 & n3992 ) | ( ~n3991 & n3994 ) | ( n3992 & n3994 ) ;
  assign n3996 = n3772 & ~n3985 ;
  assign n3997 = ( x58 & n3992 ) | ( x58 & n3996 ) | ( n3992 & n3996 ) ;
  assign n3998 = ( ~x58 & n3992 ) | ( ~x58 & n3996 ) | ( n3992 & n3996 ) ;
  assign n3999 = ( x58 & ~n3997 ) | ( x58 & n3998 ) | ( ~n3997 & n3998 ) ;
  assign n4000 = ( ~n3567 & n3995 ) | ( ~n3567 & n3999 ) | ( n3995 & n3999 ) ;
  assign n4001 = ~n3567 & n3772 ;
  assign n4002 = ( n3785 & n3985 ) | ( n3785 & n4001 ) | ( n3985 & n4001 ) ;
  assign n4003 = ( ~x59 & n3998 ) | ( ~x59 & n4002 ) | ( n3998 & n4002 ) ;
  assign n4004 = ( x59 & n3998 ) | ( x59 & n4002 ) | ( n3998 & n4002 ) ;
  assign n4005 = ( x59 & n4003 ) | ( x59 & ~n4004 ) | ( n4003 & ~n4004 ) ;
  assign n4006 = ( ~n3362 & n4000 ) | ( ~n3362 & n4005 ) | ( n4000 & n4005 ) ;
  assign n4007 = n3362 & ~n3784 ;
  assign n4008 = ( n3362 & ~n3784 ) | ( n3362 & n3985 ) | ( ~n3784 & n3985 ) ;
  assign n4009 = ( n3788 & n4007 ) | ( n3788 & n4008 ) | ( n4007 & n4008 ) ;
  assign n4010 = ( ~n3788 & n4007 ) | ( ~n3788 & n4008 ) | ( n4007 & n4008 ) ;
  assign n4011 = ( n3788 & ~n4009 ) | ( n3788 & n4010 ) | ( ~n4009 & n4010 ) ;
  assign n4012 = ( ~n3169 & n4006 ) | ( ~n3169 & n4011 ) | ( n4006 & n4011 ) ;
  assign n4013 = ~n3169 & n3789 ;
  assign n4014 = ( ~n3169 & n3789 ) | ( ~n3169 & n3985 ) | ( n3789 & n3985 ) ;
  assign n4015 = ( ~n3794 & n4013 ) | ( ~n3794 & n4014 ) | ( n4013 & n4014 ) ;
  assign n4016 = ( n3794 & n4013 ) | ( n3794 & n4014 ) | ( n4013 & n4014 ) ;
  assign n4017 = ( n3794 & n4015 ) | ( n3794 & ~n4016 ) | ( n4015 & ~n4016 ) ;
  assign n4018 = ( ~n2979 & n4012 ) | ( ~n2979 & n4017 ) | ( n4012 & n4017 ) ;
  assign n4019 = n2979 & ~n3795 ;
  assign n4020 = ( n2979 & ~n3795 ) | ( n2979 & n3985 ) | ( ~n3795 & n3985 ) ;
  assign n4021 = ( n3800 & n4019 ) | ( n3800 & n4020 ) | ( n4019 & n4020 ) ;
  assign n4022 = ( ~n3800 & n4019 ) | ( ~n3800 & n4020 ) | ( n4019 & n4020 ) ;
  assign n4023 = ( n3800 & ~n4021 ) | ( n3800 & n4022 ) | ( ~n4021 & n4022 ) ;
  assign n4024 = ( ~n2791 & n4018 ) | ( ~n2791 & n4023 ) | ( n4018 & n4023 ) ;
  assign n4025 = ~n2791 & n3801 ;
  assign n4026 = ( ~n2791 & n3801 ) | ( ~n2791 & n3985 ) | ( n3801 & n3985 ) ;
  assign n4027 = ( n3806 & n4025 ) | ( n3806 & n4026 ) | ( n4025 & n4026 ) ;
  assign n4028 = ( ~n3806 & n4025 ) | ( ~n3806 & n4026 ) | ( n4025 & n4026 ) ;
  assign n4029 = ( n3806 & ~n4027 ) | ( n3806 & n4028 ) | ( ~n4027 & n4028 ) ;
  assign n4030 = ( ~n2615 & n4024 ) | ( ~n2615 & n4029 ) | ( n4024 & n4029 ) ;
  assign n4031 = ( n2615 & ~n3807 ) | ( n2615 & n3985 ) | ( ~n3807 & n3985 ) ;
  assign n4032 = n2615 & ~n3807 ;
  assign n4033 = ( n3812 & n4031 ) | ( n3812 & n4032 ) | ( n4031 & n4032 ) ;
  assign n4034 = ( ~n3812 & n4031 ) | ( ~n3812 & n4032 ) | ( n4031 & n4032 ) ;
  assign n4035 = ( n3812 & ~n4033 ) | ( n3812 & n4034 ) | ( ~n4033 & n4034 ) ;
  assign n4036 = ( ~n2443 & n4030 ) | ( ~n2443 & n4035 ) | ( n4030 & n4035 ) ;
  assign n4037 = ( n2443 & ~n3813 ) | ( n2443 & n3985 ) | ( ~n3813 & n3985 ) ;
  assign n4038 = n2443 & ~n3813 ;
  assign n4039 = ( n3818 & n4037 ) | ( n3818 & n4038 ) | ( n4037 & n4038 ) ;
  assign n4040 = ( ~n3818 & n4037 ) | ( ~n3818 & n4038 ) | ( n4037 & n4038 ) ;
  assign n4041 = ( n3818 & ~n4039 ) | ( n3818 & n4040 ) | ( ~n4039 & n4040 ) ;
  assign n4042 = ( ~n2277 & n4036 ) | ( ~n2277 & n4041 ) | ( n4036 & n4041 ) ;
  assign n4043 = ~n2277 & n3819 ;
  assign n4044 = ( ~n2277 & n3819 ) | ( ~n2277 & n3985 ) | ( n3819 & n3985 ) ;
  assign n4045 = ( n3824 & n4043 ) | ( n3824 & n4044 ) | ( n4043 & n4044 ) ;
  assign n4046 = ( ~n3824 & n4043 ) | ( ~n3824 & n4044 ) | ( n4043 & n4044 ) ;
  assign n4047 = ( n3824 & ~n4045 ) | ( n3824 & n4046 ) | ( ~n4045 & n4046 ) ;
  assign n4048 = ( ~n2111 & n4042 ) | ( ~n2111 & n4047 ) | ( n4042 & n4047 ) ;
  assign n4049 = ( n2111 & ~n3825 ) | ( n2111 & n3985 ) | ( ~n3825 & n3985 ) ;
  assign n4050 = n2111 & ~n3825 ;
  assign n4051 = ( n3830 & n4049 ) | ( n3830 & n4050 ) | ( n4049 & n4050 ) ;
  assign n4052 = ( ~n3830 & n4049 ) | ( ~n3830 & n4050 ) | ( n4049 & n4050 ) ;
  assign n4053 = ( n3830 & ~n4051 ) | ( n3830 & n4052 ) | ( ~n4051 & n4052 ) ;
  assign n4054 = ( ~n1949 & n4048 ) | ( ~n1949 & n4053 ) | ( n4048 & n4053 ) ;
  assign n4055 = ~n1949 & n3831 ;
  assign n4056 = ( ~n1949 & n3831 ) | ( ~n1949 & n3985 ) | ( n3831 & n3985 ) ;
  assign n4057 = ( ~n3836 & n4055 ) | ( ~n3836 & n4056 ) | ( n4055 & n4056 ) ;
  assign n4058 = ( n3836 & n4055 ) | ( n3836 & n4056 ) | ( n4055 & n4056 ) ;
  assign n4059 = ( n3836 & n4057 ) | ( n3836 & ~n4058 ) | ( n4057 & ~n4058 ) ;
  assign n4060 = ( ~n1802 & n4054 ) | ( ~n1802 & n4059 ) | ( n4054 & n4059 ) ;
  assign n4061 = ( n1802 & ~n3837 ) | ( n1802 & n3985 ) | ( ~n3837 & n3985 ) ;
  assign n4062 = n1802 & ~n3837 ;
  assign n4063 = ( n3842 & n4061 ) | ( n3842 & n4062 ) | ( n4061 & n4062 ) ;
  assign n4064 = ( ~n3842 & n4061 ) | ( ~n3842 & n4062 ) | ( n4061 & n4062 ) ;
  assign n4065 = ( n3842 & ~n4063 ) | ( n3842 & n4064 ) | ( ~n4063 & n4064 ) ;
  assign n4066 = ( ~n1661 & n4060 ) | ( ~n1661 & n4065 ) | ( n4060 & n4065 ) ;
  assign n4067 = ~n1661 & n3843 ;
  assign n4068 = ( ~n1661 & n3843 ) | ( ~n1661 & n3985 ) | ( n3843 & n3985 ) ;
  assign n4069 = ( ~n3848 & n4067 ) | ( ~n3848 & n4068 ) | ( n4067 & n4068 ) ;
  assign n4070 = ( n3848 & n4067 ) | ( n3848 & n4068 ) | ( n4067 & n4068 ) ;
  assign n4071 = ( n3848 & n4069 ) | ( n3848 & ~n4070 ) | ( n4069 & ~n4070 ) ;
  assign n4072 = ( ~n1523 & n4066 ) | ( ~n1523 & n4071 ) | ( n4066 & n4071 ) ;
  assign n4073 = n1523 & ~n3849 ;
  assign n4074 = ( n1523 & ~n3849 ) | ( n1523 & n3985 ) | ( ~n3849 & n3985 ) ;
  assign n4075 = ( ~n3854 & n4073 ) | ( ~n3854 & n4074 ) | ( n4073 & n4074 ) ;
  assign n4076 = ( n3854 & n4073 ) | ( n3854 & n4074 ) | ( n4073 & n4074 ) ;
  assign n4077 = ( n3854 & n4075 ) | ( n3854 & ~n4076 ) | ( n4075 & ~n4076 ) ;
  assign n4078 = ( ~n1393 & n4072 ) | ( ~n1393 & n4077 ) | ( n4072 & n4077 ) ;
  assign n4079 = ( n1393 & ~n3855 ) | ( n1393 & n3985 ) | ( ~n3855 & n3985 ) ;
  assign n4080 = n1393 & ~n3855 ;
  assign n4081 = ( n3860 & n4079 ) | ( n3860 & n4080 ) | ( n4079 & n4080 ) ;
  assign n4082 = ( ~n3860 & n4079 ) | ( ~n3860 & n4080 ) | ( n4079 & n4080 ) ;
  assign n4083 = ( n3860 & ~n4081 ) | ( n3860 & n4082 ) | ( ~n4081 & n4082 ) ;
  assign n4084 = ( ~n1266 & n4078 ) | ( ~n1266 & n4083 ) | ( n4078 & n4083 ) ;
  assign n4085 = ( n1266 & ~n3861 ) | ( n1266 & n3985 ) | ( ~n3861 & n3985 ) ;
  assign n4086 = n1266 & ~n3861 ;
  assign n4087 = ( n3866 & n4085 ) | ( n3866 & n4086 ) | ( n4085 & n4086 ) ;
  assign n4088 = ( ~n3866 & n4085 ) | ( ~n3866 & n4086 ) | ( n4085 & n4086 ) ;
  assign n4089 = ( n3866 & ~n4087 ) | ( n3866 & n4088 ) | ( ~n4087 & n4088 ) ;
  assign n4090 = ( ~n1150 & n4084 ) | ( ~n1150 & n4089 ) | ( n4084 & n4089 ) ;
  assign n4091 = ~n1150 & n3867 ;
  assign n4092 = ( ~n1150 & n3867 ) | ( ~n1150 & n3985 ) | ( n3867 & n3985 ) ;
  assign n4093 = ( ~n3872 & n4091 ) | ( ~n3872 & n4092 ) | ( n4091 & n4092 ) ;
  assign n4094 = ( n3872 & n4091 ) | ( n3872 & n4092 ) | ( n4091 & n4092 ) ;
  assign n4095 = ( n3872 & n4093 ) | ( n3872 & ~n4094 ) | ( n4093 & ~n4094 ) ;
  assign n4096 = ( ~n1038 & n4090 ) | ( ~n1038 & n4095 ) | ( n4090 & n4095 ) ;
  assign n4097 = ~n1038 & n3873 ;
  assign n4098 = ( ~n1038 & n3873 ) | ( ~n1038 & n3985 ) | ( n3873 & n3985 ) ;
  assign n4099 = ( ~n3878 & n4097 ) | ( ~n3878 & n4098 ) | ( n4097 & n4098 ) ;
  assign n4100 = ( n3878 & n4097 ) | ( n3878 & n4098 ) | ( n4097 & n4098 ) ;
  assign n4101 = ( n3878 & n4099 ) | ( n3878 & ~n4100 ) | ( n4099 & ~n4100 ) ;
  assign n4102 = ( ~n933 & n4096 ) | ( ~n933 & n4101 ) | ( n4096 & n4101 ) ;
  assign n4103 = ( n933 & ~n3879 ) | ( n933 & n3985 ) | ( ~n3879 & n3985 ) ;
  assign n4104 = n933 & ~n3879 ;
  assign n4105 = ( n3884 & n4103 ) | ( n3884 & n4104 ) | ( n4103 & n4104 ) ;
  assign n4106 = ( ~n3884 & n4103 ) | ( ~n3884 & n4104 ) | ( n4103 & n4104 ) ;
  assign n4107 = ( n3884 & ~n4105 ) | ( n3884 & n4106 ) | ( ~n4105 & n4106 ) ;
  assign n4108 = ( ~n839 & n4102 ) | ( ~n839 & n4107 ) | ( n4102 & n4107 ) ;
  assign n4109 = ( n839 & ~n3885 ) | ( n839 & n3985 ) | ( ~n3885 & n3985 ) ;
  assign n4110 = n839 & ~n3885 ;
  assign n4111 = ( n3890 & n4109 ) | ( n3890 & n4110 ) | ( n4109 & n4110 ) ;
  assign n4112 = ( ~n3890 & n4109 ) | ( ~n3890 & n4110 ) | ( n4109 & n4110 ) ;
  assign n4113 = ( n3890 & ~n4111 ) | ( n3890 & n4112 ) | ( ~n4111 & n4112 ) ;
  assign n4114 = ( ~n746 & n4108 ) | ( ~n746 & n4113 ) | ( n4108 & n4113 ) ;
  assign n4115 = ~n746 & n3891 ;
  assign n4116 = ( ~n746 & n3891 ) | ( ~n746 & n3985 ) | ( n3891 & n3985 ) ;
  assign n4117 = ( n3896 & n4115 ) | ( n3896 & n4116 ) | ( n4115 & n4116 ) ;
  assign n4118 = ( ~n3896 & n4115 ) | ( ~n3896 & n4116 ) | ( n4115 & n4116 ) ;
  assign n4119 = ( n3896 & ~n4117 ) | ( n3896 & n4118 ) | ( ~n4117 & n4118 ) ;
  assign n4120 = ( ~n664 & n4114 ) | ( ~n664 & n4119 ) | ( n4114 & n4119 ) ;
  assign n4121 = ( n664 & ~n3897 ) | ( n664 & n3985 ) | ( ~n3897 & n3985 ) ;
  assign n4122 = n664 & ~n3897 ;
  assign n4123 = ( n3902 & n4121 ) | ( n3902 & n4122 ) | ( n4121 & n4122 ) ;
  assign n4124 = ( ~n3902 & n4121 ) | ( ~n3902 & n4122 ) | ( n4121 & n4122 ) ;
  assign n4125 = ( n3902 & ~n4123 ) | ( n3902 & n4124 ) | ( ~n4123 & n4124 ) ;
  assign n4126 = ( ~n588 & n4120 ) | ( ~n588 & n4125 ) | ( n4120 & n4125 ) ;
  assign n4127 = n588 & ~n3903 ;
  assign n4128 = ( n588 & ~n3903 ) | ( n588 & n3985 ) | ( ~n3903 & n3985 ) ;
  assign n4129 = ( n3908 & n4127 ) | ( n3908 & n4128 ) | ( n4127 & n4128 ) ;
  assign n4130 = ( ~n3908 & n4127 ) | ( ~n3908 & n4128 ) | ( n4127 & n4128 ) ;
  assign n4131 = ( n3908 & ~n4129 ) | ( n3908 & n4130 ) | ( ~n4129 & n4130 ) ;
  assign n4132 = ( ~n518 & n4126 ) | ( ~n518 & n4131 ) | ( n4126 & n4131 ) ;
  assign n4133 = ( n518 & ~n3909 ) | ( n518 & n3985 ) | ( ~n3909 & n3985 ) ;
  assign n4134 = n518 & ~n3909 ;
  assign n4135 = ( n3914 & n4133 ) | ( n3914 & n4134 ) | ( n4133 & n4134 ) ;
  assign n4136 = ( ~n3914 & n4133 ) | ( ~n3914 & n4134 ) | ( n4133 & n4134 ) ;
  assign n4137 = ( n3914 & ~n4135 ) | ( n3914 & n4136 ) | ( ~n4135 & n4136 ) ;
  assign n4138 = ( ~n454 & n4132 ) | ( ~n454 & n4137 ) | ( n4132 & n4137 ) ;
  assign n4139 = ~n454 & n3915 ;
  assign n4140 = ( ~n454 & n3915 ) | ( ~n454 & n3985 ) | ( n3915 & n3985 ) ;
  assign n4141 = ( ~n3920 & n4139 ) | ( ~n3920 & n4140 ) | ( n4139 & n4140 ) ;
  assign n4142 = ( n3920 & n4139 ) | ( n3920 & n4140 ) | ( n4139 & n4140 ) ;
  assign n4143 = ( n3920 & n4141 ) | ( n3920 & ~n4142 ) | ( n4141 & ~n4142 ) ;
  assign n4144 = ( ~n396 & n4138 ) | ( ~n396 & n4143 ) | ( n4138 & n4143 ) ;
  assign n4145 = ( n396 & ~n3921 ) | ( n396 & n3985 ) | ( ~n3921 & n3985 ) ;
  assign n4146 = n396 & ~n3921 ;
  assign n4147 = ( n3926 & n4145 ) | ( n3926 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4148 = ( ~n3926 & n4145 ) | ( ~n3926 & n4146 ) | ( n4145 & n4146 ) ;
  assign n4149 = ( n3926 & ~n4147 ) | ( n3926 & n4148 ) | ( ~n4147 & n4148 ) ;
  assign n4150 = ( ~n344 & n4144 ) | ( ~n344 & n4149 ) | ( n4144 & n4149 ) ;
  assign n4151 = ( n344 & ~n3927 ) | ( n344 & n3985 ) | ( ~n3927 & n3985 ) ;
  assign n4152 = n344 & ~n3927 ;
  assign n4153 = ( n3932 & n4151 ) | ( n3932 & n4152 ) | ( n4151 & n4152 ) ;
  assign n4154 = ( ~n3932 & n4151 ) | ( ~n3932 & n4152 ) | ( n4151 & n4152 ) ;
  assign n4155 = ( n3932 & ~n4153 ) | ( n3932 & n4154 ) | ( ~n4153 & n4154 ) ;
  assign n4156 = ( ~n298 & n4150 ) | ( ~n298 & n4155 ) | ( n4150 & n4155 ) ;
  assign n4157 = n298 & ~n3933 ;
  assign n4158 = ( n298 & ~n3933 ) | ( n298 & n3985 ) | ( ~n3933 & n3985 ) ;
  assign n4159 = ( n3938 & n4157 ) | ( n3938 & n4158 ) | ( n4157 & n4158 ) ;
  assign n4160 = ( ~n3938 & n4157 ) | ( ~n3938 & n4158 ) | ( n4157 & n4158 ) ;
  assign n4161 = ( n3938 & ~n4159 ) | ( n3938 & n4160 ) | ( ~n4159 & n4160 ) ;
  assign n4162 = ( ~n258 & n4156 ) | ( ~n258 & n4161 ) | ( n4156 & n4161 ) ;
  assign n4163 = ( n258 & ~n3939 ) | ( n258 & n3985 ) | ( ~n3939 & n3985 ) ;
  assign n4164 = n258 & ~n3939 ;
  assign n4165 = ( n3944 & n4163 ) | ( n3944 & n4164 ) | ( n4163 & n4164 ) ;
  assign n4166 = ( ~n3944 & n4163 ) | ( ~n3944 & n4164 ) | ( n4163 & n4164 ) ;
  assign n4167 = ( n3944 & ~n4165 ) | ( n3944 & n4166 ) | ( ~n4165 & n4166 ) ;
  assign n4168 = ( ~n225 & n4162 ) | ( ~n225 & n4167 ) | ( n4162 & n4167 ) ;
  assign n4169 = ( n225 & ~n3945 ) | ( n225 & n3985 ) | ( ~n3945 & n3985 ) ;
  assign n4170 = n225 & ~n3945 ;
  assign n4171 = ( n3950 & n4169 ) | ( n3950 & n4170 ) | ( n4169 & n4170 ) ;
  assign n4172 = ( ~n3950 & n4169 ) | ( ~n3950 & n4170 ) | ( n4169 & n4170 ) ;
  assign n4173 = ( n3950 & ~n4171 ) | ( n3950 & n4172 ) | ( ~n4171 & n4172 ) ;
  assign n4174 = ( ~n197 & n4168 ) | ( ~n197 & n4173 ) | ( n4168 & n4173 ) ;
  assign n4175 = ( n197 & ~n3951 ) | ( n197 & n3985 ) | ( ~n3951 & n3985 ) ;
  assign n4176 = n197 & ~n3951 ;
  assign n4177 = ( n3956 & n4175 ) | ( n3956 & n4176 ) | ( n4175 & n4176 ) ;
  assign n4178 = ( ~n3956 & n4175 ) | ( ~n3956 & n4176 ) | ( n4175 & n4176 ) ;
  assign n4179 = ( n3956 & ~n4177 ) | ( n3956 & n4178 ) | ( ~n4177 & n4178 ) ;
  assign n4180 = ( ~n170 & n4174 ) | ( ~n170 & n4179 ) | ( n4174 & n4179 ) ;
  assign n4181 = ( n170 & ~n3957 ) | ( n170 & n3985 ) | ( ~n3957 & n3985 ) ;
  assign n4182 = n170 & ~n3957 ;
  assign n4183 = ( n3962 & n4181 ) | ( n3962 & n4182 ) | ( n4181 & n4182 ) ;
  assign n4184 = ( ~n3962 & n4181 ) | ( ~n3962 & n4182 ) | ( n4181 & n4182 ) ;
  assign n4185 = ( n3962 & ~n4183 ) | ( n3962 & n4184 ) | ( ~n4183 & n4184 ) ;
  assign n4186 = ( ~n142 & n4180 ) | ( ~n142 & n4185 ) | ( n4180 & n4185 ) ;
  assign n4187 = ( n142 & ~n3963 ) | ( n142 & n3985 ) | ( ~n3963 & n3985 ) ;
  assign n4188 = n142 & ~n3963 ;
  assign n4189 = ( n3968 & n4187 ) | ( n3968 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4190 = ( ~n3968 & n4187 ) | ( ~n3968 & n4188 ) | ( n4187 & n4188 ) ;
  assign n4191 = ( n3968 & ~n4189 ) | ( n3968 & n4190 ) | ( ~n4189 & n4190 ) ;
  assign n4192 = ( ~n132 & n4186 ) | ( ~n132 & n4191 ) | ( n4186 & n4191 ) ;
  assign n4193 = ( n132 & ~n3969 ) | ( n132 & n3985 ) | ( ~n3969 & n3985 ) ;
  assign n4194 = n132 & ~n3969 ;
  assign n4195 = ( n3974 & n4193 ) | ( n3974 & n4194 ) | ( n4193 & n4194 ) ;
  assign n4196 = ( ~n3974 & n4193 ) | ( ~n3974 & n4194 ) | ( n4193 & n4194 ) ;
  assign n4197 = ( n3974 & ~n4195 ) | ( n3974 & n4196 ) | ( ~n4195 & n4196 ) ;
  assign n4198 = ( ~n131 & n4192 ) | ( ~n131 & n4197 ) | ( n4192 & n4197 ) ;
  assign n4199 = ( n3987 & ~n3988 ) | ( n3987 & n4198 ) | ( ~n3988 & n4198 ) ;
  assign n4200 = ( ~n131 & n3776 ) | ( ~n131 & n3975 ) | ( n3776 & n3975 ) ;
  assign n4201 = ~n3983 & n4200 ;
  assign n4202 = ( n131 & n3988 ) | ( n131 & n4201 ) | ( n3988 & n4201 ) ;
  assign n4203 = n4199 | n4202 ;
  assign n4204 = n4192 & n4197 ;
  assign n4205 = n4192 | n4197 ;
  assign n4206 = ~n4204 & n4205 ;
  assign n4207 = ( n131 & ~n4192 ) | ( n131 & n4202 ) | ( ~n4192 & n4202 ) ;
  assign n4208 = n4206 & n4207 ;
  assign n4209 = ( n132 & ~n4186 ) | ( n132 & n4203 ) | ( ~n4186 & n4203 ) ;
  assign n4210 = n132 & ~n4186 ;
  assign n4211 = ( n4191 & ~n4209 ) | ( n4191 & n4210 ) | ( ~n4209 & n4210 ) ;
  assign n4212 = ( n4191 & n4209 ) | ( n4191 & n4210 ) | ( n4209 & n4210 ) ;
  assign n4213 = ( n4209 & n4211 ) | ( n4209 & ~n4212 ) | ( n4211 & ~n4212 ) ;
  assign n4214 = n131 & ~n4213 ;
  assign n4215 = x55 & n4203 ;
  assign n4216 = x52 | x53 ;
  assign n4217 = x54 | n4216 ;
  assign n4218 = ( x55 & n4203 ) | ( x55 & n4217 ) | ( n4203 & n4217 ) ;
  assign n4219 = ( n3985 & n4215 ) | ( n3985 & ~n4218 ) | ( n4215 & ~n4218 ) ;
  assign n4220 = ( ~x55 & n4203 ) | ( ~x55 & n4216 ) | ( n4203 & n4216 ) ;
  assign n4221 = x54 | n4220 ;
  assign n4222 = ( x54 & x55 ) | ( x54 & n4203 ) | ( x55 & n4203 ) ;
  assign n4223 = ( x55 & n4221 ) | ( x55 & ~n4222 ) | ( n4221 & ~n4222 ) ;
  assign n4224 = ~n4219 & n4223 ;
  assign n4225 = ~n3989 & n4203 ;
  assign n4226 = n3985 & ~n4203 ;
  assign n4227 = ( x56 & n4225 ) | ( x56 & n4226 ) | ( n4225 & n4226 ) ;
  assign n4228 = ( ~x56 & n4225 ) | ( ~x56 & n4226 ) | ( n4225 & n4226 ) ;
  assign n4229 = ( x56 & ~n4227 ) | ( x56 & n4228 ) | ( ~n4227 & n4228 ) ;
  assign n4230 = ( ~n3772 & n4224 ) | ( ~n3772 & n4229 ) | ( n4224 & n4229 ) ;
  assign n4231 = ~n3772 & n3985 ;
  assign n4232 = ( n3996 & n4203 ) | ( n3996 & n4231 ) | ( n4203 & n4231 ) ;
  assign n4233 = ( ~x57 & n4228 ) | ( ~x57 & n4232 ) | ( n4228 & n4232 ) ;
  assign n4234 = ( x57 & n4228 ) | ( x57 & n4232 ) | ( n4228 & n4232 ) ;
  assign n4235 = ( x57 & n4233 ) | ( x57 & ~n4234 ) | ( n4233 & ~n4234 ) ;
  assign n4236 = ( ~n3567 & n4230 ) | ( ~n3567 & n4235 ) | ( n4230 & n4235 ) ;
  assign n4237 = n3567 & ~n3995 ;
  assign n4238 = ( n3567 & ~n3995 ) | ( n3567 & n4203 ) | ( ~n3995 & n4203 ) ;
  assign n4239 = ( ~n3999 & n4237 ) | ( ~n3999 & n4238 ) | ( n4237 & n4238 ) ;
  assign n4240 = ( n3999 & n4237 ) | ( n3999 & n4238 ) | ( n4237 & n4238 ) ;
  assign n4241 = ( n3999 & n4239 ) | ( n3999 & ~n4240 ) | ( n4239 & ~n4240 ) ;
  assign n4242 = ( ~n3362 & n4236 ) | ( ~n3362 & n4241 ) | ( n4236 & n4241 ) ;
  assign n4243 = ( n3362 & ~n4000 ) | ( n3362 & n4203 ) | ( ~n4000 & n4203 ) ;
  assign n4244 = n3362 & ~n4000 ;
  assign n4245 = ( n4005 & n4243 ) | ( n4005 & n4244 ) | ( n4243 & n4244 ) ;
  assign n4246 = ( ~n4005 & n4243 ) | ( ~n4005 & n4244 ) | ( n4243 & n4244 ) ;
  assign n4247 = ( n4005 & ~n4245 ) | ( n4005 & n4246 ) | ( ~n4245 & n4246 ) ;
  assign n4248 = ( ~n3169 & n4242 ) | ( ~n3169 & n4247 ) | ( n4242 & n4247 ) ;
  assign n4249 = ( n3169 & ~n4006 ) | ( n3169 & n4203 ) | ( ~n4006 & n4203 ) ;
  assign n4250 = n3169 & ~n4006 ;
  assign n4251 = ( n4011 & n4249 ) | ( n4011 & n4250 ) | ( n4249 & n4250 ) ;
  assign n4252 = ( ~n4011 & n4249 ) | ( ~n4011 & n4250 ) | ( n4249 & n4250 ) ;
  assign n4253 = ( n4011 & ~n4251 ) | ( n4011 & n4252 ) | ( ~n4251 & n4252 ) ;
  assign n4254 = ( ~n2979 & n4248 ) | ( ~n2979 & n4253 ) | ( n4248 & n4253 ) ;
  assign n4255 = ( n2979 & ~n4012 ) | ( n2979 & n4203 ) | ( ~n4012 & n4203 ) ;
  assign n4256 = n2979 & ~n4012 ;
  assign n4257 = ( n4017 & n4255 ) | ( n4017 & n4256 ) | ( n4255 & n4256 ) ;
  assign n4258 = ( ~n4017 & n4255 ) | ( ~n4017 & n4256 ) | ( n4255 & n4256 ) ;
  assign n4259 = ( n4017 & ~n4257 ) | ( n4017 & n4258 ) | ( ~n4257 & n4258 ) ;
  assign n4260 = ( ~n2791 & n4254 ) | ( ~n2791 & n4259 ) | ( n4254 & n4259 ) ;
  assign n4261 = n2791 & ~n4018 ;
  assign n4262 = ( n2791 & ~n4018 ) | ( n2791 & n4203 ) | ( ~n4018 & n4203 ) ;
  assign n4263 = ( ~n4023 & n4261 ) | ( ~n4023 & n4262 ) | ( n4261 & n4262 ) ;
  assign n4264 = ( n4023 & n4261 ) | ( n4023 & n4262 ) | ( n4261 & n4262 ) ;
  assign n4265 = ( n4023 & n4263 ) | ( n4023 & ~n4264 ) | ( n4263 & ~n4264 ) ;
  assign n4266 = ( ~n2615 & n4260 ) | ( ~n2615 & n4265 ) | ( n4260 & n4265 ) ;
  assign n4267 = n2615 & ~n4024 ;
  assign n4268 = ( n2615 & ~n4024 ) | ( n2615 & n4203 ) | ( ~n4024 & n4203 ) ;
  assign n4269 = ( n4029 & n4267 ) | ( n4029 & n4268 ) | ( n4267 & n4268 ) ;
  assign n4270 = ( ~n4029 & n4267 ) | ( ~n4029 & n4268 ) | ( n4267 & n4268 ) ;
  assign n4271 = ( n4029 & ~n4269 ) | ( n4029 & n4270 ) | ( ~n4269 & n4270 ) ;
  assign n4272 = ( ~n2443 & n4266 ) | ( ~n2443 & n4271 ) | ( n4266 & n4271 ) ;
  assign n4273 = ( n2443 & ~n4030 ) | ( n2443 & n4203 ) | ( ~n4030 & n4203 ) ;
  assign n4274 = n2443 & ~n4030 ;
  assign n4275 = ( n4035 & n4273 ) | ( n4035 & n4274 ) | ( n4273 & n4274 ) ;
  assign n4276 = ( ~n4035 & n4273 ) | ( ~n4035 & n4274 ) | ( n4273 & n4274 ) ;
  assign n4277 = ( n4035 & ~n4275 ) | ( n4035 & n4276 ) | ( ~n4275 & n4276 ) ;
  assign n4278 = ( ~n2277 & n4272 ) | ( ~n2277 & n4277 ) | ( n4272 & n4277 ) ;
  assign n4279 = ( n2277 & ~n4036 ) | ( n2277 & n4203 ) | ( ~n4036 & n4203 ) ;
  assign n4280 = n2277 & ~n4036 ;
  assign n4281 = ( n4041 & n4279 ) | ( n4041 & n4280 ) | ( n4279 & n4280 ) ;
  assign n4282 = ( ~n4041 & n4279 ) | ( ~n4041 & n4280 ) | ( n4279 & n4280 ) ;
  assign n4283 = ( n4041 & ~n4281 ) | ( n4041 & n4282 ) | ( ~n4281 & n4282 ) ;
  assign n4284 = ( ~n2111 & n4278 ) | ( ~n2111 & n4283 ) | ( n4278 & n4283 ) ;
  assign n4285 = ( n2111 & ~n4042 ) | ( n2111 & n4203 ) | ( ~n4042 & n4203 ) ;
  assign n4286 = n2111 & ~n4042 ;
  assign n4287 = ( n4047 & n4285 ) | ( n4047 & n4286 ) | ( n4285 & n4286 ) ;
  assign n4288 = ( ~n4047 & n4285 ) | ( ~n4047 & n4286 ) | ( n4285 & n4286 ) ;
  assign n4289 = ( n4047 & ~n4287 ) | ( n4047 & n4288 ) | ( ~n4287 & n4288 ) ;
  assign n4290 = ( ~n1949 & n4284 ) | ( ~n1949 & n4289 ) | ( n4284 & n4289 ) ;
  assign n4291 = ( n1949 & ~n4048 ) | ( n1949 & n4203 ) | ( ~n4048 & n4203 ) ;
  assign n4292 = n1949 & ~n4048 ;
  assign n4293 = ( n4053 & n4291 ) | ( n4053 & n4292 ) | ( n4291 & n4292 ) ;
  assign n4294 = ( ~n4053 & n4291 ) | ( ~n4053 & n4292 ) | ( n4291 & n4292 ) ;
  assign n4295 = ( n4053 & ~n4293 ) | ( n4053 & n4294 ) | ( ~n4293 & n4294 ) ;
  assign n4296 = ( ~n1802 & n4290 ) | ( ~n1802 & n4295 ) | ( n4290 & n4295 ) ;
  assign n4297 = ~n1802 & n4054 ;
  assign n4298 = ( ~n1802 & n4054 ) | ( ~n1802 & n4203 ) | ( n4054 & n4203 ) ;
  assign n4299 = ( n4059 & n4297 ) | ( n4059 & n4298 ) | ( n4297 & n4298 ) ;
  assign n4300 = ( ~n4059 & n4297 ) | ( ~n4059 & n4298 ) | ( n4297 & n4298 ) ;
  assign n4301 = ( n4059 & ~n4299 ) | ( n4059 & n4300 ) | ( ~n4299 & n4300 ) ;
  assign n4302 = ( ~n1661 & n4296 ) | ( ~n1661 & n4301 ) | ( n4296 & n4301 ) ;
  assign n4303 = ~n1661 & n4060 ;
  assign n4304 = ( ~n1661 & n4060 ) | ( ~n1661 & n4203 ) | ( n4060 & n4203 ) ;
  assign n4305 = ( ~n4065 & n4303 ) | ( ~n4065 & n4304 ) | ( n4303 & n4304 ) ;
  assign n4306 = ( n4065 & n4303 ) | ( n4065 & n4304 ) | ( n4303 & n4304 ) ;
  assign n4307 = ( n4065 & n4305 ) | ( n4065 & ~n4306 ) | ( n4305 & ~n4306 ) ;
  assign n4308 = ( ~n1523 & n4302 ) | ( ~n1523 & n4307 ) | ( n4302 & n4307 ) ;
  assign n4309 = ( n1523 & ~n4066 ) | ( n1523 & n4203 ) | ( ~n4066 & n4203 ) ;
  assign n4310 = n1523 & ~n4066 ;
  assign n4311 = ( n4071 & n4309 ) | ( n4071 & n4310 ) | ( n4309 & n4310 ) ;
  assign n4312 = ( ~n4071 & n4309 ) | ( ~n4071 & n4310 ) | ( n4309 & n4310 ) ;
  assign n4313 = ( n4071 & ~n4311 ) | ( n4071 & n4312 ) | ( ~n4311 & n4312 ) ;
  assign n4314 = ( ~n1393 & n4308 ) | ( ~n1393 & n4313 ) | ( n4308 & n4313 ) ;
  assign n4315 = ~n1393 & n4072 ;
  assign n4316 = ( ~n1393 & n4072 ) | ( ~n1393 & n4203 ) | ( n4072 & n4203 ) ;
  assign n4317 = ( n4077 & n4315 ) | ( n4077 & n4316 ) | ( n4315 & n4316 ) ;
  assign n4318 = ( ~n4077 & n4315 ) | ( ~n4077 & n4316 ) | ( n4315 & n4316 ) ;
  assign n4319 = ( n4077 & ~n4317 ) | ( n4077 & n4318 ) | ( ~n4317 & n4318 ) ;
  assign n4320 = ( ~n1266 & n4314 ) | ( ~n1266 & n4319 ) | ( n4314 & n4319 ) ;
  assign n4321 = ( n1266 & ~n4078 ) | ( n1266 & n4203 ) | ( ~n4078 & n4203 ) ;
  assign n4322 = n1266 & ~n4078 ;
  assign n4323 = ( n4083 & n4321 ) | ( n4083 & n4322 ) | ( n4321 & n4322 ) ;
  assign n4324 = ( ~n4083 & n4321 ) | ( ~n4083 & n4322 ) | ( n4321 & n4322 ) ;
  assign n4325 = ( n4083 & ~n4323 ) | ( n4083 & n4324 ) | ( ~n4323 & n4324 ) ;
  assign n4326 = ( ~n1150 & n4320 ) | ( ~n1150 & n4325 ) | ( n4320 & n4325 ) ;
  assign n4327 = ~n1150 & n4084 ;
  assign n4328 = ( ~n1150 & n4084 ) | ( ~n1150 & n4203 ) | ( n4084 & n4203 ) ;
  assign n4329 = ( n4089 & n4327 ) | ( n4089 & n4328 ) | ( n4327 & n4328 ) ;
  assign n4330 = ( ~n4089 & n4327 ) | ( ~n4089 & n4328 ) | ( n4327 & n4328 ) ;
  assign n4331 = ( n4089 & ~n4329 ) | ( n4089 & n4330 ) | ( ~n4329 & n4330 ) ;
  assign n4332 = ( ~n1038 & n4326 ) | ( ~n1038 & n4331 ) | ( n4326 & n4331 ) ;
  assign n4333 = ( n1038 & ~n4090 ) | ( n1038 & n4203 ) | ( ~n4090 & n4203 ) ;
  assign n4334 = n1038 & ~n4090 ;
  assign n4335 = ( n4095 & n4333 ) | ( n4095 & n4334 ) | ( n4333 & n4334 ) ;
  assign n4336 = ( ~n4095 & n4333 ) | ( ~n4095 & n4334 ) | ( n4333 & n4334 ) ;
  assign n4337 = ( n4095 & ~n4335 ) | ( n4095 & n4336 ) | ( ~n4335 & n4336 ) ;
  assign n4338 = ( ~n933 & n4332 ) | ( ~n933 & n4337 ) | ( n4332 & n4337 ) ;
  assign n4339 = ( n933 & ~n4096 ) | ( n933 & n4203 ) | ( ~n4096 & n4203 ) ;
  assign n4340 = n933 & ~n4096 ;
  assign n4341 = ( n4101 & n4339 ) | ( n4101 & n4340 ) | ( n4339 & n4340 ) ;
  assign n4342 = ( ~n4101 & n4339 ) | ( ~n4101 & n4340 ) | ( n4339 & n4340 ) ;
  assign n4343 = ( n4101 & ~n4341 ) | ( n4101 & n4342 ) | ( ~n4341 & n4342 ) ;
  assign n4344 = ( ~n839 & n4338 ) | ( ~n839 & n4343 ) | ( n4338 & n4343 ) ;
  assign n4345 = ~n839 & n4102 ;
  assign n4346 = ( ~n839 & n4102 ) | ( ~n839 & n4203 ) | ( n4102 & n4203 ) ;
  assign n4347 = ( ~n4107 & n4345 ) | ( ~n4107 & n4346 ) | ( n4345 & n4346 ) ;
  assign n4348 = ( n4107 & n4345 ) | ( n4107 & n4346 ) | ( n4345 & n4346 ) ;
  assign n4349 = ( n4107 & n4347 ) | ( n4107 & ~n4348 ) | ( n4347 & ~n4348 ) ;
  assign n4350 = ( ~n746 & n4344 ) | ( ~n746 & n4349 ) | ( n4344 & n4349 ) ;
  assign n4351 = n746 & ~n4108 ;
  assign n4352 = ( n746 & ~n4108 ) | ( n746 & n4203 ) | ( ~n4108 & n4203 ) ;
  assign n4353 = ( ~n4113 & n4351 ) | ( ~n4113 & n4352 ) | ( n4351 & n4352 ) ;
  assign n4354 = ( n4113 & n4351 ) | ( n4113 & n4352 ) | ( n4351 & n4352 ) ;
  assign n4355 = ( n4113 & n4353 ) | ( n4113 & ~n4354 ) | ( n4353 & ~n4354 ) ;
  assign n4356 = ( ~n664 & n4350 ) | ( ~n664 & n4355 ) | ( n4350 & n4355 ) ;
  assign n4357 = ( n664 & ~n4114 ) | ( n664 & n4203 ) | ( ~n4114 & n4203 ) ;
  assign n4358 = n664 & ~n4114 ;
  assign n4359 = ( n4119 & n4357 ) | ( n4119 & n4358 ) | ( n4357 & n4358 ) ;
  assign n4360 = ( ~n4119 & n4357 ) | ( ~n4119 & n4358 ) | ( n4357 & n4358 ) ;
  assign n4361 = ( n4119 & ~n4359 ) | ( n4119 & n4360 ) | ( ~n4359 & n4360 ) ;
  assign n4362 = ( ~n588 & n4356 ) | ( ~n588 & n4361 ) | ( n4356 & n4361 ) ;
  assign n4363 = ( n588 & ~n4120 ) | ( n588 & n4203 ) | ( ~n4120 & n4203 ) ;
  assign n4364 = n588 & ~n4120 ;
  assign n4365 = ( n4125 & n4363 ) | ( n4125 & n4364 ) | ( n4363 & n4364 ) ;
  assign n4366 = ( ~n4125 & n4363 ) | ( ~n4125 & n4364 ) | ( n4363 & n4364 ) ;
  assign n4367 = ( n4125 & ~n4365 ) | ( n4125 & n4366 ) | ( ~n4365 & n4366 ) ;
  assign n4368 = ( ~n518 & n4362 ) | ( ~n518 & n4367 ) | ( n4362 & n4367 ) ;
  assign n4369 = ~n518 & n4126 ;
  assign n4370 = ( ~n518 & n4126 ) | ( ~n518 & n4203 ) | ( n4126 & n4203 ) ;
  assign n4371 = ( ~n4131 & n4369 ) | ( ~n4131 & n4370 ) | ( n4369 & n4370 ) ;
  assign n4372 = ( n4131 & n4369 ) | ( n4131 & n4370 ) | ( n4369 & n4370 ) ;
  assign n4373 = ( n4131 & n4371 ) | ( n4131 & ~n4372 ) | ( n4371 & ~n4372 ) ;
  assign n4374 = ( ~n454 & n4368 ) | ( ~n454 & n4373 ) | ( n4368 & n4373 ) ;
  assign n4375 = ~n454 & n4132 ;
  assign n4376 = ( ~n454 & n4132 ) | ( ~n454 & n4203 ) | ( n4132 & n4203 ) ;
  assign n4377 = ( n4137 & n4375 ) | ( n4137 & n4376 ) | ( n4375 & n4376 ) ;
  assign n4378 = ( ~n4137 & n4375 ) | ( ~n4137 & n4376 ) | ( n4375 & n4376 ) ;
  assign n4379 = ( n4137 & ~n4377 ) | ( n4137 & n4378 ) | ( ~n4377 & n4378 ) ;
  assign n4380 = ( ~n396 & n4374 ) | ( ~n396 & n4379 ) | ( n4374 & n4379 ) ;
  assign n4381 = ~n396 & n4138 ;
  assign n4382 = ( ~n396 & n4138 ) | ( ~n396 & n4203 ) | ( n4138 & n4203 ) ;
  assign n4383 = ( ~n4143 & n4381 ) | ( ~n4143 & n4382 ) | ( n4381 & n4382 ) ;
  assign n4384 = ( n4143 & n4381 ) | ( n4143 & n4382 ) | ( n4381 & n4382 ) ;
  assign n4385 = ( n4143 & n4383 ) | ( n4143 & ~n4384 ) | ( n4383 & ~n4384 ) ;
  assign n4386 = ( ~n344 & n4380 ) | ( ~n344 & n4385 ) | ( n4380 & n4385 ) ;
  assign n4387 = ~n344 & n4144 ;
  assign n4388 = ( ~n344 & n4144 ) | ( ~n344 & n4203 ) | ( n4144 & n4203 ) ;
  assign n4389 = ( n4149 & n4387 ) | ( n4149 & n4388 ) | ( n4387 & n4388 ) ;
  assign n4390 = ( ~n4149 & n4387 ) | ( ~n4149 & n4388 ) | ( n4387 & n4388 ) ;
  assign n4391 = ( n4149 & ~n4389 ) | ( n4149 & n4390 ) | ( ~n4389 & n4390 ) ;
  assign n4392 = ( ~n298 & n4386 ) | ( ~n298 & n4391 ) | ( n4386 & n4391 ) ;
  assign n4393 = ~n298 & n4150 ;
  assign n4394 = ( ~n298 & n4150 ) | ( ~n298 & n4203 ) | ( n4150 & n4203 ) ;
  assign n4395 = ( n4155 & n4393 ) | ( n4155 & n4394 ) | ( n4393 & n4394 ) ;
  assign n4396 = ( ~n4155 & n4393 ) | ( ~n4155 & n4394 ) | ( n4393 & n4394 ) ;
  assign n4397 = ( n4155 & ~n4395 ) | ( n4155 & n4396 ) | ( ~n4395 & n4396 ) ;
  assign n4398 = ( ~n258 & n4392 ) | ( ~n258 & n4397 ) | ( n4392 & n4397 ) ;
  assign n4399 = n258 & ~n4156 ;
  assign n4400 = ( n258 & ~n4156 ) | ( n258 & n4203 ) | ( ~n4156 & n4203 ) ;
  assign n4401 = ( n4161 & n4399 ) | ( n4161 & n4400 ) | ( n4399 & n4400 ) ;
  assign n4402 = ( ~n4161 & n4399 ) | ( ~n4161 & n4400 ) | ( n4399 & n4400 ) ;
  assign n4403 = ( n4161 & ~n4401 ) | ( n4161 & n4402 ) | ( ~n4401 & n4402 ) ;
  assign n4404 = ( ~n225 & n4398 ) | ( ~n225 & n4403 ) | ( n4398 & n4403 ) ;
  assign n4405 = ( n225 & ~n4162 ) | ( n225 & n4203 ) | ( ~n4162 & n4203 ) ;
  assign n4406 = n225 & ~n4162 ;
  assign n4407 = ( n4167 & n4405 ) | ( n4167 & n4406 ) | ( n4405 & n4406 ) ;
  assign n4408 = ( ~n4167 & n4405 ) | ( ~n4167 & n4406 ) | ( n4405 & n4406 ) ;
  assign n4409 = ( n4167 & ~n4407 ) | ( n4167 & n4408 ) | ( ~n4407 & n4408 ) ;
  assign n4410 = ( ~n197 & n4404 ) | ( ~n197 & n4409 ) | ( n4404 & n4409 ) ;
  assign n4411 = ( n197 & ~n4168 ) | ( n197 & n4203 ) | ( ~n4168 & n4203 ) ;
  assign n4412 = n197 & ~n4168 ;
  assign n4413 = ( n4173 & n4411 ) | ( n4173 & n4412 ) | ( n4411 & n4412 ) ;
  assign n4414 = ( ~n4173 & n4411 ) | ( ~n4173 & n4412 ) | ( n4411 & n4412 ) ;
  assign n4415 = ( n4173 & ~n4413 ) | ( n4173 & n4414 ) | ( ~n4413 & n4414 ) ;
  assign n4416 = ( ~n170 & n4410 ) | ( ~n170 & n4415 ) | ( n4410 & n4415 ) ;
  assign n4417 = n170 & ~n4174 ;
  assign n4418 = ( n170 & ~n4174 ) | ( n170 & n4203 ) | ( ~n4174 & n4203 ) ;
  assign n4419 = ( n4179 & n4417 ) | ( n4179 & n4418 ) | ( n4417 & n4418 ) ;
  assign n4420 = ( ~n4179 & n4417 ) | ( ~n4179 & n4418 ) | ( n4417 & n4418 ) ;
  assign n4421 = ( n4179 & ~n4419 ) | ( n4179 & n4420 ) | ( ~n4419 & n4420 ) ;
  assign n4422 = ( ~n142 & n4416 ) | ( ~n142 & n4421 ) | ( n4416 & n4421 ) ;
  assign n4423 = ~n142 & n4180 ;
  assign n4424 = ( ~n142 & n4180 ) | ( ~n142 & n4203 ) | ( n4180 & n4203 ) ;
  assign n4425 = ( ~n4185 & n4423 ) | ( ~n4185 & n4424 ) | ( n4423 & n4424 ) ;
  assign n4426 = ( n4185 & n4423 ) | ( n4185 & n4424 ) | ( n4423 & n4424 ) ;
  assign n4427 = ( n4185 & n4425 ) | ( n4185 & ~n4426 ) | ( n4425 & ~n4426 ) ;
  assign n4428 = ( ~n132 & n4422 ) | ( ~n132 & n4427 ) | ( n4422 & n4427 ) ;
  assign n4429 = ( n4203 & ~n4206 ) | ( n4203 & n4213 ) | ( ~n4206 & n4213 ) ;
  assign n4430 = ~n131 & n4429 ;
  assign n4431 = ( ~n4214 & n4428 ) | ( ~n4214 & n4430 ) | ( n4428 & n4430 ) ;
  assign n4432 = n4208 | n4431 ;
  assign n4433 = n4213 | n4428 ;
  assign n4434 = n4208 & ~n4213 ;
  assign n4435 = n4428 & ~n4434 ;
  assign n4436 = ( n4430 & n4433 ) | ( n4430 & ~n4435 ) | ( n4433 & ~n4435 ) ;
  assign n4437 = ( n131 & n4213 ) | ( n131 & n4428 ) | ( n4213 & n4428 ) ;
  assign n4438 = ( ~n4433 & n4436 ) | ( ~n4433 & n4437 ) | ( n4436 & n4437 ) ;
  assign n4439 = ( n132 & ~n4422 ) | ( n132 & n4432 ) | ( ~n4422 & n4432 ) ;
  assign n4440 = n132 & ~n4422 ;
  assign n4441 = ( n4427 & n4439 ) | ( n4427 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4442 = ( n4427 & ~n4439 ) | ( n4427 & n4440 ) | ( ~n4439 & n4440 ) ;
  assign n4443 = ( n4439 & ~n4441 ) | ( n4439 & n4442 ) | ( ~n4441 & n4442 ) ;
  assign n4444 = x50 | x51 ;
  assign n4445 = x52 | n4444 ;
  assign n4446 = ~n4203 & n4445 ;
  assign n4447 = ( x53 & ~n4432 ) | ( x53 & n4446 ) | ( ~n4432 & n4446 ) ;
  assign n4448 = n4203 & ~n4445 ;
  assign n4449 = ~n4216 & n4432 ;
  assign n4450 = ( n4447 & ~n4448 ) | ( n4447 & n4449 ) | ( ~n4448 & n4449 ) ;
  assign n4451 = n4203 & ~n4432 ;
  assign n4452 = ( x54 & n4449 ) | ( x54 & n4451 ) | ( n4449 & n4451 ) ;
  assign n4453 = ( ~x54 & n4449 ) | ( ~x54 & n4451 ) | ( n4449 & n4451 ) ;
  assign n4454 = ( x54 & ~n4452 ) | ( x54 & n4453 ) | ( ~n4452 & n4453 ) ;
  assign n4455 = ( ~n3985 & n4450 ) | ( ~n3985 & n4454 ) | ( n4450 & n4454 ) ;
  assign n4456 = ~n3985 & n4203 ;
  assign n4457 = ( n4226 & n4432 ) | ( n4226 & n4456 ) | ( n4432 & n4456 ) ;
  assign n4458 = ( ~x55 & n4453 ) | ( ~x55 & n4457 ) | ( n4453 & n4457 ) ;
  assign n4459 = ( x55 & n4453 ) | ( x55 & n4457 ) | ( n4453 & n4457 ) ;
  assign n4460 = ( x55 & n4458 ) | ( x55 & ~n4459 ) | ( n4458 & ~n4459 ) ;
  assign n4461 = ( ~n3772 & n4455 ) | ( ~n3772 & n4460 ) | ( n4455 & n4460 ) ;
  assign n4462 = n3772 & ~n4224 ;
  assign n4463 = ( n3772 & ~n4224 ) | ( n3772 & n4432 ) | ( ~n4224 & n4432 ) ;
  assign n4464 = ( n4229 & n4462 ) | ( n4229 & n4463 ) | ( n4462 & n4463 ) ;
  assign n4465 = ( ~n4229 & n4462 ) | ( ~n4229 & n4463 ) | ( n4462 & n4463 ) ;
  assign n4466 = ( n4229 & ~n4464 ) | ( n4229 & n4465 ) | ( ~n4464 & n4465 ) ;
  assign n4467 = ( ~n3567 & n4461 ) | ( ~n3567 & n4466 ) | ( n4461 & n4466 ) ;
  assign n4468 = n3567 & ~n4230 ;
  assign n4469 = ( n3567 & ~n4230 ) | ( n3567 & n4432 ) | ( ~n4230 & n4432 ) ;
  assign n4470 = ( n4235 & n4468 ) | ( n4235 & n4469 ) | ( n4468 & n4469 ) ;
  assign n4471 = ( ~n4235 & n4468 ) | ( ~n4235 & n4469 ) | ( n4468 & n4469 ) ;
  assign n4472 = ( n4235 & ~n4470 ) | ( n4235 & n4471 ) | ( ~n4470 & n4471 ) ;
  assign n4473 = ( ~n3362 & n4467 ) | ( ~n3362 & n4472 ) | ( n4467 & n4472 ) ;
  assign n4474 = n3362 & ~n4236 ;
  assign n4475 = ( n3362 & ~n4236 ) | ( n3362 & n4432 ) | ( ~n4236 & n4432 ) ;
  assign n4476 = ( ~n4241 & n4474 ) | ( ~n4241 & n4475 ) | ( n4474 & n4475 ) ;
  assign n4477 = ( n4241 & n4474 ) | ( n4241 & n4475 ) | ( n4474 & n4475 ) ;
  assign n4478 = ( n4241 & n4476 ) | ( n4241 & ~n4477 ) | ( n4476 & ~n4477 ) ;
  assign n4479 = ( ~n3169 & n4473 ) | ( ~n3169 & n4478 ) | ( n4473 & n4478 ) ;
  assign n4480 = ~n3169 & n4242 ;
  assign n4481 = ( ~n3169 & n4242 ) | ( ~n3169 & n4432 ) | ( n4242 & n4432 ) ;
  assign n4482 = ( n4247 & n4480 ) | ( n4247 & n4481 ) | ( n4480 & n4481 ) ;
  assign n4483 = ( ~n4247 & n4480 ) | ( ~n4247 & n4481 ) | ( n4480 & n4481 ) ;
  assign n4484 = ( n4247 & ~n4482 ) | ( n4247 & n4483 ) | ( ~n4482 & n4483 ) ;
  assign n4485 = ( ~n2979 & n4479 ) | ( ~n2979 & n4484 ) | ( n4479 & n4484 ) ;
  assign n4486 = ~n2979 & n4248 ;
  assign n4487 = ( ~n2979 & n4248 ) | ( ~n2979 & n4432 ) | ( n4248 & n4432 ) ;
  assign n4488 = ( ~n4253 & n4486 ) | ( ~n4253 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4489 = ( n4253 & n4486 ) | ( n4253 & n4487 ) | ( n4486 & n4487 ) ;
  assign n4490 = ( n4253 & n4488 ) | ( n4253 & ~n4489 ) | ( n4488 & ~n4489 ) ;
  assign n4491 = ( ~n2791 & n4485 ) | ( ~n2791 & n4490 ) | ( n4485 & n4490 ) ;
  assign n4492 = ( n2791 & ~n4254 ) | ( n2791 & n4432 ) | ( ~n4254 & n4432 ) ;
  assign n4493 = n2791 & ~n4254 ;
  assign n4494 = ( n4259 & n4492 ) | ( n4259 & n4493 ) | ( n4492 & n4493 ) ;
  assign n4495 = ( ~n4259 & n4492 ) | ( ~n4259 & n4493 ) | ( n4492 & n4493 ) ;
  assign n4496 = ( n4259 & ~n4494 ) | ( n4259 & n4495 ) | ( ~n4494 & n4495 ) ;
  assign n4497 = ( ~n2615 & n4491 ) | ( ~n2615 & n4496 ) | ( n4491 & n4496 ) ;
  assign n4498 = n2615 & ~n4260 ;
  assign n4499 = ( n2615 & ~n4260 ) | ( n2615 & n4432 ) | ( ~n4260 & n4432 ) ;
  assign n4500 = ( ~n4265 & n4498 ) | ( ~n4265 & n4499 ) | ( n4498 & n4499 ) ;
  assign n4501 = ( n4265 & n4498 ) | ( n4265 & n4499 ) | ( n4498 & n4499 ) ;
  assign n4502 = ( n4265 & n4500 ) | ( n4265 & ~n4501 ) | ( n4500 & ~n4501 ) ;
  assign n4503 = ( ~n2443 & n4497 ) | ( ~n2443 & n4502 ) | ( n4497 & n4502 ) ;
  assign n4504 = ( n2443 & ~n4266 ) | ( n2443 & n4432 ) | ( ~n4266 & n4432 ) ;
  assign n4505 = n2443 & ~n4266 ;
  assign n4506 = ( n4271 & n4504 ) | ( n4271 & n4505 ) | ( n4504 & n4505 ) ;
  assign n4507 = ( ~n4271 & n4504 ) | ( ~n4271 & n4505 ) | ( n4504 & n4505 ) ;
  assign n4508 = ( n4271 & ~n4506 ) | ( n4271 & n4507 ) | ( ~n4506 & n4507 ) ;
  assign n4509 = ( ~n2277 & n4503 ) | ( ~n2277 & n4508 ) | ( n4503 & n4508 ) ;
  assign n4510 = ( n2277 & ~n4272 ) | ( n2277 & n4432 ) | ( ~n4272 & n4432 ) ;
  assign n4511 = n2277 & ~n4272 ;
  assign n4512 = ( n4277 & n4510 ) | ( n4277 & n4511 ) | ( n4510 & n4511 ) ;
  assign n4513 = ( ~n4277 & n4510 ) | ( ~n4277 & n4511 ) | ( n4510 & n4511 ) ;
  assign n4514 = ( n4277 & ~n4512 ) | ( n4277 & n4513 ) | ( ~n4512 & n4513 ) ;
  assign n4515 = ( ~n2111 & n4509 ) | ( ~n2111 & n4514 ) | ( n4509 & n4514 ) ;
  assign n4516 = ( n2111 & ~n4278 ) | ( n2111 & n4432 ) | ( ~n4278 & n4432 ) ;
  assign n4517 = n2111 & ~n4278 ;
  assign n4518 = ( n4283 & n4516 ) | ( n4283 & n4517 ) | ( n4516 & n4517 ) ;
  assign n4519 = ( ~n4283 & n4516 ) | ( ~n4283 & n4517 ) | ( n4516 & n4517 ) ;
  assign n4520 = ( n4283 & ~n4518 ) | ( n4283 & n4519 ) | ( ~n4518 & n4519 ) ;
  assign n4521 = ( ~n1949 & n4515 ) | ( ~n1949 & n4520 ) | ( n4515 & n4520 ) ;
  assign n4522 = ~n1949 & n4284 ;
  assign n4523 = ( ~n1949 & n4284 ) | ( ~n1949 & n4432 ) | ( n4284 & n4432 ) ;
  assign n4524 = ( ~n4289 & n4522 ) | ( ~n4289 & n4523 ) | ( n4522 & n4523 ) ;
  assign n4525 = ( n4289 & n4522 ) | ( n4289 & n4523 ) | ( n4522 & n4523 ) ;
  assign n4526 = ( n4289 & n4524 ) | ( n4289 & ~n4525 ) | ( n4524 & ~n4525 ) ;
  assign n4527 = ( ~n1802 & n4521 ) | ( ~n1802 & n4526 ) | ( n4521 & n4526 ) ;
  assign n4528 = ~n1802 & n4290 ;
  assign n4529 = ( ~n1802 & n4290 ) | ( ~n1802 & n4432 ) | ( n4290 & n4432 ) ;
  assign n4530 = ( ~n4295 & n4528 ) | ( ~n4295 & n4529 ) | ( n4528 & n4529 ) ;
  assign n4531 = ( n4295 & n4528 ) | ( n4295 & n4529 ) | ( n4528 & n4529 ) ;
  assign n4532 = ( n4295 & n4530 ) | ( n4295 & ~n4531 ) | ( n4530 & ~n4531 ) ;
  assign n4533 = ( ~n1661 & n4527 ) | ( ~n1661 & n4532 ) | ( n4527 & n4532 ) ;
  assign n4534 = ( n1661 & ~n4296 ) | ( n1661 & n4432 ) | ( ~n4296 & n4432 ) ;
  assign n4535 = n1661 & ~n4296 ;
  assign n4536 = ( n4301 & n4534 ) | ( n4301 & n4535 ) | ( n4534 & n4535 ) ;
  assign n4537 = ( ~n4301 & n4534 ) | ( ~n4301 & n4535 ) | ( n4534 & n4535 ) ;
  assign n4538 = ( n4301 & ~n4536 ) | ( n4301 & n4537 ) | ( ~n4536 & n4537 ) ;
  assign n4539 = ( ~n1523 & n4533 ) | ( ~n1523 & n4538 ) | ( n4533 & n4538 ) ;
  assign n4540 = ( n1523 & ~n4302 ) | ( n1523 & n4432 ) | ( ~n4302 & n4432 ) ;
  assign n4541 = n1523 & ~n4302 ;
  assign n4542 = ( n4307 & n4540 ) | ( n4307 & n4541 ) | ( n4540 & n4541 ) ;
  assign n4543 = ( ~n4307 & n4540 ) | ( ~n4307 & n4541 ) | ( n4540 & n4541 ) ;
  assign n4544 = ( n4307 & ~n4542 ) | ( n4307 & n4543 ) | ( ~n4542 & n4543 ) ;
  assign n4545 = ( ~n1393 & n4539 ) | ( ~n1393 & n4544 ) | ( n4539 & n4544 ) ;
  assign n4546 = ~n1393 & n4308 ;
  assign n4547 = ( ~n1393 & n4308 ) | ( ~n1393 & n4432 ) | ( n4308 & n4432 ) ;
  assign n4548 = ( n4313 & n4546 ) | ( n4313 & n4547 ) | ( n4546 & n4547 ) ;
  assign n4549 = ( ~n4313 & n4546 ) | ( ~n4313 & n4547 ) | ( n4546 & n4547 ) ;
  assign n4550 = ( n4313 & ~n4548 ) | ( n4313 & n4549 ) | ( ~n4548 & n4549 ) ;
  assign n4551 = ( ~n1266 & n4545 ) | ( ~n1266 & n4550 ) | ( n4545 & n4550 ) ;
  assign n4552 = ( n1266 & ~n4314 ) | ( n1266 & n4432 ) | ( ~n4314 & n4432 ) ;
  assign n4553 = n1266 & ~n4314 ;
  assign n4554 = ( n4319 & n4552 ) | ( n4319 & n4553 ) | ( n4552 & n4553 ) ;
  assign n4555 = ( ~n4319 & n4552 ) | ( ~n4319 & n4553 ) | ( n4552 & n4553 ) ;
  assign n4556 = ( n4319 & ~n4554 ) | ( n4319 & n4555 ) | ( ~n4554 & n4555 ) ;
  assign n4557 = ( ~n1150 & n4551 ) | ( ~n1150 & n4556 ) | ( n4551 & n4556 ) ;
  assign n4558 = n1150 & ~n4320 ;
  assign n4559 = ( n1150 & ~n4320 ) | ( n1150 & n4432 ) | ( ~n4320 & n4432 ) ;
  assign n4560 = ( ~n4325 & n4558 ) | ( ~n4325 & n4559 ) | ( n4558 & n4559 ) ;
  assign n4561 = ( n4325 & n4558 ) | ( n4325 & n4559 ) | ( n4558 & n4559 ) ;
  assign n4562 = ( n4325 & n4560 ) | ( n4325 & ~n4561 ) | ( n4560 & ~n4561 ) ;
  assign n4563 = ( ~n1038 & n4557 ) | ( ~n1038 & n4562 ) | ( n4557 & n4562 ) ;
  assign n4564 = ( n1038 & ~n4326 ) | ( n1038 & n4432 ) | ( ~n4326 & n4432 ) ;
  assign n4565 = n1038 & ~n4326 ;
  assign n4566 = ( n4331 & n4564 ) | ( n4331 & n4565 ) | ( n4564 & n4565 ) ;
  assign n4567 = ( ~n4331 & n4564 ) | ( ~n4331 & n4565 ) | ( n4564 & n4565 ) ;
  assign n4568 = ( n4331 & ~n4566 ) | ( n4331 & n4567 ) | ( ~n4566 & n4567 ) ;
  assign n4569 = ( ~n933 & n4563 ) | ( ~n933 & n4568 ) | ( n4563 & n4568 ) ;
  assign n4570 = ( n933 & ~n4332 ) | ( n933 & n4432 ) | ( ~n4332 & n4432 ) ;
  assign n4571 = n933 & ~n4332 ;
  assign n4572 = ( n4337 & n4570 ) | ( n4337 & n4571 ) | ( n4570 & n4571 ) ;
  assign n4573 = ( ~n4337 & n4570 ) | ( ~n4337 & n4571 ) | ( n4570 & n4571 ) ;
  assign n4574 = ( n4337 & ~n4572 ) | ( n4337 & n4573 ) | ( ~n4572 & n4573 ) ;
  assign n4575 = ( ~n839 & n4569 ) | ( ~n839 & n4574 ) | ( n4569 & n4574 ) ;
  assign n4576 = ~n839 & n4338 ;
  assign n4577 = ( ~n839 & n4338 ) | ( ~n839 & n4432 ) | ( n4338 & n4432 ) ;
  assign n4578 = ( ~n4343 & n4576 ) | ( ~n4343 & n4577 ) | ( n4576 & n4577 ) ;
  assign n4579 = ( n4343 & n4576 ) | ( n4343 & n4577 ) | ( n4576 & n4577 ) ;
  assign n4580 = ( n4343 & n4578 ) | ( n4343 & ~n4579 ) | ( n4578 & ~n4579 ) ;
  assign n4581 = ( ~n746 & n4575 ) | ( ~n746 & n4580 ) | ( n4575 & n4580 ) ;
  assign n4582 = ~n746 & n4344 ;
  assign n4583 = ( ~n746 & n4344 ) | ( ~n746 & n4432 ) | ( n4344 & n4432 ) ;
  assign n4584 = ( ~n4349 & n4582 ) | ( ~n4349 & n4583 ) | ( n4582 & n4583 ) ;
  assign n4585 = ( n4349 & n4582 ) | ( n4349 & n4583 ) | ( n4582 & n4583 ) ;
  assign n4586 = ( n4349 & n4584 ) | ( n4349 & ~n4585 ) | ( n4584 & ~n4585 ) ;
  assign n4587 = ( ~n664 & n4581 ) | ( ~n664 & n4586 ) | ( n4581 & n4586 ) ;
  assign n4588 = ( n664 & ~n4350 ) | ( n664 & n4432 ) | ( ~n4350 & n4432 ) ;
  assign n4589 = n664 & ~n4350 ;
  assign n4590 = ( n4355 & n4588 ) | ( n4355 & n4589 ) | ( n4588 & n4589 ) ;
  assign n4591 = ( ~n4355 & n4588 ) | ( ~n4355 & n4589 ) | ( n4588 & n4589 ) ;
  assign n4592 = ( n4355 & ~n4590 ) | ( n4355 & n4591 ) | ( ~n4590 & n4591 ) ;
  assign n4593 = ( ~n588 & n4587 ) | ( ~n588 & n4592 ) | ( n4587 & n4592 ) ;
  assign n4594 = ( n588 & ~n4356 ) | ( n588 & n4432 ) | ( ~n4356 & n4432 ) ;
  assign n4595 = n588 & ~n4356 ;
  assign n4596 = ( n4361 & n4594 ) | ( n4361 & n4595 ) | ( n4594 & n4595 ) ;
  assign n4597 = ( ~n4361 & n4594 ) | ( ~n4361 & n4595 ) | ( n4594 & n4595 ) ;
  assign n4598 = ( n4361 & ~n4596 ) | ( n4361 & n4597 ) | ( ~n4596 & n4597 ) ;
  assign n4599 = ( ~n518 & n4593 ) | ( ~n518 & n4598 ) | ( n4593 & n4598 ) ;
  assign n4600 = ~n518 & n4362 ;
  assign n4601 = ( ~n518 & n4362 ) | ( ~n518 & n4432 ) | ( n4362 & n4432 ) ;
  assign n4602 = ( n4367 & n4600 ) | ( n4367 & n4601 ) | ( n4600 & n4601 ) ;
  assign n4603 = ( ~n4367 & n4600 ) | ( ~n4367 & n4601 ) | ( n4600 & n4601 ) ;
  assign n4604 = ( n4367 & ~n4602 ) | ( n4367 & n4603 ) | ( ~n4602 & n4603 ) ;
  assign n4605 = ( ~n454 & n4599 ) | ( ~n454 & n4604 ) | ( n4599 & n4604 ) ;
  assign n4606 = ( n454 & ~n4368 ) | ( n454 & n4432 ) | ( ~n4368 & n4432 ) ;
  assign n4607 = n454 & ~n4368 ;
  assign n4608 = ( n4373 & n4606 ) | ( n4373 & n4607 ) | ( n4606 & n4607 ) ;
  assign n4609 = ( ~n4373 & n4606 ) | ( ~n4373 & n4607 ) | ( n4606 & n4607 ) ;
  assign n4610 = ( n4373 & ~n4608 ) | ( n4373 & n4609 ) | ( ~n4608 & n4609 ) ;
  assign n4611 = ( ~n396 & n4605 ) | ( ~n396 & n4610 ) | ( n4605 & n4610 ) ;
  assign n4612 = ~n396 & n4374 ;
  assign n4613 = ( ~n396 & n4374 ) | ( ~n396 & n4432 ) | ( n4374 & n4432 ) ;
  assign n4614 = ( ~n4379 & n4612 ) | ( ~n4379 & n4613 ) | ( n4612 & n4613 ) ;
  assign n4615 = ( n4379 & n4612 ) | ( n4379 & n4613 ) | ( n4612 & n4613 ) ;
  assign n4616 = ( n4379 & n4614 ) | ( n4379 & ~n4615 ) | ( n4614 & ~n4615 ) ;
  assign n4617 = ( ~n344 & n4611 ) | ( ~n344 & n4616 ) | ( n4611 & n4616 ) ;
  assign n4618 = ( n344 & ~n4380 ) | ( n344 & n4432 ) | ( ~n4380 & n4432 ) ;
  assign n4619 = n344 & ~n4380 ;
  assign n4620 = ( n4385 & n4618 ) | ( n4385 & n4619 ) | ( n4618 & n4619 ) ;
  assign n4621 = ( ~n4385 & n4618 ) | ( ~n4385 & n4619 ) | ( n4618 & n4619 ) ;
  assign n4622 = ( n4385 & ~n4620 ) | ( n4385 & n4621 ) | ( ~n4620 & n4621 ) ;
  assign n4623 = ( ~n298 & n4617 ) | ( ~n298 & n4622 ) | ( n4617 & n4622 ) ;
  assign n4624 = n298 & ~n4386 ;
  assign n4625 = ( n298 & ~n4386 ) | ( n298 & n4432 ) | ( ~n4386 & n4432 ) ;
  assign n4626 = ( n4391 & n4624 ) | ( n4391 & n4625 ) | ( n4624 & n4625 ) ;
  assign n4627 = ( ~n4391 & n4624 ) | ( ~n4391 & n4625 ) | ( n4624 & n4625 ) ;
  assign n4628 = ( n4391 & ~n4626 ) | ( n4391 & n4627 ) | ( ~n4626 & n4627 ) ;
  assign n4629 = ( ~n258 & n4623 ) | ( ~n258 & n4628 ) | ( n4623 & n4628 ) ;
  assign n4630 = ~n258 & n4392 ;
  assign n4631 = ( ~n258 & n4392 ) | ( ~n258 & n4432 ) | ( n4392 & n4432 ) ;
  assign n4632 = ( n4397 & n4630 ) | ( n4397 & n4631 ) | ( n4630 & n4631 ) ;
  assign n4633 = ( ~n4397 & n4630 ) | ( ~n4397 & n4631 ) | ( n4630 & n4631 ) ;
  assign n4634 = ( n4397 & ~n4632 ) | ( n4397 & n4633 ) | ( ~n4632 & n4633 ) ;
  assign n4635 = ( ~n225 & n4629 ) | ( ~n225 & n4634 ) | ( n4629 & n4634 ) ;
  assign n4636 = ( n225 & ~n4398 ) | ( n225 & n4432 ) | ( ~n4398 & n4432 ) ;
  assign n4637 = n225 & ~n4398 ;
  assign n4638 = ( n4403 & n4636 ) | ( n4403 & n4637 ) | ( n4636 & n4637 ) ;
  assign n4639 = ( ~n4403 & n4636 ) | ( ~n4403 & n4637 ) | ( n4636 & n4637 ) ;
  assign n4640 = ( n4403 & ~n4638 ) | ( n4403 & n4639 ) | ( ~n4638 & n4639 ) ;
  assign n4641 = ( ~n197 & n4635 ) | ( ~n197 & n4640 ) | ( n4635 & n4640 ) ;
  assign n4642 = ~n197 & n4404 ;
  assign n4643 = ( ~n197 & n4404 ) | ( ~n197 & n4432 ) | ( n4404 & n4432 ) ;
  assign n4644 = ( ~n4409 & n4642 ) | ( ~n4409 & n4643 ) | ( n4642 & n4643 ) ;
  assign n4645 = ( n4409 & n4642 ) | ( n4409 & n4643 ) | ( n4642 & n4643 ) ;
  assign n4646 = ( n4409 & n4644 ) | ( n4409 & ~n4645 ) | ( n4644 & ~n4645 ) ;
  assign n4647 = ( ~n170 & n4641 ) | ( ~n170 & n4646 ) | ( n4641 & n4646 ) ;
  assign n4648 = ( n170 & ~n4410 ) | ( n170 & n4432 ) | ( ~n4410 & n4432 ) ;
  assign n4649 = n170 & ~n4410 ;
  assign n4650 = ( n4415 & n4648 ) | ( n4415 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4651 = ( ~n4415 & n4648 ) | ( ~n4415 & n4649 ) | ( n4648 & n4649 ) ;
  assign n4652 = ( n4415 & ~n4650 ) | ( n4415 & n4651 ) | ( ~n4650 & n4651 ) ;
  assign n4653 = ( ~n142 & n4647 ) | ( ~n142 & n4652 ) | ( n4647 & n4652 ) ;
  assign n4654 = ( n142 & ~n4416 ) | ( n142 & n4432 ) | ( ~n4416 & n4432 ) ;
  assign n4655 = n142 & ~n4416 ;
  assign n4656 = ( n4421 & n4654 ) | ( n4421 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4657 = ( ~n4421 & n4654 ) | ( ~n4421 & n4655 ) | ( n4654 & n4655 ) ;
  assign n4658 = ( n4421 & ~n4656 ) | ( n4421 & n4657 ) | ( ~n4656 & n4657 ) ;
  assign n4659 = ( ~n132 & n4653 ) | ( ~n132 & n4658 ) | ( n4653 & n4658 ) ;
  assign n4660 = ( ~n131 & n4443 ) | ( ~n131 & n4659 ) | ( n4443 & n4659 ) ;
  assign n4661 = n4438 | n4660 ;
  assign n4662 = ( n4433 & ~n4435 ) | ( n4433 & n4443 ) | ( ~n4435 & n4443 ) ;
  assign n4663 = ( n4443 & n4659 ) | ( n4443 & n4662 ) | ( n4659 & n4662 ) ;
  assign n4664 = ~n4660 & n4663 ;
  assign n4665 = ( n132 & ~n4653 ) | ( n132 & n4661 ) | ( ~n4653 & n4661 ) ;
  assign n4666 = n132 & ~n4653 ;
  assign n4667 = ( n4658 & n4665 ) | ( n4658 & n4666 ) | ( n4665 & n4666 ) ;
  assign n4668 = ( n4658 & ~n4665 ) | ( n4658 & n4666 ) | ( ~n4665 & n4666 ) ;
  assign n4669 = ( n4665 & ~n4667 ) | ( n4665 & n4668 ) | ( ~n4667 & n4668 ) ;
  assign n4670 = x48 | x49 ;
  assign n4671 = x50 | n4670 ;
  assign n4672 = n4432 & ~n4671 ;
  assign n4673 = ~n4444 & n4661 ;
  assign n4674 = ~n4432 & n4671 ;
  assign n4675 = ( x51 & ~n4661 ) | ( x51 & n4674 ) | ( ~n4661 & n4674 ) ;
  assign n4676 = ( ~n4672 & n4673 ) | ( ~n4672 & n4675 ) | ( n4673 & n4675 ) ;
  assign n4677 = n4432 & ~n4661 ;
  assign n4678 = ( x52 & n4673 ) | ( x52 & n4677 ) | ( n4673 & n4677 ) ;
  assign n4679 = ( ~x52 & n4673 ) | ( ~x52 & n4677 ) | ( n4673 & n4677 ) ;
  assign n4680 = ( x52 & ~n4678 ) | ( x52 & n4679 ) | ( ~n4678 & n4679 ) ;
  assign n4681 = ( ~n4203 & n4676 ) | ( ~n4203 & n4680 ) | ( n4676 & n4680 ) ;
  assign n4682 = ~n4203 & n4432 ;
  assign n4683 = ( n4451 & n4661 ) | ( n4451 & n4682 ) | ( n4661 & n4682 ) ;
  assign n4684 = ( ~x53 & n4679 ) | ( ~x53 & n4683 ) | ( n4679 & n4683 ) ;
  assign n4685 = ( x53 & n4679 ) | ( x53 & n4683 ) | ( n4679 & n4683 ) ;
  assign n4686 = ( x53 & n4684 ) | ( x53 & ~n4685 ) | ( n4684 & ~n4685 ) ;
  assign n4687 = ( ~n3985 & n4681 ) | ( ~n3985 & n4686 ) | ( n4681 & n4686 ) ;
  assign n4688 = n3985 & ~n4450 ;
  assign n4689 = ( n3985 & ~n4450 ) | ( n3985 & n4661 ) | ( ~n4450 & n4661 ) ;
  assign n4690 = ( n4454 & n4688 ) | ( n4454 & n4689 ) | ( n4688 & n4689 ) ;
  assign n4691 = ( ~n4454 & n4688 ) | ( ~n4454 & n4689 ) | ( n4688 & n4689 ) ;
  assign n4692 = ( n4454 & ~n4690 ) | ( n4454 & n4691 ) | ( ~n4690 & n4691 ) ;
  assign n4693 = ( ~n3772 & n4687 ) | ( ~n3772 & n4692 ) | ( n4687 & n4692 ) ;
  assign n4694 = ( n3772 & ~n4455 ) | ( n3772 & n4661 ) | ( ~n4455 & n4661 ) ;
  assign n4695 = n3772 & ~n4455 ;
  assign n4696 = ( n4460 & n4694 ) | ( n4460 & n4695 ) | ( n4694 & n4695 ) ;
  assign n4697 = ( ~n4460 & n4694 ) | ( ~n4460 & n4695 ) | ( n4694 & n4695 ) ;
  assign n4698 = ( n4460 & ~n4696 ) | ( n4460 & n4697 ) | ( ~n4696 & n4697 ) ;
  assign n4699 = ( ~n3567 & n4693 ) | ( ~n3567 & n4698 ) | ( n4693 & n4698 ) ;
  assign n4700 = ~n3567 & n4461 ;
  assign n4701 = ( ~n3567 & n4461 ) | ( ~n3567 & n4661 ) | ( n4461 & n4661 ) ;
  assign n4702 = ( ~n4466 & n4700 ) | ( ~n4466 & n4701 ) | ( n4700 & n4701 ) ;
  assign n4703 = ( n4466 & n4700 ) | ( n4466 & n4701 ) | ( n4700 & n4701 ) ;
  assign n4704 = ( n4466 & n4702 ) | ( n4466 & ~n4703 ) | ( n4702 & ~n4703 ) ;
  assign n4705 = ( ~n3362 & n4699 ) | ( ~n3362 & n4704 ) | ( n4699 & n4704 ) ;
  assign n4706 = ( n3362 & ~n4467 ) | ( n3362 & n4661 ) | ( ~n4467 & n4661 ) ;
  assign n4707 = n3362 & ~n4467 ;
  assign n4708 = ( n4472 & n4706 ) | ( n4472 & n4707 ) | ( n4706 & n4707 ) ;
  assign n4709 = ( ~n4472 & n4706 ) | ( ~n4472 & n4707 ) | ( n4706 & n4707 ) ;
  assign n4710 = ( n4472 & ~n4708 ) | ( n4472 & n4709 ) | ( ~n4708 & n4709 ) ;
  assign n4711 = ( ~n3169 & n4705 ) | ( ~n3169 & n4710 ) | ( n4705 & n4710 ) ;
  assign n4712 = ( n3169 & ~n4473 ) | ( n3169 & n4661 ) | ( ~n4473 & n4661 ) ;
  assign n4713 = n3169 & ~n4473 ;
  assign n4714 = ( n4478 & n4712 ) | ( n4478 & n4713 ) | ( n4712 & n4713 ) ;
  assign n4715 = ( ~n4478 & n4712 ) | ( ~n4478 & n4713 ) | ( n4712 & n4713 ) ;
  assign n4716 = ( n4478 & ~n4714 ) | ( n4478 & n4715 ) | ( ~n4714 & n4715 ) ;
  assign n4717 = ( ~n2979 & n4711 ) | ( ~n2979 & n4716 ) | ( n4711 & n4716 ) ;
  assign n4718 = ( n2979 & ~n4479 ) | ( n2979 & n4661 ) | ( ~n4479 & n4661 ) ;
  assign n4719 = n2979 & ~n4479 ;
  assign n4720 = ( n4484 & n4718 ) | ( n4484 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4721 = ( ~n4484 & n4718 ) | ( ~n4484 & n4719 ) | ( n4718 & n4719 ) ;
  assign n4722 = ( n4484 & ~n4720 ) | ( n4484 & n4721 ) | ( ~n4720 & n4721 ) ;
  assign n4723 = ( ~n2791 & n4717 ) | ( ~n2791 & n4722 ) | ( n4717 & n4722 ) ;
  assign n4724 = ~n2791 & n4485 ;
  assign n4725 = ( ~n2791 & n4485 ) | ( ~n2791 & n4661 ) | ( n4485 & n4661 ) ;
  assign n4726 = ( n4490 & n4724 ) | ( n4490 & n4725 ) | ( n4724 & n4725 ) ;
  assign n4727 = ( ~n4490 & n4724 ) | ( ~n4490 & n4725 ) | ( n4724 & n4725 ) ;
  assign n4728 = ( n4490 & ~n4726 ) | ( n4490 & n4727 ) | ( ~n4726 & n4727 ) ;
  assign n4729 = ( ~n2615 & n4723 ) | ( ~n2615 & n4728 ) | ( n4723 & n4728 ) ;
  assign n4730 = ~n2615 & n4491 ;
  assign n4731 = ( ~n2615 & n4491 ) | ( ~n2615 & n4661 ) | ( n4491 & n4661 ) ;
  assign n4732 = ( ~n4496 & n4730 ) | ( ~n4496 & n4731 ) | ( n4730 & n4731 ) ;
  assign n4733 = ( n4496 & n4730 ) | ( n4496 & n4731 ) | ( n4730 & n4731 ) ;
  assign n4734 = ( n4496 & n4732 ) | ( n4496 & ~n4733 ) | ( n4732 & ~n4733 ) ;
  assign n4735 = ( ~n2443 & n4729 ) | ( ~n2443 & n4734 ) | ( n4729 & n4734 ) ;
  assign n4736 = ( n2443 & ~n4497 ) | ( n2443 & n4661 ) | ( ~n4497 & n4661 ) ;
  assign n4737 = n2443 & ~n4497 ;
  assign n4738 = ( n4502 & n4736 ) | ( n4502 & n4737 ) | ( n4736 & n4737 ) ;
  assign n4739 = ( ~n4502 & n4736 ) | ( ~n4502 & n4737 ) | ( n4736 & n4737 ) ;
  assign n4740 = ( n4502 & ~n4738 ) | ( n4502 & n4739 ) | ( ~n4738 & n4739 ) ;
  assign n4741 = ( ~n2277 & n4735 ) | ( ~n2277 & n4740 ) | ( n4735 & n4740 ) ;
  assign n4742 = ~n2277 & n4503 ;
  assign n4743 = ( ~n2277 & n4503 ) | ( ~n2277 & n4661 ) | ( n4503 & n4661 ) ;
  assign n4744 = ( ~n4508 & n4742 ) | ( ~n4508 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4745 = ( n4508 & n4742 ) | ( n4508 & n4743 ) | ( n4742 & n4743 ) ;
  assign n4746 = ( n4508 & n4744 ) | ( n4508 & ~n4745 ) | ( n4744 & ~n4745 ) ;
  assign n4747 = ( ~n2111 & n4741 ) | ( ~n2111 & n4746 ) | ( n4741 & n4746 ) ;
  assign n4748 = ~n2111 & n4509 ;
  assign n4749 = ( ~n2111 & n4509 ) | ( ~n2111 & n4661 ) | ( n4509 & n4661 ) ;
  assign n4750 = ( ~n4514 & n4748 ) | ( ~n4514 & n4749 ) | ( n4748 & n4749 ) ;
  assign n4751 = ( n4514 & n4748 ) | ( n4514 & n4749 ) | ( n4748 & n4749 ) ;
  assign n4752 = ( n4514 & n4750 ) | ( n4514 & ~n4751 ) | ( n4750 & ~n4751 ) ;
  assign n4753 = ( ~n1949 & n4747 ) | ( ~n1949 & n4752 ) | ( n4747 & n4752 ) ;
  assign n4754 = ( n1949 & ~n4515 ) | ( n1949 & n4661 ) | ( ~n4515 & n4661 ) ;
  assign n4755 = n1949 & ~n4515 ;
  assign n4756 = ( n4520 & n4754 ) | ( n4520 & n4755 ) | ( n4754 & n4755 ) ;
  assign n4757 = ( ~n4520 & n4754 ) | ( ~n4520 & n4755 ) | ( n4754 & n4755 ) ;
  assign n4758 = ( n4520 & ~n4756 ) | ( n4520 & n4757 ) | ( ~n4756 & n4757 ) ;
  assign n4759 = ( ~n1802 & n4753 ) | ( ~n1802 & n4758 ) | ( n4753 & n4758 ) ;
  assign n4760 = ( n1802 & ~n4521 ) | ( n1802 & n4661 ) | ( ~n4521 & n4661 ) ;
  assign n4761 = n1802 & ~n4521 ;
  assign n4762 = ( n4526 & n4760 ) | ( n4526 & n4761 ) | ( n4760 & n4761 ) ;
  assign n4763 = ( ~n4526 & n4760 ) | ( ~n4526 & n4761 ) | ( n4760 & n4761 ) ;
  assign n4764 = ( n4526 & ~n4762 ) | ( n4526 & n4763 ) | ( ~n4762 & n4763 ) ;
  assign n4765 = ( ~n1661 & n4759 ) | ( ~n1661 & n4764 ) | ( n4759 & n4764 ) ;
  assign n4766 = ( n1661 & ~n4527 ) | ( n1661 & n4661 ) | ( ~n4527 & n4661 ) ;
  assign n4767 = n1661 & ~n4527 ;
  assign n4768 = ( n4532 & n4766 ) | ( n4532 & n4767 ) | ( n4766 & n4767 ) ;
  assign n4769 = ( ~n4532 & n4766 ) | ( ~n4532 & n4767 ) | ( n4766 & n4767 ) ;
  assign n4770 = ( n4532 & ~n4768 ) | ( n4532 & n4769 ) | ( ~n4768 & n4769 ) ;
  assign n4771 = ( ~n1523 & n4765 ) | ( ~n1523 & n4770 ) | ( n4765 & n4770 ) ;
  assign n4772 = ( n1523 & ~n4533 ) | ( n1523 & n4661 ) | ( ~n4533 & n4661 ) ;
  assign n4773 = n1523 & ~n4533 ;
  assign n4774 = ( n4538 & n4772 ) | ( n4538 & n4773 ) | ( n4772 & n4773 ) ;
  assign n4775 = ( ~n4538 & n4772 ) | ( ~n4538 & n4773 ) | ( n4772 & n4773 ) ;
  assign n4776 = ( n4538 & ~n4774 ) | ( n4538 & n4775 ) | ( ~n4774 & n4775 ) ;
  assign n4777 = ( ~n1393 & n4771 ) | ( ~n1393 & n4776 ) | ( n4771 & n4776 ) ;
  assign n4778 = ~n1393 & n4539 ;
  assign n4779 = ( ~n1393 & n4539 ) | ( ~n1393 & n4661 ) | ( n4539 & n4661 ) ;
  assign n4780 = ( ~n4544 & n4778 ) | ( ~n4544 & n4779 ) | ( n4778 & n4779 ) ;
  assign n4781 = ( n4544 & n4778 ) | ( n4544 & n4779 ) | ( n4778 & n4779 ) ;
  assign n4782 = ( n4544 & n4780 ) | ( n4544 & ~n4781 ) | ( n4780 & ~n4781 ) ;
  assign n4783 = ( ~n1266 & n4777 ) | ( ~n1266 & n4782 ) | ( n4777 & n4782 ) ;
  assign n4784 = ( n1266 & ~n4545 ) | ( n1266 & n4661 ) | ( ~n4545 & n4661 ) ;
  assign n4785 = n1266 & ~n4545 ;
  assign n4786 = ( n4550 & n4784 ) | ( n4550 & n4785 ) | ( n4784 & n4785 ) ;
  assign n4787 = ( ~n4550 & n4784 ) | ( ~n4550 & n4785 ) | ( n4784 & n4785 ) ;
  assign n4788 = ( n4550 & ~n4786 ) | ( n4550 & n4787 ) | ( ~n4786 & n4787 ) ;
  assign n4789 = ( ~n1150 & n4783 ) | ( ~n1150 & n4788 ) | ( n4783 & n4788 ) ;
  assign n4790 = ( n1150 & ~n4551 ) | ( n1150 & n4661 ) | ( ~n4551 & n4661 ) ;
  assign n4791 = n1150 & ~n4551 ;
  assign n4792 = ( n4556 & n4790 ) | ( n4556 & n4791 ) | ( n4790 & n4791 ) ;
  assign n4793 = ( ~n4556 & n4790 ) | ( ~n4556 & n4791 ) | ( n4790 & n4791 ) ;
  assign n4794 = ( n4556 & ~n4792 ) | ( n4556 & n4793 ) | ( ~n4792 & n4793 ) ;
  assign n4795 = ( ~n1038 & n4789 ) | ( ~n1038 & n4794 ) | ( n4789 & n4794 ) ;
  assign n4796 = ~n1038 & n4557 ;
  assign n4797 = ( ~n1038 & n4557 ) | ( ~n1038 & n4661 ) | ( n4557 & n4661 ) ;
  assign n4798 = ( ~n4562 & n4796 ) | ( ~n4562 & n4797 ) | ( n4796 & n4797 ) ;
  assign n4799 = ( n4562 & n4796 ) | ( n4562 & n4797 ) | ( n4796 & n4797 ) ;
  assign n4800 = ( n4562 & n4798 ) | ( n4562 & ~n4799 ) | ( n4798 & ~n4799 ) ;
  assign n4801 = ( ~n933 & n4795 ) | ( ~n933 & n4800 ) | ( n4795 & n4800 ) ;
  assign n4802 = ( n933 & ~n4563 ) | ( n933 & n4661 ) | ( ~n4563 & n4661 ) ;
  assign n4803 = n933 & ~n4563 ;
  assign n4804 = ( n4568 & n4802 ) | ( n4568 & n4803 ) | ( n4802 & n4803 ) ;
  assign n4805 = ( ~n4568 & n4802 ) | ( ~n4568 & n4803 ) | ( n4802 & n4803 ) ;
  assign n4806 = ( n4568 & ~n4804 ) | ( n4568 & n4805 ) | ( ~n4804 & n4805 ) ;
  assign n4807 = ( ~n839 & n4801 ) | ( ~n839 & n4806 ) | ( n4801 & n4806 ) ;
  assign n4808 = ( n839 & ~n4569 ) | ( n839 & n4661 ) | ( ~n4569 & n4661 ) ;
  assign n4809 = n839 & ~n4569 ;
  assign n4810 = ( n4574 & n4808 ) | ( n4574 & n4809 ) | ( n4808 & n4809 ) ;
  assign n4811 = ( ~n4574 & n4808 ) | ( ~n4574 & n4809 ) | ( n4808 & n4809 ) ;
  assign n4812 = ( n4574 & ~n4810 ) | ( n4574 & n4811 ) | ( ~n4810 & n4811 ) ;
  assign n4813 = ( ~n746 & n4807 ) | ( ~n746 & n4812 ) | ( n4807 & n4812 ) ;
  assign n4814 = ~n746 & n4575 ;
  assign n4815 = ( ~n746 & n4575 ) | ( ~n746 & n4661 ) | ( n4575 & n4661 ) ;
  assign n4816 = ( ~n4580 & n4814 ) | ( ~n4580 & n4815 ) | ( n4814 & n4815 ) ;
  assign n4817 = ( n4580 & n4814 ) | ( n4580 & n4815 ) | ( n4814 & n4815 ) ;
  assign n4818 = ( n4580 & n4816 ) | ( n4580 & ~n4817 ) | ( n4816 & ~n4817 ) ;
  assign n4819 = ( ~n664 & n4813 ) | ( ~n664 & n4818 ) | ( n4813 & n4818 ) ;
  assign n4820 = ~n664 & n4581 ;
  assign n4821 = ( ~n664 & n4581 ) | ( ~n664 & n4661 ) | ( n4581 & n4661 ) ;
  assign n4822 = ( n4586 & n4820 ) | ( n4586 & n4821 ) | ( n4820 & n4821 ) ;
  assign n4823 = ( ~n4586 & n4820 ) | ( ~n4586 & n4821 ) | ( n4820 & n4821 ) ;
  assign n4824 = ( n4586 & ~n4822 ) | ( n4586 & n4823 ) | ( ~n4822 & n4823 ) ;
  assign n4825 = ( ~n588 & n4819 ) | ( ~n588 & n4824 ) | ( n4819 & n4824 ) ;
  assign n4826 = ( n588 & ~n4587 ) | ( n588 & n4661 ) | ( ~n4587 & n4661 ) ;
  assign n4827 = n588 & ~n4587 ;
  assign n4828 = ( n4592 & n4826 ) | ( n4592 & n4827 ) | ( n4826 & n4827 ) ;
  assign n4829 = ( ~n4592 & n4826 ) | ( ~n4592 & n4827 ) | ( n4826 & n4827 ) ;
  assign n4830 = ( n4592 & ~n4828 ) | ( n4592 & n4829 ) | ( ~n4828 & n4829 ) ;
  assign n4831 = ( ~n518 & n4825 ) | ( ~n518 & n4830 ) | ( n4825 & n4830 ) ;
  assign n4832 = ( n518 & ~n4593 ) | ( n518 & n4661 ) | ( ~n4593 & n4661 ) ;
  assign n4833 = n518 & ~n4593 ;
  assign n4834 = ( n4598 & n4832 ) | ( n4598 & n4833 ) | ( n4832 & n4833 ) ;
  assign n4835 = ( ~n4598 & n4832 ) | ( ~n4598 & n4833 ) | ( n4832 & n4833 ) ;
  assign n4836 = ( n4598 & ~n4834 ) | ( n4598 & n4835 ) | ( ~n4834 & n4835 ) ;
  assign n4837 = ( ~n454 & n4831 ) | ( ~n454 & n4836 ) | ( n4831 & n4836 ) ;
  assign n4838 = ( n454 & ~n4599 ) | ( n454 & n4661 ) | ( ~n4599 & n4661 ) ;
  assign n4839 = n454 & ~n4599 ;
  assign n4840 = ( n4604 & n4838 ) | ( n4604 & n4839 ) | ( n4838 & n4839 ) ;
  assign n4841 = ( ~n4604 & n4838 ) | ( ~n4604 & n4839 ) | ( n4838 & n4839 ) ;
  assign n4842 = ( n4604 & ~n4840 ) | ( n4604 & n4841 ) | ( ~n4840 & n4841 ) ;
  assign n4843 = ( ~n396 & n4837 ) | ( ~n396 & n4842 ) | ( n4837 & n4842 ) ;
  assign n4844 = ( n396 & ~n4605 ) | ( n396 & n4661 ) | ( ~n4605 & n4661 ) ;
  assign n4845 = n396 & ~n4605 ;
  assign n4846 = ( n4610 & n4844 ) | ( n4610 & n4845 ) | ( n4844 & n4845 ) ;
  assign n4847 = ( ~n4610 & n4844 ) | ( ~n4610 & n4845 ) | ( n4844 & n4845 ) ;
  assign n4848 = ( n4610 & ~n4846 ) | ( n4610 & n4847 ) | ( ~n4846 & n4847 ) ;
  assign n4849 = ( ~n344 & n4843 ) | ( ~n344 & n4848 ) | ( n4843 & n4848 ) ;
  assign n4850 = ( n344 & ~n4611 ) | ( n344 & n4661 ) | ( ~n4611 & n4661 ) ;
  assign n4851 = n344 & ~n4611 ;
  assign n4852 = ( n4616 & n4850 ) | ( n4616 & n4851 ) | ( n4850 & n4851 ) ;
  assign n4853 = ( ~n4616 & n4850 ) | ( ~n4616 & n4851 ) | ( n4850 & n4851 ) ;
  assign n4854 = ( n4616 & ~n4852 ) | ( n4616 & n4853 ) | ( ~n4852 & n4853 ) ;
  assign n4855 = ( ~n298 & n4849 ) | ( ~n298 & n4854 ) | ( n4849 & n4854 ) ;
  assign n4856 = ( n298 & ~n4617 ) | ( n298 & n4661 ) | ( ~n4617 & n4661 ) ;
  assign n4857 = n298 & ~n4617 ;
  assign n4858 = ( ~n4622 & n4856 ) | ( ~n4622 & n4857 ) | ( n4856 & n4857 ) ;
  assign n4859 = ( n4622 & n4856 ) | ( n4622 & n4857 ) | ( n4856 & n4857 ) ;
  assign n4860 = ( n4622 & n4858 ) | ( n4622 & ~n4859 ) | ( n4858 & ~n4859 ) ;
  assign n4861 = ( ~n258 & n4855 ) | ( ~n258 & n4860 ) | ( n4855 & n4860 ) ;
  assign n4862 = ( n258 & ~n4623 ) | ( n258 & n4661 ) | ( ~n4623 & n4661 ) ;
  assign n4863 = n258 & ~n4623 ;
  assign n4864 = ( n4628 & n4862 ) | ( n4628 & n4863 ) | ( n4862 & n4863 ) ;
  assign n4865 = ( ~n4628 & n4862 ) | ( ~n4628 & n4863 ) | ( n4862 & n4863 ) ;
  assign n4866 = ( n4628 & ~n4864 ) | ( n4628 & n4865 ) | ( ~n4864 & n4865 ) ;
  assign n4867 = ( ~n225 & n4861 ) | ( ~n225 & n4866 ) | ( n4861 & n4866 ) ;
  assign n4868 = ( n225 & ~n4629 ) | ( n225 & n4661 ) | ( ~n4629 & n4661 ) ;
  assign n4869 = n225 & ~n4629 ;
  assign n4870 = ( n4634 & n4868 ) | ( n4634 & n4869 ) | ( n4868 & n4869 ) ;
  assign n4871 = ( ~n4634 & n4868 ) | ( ~n4634 & n4869 ) | ( n4868 & n4869 ) ;
  assign n4872 = ( n4634 & ~n4870 ) | ( n4634 & n4871 ) | ( ~n4870 & n4871 ) ;
  assign n4873 = ( ~n197 & n4867 ) | ( ~n197 & n4872 ) | ( n4867 & n4872 ) ;
  assign n4874 = ~n197 & n4635 ;
  assign n4875 = ( ~n197 & n4635 ) | ( ~n197 & n4661 ) | ( n4635 & n4661 ) ;
  assign n4876 = ( ~n4640 & n4874 ) | ( ~n4640 & n4875 ) | ( n4874 & n4875 ) ;
  assign n4877 = ( n4640 & n4874 ) | ( n4640 & n4875 ) | ( n4874 & n4875 ) ;
  assign n4878 = ( n4640 & n4876 ) | ( n4640 & ~n4877 ) | ( n4876 & ~n4877 ) ;
  assign n4879 = ( ~n170 & n4873 ) | ( ~n170 & n4878 ) | ( n4873 & n4878 ) ;
  assign n4880 = ( n170 & ~n4641 ) | ( n170 & n4661 ) | ( ~n4641 & n4661 ) ;
  assign n4881 = n170 & ~n4641 ;
  assign n4882 = ( n4646 & n4880 ) | ( n4646 & n4881 ) | ( n4880 & n4881 ) ;
  assign n4883 = ( ~n4646 & n4880 ) | ( ~n4646 & n4881 ) | ( n4880 & n4881 ) ;
  assign n4884 = ( n4646 & ~n4882 ) | ( n4646 & n4883 ) | ( ~n4882 & n4883 ) ;
  assign n4885 = ( ~n142 & n4879 ) | ( ~n142 & n4884 ) | ( n4879 & n4884 ) ;
  assign n4886 = ( n142 & ~n4647 ) | ( n142 & n4661 ) | ( ~n4647 & n4661 ) ;
  assign n4887 = n142 & ~n4647 ;
  assign n4888 = ( n4652 & n4886 ) | ( n4652 & n4887 ) | ( n4886 & n4887 ) ;
  assign n4889 = ( ~n4652 & n4886 ) | ( ~n4652 & n4887 ) | ( n4886 & n4887 ) ;
  assign n4890 = ( n4652 & ~n4888 ) | ( n4652 & n4889 ) | ( ~n4888 & n4889 ) ;
  assign n4891 = ( ~n132 & n4885 ) | ( ~n132 & n4890 ) | ( n4885 & n4890 ) ;
  assign n4892 = n4443 & n4659 ;
  assign n4893 = n4438 & ~n4443 ;
  assign n4894 = ~n4659 & n4893 ;
  assign n4895 = ( ~n4669 & n4892 ) | ( ~n4669 & n4894 ) | ( n4892 & n4894 ) ;
  assign n4896 = n4891 | n4895 ;
  assign n4897 = ( ~n131 & n4669 ) | ( ~n131 & n4896 ) | ( n4669 & n4896 ) ;
  assign n4898 = n4664 | n4897 ;
  assign n4899 = ~n4670 & n4898 ;
  assign n4900 = x46 | x47 ;
  assign n4901 = x48 | n4900 ;
  assign n4902 = n4661 & ~n4901 ;
  assign n4903 = ~n4661 & n4901 ;
  assign n4904 = ( x49 & ~n4898 ) | ( x49 & n4903 ) | ( ~n4898 & n4903 ) ;
  assign n4905 = ( n4899 & ~n4902 ) | ( n4899 & n4904 ) | ( ~n4902 & n4904 ) ;
  assign n4906 = n4661 & ~n4898 ;
  assign n4907 = ( x50 & n4899 ) | ( x50 & n4906 ) | ( n4899 & n4906 ) ;
  assign n4908 = ( ~x50 & n4899 ) | ( ~x50 & n4906 ) | ( n4899 & n4906 ) ;
  assign n4909 = ( x50 & ~n4907 ) | ( x50 & n4908 ) | ( ~n4907 & n4908 ) ;
  assign n4910 = ( ~n4432 & n4905 ) | ( ~n4432 & n4909 ) | ( n4905 & n4909 ) ;
  assign n4911 = ~n4432 & n4661 ;
  assign n4912 = ( n4677 & n4898 ) | ( n4677 & n4911 ) | ( n4898 & n4911 ) ;
  assign n4913 = ( x51 & n4908 ) | ( x51 & n4912 ) | ( n4908 & n4912 ) ;
  assign n4914 = ( ~x51 & n4908 ) | ( ~x51 & n4912 ) | ( n4908 & n4912 ) ;
  assign n4915 = ( x51 & ~n4913 ) | ( x51 & n4914 ) | ( ~n4913 & n4914 ) ;
  assign n4916 = ( ~n4203 & n4910 ) | ( ~n4203 & n4915 ) | ( n4910 & n4915 ) ;
  assign n4917 = ( n4203 & ~n4676 ) | ( n4203 & n4898 ) | ( ~n4676 & n4898 ) ;
  assign n4918 = n4203 & ~n4676 ;
  assign n4919 = ( n4680 & n4917 ) | ( n4680 & n4918 ) | ( n4917 & n4918 ) ;
  assign n4920 = ( ~n4680 & n4917 ) | ( ~n4680 & n4918 ) | ( n4917 & n4918 ) ;
  assign n4921 = ( n4680 & ~n4919 ) | ( n4680 & n4920 ) | ( ~n4919 & n4920 ) ;
  assign n4922 = ( ~n3985 & n4916 ) | ( ~n3985 & n4921 ) | ( n4916 & n4921 ) ;
  assign n4923 = ~n3985 & n4681 ;
  assign n4924 = ( ~n3985 & n4681 ) | ( ~n3985 & n4898 ) | ( n4681 & n4898 ) ;
  assign n4925 = ( n4686 & n4923 ) | ( n4686 & n4924 ) | ( n4923 & n4924 ) ;
  assign n4926 = ( ~n4686 & n4923 ) | ( ~n4686 & n4924 ) | ( n4923 & n4924 ) ;
  assign n4927 = ( n4686 & ~n4925 ) | ( n4686 & n4926 ) | ( ~n4925 & n4926 ) ;
  assign n4928 = ( ~n3772 & n4922 ) | ( ~n3772 & n4927 ) | ( n4922 & n4927 ) ;
  assign n4929 = ( n3772 & ~n4687 ) | ( n3772 & n4898 ) | ( ~n4687 & n4898 ) ;
  assign n4930 = n3772 & ~n4687 ;
  assign n4931 = ( n4692 & n4929 ) | ( n4692 & n4930 ) | ( n4929 & n4930 ) ;
  assign n4932 = ( ~n4692 & n4929 ) | ( ~n4692 & n4930 ) | ( n4929 & n4930 ) ;
  assign n4933 = ( n4692 & ~n4931 ) | ( n4692 & n4932 ) | ( ~n4931 & n4932 ) ;
  assign n4934 = ( ~n3567 & n4928 ) | ( ~n3567 & n4933 ) | ( n4928 & n4933 ) ;
  assign n4935 = ~n3567 & n4693 ;
  assign n4936 = ( ~n3567 & n4693 ) | ( ~n3567 & n4898 ) | ( n4693 & n4898 ) ;
  assign n4937 = ( ~n4698 & n4935 ) | ( ~n4698 & n4936 ) | ( n4935 & n4936 ) ;
  assign n4938 = ( n4698 & n4935 ) | ( n4698 & n4936 ) | ( n4935 & n4936 ) ;
  assign n4939 = ( n4698 & n4937 ) | ( n4698 & ~n4938 ) | ( n4937 & ~n4938 ) ;
  assign n4940 = ( ~n3362 & n4934 ) | ( ~n3362 & n4939 ) | ( n4934 & n4939 ) ;
  assign n4941 = ~n3362 & n4699 ;
  assign n4942 = ( ~n3362 & n4699 ) | ( ~n3362 & n4898 ) | ( n4699 & n4898 ) ;
  assign n4943 = ( ~n4704 & n4941 ) | ( ~n4704 & n4942 ) | ( n4941 & n4942 ) ;
  assign n4944 = ( n4704 & n4941 ) | ( n4704 & n4942 ) | ( n4941 & n4942 ) ;
  assign n4945 = ( n4704 & n4943 ) | ( n4704 & ~n4944 ) | ( n4943 & ~n4944 ) ;
  assign n4946 = ( ~n3169 & n4940 ) | ( ~n3169 & n4945 ) | ( n4940 & n4945 ) ;
  assign n4947 = ( n3169 & ~n4705 ) | ( n3169 & n4898 ) | ( ~n4705 & n4898 ) ;
  assign n4948 = n3169 & ~n4705 ;
  assign n4949 = ( n4710 & n4947 ) | ( n4710 & n4948 ) | ( n4947 & n4948 ) ;
  assign n4950 = ( ~n4710 & n4947 ) | ( ~n4710 & n4948 ) | ( n4947 & n4948 ) ;
  assign n4951 = ( n4710 & ~n4949 ) | ( n4710 & n4950 ) | ( ~n4949 & n4950 ) ;
  assign n4952 = ( ~n2979 & n4946 ) | ( ~n2979 & n4951 ) | ( n4946 & n4951 ) ;
  assign n4953 = ( n2979 & ~n4711 ) | ( n2979 & n4898 ) | ( ~n4711 & n4898 ) ;
  assign n4954 = n2979 & ~n4711 ;
  assign n4955 = ( ~n4716 & n4953 ) | ( ~n4716 & n4954 ) | ( n4953 & n4954 ) ;
  assign n4956 = ( n4716 & n4953 ) | ( n4716 & n4954 ) | ( n4953 & n4954 ) ;
  assign n4957 = ( n4716 & n4955 ) | ( n4716 & ~n4956 ) | ( n4955 & ~n4956 ) ;
  assign n4958 = ( ~n2791 & n4952 ) | ( ~n2791 & n4957 ) | ( n4952 & n4957 ) ;
  assign n4959 = ( n2791 & ~n4717 ) | ( n2791 & n4898 ) | ( ~n4717 & n4898 ) ;
  assign n4960 = n2791 & ~n4717 ;
  assign n4961 = ( n4722 & n4959 ) | ( n4722 & n4960 ) | ( n4959 & n4960 ) ;
  assign n4962 = ( ~n4722 & n4959 ) | ( ~n4722 & n4960 ) | ( n4959 & n4960 ) ;
  assign n4963 = ( n4722 & ~n4961 ) | ( n4722 & n4962 ) | ( ~n4961 & n4962 ) ;
  assign n4964 = ( ~n2615 & n4958 ) | ( ~n2615 & n4963 ) | ( n4958 & n4963 ) ;
  assign n4965 = ( n2615 & ~n4723 ) | ( n2615 & n4898 ) | ( ~n4723 & n4898 ) ;
  assign n4966 = n2615 & ~n4723 ;
  assign n4967 = ( n4728 & n4965 ) | ( n4728 & n4966 ) | ( n4965 & n4966 ) ;
  assign n4968 = ( ~n4728 & n4965 ) | ( ~n4728 & n4966 ) | ( n4965 & n4966 ) ;
  assign n4969 = ( n4728 & ~n4967 ) | ( n4728 & n4968 ) | ( ~n4967 & n4968 ) ;
  assign n4970 = ( ~n2443 & n4964 ) | ( ~n2443 & n4969 ) | ( n4964 & n4969 ) ;
  assign n4971 = ( ~n2443 & n4729 ) | ( ~n2443 & n4898 ) | ( n4729 & n4898 ) ;
  assign n4972 = ~n2443 & n4729 ;
  assign n4973 = ( ~n4734 & n4971 ) | ( ~n4734 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4974 = ( n4734 & n4971 ) | ( n4734 & n4972 ) | ( n4971 & n4972 ) ;
  assign n4975 = ( n4734 & n4973 ) | ( n4734 & ~n4974 ) | ( n4973 & ~n4974 ) ;
  assign n4976 = ( ~n2277 & n4970 ) | ( ~n2277 & n4975 ) | ( n4970 & n4975 ) ;
  assign n4977 = ~n2277 & n4735 ;
  assign n4978 = ( ~n2277 & n4735 ) | ( ~n2277 & n4898 ) | ( n4735 & n4898 ) ;
  assign n4979 = ( ~n4740 & n4977 ) | ( ~n4740 & n4978 ) | ( n4977 & n4978 ) ;
  assign n4980 = ( n4740 & n4977 ) | ( n4740 & n4978 ) | ( n4977 & n4978 ) ;
  assign n4981 = ( n4740 & n4979 ) | ( n4740 & ~n4980 ) | ( n4979 & ~n4980 ) ;
  assign n4982 = ( ~n2111 & n4976 ) | ( ~n2111 & n4981 ) | ( n4976 & n4981 ) ;
  assign n4983 = ~n2111 & n4741 ;
  assign n4984 = ( ~n2111 & n4741 ) | ( ~n2111 & n4898 ) | ( n4741 & n4898 ) ;
  assign n4985 = ( n4746 & n4983 ) | ( n4746 & n4984 ) | ( n4983 & n4984 ) ;
  assign n4986 = ( ~n4746 & n4983 ) | ( ~n4746 & n4984 ) | ( n4983 & n4984 ) ;
  assign n4987 = ( n4746 & ~n4985 ) | ( n4746 & n4986 ) | ( ~n4985 & n4986 ) ;
  assign n4988 = ( ~n1949 & n4982 ) | ( ~n1949 & n4987 ) | ( n4982 & n4987 ) ;
  assign n4989 = ( n1949 & ~n4747 ) | ( n1949 & n4898 ) | ( ~n4747 & n4898 ) ;
  assign n4990 = n1949 & ~n4747 ;
  assign n4991 = ( n4752 & n4989 ) | ( n4752 & n4990 ) | ( n4989 & n4990 ) ;
  assign n4992 = ( ~n4752 & n4989 ) | ( ~n4752 & n4990 ) | ( n4989 & n4990 ) ;
  assign n4993 = ( n4752 & ~n4991 ) | ( n4752 & n4992 ) | ( ~n4991 & n4992 ) ;
  assign n4994 = ( ~n1802 & n4988 ) | ( ~n1802 & n4993 ) | ( n4988 & n4993 ) ;
  assign n4995 = ~n1802 & n4753 ;
  assign n4996 = ( ~n1802 & n4753 ) | ( ~n1802 & n4898 ) | ( n4753 & n4898 ) ;
  assign n4997 = ( n4758 & n4995 ) | ( n4758 & n4996 ) | ( n4995 & n4996 ) ;
  assign n4998 = ( ~n4758 & n4995 ) | ( ~n4758 & n4996 ) | ( n4995 & n4996 ) ;
  assign n4999 = ( n4758 & ~n4997 ) | ( n4758 & n4998 ) | ( ~n4997 & n4998 ) ;
  assign n5000 = ( ~n1661 & n4994 ) | ( ~n1661 & n4999 ) | ( n4994 & n4999 ) ;
  assign n5001 = ( n1661 & ~n4759 ) | ( n1661 & n4898 ) | ( ~n4759 & n4898 ) ;
  assign n5002 = n1661 & ~n4759 ;
  assign n5003 = ( n4764 & n5001 ) | ( n4764 & n5002 ) | ( n5001 & n5002 ) ;
  assign n5004 = ( ~n4764 & n5001 ) | ( ~n4764 & n5002 ) | ( n5001 & n5002 ) ;
  assign n5005 = ( n4764 & ~n5003 ) | ( n4764 & n5004 ) | ( ~n5003 & n5004 ) ;
  assign n5006 = ( ~n1523 & n5000 ) | ( ~n1523 & n5005 ) | ( n5000 & n5005 ) ;
  assign n5007 = ~n1523 & n4765 ;
  assign n5008 = ( ~n1523 & n4765 ) | ( ~n1523 & n4898 ) | ( n4765 & n4898 ) ;
  assign n5009 = ( n4770 & n5007 ) | ( n4770 & n5008 ) | ( n5007 & n5008 ) ;
  assign n5010 = ( ~n4770 & n5007 ) | ( ~n4770 & n5008 ) | ( n5007 & n5008 ) ;
  assign n5011 = ( n4770 & ~n5009 ) | ( n4770 & n5010 ) | ( ~n5009 & n5010 ) ;
  assign n5012 = ( ~n1393 & n5006 ) | ( ~n1393 & n5011 ) | ( n5006 & n5011 ) ;
  assign n5013 = ~n1393 & n4771 ;
  assign n5014 = ( ~n1393 & n4771 ) | ( ~n1393 & n4898 ) | ( n4771 & n4898 ) ;
  assign n5015 = ( n4776 & n5013 ) | ( n4776 & n5014 ) | ( n5013 & n5014 ) ;
  assign n5016 = ( ~n4776 & n5013 ) | ( ~n4776 & n5014 ) | ( n5013 & n5014 ) ;
  assign n5017 = ( n4776 & ~n5015 ) | ( n4776 & n5016 ) | ( ~n5015 & n5016 ) ;
  assign n5018 = ( ~n1266 & n5012 ) | ( ~n1266 & n5017 ) | ( n5012 & n5017 ) ;
  assign n5019 = ~n1266 & n4777 ;
  assign n5020 = ( ~n1266 & n4777 ) | ( ~n1266 & n4898 ) | ( n4777 & n4898 ) ;
  assign n5021 = ( ~n4782 & n5019 ) | ( ~n4782 & n5020 ) | ( n5019 & n5020 ) ;
  assign n5022 = ( n4782 & n5019 ) | ( n4782 & n5020 ) | ( n5019 & n5020 ) ;
  assign n5023 = ( n4782 & n5021 ) | ( n4782 & ~n5022 ) | ( n5021 & ~n5022 ) ;
  assign n5024 = ( ~n1150 & n5018 ) | ( ~n1150 & n5023 ) | ( n5018 & n5023 ) ;
  assign n5025 = ~n1150 & n4783 ;
  assign n5026 = ( ~n1150 & n4783 ) | ( ~n1150 & n4898 ) | ( n4783 & n4898 ) ;
  assign n5027 = ( n4788 & n5025 ) | ( n4788 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5028 = ( ~n4788 & n5025 ) | ( ~n4788 & n5026 ) | ( n5025 & n5026 ) ;
  assign n5029 = ( n4788 & ~n5027 ) | ( n4788 & n5028 ) | ( ~n5027 & n5028 ) ;
  assign n5030 = ( ~n1038 & n5024 ) | ( ~n1038 & n5029 ) | ( n5024 & n5029 ) ;
  assign n5031 = ( n1038 & ~n4789 ) | ( n1038 & n4898 ) | ( ~n4789 & n4898 ) ;
  assign n5032 = n1038 & ~n4789 ;
  assign n5033 = ( n4794 & n5031 ) | ( n4794 & n5032 ) | ( n5031 & n5032 ) ;
  assign n5034 = ( ~n4794 & n5031 ) | ( ~n4794 & n5032 ) | ( n5031 & n5032 ) ;
  assign n5035 = ( n4794 & ~n5033 ) | ( n4794 & n5034 ) | ( ~n5033 & n5034 ) ;
  assign n5036 = ( ~n933 & n5030 ) | ( ~n933 & n5035 ) | ( n5030 & n5035 ) ;
  assign n5037 = ( n933 & ~n4795 ) | ( n933 & n4898 ) | ( ~n4795 & n4898 ) ;
  assign n5038 = n933 & ~n4795 ;
  assign n5039 = ( n4800 & n5037 ) | ( n4800 & n5038 ) | ( n5037 & n5038 ) ;
  assign n5040 = ( ~n4800 & n5037 ) | ( ~n4800 & n5038 ) | ( n5037 & n5038 ) ;
  assign n5041 = ( n4800 & ~n5039 ) | ( n4800 & n5040 ) | ( ~n5039 & n5040 ) ;
  assign n5042 = ( ~n839 & n5036 ) | ( ~n839 & n5041 ) | ( n5036 & n5041 ) ;
  assign n5043 = ( n839 & ~n4801 ) | ( n839 & n4898 ) | ( ~n4801 & n4898 ) ;
  assign n5044 = n839 & ~n4801 ;
  assign n5045 = ( n4806 & n5043 ) | ( n4806 & n5044 ) | ( n5043 & n5044 ) ;
  assign n5046 = ( ~n4806 & n5043 ) | ( ~n4806 & n5044 ) | ( n5043 & n5044 ) ;
  assign n5047 = ( n4806 & ~n5045 ) | ( n4806 & n5046 ) | ( ~n5045 & n5046 ) ;
  assign n5048 = ( ~n746 & n5042 ) | ( ~n746 & n5047 ) | ( n5042 & n5047 ) ;
  assign n5049 = n746 & ~n4807 ;
  assign n5050 = ( n746 & ~n4807 ) | ( n746 & n4898 ) | ( ~n4807 & n4898 ) ;
  assign n5051 = ( ~n4812 & n5049 ) | ( ~n4812 & n5050 ) | ( n5049 & n5050 ) ;
  assign n5052 = ( n4812 & n5049 ) | ( n4812 & n5050 ) | ( n5049 & n5050 ) ;
  assign n5053 = ( n4812 & n5051 ) | ( n4812 & ~n5052 ) | ( n5051 & ~n5052 ) ;
  assign n5054 = ( ~n664 & n5048 ) | ( ~n664 & n5053 ) | ( n5048 & n5053 ) ;
  assign n5055 = ( n664 & ~n4813 ) | ( n664 & n4898 ) | ( ~n4813 & n4898 ) ;
  assign n5056 = n664 & ~n4813 ;
  assign n5057 = ( n4818 & n5055 ) | ( n4818 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5058 = ( ~n4818 & n5055 ) | ( ~n4818 & n5056 ) | ( n5055 & n5056 ) ;
  assign n5059 = ( n4818 & ~n5057 ) | ( n4818 & n5058 ) | ( ~n5057 & n5058 ) ;
  assign n5060 = ( ~n588 & n5054 ) | ( ~n588 & n5059 ) | ( n5054 & n5059 ) ;
  assign n5061 = ( n588 & ~n4819 ) | ( n588 & n4898 ) | ( ~n4819 & n4898 ) ;
  assign n5062 = n588 & ~n4819 ;
  assign n5063 = ( n4824 & n5061 ) | ( n4824 & n5062 ) | ( n5061 & n5062 ) ;
  assign n5064 = ( ~n4824 & n5061 ) | ( ~n4824 & n5062 ) | ( n5061 & n5062 ) ;
  assign n5065 = ( n4824 & ~n5063 ) | ( n4824 & n5064 ) | ( ~n5063 & n5064 ) ;
  assign n5066 = ( ~n518 & n5060 ) | ( ~n518 & n5065 ) | ( n5060 & n5065 ) ;
  assign n5067 = ~n518 & n4825 ;
  assign n5068 = ( ~n518 & n4825 ) | ( ~n518 & n4898 ) | ( n4825 & n4898 ) ;
  assign n5069 = ( ~n4830 & n5067 ) | ( ~n4830 & n5068 ) | ( n5067 & n5068 ) ;
  assign n5070 = ( n4830 & n5067 ) | ( n4830 & n5068 ) | ( n5067 & n5068 ) ;
  assign n5071 = ( n4830 & n5069 ) | ( n4830 & ~n5070 ) | ( n5069 & ~n5070 ) ;
  assign n5072 = ( ~n454 & n5066 ) | ( ~n454 & n5071 ) | ( n5066 & n5071 ) ;
  assign n5073 = ~n454 & n4831 ;
  assign n5074 = ( ~n454 & n4831 ) | ( ~n454 & n4898 ) | ( n4831 & n4898 ) ;
  assign n5075 = ( n4836 & n5073 ) | ( n4836 & n5074 ) | ( n5073 & n5074 ) ;
  assign n5076 = ( ~n4836 & n5073 ) | ( ~n4836 & n5074 ) | ( n5073 & n5074 ) ;
  assign n5077 = ( n4836 & ~n5075 ) | ( n4836 & n5076 ) | ( ~n5075 & n5076 ) ;
  assign n5078 = ( ~n396 & n5072 ) | ( ~n396 & n5077 ) | ( n5072 & n5077 ) ;
  assign n5079 = ( n396 & ~n4837 ) | ( n396 & n4898 ) | ( ~n4837 & n4898 ) ;
  assign n5080 = n396 & ~n4837 ;
  assign n5081 = ( n4842 & n5079 ) | ( n4842 & n5080 ) | ( n5079 & n5080 ) ;
  assign n5082 = ( ~n4842 & n5079 ) | ( ~n4842 & n5080 ) | ( n5079 & n5080 ) ;
  assign n5083 = ( n4842 & ~n5081 ) | ( n4842 & n5082 ) | ( ~n5081 & n5082 ) ;
  assign n5084 = ( ~n344 & n5078 ) | ( ~n344 & n5083 ) | ( n5078 & n5083 ) ;
  assign n5085 = ( n344 & ~n4843 ) | ( n344 & n4898 ) | ( ~n4843 & n4898 ) ;
  assign n5086 = n344 & ~n4843 ;
  assign n5087 = ( n4848 & n5085 ) | ( n4848 & n5086 ) | ( n5085 & n5086 ) ;
  assign n5088 = ( ~n4848 & n5085 ) | ( ~n4848 & n5086 ) | ( n5085 & n5086 ) ;
  assign n5089 = ( n4848 & ~n5087 ) | ( n4848 & n5088 ) | ( ~n5087 & n5088 ) ;
  assign n5090 = ( ~n298 & n5084 ) | ( ~n298 & n5089 ) | ( n5084 & n5089 ) ;
  assign n5091 = n298 & ~n4849 ;
  assign n5092 = ( n298 & ~n4849 ) | ( n298 & n4898 ) | ( ~n4849 & n4898 ) ;
  assign n5093 = ( ~n4854 & n5091 ) | ( ~n4854 & n5092 ) | ( n5091 & n5092 ) ;
  assign n5094 = ( n4854 & n5091 ) | ( n4854 & n5092 ) | ( n5091 & n5092 ) ;
  assign n5095 = ( n4854 & n5093 ) | ( n4854 & ~n5094 ) | ( n5093 & ~n5094 ) ;
  assign n5096 = ( ~n258 & n5090 ) | ( ~n258 & n5095 ) | ( n5090 & n5095 ) ;
  assign n5097 = ( n258 & ~n4855 ) | ( n258 & n4898 ) | ( ~n4855 & n4898 ) ;
  assign n5098 = n258 & ~n4855 ;
  assign n5099 = ( n4860 & n5097 ) | ( n4860 & n5098 ) | ( n5097 & n5098 ) ;
  assign n5100 = ( ~n4860 & n5097 ) | ( ~n4860 & n5098 ) | ( n5097 & n5098 ) ;
  assign n5101 = ( n4860 & ~n5099 ) | ( n4860 & n5100 ) | ( ~n5099 & n5100 ) ;
  assign n5102 = ( ~n225 & n5096 ) | ( ~n225 & n5101 ) | ( n5096 & n5101 ) ;
  assign n5103 = ~n225 & n4861 ;
  assign n5104 = ( ~n225 & n4861 ) | ( ~n225 & n4898 ) | ( n4861 & n4898 ) ;
  assign n5105 = ( ~n4866 & n5103 ) | ( ~n4866 & n5104 ) | ( n5103 & n5104 ) ;
  assign n5106 = ( n4866 & n5103 ) | ( n4866 & n5104 ) | ( n5103 & n5104 ) ;
  assign n5107 = ( n4866 & n5105 ) | ( n4866 & ~n5106 ) | ( n5105 & ~n5106 ) ;
  assign n5108 = ( ~n197 & n5102 ) | ( ~n197 & n5107 ) | ( n5102 & n5107 ) ;
  assign n5109 = ( n197 & ~n4867 ) | ( n197 & n4898 ) | ( ~n4867 & n4898 ) ;
  assign n5110 = n197 & ~n4867 ;
  assign n5111 = ( n4872 & n5109 ) | ( n4872 & n5110 ) | ( n5109 & n5110 ) ;
  assign n5112 = ( ~n4872 & n5109 ) | ( ~n4872 & n5110 ) | ( n5109 & n5110 ) ;
  assign n5113 = ( n4872 & ~n5111 ) | ( n4872 & n5112 ) | ( ~n5111 & n5112 ) ;
  assign n5114 = ( ~n170 & n5108 ) | ( ~n170 & n5113 ) | ( n5108 & n5113 ) ;
  assign n5115 = ( n170 & ~n4873 ) | ( n170 & n4898 ) | ( ~n4873 & n4898 ) ;
  assign n5116 = n170 & ~n4873 ;
  assign n5117 = ( n4878 & n5115 ) | ( n4878 & n5116 ) | ( n5115 & n5116 ) ;
  assign n5118 = ( ~n4878 & n5115 ) | ( ~n4878 & n5116 ) | ( n5115 & n5116 ) ;
  assign n5119 = ( n4878 & ~n5117 ) | ( n4878 & n5118 ) | ( ~n5117 & n5118 ) ;
  assign n5120 = ( ~n142 & n5114 ) | ( ~n142 & n5119 ) | ( n5114 & n5119 ) ;
  assign n5121 = ~n142 & n4879 ;
  assign n5122 = ( ~n142 & n4879 ) | ( ~n142 & n4898 ) | ( n4879 & n4898 ) ;
  assign n5123 = ( ~n4884 & n5121 ) | ( ~n4884 & n5122 ) | ( n5121 & n5122 ) ;
  assign n5124 = ( n4884 & n5121 ) | ( n4884 & n5122 ) | ( n5121 & n5122 ) ;
  assign n5125 = ( n4884 & n5123 ) | ( n4884 & ~n5124 ) | ( n5123 & ~n5124 ) ;
  assign n5126 = ( ~n132 & n5120 ) | ( ~n132 & n5125 ) | ( n5120 & n5125 ) ;
  assign n5127 = n132 & ~n4885 ;
  assign n5128 = ( n132 & ~n4885 ) | ( n132 & n4898 ) | ( ~n4885 & n4898 ) ;
  assign n5129 = ( n4890 & n5127 ) | ( n4890 & n5128 ) | ( n5127 & n5128 ) ;
  assign n5130 = ( ~n4890 & n5127 ) | ( ~n4890 & n5128 ) | ( n5127 & n5128 ) ;
  assign n5131 = ( n4890 & ~n5129 ) | ( n4890 & n5130 ) | ( ~n5129 & n5130 ) ;
  assign n5132 = ( ~n131 & n5126 ) | ( ~n131 & n5131 ) | ( n5126 & n5131 ) ;
  assign n5133 = ~n4891 & n4895 ;
  assign n5134 = n4669 & n4891 ;
  assign n5135 = ( ~n131 & n5133 ) | ( ~n131 & n5134 ) | ( n5133 & n5134 ) ;
  assign n5136 = ( n131 & n4669 ) | ( n131 & n4891 ) | ( n4669 & n4891 ) ;
  assign n5137 = ( ~n4664 & n4891 ) | ( ~n4664 & n5134 ) | ( n4891 & n5134 ) ;
  assign n5138 = ( n5135 & n5136 ) | ( n5135 & ~n5137 ) | ( n5136 & ~n5137 ) ;
  assign n5139 = n5132 | n5138 ;
  assign n5140 = ~n5132 & n5135 ;
  assign n5141 = ( ~n5131 & n5136 ) | ( ~n5131 & n5137 ) | ( n5136 & n5137 ) ;
  assign n5142 = ~n5137 & n5141 ;
  assign n5143 = ( ~n131 & n5126 ) | ( ~n131 & n5142 ) | ( n5126 & n5142 ) ;
  assign n5144 = ( n5131 & ~n5132 ) | ( n5131 & n5143 ) | ( ~n5132 & n5143 ) ;
  assign n5145 = n5140 | n5144 ;
  assign n5146 = x44 | x45 ;
  assign n5147 = x46 | n5146 ;
  assign n5148 = ~n4898 & n5147 ;
  assign n5149 = ( x47 & ~n5139 ) | ( x47 & n5148 ) | ( ~n5139 & n5148 ) ;
  assign n5150 = n4898 & ~n5147 ;
  assign n5151 = ~n4900 & n5139 ;
  assign n5152 = ( n5149 & ~n5150 ) | ( n5149 & n5151 ) | ( ~n5150 & n5151 ) ;
  assign n5153 = n4898 & ~n5139 ;
  assign n5154 = ( x48 & n5151 ) | ( x48 & n5153 ) | ( n5151 & n5153 ) ;
  assign n5155 = ( ~x48 & n5151 ) | ( ~x48 & n5153 ) | ( n5151 & n5153 ) ;
  assign n5156 = ( x48 & ~n5154 ) | ( x48 & n5155 ) | ( ~n5154 & n5155 ) ;
  assign n5157 = ( ~n4661 & n5152 ) | ( ~n4661 & n5156 ) | ( n5152 & n5156 ) ;
  assign n5158 = ~n4661 & n4898 ;
  assign n5159 = ( n4906 & n5139 ) | ( n4906 & n5158 ) | ( n5139 & n5158 ) ;
  assign n5160 = ( ~x49 & n5155 ) | ( ~x49 & n5159 ) | ( n5155 & n5159 ) ;
  assign n5161 = ( x49 & n5155 ) | ( x49 & n5159 ) | ( n5155 & n5159 ) ;
  assign n5162 = ( x49 & n5160 ) | ( x49 & ~n5161 ) | ( n5160 & ~n5161 ) ;
  assign n5163 = ( ~n4432 & n5157 ) | ( ~n4432 & n5162 ) | ( n5157 & n5162 ) ;
  assign n5164 = n4432 & ~n4905 ;
  assign n5165 = ( n4432 & ~n4905 ) | ( n4432 & n5139 ) | ( ~n4905 & n5139 ) ;
  assign n5166 = ( n4909 & n5164 ) | ( n4909 & n5165 ) | ( n5164 & n5165 ) ;
  assign n5167 = ( ~n4909 & n5164 ) | ( ~n4909 & n5165 ) | ( n5164 & n5165 ) ;
  assign n5168 = ( n4909 & ~n5166 ) | ( n4909 & n5167 ) | ( ~n5166 & n5167 ) ;
  assign n5169 = ( ~n4203 & n5163 ) | ( ~n4203 & n5168 ) | ( n5163 & n5168 ) ;
  assign n5170 = ~n4203 & n4910 ;
  assign n5171 = ( ~n4203 & n4910 ) | ( ~n4203 & n5139 ) | ( n4910 & n5139 ) ;
  assign n5172 = ( ~n4915 & n5170 ) | ( ~n4915 & n5171 ) | ( n5170 & n5171 ) ;
  assign n5173 = ( n4915 & n5170 ) | ( n4915 & n5171 ) | ( n5170 & n5171 ) ;
  assign n5174 = ( n4915 & n5172 ) | ( n4915 & ~n5173 ) | ( n5172 & ~n5173 ) ;
  assign n5175 = ( ~n3985 & n5169 ) | ( ~n3985 & n5174 ) | ( n5169 & n5174 ) ;
  assign n5176 = n3985 & ~n4916 ;
  assign n5177 = ( n3985 & ~n4916 ) | ( n3985 & n5139 ) | ( ~n4916 & n5139 ) ;
  assign n5178 = ( n4921 & n5176 ) | ( n4921 & n5177 ) | ( n5176 & n5177 ) ;
  assign n5179 = ( ~n4921 & n5176 ) | ( ~n4921 & n5177 ) | ( n5176 & n5177 ) ;
  assign n5180 = ( n4921 & ~n5178 ) | ( n4921 & n5179 ) | ( ~n5178 & n5179 ) ;
  assign n5181 = ( ~n3772 & n5175 ) | ( ~n3772 & n5180 ) | ( n5175 & n5180 ) ;
  assign n5182 = ~n3772 & n4922 ;
  assign n5183 = ( ~n3772 & n4922 ) | ( ~n3772 & n5139 ) | ( n4922 & n5139 ) ;
  assign n5184 = ( n4927 & n5182 ) | ( n4927 & n5183 ) | ( n5182 & n5183 ) ;
  assign n5185 = ( ~n4927 & n5182 ) | ( ~n4927 & n5183 ) | ( n5182 & n5183 ) ;
  assign n5186 = ( n4927 & ~n5184 ) | ( n4927 & n5185 ) | ( ~n5184 & n5185 ) ;
  assign n5187 = ( ~n3567 & n5181 ) | ( ~n3567 & n5186 ) | ( n5181 & n5186 ) ;
  assign n5188 = n3567 & ~n4928 ;
  assign n5189 = ( n3567 & ~n4928 ) | ( n3567 & n5139 ) | ( ~n4928 & n5139 ) ;
  assign n5190 = ( n4933 & n5188 ) | ( n4933 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5191 = ( ~n4933 & n5188 ) | ( ~n4933 & n5189 ) | ( n5188 & n5189 ) ;
  assign n5192 = ( n4933 & ~n5190 ) | ( n4933 & n5191 ) | ( ~n5190 & n5191 ) ;
  assign n5193 = ( ~n3362 & n5187 ) | ( ~n3362 & n5192 ) | ( n5187 & n5192 ) ;
  assign n5194 = ( n3362 & ~n4934 ) | ( n3362 & n5139 ) | ( ~n4934 & n5139 ) ;
  assign n5195 = n3362 & ~n4934 ;
  assign n5196 = ( n4939 & n5194 ) | ( n4939 & n5195 ) | ( n5194 & n5195 ) ;
  assign n5197 = ( ~n4939 & n5194 ) | ( ~n4939 & n5195 ) | ( n5194 & n5195 ) ;
  assign n5198 = ( n4939 & ~n5196 ) | ( n4939 & n5197 ) | ( ~n5196 & n5197 ) ;
  assign n5199 = ( ~n3169 & n5193 ) | ( ~n3169 & n5198 ) | ( n5193 & n5198 ) ;
  assign n5200 = ( n3169 & ~n4940 ) | ( n3169 & n5139 ) | ( ~n4940 & n5139 ) ;
  assign n5201 = n3169 & ~n4940 ;
  assign n5202 = ( n4945 & n5200 ) | ( n4945 & n5201 ) | ( n5200 & n5201 ) ;
  assign n5203 = ( ~n4945 & n5200 ) | ( ~n4945 & n5201 ) | ( n5200 & n5201 ) ;
  assign n5204 = ( n4945 & ~n5202 ) | ( n4945 & n5203 ) | ( ~n5202 & n5203 ) ;
  assign n5205 = ( ~n2979 & n5199 ) | ( ~n2979 & n5204 ) | ( n5199 & n5204 ) ;
  assign n5206 = ( n2979 & ~n4946 ) | ( n2979 & n5139 ) | ( ~n4946 & n5139 ) ;
  assign n5207 = n2979 & ~n4946 ;
  assign n5208 = ( n4951 & n5206 ) | ( n4951 & n5207 ) | ( n5206 & n5207 ) ;
  assign n5209 = ( ~n4951 & n5206 ) | ( ~n4951 & n5207 ) | ( n5206 & n5207 ) ;
  assign n5210 = ( n4951 & ~n5208 ) | ( n4951 & n5209 ) | ( ~n5208 & n5209 ) ;
  assign n5211 = ( ~n2791 & n5205 ) | ( ~n2791 & n5210 ) | ( n5205 & n5210 ) ;
  assign n5212 = ( n2791 & ~n4952 ) | ( n2791 & n5139 ) | ( ~n4952 & n5139 ) ;
  assign n5213 = n2791 & ~n4952 ;
  assign n5214 = ( n4957 & n5212 ) | ( n4957 & n5213 ) | ( n5212 & n5213 ) ;
  assign n5215 = ( ~n4957 & n5212 ) | ( ~n4957 & n5213 ) | ( n5212 & n5213 ) ;
  assign n5216 = ( n4957 & ~n5214 ) | ( n4957 & n5215 ) | ( ~n5214 & n5215 ) ;
  assign n5217 = ( ~n2615 & n5211 ) | ( ~n2615 & n5216 ) | ( n5211 & n5216 ) ;
  assign n5218 = ( n2615 & ~n4958 ) | ( n2615 & n5139 ) | ( ~n4958 & n5139 ) ;
  assign n5219 = n2615 & ~n4958 ;
  assign n5220 = ( n4963 & n5218 ) | ( n4963 & n5219 ) | ( n5218 & n5219 ) ;
  assign n5221 = ( ~n4963 & n5218 ) | ( ~n4963 & n5219 ) | ( n5218 & n5219 ) ;
  assign n5222 = ( n4963 & ~n5220 ) | ( n4963 & n5221 ) | ( ~n5220 & n5221 ) ;
  assign n5223 = ( ~n2443 & n5217 ) | ( ~n2443 & n5222 ) | ( n5217 & n5222 ) ;
  assign n5224 = ~n2443 & n4964 ;
  assign n5225 = ( ~n2443 & n4964 ) | ( ~n2443 & n5139 ) | ( n4964 & n5139 ) ;
  assign n5226 = ( n4969 & n5224 ) | ( n4969 & n5225 ) | ( n5224 & n5225 ) ;
  assign n5227 = ( ~n4969 & n5224 ) | ( ~n4969 & n5225 ) | ( n5224 & n5225 ) ;
  assign n5228 = ( n4969 & ~n5226 ) | ( n4969 & n5227 ) | ( ~n5226 & n5227 ) ;
  assign n5229 = ( ~n2277 & n5223 ) | ( ~n2277 & n5228 ) | ( n5223 & n5228 ) ;
  assign n5230 = ( n2277 & ~n4970 ) | ( n2277 & n5139 ) | ( ~n4970 & n5139 ) ;
  assign n5231 = n2277 & ~n4970 ;
  assign n5232 = ( n4975 & n5230 ) | ( n4975 & n5231 ) | ( n5230 & n5231 ) ;
  assign n5233 = ( ~n4975 & n5230 ) | ( ~n4975 & n5231 ) | ( n5230 & n5231 ) ;
  assign n5234 = ( n4975 & ~n5232 ) | ( n4975 & n5233 ) | ( ~n5232 & n5233 ) ;
  assign n5235 = ( ~n2111 & n5229 ) | ( ~n2111 & n5234 ) | ( n5229 & n5234 ) ;
  assign n5236 = ~n2111 & n4976 ;
  assign n5237 = ( ~n2111 & n4976 ) | ( ~n2111 & n5139 ) | ( n4976 & n5139 ) ;
  assign n5238 = ( ~n4981 & n5236 ) | ( ~n4981 & n5237 ) | ( n5236 & n5237 ) ;
  assign n5239 = ( n4981 & n5236 ) | ( n4981 & n5237 ) | ( n5236 & n5237 ) ;
  assign n5240 = ( n4981 & n5238 ) | ( n4981 & ~n5239 ) | ( n5238 & ~n5239 ) ;
  assign n5241 = ( ~n1949 & n5235 ) | ( ~n1949 & n5240 ) | ( n5235 & n5240 ) ;
  assign n5242 = ( n1949 & ~n4982 ) | ( n1949 & n5139 ) | ( ~n4982 & n5139 ) ;
  assign n5243 = n1949 & ~n4982 ;
  assign n5244 = ( n4987 & n5242 ) | ( n4987 & n5243 ) | ( n5242 & n5243 ) ;
  assign n5245 = ( ~n4987 & n5242 ) | ( ~n4987 & n5243 ) | ( n5242 & n5243 ) ;
  assign n5246 = ( n4987 & ~n5244 ) | ( n4987 & n5245 ) | ( ~n5244 & n5245 ) ;
  assign n5247 = ( ~n1802 & n5241 ) | ( ~n1802 & n5246 ) | ( n5241 & n5246 ) ;
  assign n5248 = ~n1802 & n4988 ;
  assign n5249 = ( ~n1802 & n4988 ) | ( ~n1802 & n5139 ) | ( n4988 & n5139 ) ;
  assign n5250 = ( n4993 & n5248 ) | ( n4993 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5251 = ( ~n4993 & n5248 ) | ( ~n4993 & n5249 ) | ( n5248 & n5249 ) ;
  assign n5252 = ( n4993 & ~n5250 ) | ( n4993 & n5251 ) | ( ~n5250 & n5251 ) ;
  assign n5253 = ( ~n1661 & n5247 ) | ( ~n1661 & n5252 ) | ( n5247 & n5252 ) ;
  assign n5254 = ~n1661 & n4994 ;
  assign n5255 = ( ~n1661 & n4994 ) | ( ~n1661 & n5139 ) | ( n4994 & n5139 ) ;
  assign n5256 = ( ~n4999 & n5254 ) | ( ~n4999 & n5255 ) | ( n5254 & n5255 ) ;
  assign n5257 = ( n4999 & n5254 ) | ( n4999 & n5255 ) | ( n5254 & n5255 ) ;
  assign n5258 = ( n4999 & n5256 ) | ( n4999 & ~n5257 ) | ( n5256 & ~n5257 ) ;
  assign n5259 = ( ~n1523 & n5253 ) | ( ~n1523 & n5258 ) | ( n5253 & n5258 ) ;
  assign n5260 = ( n1523 & ~n5000 ) | ( n1523 & n5139 ) | ( ~n5000 & n5139 ) ;
  assign n5261 = n1523 & ~n5000 ;
  assign n5262 = ( n5005 & n5260 ) | ( n5005 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5263 = ( ~n5005 & n5260 ) | ( ~n5005 & n5261 ) | ( n5260 & n5261 ) ;
  assign n5264 = ( n5005 & ~n5262 ) | ( n5005 & n5263 ) | ( ~n5262 & n5263 ) ;
  assign n5265 = ( ~n1393 & n5259 ) | ( ~n1393 & n5264 ) | ( n5259 & n5264 ) ;
  assign n5266 = ( n1393 & ~n5006 ) | ( n1393 & n5139 ) | ( ~n5006 & n5139 ) ;
  assign n5267 = n1393 & ~n5006 ;
  assign n5268 = ( n5011 & n5266 ) | ( n5011 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5269 = ( ~n5011 & n5266 ) | ( ~n5011 & n5267 ) | ( n5266 & n5267 ) ;
  assign n5270 = ( n5011 & ~n5268 ) | ( n5011 & n5269 ) | ( ~n5268 & n5269 ) ;
  assign n5271 = ( ~n1266 & n5265 ) | ( ~n1266 & n5270 ) | ( n5265 & n5270 ) ;
  assign n5272 = ( n1266 & ~n5012 ) | ( n1266 & n5139 ) | ( ~n5012 & n5139 ) ;
  assign n5273 = n1266 & ~n5012 ;
  assign n5274 = ( n5017 & n5272 ) | ( n5017 & n5273 ) | ( n5272 & n5273 ) ;
  assign n5275 = ( ~n5017 & n5272 ) | ( ~n5017 & n5273 ) | ( n5272 & n5273 ) ;
  assign n5276 = ( n5017 & ~n5274 ) | ( n5017 & n5275 ) | ( ~n5274 & n5275 ) ;
  assign n5277 = ( ~n1150 & n5271 ) | ( ~n1150 & n5276 ) | ( n5271 & n5276 ) ;
  assign n5278 = ( n1150 & ~n5018 ) | ( n1150 & n5139 ) | ( ~n5018 & n5139 ) ;
  assign n5279 = n1150 & ~n5018 ;
  assign n5280 = ( n5023 & n5278 ) | ( n5023 & n5279 ) | ( n5278 & n5279 ) ;
  assign n5281 = ( ~n5023 & n5278 ) | ( ~n5023 & n5279 ) | ( n5278 & n5279 ) ;
  assign n5282 = ( n5023 & ~n5280 ) | ( n5023 & n5281 ) | ( ~n5280 & n5281 ) ;
  assign n5283 = ( ~n1038 & n5277 ) | ( ~n1038 & n5282 ) | ( n5277 & n5282 ) ;
  assign n5284 = ( n1038 & ~n5024 ) | ( n1038 & n5139 ) | ( ~n5024 & n5139 ) ;
  assign n5285 = n1038 & ~n5024 ;
  assign n5286 = ( n5029 & n5284 ) | ( n5029 & n5285 ) | ( n5284 & n5285 ) ;
  assign n5287 = ( ~n5029 & n5284 ) | ( ~n5029 & n5285 ) | ( n5284 & n5285 ) ;
  assign n5288 = ( n5029 & ~n5286 ) | ( n5029 & n5287 ) | ( ~n5286 & n5287 ) ;
  assign n5289 = ( ~n933 & n5283 ) | ( ~n933 & n5288 ) | ( n5283 & n5288 ) ;
  assign n5290 = ~n933 & n5030 ;
  assign n5291 = ( ~n933 & n5030 ) | ( ~n933 & n5139 ) | ( n5030 & n5139 ) ;
  assign n5292 = ( n5035 & n5290 ) | ( n5035 & n5291 ) | ( n5290 & n5291 ) ;
  assign n5293 = ( ~n5035 & n5290 ) | ( ~n5035 & n5291 ) | ( n5290 & n5291 ) ;
  assign n5294 = ( n5035 & ~n5292 ) | ( n5035 & n5293 ) | ( ~n5292 & n5293 ) ;
  assign n5295 = ( ~n839 & n5289 ) | ( ~n839 & n5294 ) | ( n5289 & n5294 ) ;
  assign n5296 = ( n839 & ~n5036 ) | ( n839 & n5139 ) | ( ~n5036 & n5139 ) ;
  assign n5297 = n839 & ~n5036 ;
  assign n5298 = ( n5041 & n5296 ) | ( n5041 & n5297 ) | ( n5296 & n5297 ) ;
  assign n5299 = ( ~n5041 & n5296 ) | ( ~n5041 & n5297 ) | ( n5296 & n5297 ) ;
  assign n5300 = ( n5041 & ~n5298 ) | ( n5041 & n5299 ) | ( ~n5298 & n5299 ) ;
  assign n5301 = ( ~n746 & n5295 ) | ( ~n746 & n5300 ) | ( n5295 & n5300 ) ;
  assign n5302 = ( n746 & ~n5042 ) | ( n746 & n5139 ) | ( ~n5042 & n5139 ) ;
  assign n5303 = n746 & ~n5042 ;
  assign n5304 = ( n5047 & n5302 ) | ( n5047 & n5303 ) | ( n5302 & n5303 ) ;
  assign n5305 = ( ~n5047 & n5302 ) | ( ~n5047 & n5303 ) | ( n5302 & n5303 ) ;
  assign n5306 = ( n5047 & ~n5304 ) | ( n5047 & n5305 ) | ( ~n5304 & n5305 ) ;
  assign n5307 = ( ~n664 & n5301 ) | ( ~n664 & n5306 ) | ( n5301 & n5306 ) ;
  assign n5308 = ( n664 & ~n5048 ) | ( n664 & n5139 ) | ( ~n5048 & n5139 ) ;
  assign n5309 = n664 & ~n5048 ;
  assign n5310 = ( n5053 & n5308 ) | ( n5053 & n5309 ) | ( n5308 & n5309 ) ;
  assign n5311 = ( ~n5053 & n5308 ) | ( ~n5053 & n5309 ) | ( n5308 & n5309 ) ;
  assign n5312 = ( n5053 & ~n5310 ) | ( n5053 & n5311 ) | ( ~n5310 & n5311 ) ;
  assign n5313 = ( ~n588 & n5307 ) | ( ~n588 & n5312 ) | ( n5307 & n5312 ) ;
  assign n5314 = ~n588 & n5054 ;
  assign n5315 = ( ~n588 & n5054 ) | ( ~n588 & n5139 ) | ( n5054 & n5139 ) ;
  assign n5316 = ( ~n5059 & n5314 ) | ( ~n5059 & n5315 ) | ( n5314 & n5315 ) ;
  assign n5317 = ( n5059 & n5314 ) | ( n5059 & n5315 ) | ( n5314 & n5315 ) ;
  assign n5318 = ( n5059 & n5316 ) | ( n5059 & ~n5317 ) | ( n5316 & ~n5317 ) ;
  assign n5319 = ( ~n518 & n5313 ) | ( ~n518 & n5318 ) | ( n5313 & n5318 ) ;
  assign n5320 = ( n518 & ~n5060 ) | ( n518 & n5139 ) | ( ~n5060 & n5139 ) ;
  assign n5321 = n518 & ~n5060 ;
  assign n5322 = ( n5065 & n5320 ) | ( n5065 & n5321 ) | ( n5320 & n5321 ) ;
  assign n5323 = ( ~n5065 & n5320 ) | ( ~n5065 & n5321 ) | ( n5320 & n5321 ) ;
  assign n5324 = ( n5065 & ~n5322 ) | ( n5065 & n5323 ) | ( ~n5322 & n5323 ) ;
  assign n5325 = ( ~n454 & n5319 ) | ( ~n454 & n5324 ) | ( n5319 & n5324 ) ;
  assign n5326 = ( n454 & ~n5066 ) | ( n454 & n5139 ) | ( ~n5066 & n5139 ) ;
  assign n5327 = n454 & ~n5066 ;
  assign n5328 = ( ~n5071 & n5326 ) | ( ~n5071 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5329 = ( n5071 & n5326 ) | ( n5071 & n5327 ) | ( n5326 & n5327 ) ;
  assign n5330 = ( n5071 & n5328 ) | ( n5071 & ~n5329 ) | ( n5328 & ~n5329 ) ;
  assign n5331 = ( ~n396 & n5325 ) | ( ~n396 & n5330 ) | ( n5325 & n5330 ) ;
  assign n5332 = ( n396 & ~n5072 ) | ( n396 & n5139 ) | ( ~n5072 & n5139 ) ;
  assign n5333 = n396 & ~n5072 ;
  assign n5334 = ( n5077 & n5332 ) | ( n5077 & n5333 ) | ( n5332 & n5333 ) ;
  assign n5335 = ( ~n5077 & n5332 ) | ( ~n5077 & n5333 ) | ( n5332 & n5333 ) ;
  assign n5336 = ( n5077 & ~n5334 ) | ( n5077 & n5335 ) | ( ~n5334 & n5335 ) ;
  assign n5337 = ( ~n344 & n5331 ) | ( ~n344 & n5336 ) | ( n5331 & n5336 ) ;
  assign n5338 = ~n344 & n5078 ;
  assign n5339 = ( ~n344 & n5078 ) | ( ~n344 & n5139 ) | ( n5078 & n5139 ) ;
  assign n5340 = ( ~n5083 & n5338 ) | ( ~n5083 & n5339 ) | ( n5338 & n5339 ) ;
  assign n5341 = ( n5083 & n5338 ) | ( n5083 & n5339 ) | ( n5338 & n5339 ) ;
  assign n5342 = ( n5083 & n5340 ) | ( n5083 & ~n5341 ) | ( n5340 & ~n5341 ) ;
  assign n5343 = ( ~n298 & n5337 ) | ( ~n298 & n5342 ) | ( n5337 & n5342 ) ;
  assign n5344 = ( n298 & ~n5084 ) | ( n298 & n5139 ) | ( ~n5084 & n5139 ) ;
  assign n5345 = n298 & ~n5084 ;
  assign n5346 = ( n5089 & n5344 ) | ( n5089 & n5345 ) | ( n5344 & n5345 ) ;
  assign n5347 = ( ~n5089 & n5344 ) | ( ~n5089 & n5345 ) | ( n5344 & n5345 ) ;
  assign n5348 = ( n5089 & ~n5346 ) | ( n5089 & n5347 ) | ( ~n5346 & n5347 ) ;
  assign n5349 = ( ~n258 & n5343 ) | ( ~n258 & n5348 ) | ( n5343 & n5348 ) ;
  assign n5350 = ~n258 & n5090 ;
  assign n5351 = ( ~n258 & n5090 ) | ( ~n258 & n5139 ) | ( n5090 & n5139 ) ;
  assign n5352 = ( n5095 & n5350 ) | ( n5095 & n5351 ) | ( n5350 & n5351 ) ;
  assign n5353 = ( ~n5095 & n5350 ) | ( ~n5095 & n5351 ) | ( n5350 & n5351 ) ;
  assign n5354 = ( n5095 & ~n5352 ) | ( n5095 & n5353 ) | ( ~n5352 & n5353 ) ;
  assign n5355 = ( ~n225 & n5349 ) | ( ~n225 & n5354 ) | ( n5349 & n5354 ) ;
  assign n5356 = ( n225 & ~n5096 ) | ( n225 & n5139 ) | ( ~n5096 & n5139 ) ;
  assign n5357 = n225 & ~n5096 ;
  assign n5358 = ( n5101 & n5356 ) | ( n5101 & n5357 ) | ( n5356 & n5357 ) ;
  assign n5359 = ( ~n5101 & n5356 ) | ( ~n5101 & n5357 ) | ( n5356 & n5357 ) ;
  assign n5360 = ( n5101 & ~n5358 ) | ( n5101 & n5359 ) | ( ~n5358 & n5359 ) ;
  assign n5361 = ( ~n197 & n5355 ) | ( ~n197 & n5360 ) | ( n5355 & n5360 ) ;
  assign n5362 = ~n197 & n5102 ;
  assign n5363 = ( ~n197 & n5102 ) | ( ~n197 & n5139 ) | ( n5102 & n5139 ) ;
  assign n5364 = ( n5107 & n5362 ) | ( n5107 & n5363 ) | ( n5362 & n5363 ) ;
  assign n5365 = ( ~n5107 & n5362 ) | ( ~n5107 & n5363 ) | ( n5362 & n5363 ) ;
  assign n5366 = ( n5107 & ~n5364 ) | ( n5107 & n5365 ) | ( ~n5364 & n5365 ) ;
  assign n5367 = ( ~n170 & n5361 ) | ( ~n170 & n5366 ) | ( n5361 & n5366 ) ;
  assign n5368 = ( n170 & ~n5108 ) | ( n170 & n5139 ) | ( ~n5108 & n5139 ) ;
  assign n5369 = n170 & ~n5108 ;
  assign n5370 = ( n5113 & n5368 ) | ( n5113 & n5369 ) | ( n5368 & n5369 ) ;
  assign n5371 = ( ~n5113 & n5368 ) | ( ~n5113 & n5369 ) | ( n5368 & n5369 ) ;
  assign n5372 = ( n5113 & ~n5370 ) | ( n5113 & n5371 ) | ( ~n5370 & n5371 ) ;
  assign n5373 = ( ~n142 & n5367 ) | ( ~n142 & n5372 ) | ( n5367 & n5372 ) ;
  assign n5374 = ( n142 & ~n5114 ) | ( n142 & n5139 ) | ( ~n5114 & n5139 ) ;
  assign n5375 = n142 & ~n5114 ;
  assign n5376 = ( n5119 & n5374 ) | ( n5119 & n5375 ) | ( n5374 & n5375 ) ;
  assign n5377 = ( ~n5119 & n5374 ) | ( ~n5119 & n5375 ) | ( n5374 & n5375 ) ;
  assign n5378 = ( n5119 & ~n5376 ) | ( n5119 & n5377 ) | ( ~n5376 & n5377 ) ;
  assign n5379 = ( ~n132 & n5373 ) | ( ~n132 & n5378 ) | ( n5373 & n5378 ) ;
  assign n5380 = ( n132 & ~n5120 ) | ( n132 & n5139 ) | ( ~n5120 & n5139 ) ;
  assign n5381 = n132 & ~n5120 ;
  assign n5382 = ( n5125 & n5380 ) | ( n5125 & n5381 ) | ( n5380 & n5381 ) ;
  assign n5383 = ( ~n5125 & n5380 ) | ( ~n5125 & n5381 ) | ( n5380 & n5381 ) ;
  assign n5384 = ( n5125 & ~n5382 ) | ( n5125 & n5383 ) | ( ~n5382 & n5383 ) ;
  assign n5385 = ( ~n131 & n5379 ) | ( ~n131 & n5384 ) | ( n5379 & n5384 ) ;
  assign n5386 = n5145 | n5385 ;
  assign n5387 = x42 | x43 ;
  assign n5388 = x44 | n5387 ;
  assign n5389 = ~n5139 & n5388 ;
  assign n5390 = ( x45 & ~n5386 ) | ( x45 & n5389 ) | ( ~n5386 & n5389 ) ;
  assign n5391 = ~n5146 & n5386 ;
  assign n5392 = n5139 & ~n5388 ;
  assign n5393 = ( n5390 & n5391 ) | ( n5390 & ~n5392 ) | ( n5391 & ~n5392 ) ;
  assign n5394 = n5139 & ~n5386 ;
  assign n5395 = ( x46 & n5391 ) | ( x46 & n5394 ) | ( n5391 & n5394 ) ;
  assign n5396 = ( ~x46 & n5391 ) | ( ~x46 & n5394 ) | ( n5391 & n5394 ) ;
  assign n5397 = ( x46 & ~n5395 ) | ( x46 & n5396 ) | ( ~n5395 & n5396 ) ;
  assign n5398 = ( ~n4898 & n5393 ) | ( ~n4898 & n5397 ) | ( n5393 & n5397 ) ;
  assign n5399 = ~n4898 & n5139 ;
  assign n5400 = ( n5153 & n5386 ) | ( n5153 & n5399 ) | ( n5386 & n5399 ) ;
  assign n5401 = ( ~x47 & n5396 ) | ( ~x47 & n5400 ) | ( n5396 & n5400 ) ;
  assign n5402 = ( x47 & n5396 ) | ( x47 & n5400 ) | ( n5396 & n5400 ) ;
  assign n5403 = ( x47 & n5401 ) | ( x47 & ~n5402 ) | ( n5401 & ~n5402 ) ;
  assign n5404 = ( ~n4661 & n5398 ) | ( ~n4661 & n5403 ) | ( n5398 & n5403 ) ;
  assign n5405 = ( n4661 & ~n5152 ) | ( n4661 & n5386 ) | ( ~n5152 & n5386 ) ;
  assign n5406 = n4661 & ~n5152 ;
  assign n5407 = ( n5156 & n5405 ) | ( n5156 & n5406 ) | ( n5405 & n5406 ) ;
  assign n5408 = ( ~n5156 & n5405 ) | ( ~n5156 & n5406 ) | ( n5405 & n5406 ) ;
  assign n5409 = ( n5156 & ~n5407 ) | ( n5156 & n5408 ) | ( ~n5407 & n5408 ) ;
  assign n5410 = ( ~n4432 & n5404 ) | ( ~n4432 & n5409 ) | ( n5404 & n5409 ) ;
  assign n5411 = ( n4432 & ~n5157 ) | ( n4432 & n5386 ) | ( ~n5157 & n5386 ) ;
  assign n5412 = n4432 & ~n5157 ;
  assign n5413 = ( n5162 & n5411 ) | ( n5162 & n5412 ) | ( n5411 & n5412 ) ;
  assign n5414 = ( ~n5162 & n5411 ) | ( ~n5162 & n5412 ) | ( n5411 & n5412 ) ;
  assign n5415 = ( n5162 & ~n5413 ) | ( n5162 & n5414 ) | ( ~n5413 & n5414 ) ;
  assign n5416 = ( ~n4203 & n5410 ) | ( ~n4203 & n5415 ) | ( n5410 & n5415 ) ;
  assign n5417 = n4203 & ~n5163 ;
  assign n5418 = ( n4203 & ~n5163 ) | ( n4203 & n5386 ) | ( ~n5163 & n5386 ) ;
  assign n5419 = ( n5168 & n5417 ) | ( n5168 & n5418 ) | ( n5417 & n5418 ) ;
  assign n5420 = ( ~n5168 & n5417 ) | ( ~n5168 & n5418 ) | ( n5417 & n5418 ) ;
  assign n5421 = ( n5168 & ~n5419 ) | ( n5168 & n5420 ) | ( ~n5419 & n5420 ) ;
  assign n5422 = ( ~n3985 & n5416 ) | ( ~n3985 & n5421 ) | ( n5416 & n5421 ) ;
  assign n5423 = ( n3985 & ~n5169 ) | ( n3985 & n5386 ) | ( ~n5169 & n5386 ) ;
  assign n5424 = n3985 & ~n5169 ;
  assign n5425 = ( n5174 & n5423 ) | ( n5174 & n5424 ) | ( n5423 & n5424 ) ;
  assign n5426 = ( ~n5174 & n5423 ) | ( ~n5174 & n5424 ) | ( n5423 & n5424 ) ;
  assign n5427 = ( n5174 & ~n5425 ) | ( n5174 & n5426 ) | ( ~n5425 & n5426 ) ;
  assign n5428 = ( ~n3772 & n5422 ) | ( ~n3772 & n5427 ) | ( n5422 & n5427 ) ;
  assign n5429 = n3772 & ~n5175 ;
  assign n5430 = ( n3772 & ~n5175 ) | ( n3772 & n5386 ) | ( ~n5175 & n5386 ) ;
  assign n5431 = ( ~n5180 & n5429 ) | ( ~n5180 & n5430 ) | ( n5429 & n5430 ) ;
  assign n5432 = ( n5180 & n5429 ) | ( n5180 & n5430 ) | ( n5429 & n5430 ) ;
  assign n5433 = ( n5180 & n5431 ) | ( n5180 & ~n5432 ) | ( n5431 & ~n5432 ) ;
  assign n5434 = ( ~n3567 & n5428 ) | ( ~n3567 & n5433 ) | ( n5428 & n5433 ) ;
  assign n5435 = ( n3567 & ~n5181 ) | ( n3567 & n5386 ) | ( ~n5181 & n5386 ) ;
  assign n5436 = n3567 & ~n5181 ;
  assign n5437 = ( n5186 & n5435 ) | ( n5186 & n5436 ) | ( n5435 & n5436 ) ;
  assign n5438 = ( ~n5186 & n5435 ) | ( ~n5186 & n5436 ) | ( n5435 & n5436 ) ;
  assign n5439 = ( n5186 & ~n5437 ) | ( n5186 & n5438 ) | ( ~n5437 & n5438 ) ;
  assign n5440 = ( ~n3362 & n5434 ) | ( ~n3362 & n5439 ) | ( n5434 & n5439 ) ;
  assign n5441 = ( n3362 & ~n5187 ) | ( n3362 & n5386 ) | ( ~n5187 & n5386 ) ;
  assign n5442 = n3362 & ~n5187 ;
  assign n5443 = ( n5192 & n5441 ) | ( n5192 & n5442 ) | ( n5441 & n5442 ) ;
  assign n5444 = ( ~n5192 & n5441 ) | ( ~n5192 & n5442 ) | ( n5441 & n5442 ) ;
  assign n5445 = ( n5192 & ~n5443 ) | ( n5192 & n5444 ) | ( ~n5443 & n5444 ) ;
  assign n5446 = ( ~n3169 & n5440 ) | ( ~n3169 & n5445 ) | ( n5440 & n5445 ) ;
  assign n5447 = ( n3169 & ~n5193 ) | ( n3169 & n5386 ) | ( ~n5193 & n5386 ) ;
  assign n5448 = n3169 & ~n5193 ;
  assign n5449 = ( n5198 & n5447 ) | ( n5198 & n5448 ) | ( n5447 & n5448 ) ;
  assign n5450 = ( ~n5198 & n5447 ) | ( ~n5198 & n5448 ) | ( n5447 & n5448 ) ;
  assign n5451 = ( n5198 & ~n5449 ) | ( n5198 & n5450 ) | ( ~n5449 & n5450 ) ;
  assign n5452 = ( ~n2979 & n5446 ) | ( ~n2979 & n5451 ) | ( n5446 & n5451 ) ;
  assign n5453 = ( n2979 & ~n5199 ) | ( n2979 & n5386 ) | ( ~n5199 & n5386 ) ;
  assign n5454 = n2979 & ~n5199 ;
  assign n5455 = ( n5204 & n5453 ) | ( n5204 & n5454 ) | ( n5453 & n5454 ) ;
  assign n5456 = ( ~n5204 & n5453 ) | ( ~n5204 & n5454 ) | ( n5453 & n5454 ) ;
  assign n5457 = ( n5204 & ~n5455 ) | ( n5204 & n5456 ) | ( ~n5455 & n5456 ) ;
  assign n5458 = ( ~n2791 & n5452 ) | ( ~n2791 & n5457 ) | ( n5452 & n5457 ) ;
  assign n5459 = ~n2791 & n5205 ;
  assign n5460 = ( ~n2791 & n5205 ) | ( ~n2791 & n5386 ) | ( n5205 & n5386 ) ;
  assign n5461 = ( ~n5210 & n5459 ) | ( ~n5210 & n5460 ) | ( n5459 & n5460 ) ;
  assign n5462 = ( n5210 & n5459 ) | ( n5210 & n5460 ) | ( n5459 & n5460 ) ;
  assign n5463 = ( n5210 & n5461 ) | ( n5210 & ~n5462 ) | ( n5461 & ~n5462 ) ;
  assign n5464 = ( ~n2615 & n5458 ) | ( ~n2615 & n5463 ) | ( n5458 & n5463 ) ;
  assign n5465 = ( n2615 & ~n5211 ) | ( n2615 & n5386 ) | ( ~n5211 & n5386 ) ;
  assign n5466 = n2615 & ~n5211 ;
  assign n5467 = ( n5216 & n5465 ) | ( n5216 & n5466 ) | ( n5465 & n5466 ) ;
  assign n5468 = ( ~n5216 & n5465 ) | ( ~n5216 & n5466 ) | ( n5465 & n5466 ) ;
  assign n5469 = ( n5216 & ~n5467 ) | ( n5216 & n5468 ) | ( ~n5467 & n5468 ) ;
  assign n5470 = ( ~n2443 & n5464 ) | ( ~n2443 & n5469 ) | ( n5464 & n5469 ) ;
  assign n5471 = ( n2443 & ~n5217 ) | ( n2443 & n5386 ) | ( ~n5217 & n5386 ) ;
  assign n5472 = n2443 & ~n5217 ;
  assign n5473 = ( n5222 & n5471 ) | ( n5222 & n5472 ) | ( n5471 & n5472 ) ;
  assign n5474 = ( ~n5222 & n5471 ) | ( ~n5222 & n5472 ) | ( n5471 & n5472 ) ;
  assign n5475 = ( n5222 & ~n5473 ) | ( n5222 & n5474 ) | ( ~n5473 & n5474 ) ;
  assign n5476 = ( ~n2277 & n5470 ) | ( ~n2277 & n5475 ) | ( n5470 & n5475 ) ;
  assign n5477 = ( n2277 & ~n5223 ) | ( n2277 & n5386 ) | ( ~n5223 & n5386 ) ;
  assign n5478 = n2277 & ~n5223 ;
  assign n5479 = ( n5228 & n5477 ) | ( n5228 & n5478 ) | ( n5477 & n5478 ) ;
  assign n5480 = ( ~n5228 & n5477 ) | ( ~n5228 & n5478 ) | ( n5477 & n5478 ) ;
  assign n5481 = ( n5228 & ~n5479 ) | ( n5228 & n5480 ) | ( ~n5479 & n5480 ) ;
  assign n5482 = ( ~n2111 & n5476 ) | ( ~n2111 & n5481 ) | ( n5476 & n5481 ) ;
  assign n5483 = ~n2111 & n5229 ;
  assign n5484 = ( ~n2111 & n5229 ) | ( ~n2111 & n5386 ) | ( n5229 & n5386 ) ;
  assign n5485 = ( ~n5234 & n5483 ) | ( ~n5234 & n5484 ) | ( n5483 & n5484 ) ;
  assign n5486 = ( n5234 & n5483 ) | ( n5234 & n5484 ) | ( n5483 & n5484 ) ;
  assign n5487 = ( n5234 & n5485 ) | ( n5234 & ~n5486 ) | ( n5485 & ~n5486 ) ;
  assign n5488 = ( ~n1949 & n5482 ) | ( ~n1949 & n5487 ) | ( n5482 & n5487 ) ;
  assign n5489 = ( n1949 & ~n5235 ) | ( n1949 & n5386 ) | ( ~n5235 & n5386 ) ;
  assign n5490 = n1949 & ~n5235 ;
  assign n5491 = ( n5240 & n5489 ) | ( n5240 & n5490 ) | ( n5489 & n5490 ) ;
  assign n5492 = ( ~n5240 & n5489 ) | ( ~n5240 & n5490 ) | ( n5489 & n5490 ) ;
  assign n5493 = ( n5240 & ~n5491 ) | ( n5240 & n5492 ) | ( ~n5491 & n5492 ) ;
  assign n5494 = ( ~n1802 & n5488 ) | ( ~n1802 & n5493 ) | ( n5488 & n5493 ) ;
  assign n5495 = ( n1802 & ~n5241 ) | ( n1802 & n5386 ) | ( ~n5241 & n5386 ) ;
  assign n5496 = n1802 & ~n5241 ;
  assign n5497 = ( n5246 & n5495 ) | ( n5246 & n5496 ) | ( n5495 & n5496 ) ;
  assign n5498 = ( ~n5246 & n5495 ) | ( ~n5246 & n5496 ) | ( n5495 & n5496 ) ;
  assign n5499 = ( n5246 & ~n5497 ) | ( n5246 & n5498 ) | ( ~n5497 & n5498 ) ;
  assign n5500 = ( ~n1661 & n5494 ) | ( ~n1661 & n5499 ) | ( n5494 & n5499 ) ;
  assign n5501 = ( n1661 & ~n5247 ) | ( n1661 & n5386 ) | ( ~n5247 & n5386 ) ;
  assign n5502 = n1661 & ~n5247 ;
  assign n5503 = ( n5252 & n5501 ) | ( n5252 & n5502 ) | ( n5501 & n5502 ) ;
  assign n5504 = ( ~n5252 & n5501 ) | ( ~n5252 & n5502 ) | ( n5501 & n5502 ) ;
  assign n5505 = ( n5252 & ~n5503 ) | ( n5252 & n5504 ) | ( ~n5503 & n5504 ) ;
  assign n5506 = ( ~n1523 & n5500 ) | ( ~n1523 & n5505 ) | ( n5500 & n5505 ) ;
  assign n5507 = ( n1523 & ~n5253 ) | ( n1523 & n5386 ) | ( ~n5253 & n5386 ) ;
  assign n5508 = n1523 & ~n5253 ;
  assign n5509 = ( n5258 & n5507 ) | ( n5258 & n5508 ) | ( n5507 & n5508 ) ;
  assign n5510 = ( ~n5258 & n5507 ) | ( ~n5258 & n5508 ) | ( n5507 & n5508 ) ;
  assign n5511 = ( n5258 & ~n5509 ) | ( n5258 & n5510 ) | ( ~n5509 & n5510 ) ;
  assign n5512 = ( ~n1393 & n5506 ) | ( ~n1393 & n5511 ) | ( n5506 & n5511 ) ;
  assign n5513 = ~n1393 & n5259 ;
  assign n5514 = ( ~n1393 & n5259 ) | ( ~n1393 & n5386 ) | ( n5259 & n5386 ) ;
  assign n5515 = ( n5264 & n5513 ) | ( n5264 & n5514 ) | ( n5513 & n5514 ) ;
  assign n5516 = ( ~n5264 & n5513 ) | ( ~n5264 & n5514 ) | ( n5513 & n5514 ) ;
  assign n5517 = ( n5264 & ~n5515 ) | ( n5264 & n5516 ) | ( ~n5515 & n5516 ) ;
  assign n5518 = ( ~n1266 & n5512 ) | ( ~n1266 & n5517 ) | ( n5512 & n5517 ) ;
  assign n5519 = ( n1266 & ~n5265 ) | ( n1266 & n5386 ) | ( ~n5265 & n5386 ) ;
  assign n5520 = n1266 & ~n5265 ;
  assign n5521 = ( n5270 & n5519 ) | ( n5270 & n5520 ) | ( n5519 & n5520 ) ;
  assign n5522 = ( ~n5270 & n5519 ) | ( ~n5270 & n5520 ) | ( n5519 & n5520 ) ;
  assign n5523 = ( n5270 & ~n5521 ) | ( n5270 & n5522 ) | ( ~n5521 & n5522 ) ;
  assign n5524 = ( ~n1150 & n5518 ) | ( ~n1150 & n5523 ) | ( n5518 & n5523 ) ;
  assign n5525 = ( n1150 & ~n5271 ) | ( n1150 & n5386 ) | ( ~n5271 & n5386 ) ;
  assign n5526 = n1150 & ~n5271 ;
  assign n5527 = ( n5276 & n5525 ) | ( n5276 & n5526 ) | ( n5525 & n5526 ) ;
  assign n5528 = ( ~n5276 & n5525 ) | ( ~n5276 & n5526 ) | ( n5525 & n5526 ) ;
  assign n5529 = ( n5276 & ~n5527 ) | ( n5276 & n5528 ) | ( ~n5527 & n5528 ) ;
  assign n5530 = ( ~n1038 & n5524 ) | ( ~n1038 & n5529 ) | ( n5524 & n5529 ) ;
  assign n5531 = ( n1038 & ~n5277 ) | ( n1038 & n5386 ) | ( ~n5277 & n5386 ) ;
  assign n5532 = n1038 & ~n5277 ;
  assign n5533 = ( n5282 & n5531 ) | ( n5282 & n5532 ) | ( n5531 & n5532 ) ;
  assign n5534 = ( ~n5282 & n5531 ) | ( ~n5282 & n5532 ) | ( n5531 & n5532 ) ;
  assign n5535 = ( n5282 & ~n5533 ) | ( n5282 & n5534 ) | ( ~n5533 & n5534 ) ;
  assign n5536 = ( ~n933 & n5530 ) | ( ~n933 & n5535 ) | ( n5530 & n5535 ) ;
  assign n5537 = ( n933 & ~n5283 ) | ( n933 & n5386 ) | ( ~n5283 & n5386 ) ;
  assign n5538 = n933 & ~n5283 ;
  assign n5539 = ( n5288 & n5537 ) | ( n5288 & n5538 ) | ( n5537 & n5538 ) ;
  assign n5540 = ( ~n5288 & n5537 ) | ( ~n5288 & n5538 ) | ( n5537 & n5538 ) ;
  assign n5541 = ( n5288 & ~n5539 ) | ( n5288 & n5540 ) | ( ~n5539 & n5540 ) ;
  assign n5542 = ( ~n839 & n5536 ) | ( ~n839 & n5541 ) | ( n5536 & n5541 ) ;
  assign n5543 = ( n839 & ~n5289 ) | ( n839 & n5386 ) | ( ~n5289 & n5386 ) ;
  assign n5544 = n839 & ~n5289 ;
  assign n5545 = ( n5294 & n5543 ) | ( n5294 & n5544 ) | ( n5543 & n5544 ) ;
  assign n5546 = ( ~n5294 & n5543 ) | ( ~n5294 & n5544 ) | ( n5543 & n5544 ) ;
  assign n5547 = ( n5294 & ~n5545 ) | ( n5294 & n5546 ) | ( ~n5545 & n5546 ) ;
  assign n5548 = ( ~n746 & n5542 ) | ( ~n746 & n5547 ) | ( n5542 & n5547 ) ;
  assign n5549 = ( n746 & ~n5295 ) | ( n746 & n5386 ) | ( ~n5295 & n5386 ) ;
  assign n5550 = n746 & ~n5295 ;
  assign n5551 = ( n5300 & n5549 ) | ( n5300 & n5550 ) | ( n5549 & n5550 ) ;
  assign n5552 = ( ~n5300 & n5549 ) | ( ~n5300 & n5550 ) | ( n5549 & n5550 ) ;
  assign n5553 = ( n5300 & ~n5551 ) | ( n5300 & n5552 ) | ( ~n5551 & n5552 ) ;
  assign n5554 = ( ~n664 & n5548 ) | ( ~n664 & n5553 ) | ( n5548 & n5553 ) ;
  assign n5555 = ( n664 & ~n5301 ) | ( n664 & n5386 ) | ( ~n5301 & n5386 ) ;
  assign n5556 = n664 & ~n5301 ;
  assign n5557 = ( n5306 & n5555 ) | ( n5306 & n5556 ) | ( n5555 & n5556 ) ;
  assign n5558 = ( ~n5306 & n5555 ) | ( ~n5306 & n5556 ) | ( n5555 & n5556 ) ;
  assign n5559 = ( n5306 & ~n5557 ) | ( n5306 & n5558 ) | ( ~n5557 & n5558 ) ;
  assign n5560 = ( ~n588 & n5554 ) | ( ~n588 & n5559 ) | ( n5554 & n5559 ) ;
  assign n5561 = ( n588 & ~n5307 ) | ( n588 & n5386 ) | ( ~n5307 & n5386 ) ;
  assign n5562 = n588 & ~n5307 ;
  assign n5563 = ( n5312 & n5561 ) | ( n5312 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5564 = ( ~n5312 & n5561 ) | ( ~n5312 & n5562 ) | ( n5561 & n5562 ) ;
  assign n5565 = ( n5312 & ~n5563 ) | ( n5312 & n5564 ) | ( ~n5563 & n5564 ) ;
  assign n5566 = ( ~n518 & n5560 ) | ( ~n518 & n5565 ) | ( n5560 & n5565 ) ;
  assign n5567 = ~n518 & n5313 ;
  assign n5568 = ( ~n518 & n5313 ) | ( ~n518 & n5386 ) | ( n5313 & n5386 ) ;
  assign n5569 = ( ~n5318 & n5567 ) | ( ~n5318 & n5568 ) | ( n5567 & n5568 ) ;
  assign n5570 = ( n5318 & n5567 ) | ( n5318 & n5568 ) | ( n5567 & n5568 ) ;
  assign n5571 = ( n5318 & n5569 ) | ( n5318 & ~n5570 ) | ( n5569 & ~n5570 ) ;
  assign n5572 = ( ~n454 & n5566 ) | ( ~n454 & n5571 ) | ( n5566 & n5571 ) ;
  assign n5573 = ( n454 & ~n5319 ) | ( n454 & n5386 ) | ( ~n5319 & n5386 ) ;
  assign n5574 = n454 & ~n5319 ;
  assign n5575 = ( n5324 & n5573 ) | ( n5324 & n5574 ) | ( n5573 & n5574 ) ;
  assign n5576 = ( ~n5324 & n5573 ) | ( ~n5324 & n5574 ) | ( n5573 & n5574 ) ;
  assign n5577 = ( n5324 & ~n5575 ) | ( n5324 & n5576 ) | ( ~n5575 & n5576 ) ;
  assign n5578 = ( ~n396 & n5572 ) | ( ~n396 & n5577 ) | ( n5572 & n5577 ) ;
  assign n5579 = ( n396 & ~n5325 ) | ( n396 & n5386 ) | ( ~n5325 & n5386 ) ;
  assign n5580 = n396 & ~n5325 ;
  assign n5581 = ( n5330 & n5579 ) | ( n5330 & n5580 ) | ( n5579 & n5580 ) ;
  assign n5582 = ( ~n5330 & n5579 ) | ( ~n5330 & n5580 ) | ( n5579 & n5580 ) ;
  assign n5583 = ( n5330 & ~n5581 ) | ( n5330 & n5582 ) | ( ~n5581 & n5582 ) ;
  assign n5584 = ( ~n344 & n5578 ) | ( ~n344 & n5583 ) | ( n5578 & n5583 ) ;
  assign n5585 = ( n344 & ~n5331 ) | ( n344 & n5386 ) | ( ~n5331 & n5386 ) ;
  assign n5586 = n344 & ~n5331 ;
  assign n5587 = ( n5336 & n5585 ) | ( n5336 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5588 = ( ~n5336 & n5585 ) | ( ~n5336 & n5586 ) | ( n5585 & n5586 ) ;
  assign n5589 = ( n5336 & ~n5587 ) | ( n5336 & n5588 ) | ( ~n5587 & n5588 ) ;
  assign n5590 = ( ~n298 & n5584 ) | ( ~n298 & n5589 ) | ( n5584 & n5589 ) ;
  assign n5591 = ~n298 & n5337 ;
  assign n5592 = ( ~n298 & n5337 ) | ( ~n298 & n5386 ) | ( n5337 & n5386 ) ;
  assign n5593 = ( ~n5342 & n5591 ) | ( ~n5342 & n5592 ) | ( n5591 & n5592 ) ;
  assign n5594 = ( n5342 & n5591 ) | ( n5342 & n5592 ) | ( n5591 & n5592 ) ;
  assign n5595 = ( n5342 & n5593 ) | ( n5342 & ~n5594 ) | ( n5593 & ~n5594 ) ;
  assign n5596 = ( ~n258 & n5590 ) | ( ~n258 & n5595 ) | ( n5590 & n5595 ) ;
  assign n5597 = ( n258 & ~n5343 ) | ( n258 & n5386 ) | ( ~n5343 & n5386 ) ;
  assign n5598 = n258 & ~n5343 ;
  assign n5599 = ( n5348 & n5597 ) | ( n5348 & n5598 ) | ( n5597 & n5598 ) ;
  assign n5600 = ( ~n5348 & n5597 ) | ( ~n5348 & n5598 ) | ( n5597 & n5598 ) ;
  assign n5601 = ( n5348 & ~n5599 ) | ( n5348 & n5600 ) | ( ~n5599 & n5600 ) ;
  assign n5602 = ( ~n225 & n5596 ) | ( ~n225 & n5601 ) | ( n5596 & n5601 ) ;
  assign n5603 = ( n225 & ~n5349 ) | ( n225 & n5386 ) | ( ~n5349 & n5386 ) ;
  assign n5604 = n225 & ~n5349 ;
  assign n5605 = ( n5354 & n5603 ) | ( n5354 & n5604 ) | ( n5603 & n5604 ) ;
  assign n5606 = ( ~n5354 & n5603 ) | ( ~n5354 & n5604 ) | ( n5603 & n5604 ) ;
  assign n5607 = ( n5354 & ~n5605 ) | ( n5354 & n5606 ) | ( ~n5605 & n5606 ) ;
  assign n5608 = ( ~n197 & n5602 ) | ( ~n197 & n5607 ) | ( n5602 & n5607 ) ;
  assign n5609 = ( n197 & ~n5355 ) | ( n197 & n5386 ) | ( ~n5355 & n5386 ) ;
  assign n5610 = n197 & ~n5355 ;
  assign n5611 = ( n5360 & n5609 ) | ( n5360 & n5610 ) | ( n5609 & n5610 ) ;
  assign n5612 = ( ~n5360 & n5609 ) | ( ~n5360 & n5610 ) | ( n5609 & n5610 ) ;
  assign n5613 = ( n5360 & ~n5611 ) | ( n5360 & n5612 ) | ( ~n5611 & n5612 ) ;
  assign n5614 = ( ~n170 & n5608 ) | ( ~n170 & n5613 ) | ( n5608 & n5613 ) ;
  assign n5615 = ( n170 & ~n5361 ) | ( n170 & n5386 ) | ( ~n5361 & n5386 ) ;
  assign n5616 = n170 & ~n5361 ;
  assign n5617 = ( n5366 & n5615 ) | ( n5366 & n5616 ) | ( n5615 & n5616 ) ;
  assign n5618 = ( ~n5366 & n5615 ) | ( ~n5366 & n5616 ) | ( n5615 & n5616 ) ;
  assign n5619 = ( n5366 & ~n5617 ) | ( n5366 & n5618 ) | ( ~n5617 & n5618 ) ;
  assign n5620 = ( ~n142 & n5614 ) | ( ~n142 & n5619 ) | ( n5614 & n5619 ) ;
  assign n5621 = ~n142 & n5367 ;
  assign n5622 = ( ~n142 & n5367 ) | ( ~n142 & n5386 ) | ( n5367 & n5386 ) ;
  assign n5623 = ( ~n5372 & n5621 ) | ( ~n5372 & n5622 ) | ( n5621 & n5622 ) ;
  assign n5624 = ( n5372 & n5621 ) | ( n5372 & n5622 ) | ( n5621 & n5622 ) ;
  assign n5625 = ( n5372 & n5623 ) | ( n5372 & ~n5624 ) | ( n5623 & ~n5624 ) ;
  assign n5626 = ( ~n132 & n5620 ) | ( ~n132 & n5625 ) | ( n5620 & n5625 ) ;
  assign n5627 = ( n132 & ~n5373 ) | ( n132 & n5386 ) | ( ~n5373 & n5386 ) ;
  assign n5628 = n132 & ~n5373 ;
  assign n5629 = ( n5378 & n5627 ) | ( n5378 & n5628 ) | ( n5627 & n5628 ) ;
  assign n5630 = ( ~n5378 & n5627 ) | ( ~n5378 & n5628 ) | ( n5627 & n5628 ) ;
  assign n5631 = ( n5378 & ~n5629 ) | ( n5378 & n5630 ) | ( ~n5629 & n5630 ) ;
  assign n5632 = ( ~n131 & n5626 ) | ( ~n131 & n5631 ) | ( n5626 & n5631 ) ;
  assign n5633 = n5144 & ~n5384 ;
  assign n5634 = n5379 & ~n5633 ;
  assign n5635 = n5379 & n5384 ;
  assign n5636 = ( n131 & n5145 ) | ( n131 & ~n5384 ) | ( n5145 & ~n5384 ) ;
  assign n5637 = ~n5379 & n5636 ;
  assign n5638 = ( ~n131 & n5635 ) | ( ~n131 & n5637 ) | ( n5635 & n5637 ) ;
  assign n5639 = n5379 | n5384 ;
  assign n5640 = ( n131 & n5634 ) | ( n131 & n5639 ) | ( n5634 & n5639 ) ;
  assign n5641 = ( ~n5634 & n5638 ) | ( ~n5634 & n5640 ) | ( n5638 & n5640 ) ;
  assign n5642 = n5632 | n5641 ;
  assign n5643 = n5626 | n5631 ;
  assign n5644 = ( ~n5631 & n5634 ) | ( ~n5631 & n5639 ) | ( n5634 & n5639 ) ;
  assign n5645 = ~n5634 & n5644 ;
  assign n5646 = n5626 & ~n5645 ;
  assign n5647 = ( n131 & ~n5643 ) | ( n131 & n5646 ) | ( ~n5643 & n5646 ) ;
  assign n5648 = ( n1802 & ~n5488 ) | ( n1802 & n5642 ) | ( ~n5488 & n5642 ) ;
  assign n5649 = n1802 & ~n5488 ;
  assign n5650 = ( n5493 & n5648 ) | ( n5493 & n5649 ) | ( n5648 & n5649 ) ;
  assign n5651 = ( n5493 & ~n5648 ) | ( n5493 & n5649 ) | ( ~n5648 & n5649 ) ;
  assign n5652 = ( n5648 & ~n5650 ) | ( n5648 & n5651 ) | ( ~n5650 & n5651 ) ;
  assign n5653 = ~n5387 & n5642 ;
  assign n5654 = x40 | x41 ;
  assign n5655 = x42 | n5654 ;
  assign n5656 = n5386 & ~n5655 ;
  assign n5657 = ~n5386 & n5655 ;
  assign n5658 = ( x43 & ~n5642 ) | ( x43 & n5657 ) | ( ~n5642 & n5657 ) ;
  assign n5659 = ( n5653 & ~n5656 ) | ( n5653 & n5658 ) | ( ~n5656 & n5658 ) ;
  assign n5660 = n5386 & ~n5642 ;
  assign n5661 = ( ~x44 & n5653 ) | ( ~x44 & n5660 ) | ( n5653 & n5660 ) ;
  assign n5662 = ( x44 & n5653 ) | ( x44 & n5660 ) | ( n5653 & n5660 ) ;
  assign n5663 = ( x44 & n5661 ) | ( x44 & ~n5662 ) | ( n5661 & ~n5662 ) ;
  assign n5664 = ( ~n5139 & n5659 ) | ( ~n5139 & n5663 ) | ( n5659 & n5663 ) ;
  assign n5665 = ~n5139 & n5386 ;
  assign n5666 = ( n5394 & n5642 ) | ( n5394 & n5665 ) | ( n5642 & n5665 ) ;
  assign n5667 = ( x45 & n5661 ) | ( x45 & n5666 ) | ( n5661 & n5666 ) ;
  assign n5668 = ( ~x45 & n5661 ) | ( ~x45 & n5666 ) | ( n5661 & n5666 ) ;
  assign n5669 = ( x45 & ~n5667 ) | ( x45 & n5668 ) | ( ~n5667 & n5668 ) ;
  assign n5670 = ( ~n4898 & n5664 ) | ( ~n4898 & n5669 ) | ( n5664 & n5669 ) ;
  assign n5671 = ( n4898 & ~n5393 ) | ( n4898 & n5642 ) | ( ~n5393 & n5642 ) ;
  assign n5672 = n4898 & ~n5393 ;
  assign n5673 = ( n5397 & n5671 ) | ( n5397 & n5672 ) | ( n5671 & n5672 ) ;
  assign n5674 = ( ~n5397 & n5671 ) | ( ~n5397 & n5672 ) | ( n5671 & n5672 ) ;
  assign n5675 = ( n5397 & ~n5673 ) | ( n5397 & n5674 ) | ( ~n5673 & n5674 ) ;
  assign n5676 = ( ~n4661 & n5670 ) | ( ~n4661 & n5675 ) | ( n5670 & n5675 ) ;
  assign n5677 = ( n4661 & ~n5398 ) | ( n4661 & n5642 ) | ( ~n5398 & n5642 ) ;
  assign n5678 = n4661 & ~n5398 ;
  assign n5679 = ( n5403 & n5677 ) | ( n5403 & n5678 ) | ( n5677 & n5678 ) ;
  assign n5680 = ( ~n5403 & n5677 ) | ( ~n5403 & n5678 ) | ( n5677 & n5678 ) ;
  assign n5681 = ( n5403 & ~n5679 ) | ( n5403 & n5680 ) | ( ~n5679 & n5680 ) ;
  assign n5682 = ( ~n4432 & n5676 ) | ( ~n4432 & n5681 ) | ( n5676 & n5681 ) ;
  assign n5683 = n4432 & ~n5404 ;
  assign n5684 = ( n4432 & ~n5404 ) | ( n4432 & n5642 ) | ( ~n5404 & n5642 ) ;
  assign n5685 = ( n5409 & n5683 ) | ( n5409 & n5684 ) | ( n5683 & n5684 ) ;
  assign n5686 = ( ~n5409 & n5683 ) | ( ~n5409 & n5684 ) | ( n5683 & n5684 ) ;
  assign n5687 = ( n5409 & ~n5685 ) | ( n5409 & n5686 ) | ( ~n5685 & n5686 ) ;
  assign n5688 = ( ~n4203 & n5682 ) | ( ~n4203 & n5687 ) | ( n5682 & n5687 ) ;
  assign n5689 = ~n4203 & n5410 ;
  assign n5690 = ( ~n4203 & n5410 ) | ( ~n4203 & n5642 ) | ( n5410 & n5642 ) ;
  assign n5691 = ( n5415 & n5689 ) | ( n5415 & n5690 ) | ( n5689 & n5690 ) ;
  assign n5692 = ( ~n5415 & n5689 ) | ( ~n5415 & n5690 ) | ( n5689 & n5690 ) ;
  assign n5693 = ( n5415 & ~n5691 ) | ( n5415 & n5692 ) | ( ~n5691 & n5692 ) ;
  assign n5694 = ( ~n3985 & n5688 ) | ( ~n3985 & n5693 ) | ( n5688 & n5693 ) ;
  assign n5695 = ~n3985 & n5416 ;
  assign n5696 = ( ~n3985 & n5416 ) | ( ~n3985 & n5642 ) | ( n5416 & n5642 ) ;
  assign n5697 = ( ~n5421 & n5695 ) | ( ~n5421 & n5696 ) | ( n5695 & n5696 ) ;
  assign n5698 = ( n5421 & n5695 ) | ( n5421 & n5696 ) | ( n5695 & n5696 ) ;
  assign n5699 = ( n5421 & n5697 ) | ( n5421 & ~n5698 ) | ( n5697 & ~n5698 ) ;
  assign n5700 = ( ~n3772 & n5694 ) | ( ~n3772 & n5699 ) | ( n5694 & n5699 ) ;
  assign n5701 = ( n3772 & ~n5422 ) | ( n3772 & n5642 ) | ( ~n5422 & n5642 ) ;
  assign n5702 = n3772 & ~n5422 ;
  assign n5703 = ( n5427 & n5701 ) | ( n5427 & n5702 ) | ( n5701 & n5702 ) ;
  assign n5704 = ( ~n5427 & n5701 ) | ( ~n5427 & n5702 ) | ( n5701 & n5702 ) ;
  assign n5705 = ( n5427 & ~n5703 ) | ( n5427 & n5704 ) | ( ~n5703 & n5704 ) ;
  assign n5706 = ( ~n3567 & n5700 ) | ( ~n3567 & n5705 ) | ( n5700 & n5705 ) ;
  assign n5707 = ( n3567 & ~n5428 ) | ( n3567 & n5642 ) | ( ~n5428 & n5642 ) ;
  assign n5708 = n3567 & ~n5428 ;
  assign n5709 = ( n5433 & n5707 ) | ( n5433 & n5708 ) | ( n5707 & n5708 ) ;
  assign n5710 = ( ~n5433 & n5707 ) | ( ~n5433 & n5708 ) | ( n5707 & n5708 ) ;
  assign n5711 = ( n5433 & ~n5709 ) | ( n5433 & n5710 ) | ( ~n5709 & n5710 ) ;
  assign n5712 = ( ~n3362 & n5706 ) | ( ~n3362 & n5711 ) | ( n5706 & n5711 ) ;
  assign n5713 = ~n3362 & n5434 ;
  assign n5714 = ( ~n3362 & n5434 ) | ( ~n3362 & n5642 ) | ( n5434 & n5642 ) ;
  assign n5715 = ( ~n5439 & n5713 ) | ( ~n5439 & n5714 ) | ( n5713 & n5714 ) ;
  assign n5716 = ( n5439 & n5713 ) | ( n5439 & n5714 ) | ( n5713 & n5714 ) ;
  assign n5717 = ( n5439 & n5715 ) | ( n5439 & ~n5716 ) | ( n5715 & ~n5716 ) ;
  assign n5718 = ( ~n3169 & n5712 ) | ( ~n3169 & n5717 ) | ( n5712 & n5717 ) ;
  assign n5719 = ( n3169 & ~n5440 ) | ( n3169 & n5642 ) | ( ~n5440 & n5642 ) ;
  assign n5720 = n3169 & ~n5440 ;
  assign n5721 = ( n5445 & n5719 ) | ( n5445 & n5720 ) | ( n5719 & n5720 ) ;
  assign n5722 = ( ~n5445 & n5719 ) | ( ~n5445 & n5720 ) | ( n5719 & n5720 ) ;
  assign n5723 = ( n5445 & ~n5721 ) | ( n5445 & n5722 ) | ( ~n5721 & n5722 ) ;
  assign n5724 = ( ~n2979 & n5718 ) | ( ~n2979 & n5723 ) | ( n5718 & n5723 ) ;
  assign n5725 = ~n2979 & n5446 ;
  assign n5726 = ( ~n2979 & n5446 ) | ( ~n2979 & n5642 ) | ( n5446 & n5642 ) ;
  assign n5727 = ( ~n5451 & n5725 ) | ( ~n5451 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5728 = ( n5451 & n5725 ) | ( n5451 & n5726 ) | ( n5725 & n5726 ) ;
  assign n5729 = ( n5451 & n5727 ) | ( n5451 & ~n5728 ) | ( n5727 & ~n5728 ) ;
  assign n5730 = ( ~n2791 & n5724 ) | ( ~n2791 & n5729 ) | ( n5724 & n5729 ) ;
  assign n5731 = ( n2791 & ~n5452 ) | ( n2791 & n5642 ) | ( ~n5452 & n5642 ) ;
  assign n5732 = n2791 & ~n5452 ;
  assign n5733 = ( n5457 & n5731 ) | ( n5457 & n5732 ) | ( n5731 & n5732 ) ;
  assign n5734 = ( ~n5457 & n5731 ) | ( ~n5457 & n5732 ) | ( n5731 & n5732 ) ;
  assign n5735 = ( n5457 & ~n5733 ) | ( n5457 & n5734 ) | ( ~n5733 & n5734 ) ;
  assign n5736 = ( ~n2615 & n5730 ) | ( ~n2615 & n5735 ) | ( n5730 & n5735 ) ;
  assign n5737 = ( n2615 & ~n5458 ) | ( n2615 & n5642 ) | ( ~n5458 & n5642 ) ;
  assign n5738 = n2615 & ~n5458 ;
  assign n5739 = ( n5463 & n5737 ) | ( n5463 & n5738 ) | ( n5737 & n5738 ) ;
  assign n5740 = ( ~n5463 & n5737 ) | ( ~n5463 & n5738 ) | ( n5737 & n5738 ) ;
  assign n5741 = ( n5463 & ~n5739 ) | ( n5463 & n5740 ) | ( ~n5739 & n5740 ) ;
  assign n5742 = ( ~n2443 & n5736 ) | ( ~n2443 & n5741 ) | ( n5736 & n5741 ) ;
  assign n5743 = ( n2443 & ~n5464 ) | ( n2443 & n5642 ) | ( ~n5464 & n5642 ) ;
  assign n5744 = n2443 & ~n5464 ;
  assign n5745 = ( n5469 & n5743 ) | ( n5469 & n5744 ) | ( n5743 & n5744 ) ;
  assign n5746 = ( ~n5469 & n5743 ) | ( ~n5469 & n5744 ) | ( n5743 & n5744 ) ;
  assign n5747 = ( n5469 & ~n5745 ) | ( n5469 & n5746 ) | ( ~n5745 & n5746 ) ;
  assign n5748 = ( ~n2277 & n5742 ) | ( ~n2277 & n5747 ) | ( n5742 & n5747 ) ;
  assign n5749 = ( n2277 & ~n5470 ) | ( n2277 & n5642 ) | ( ~n5470 & n5642 ) ;
  assign n5750 = n2277 & ~n5470 ;
  assign n5751 = ( n5475 & n5749 ) | ( n5475 & n5750 ) | ( n5749 & n5750 ) ;
  assign n5752 = ( ~n5475 & n5749 ) | ( ~n5475 & n5750 ) | ( n5749 & n5750 ) ;
  assign n5753 = ( n5475 & ~n5751 ) | ( n5475 & n5752 ) | ( ~n5751 & n5752 ) ;
  assign n5754 = ( ~n2111 & n5748 ) | ( ~n2111 & n5753 ) | ( n5748 & n5753 ) ;
  assign n5755 = n2111 & ~n5476 ;
  assign n5756 = ( n2111 & ~n5476 ) | ( n2111 & n5642 ) | ( ~n5476 & n5642 ) ;
  assign n5757 = ( n5481 & n5755 ) | ( n5481 & n5756 ) | ( n5755 & n5756 ) ;
  assign n5758 = ( ~n5481 & n5755 ) | ( ~n5481 & n5756 ) | ( n5755 & n5756 ) ;
  assign n5759 = ( n5481 & ~n5757 ) | ( n5481 & n5758 ) | ( ~n5757 & n5758 ) ;
  assign n5760 = ( ~n1949 & n5754 ) | ( ~n1949 & n5759 ) | ( n5754 & n5759 ) ;
  assign n5761 = ( n1949 & ~n5482 ) | ( n1949 & n5642 ) | ( ~n5482 & n5642 ) ;
  assign n5762 = n1949 & ~n5482 ;
  assign n5763 = ( n5487 & n5761 ) | ( n5487 & n5762 ) | ( n5761 & n5762 ) ;
  assign n5764 = ( ~n5487 & n5761 ) | ( ~n5487 & n5762 ) | ( n5761 & n5762 ) ;
  assign n5765 = ( n5487 & ~n5763 ) | ( n5487 & n5764 ) | ( ~n5763 & n5764 ) ;
  assign n5766 = ( ~n1802 & n5760 ) | ( ~n1802 & n5765 ) | ( n5760 & n5765 ) ;
  assign n5767 = ( ~n1661 & n5652 ) | ( ~n1661 & n5766 ) | ( n5652 & n5766 ) ;
  assign n5768 = ( n1661 & ~n5494 ) | ( n1661 & n5642 ) | ( ~n5494 & n5642 ) ;
  assign n5769 = n1661 & ~n5494 ;
  assign n5770 = ( n5499 & n5768 ) | ( n5499 & n5769 ) | ( n5768 & n5769 ) ;
  assign n5771 = ( ~n5499 & n5768 ) | ( ~n5499 & n5769 ) | ( n5768 & n5769 ) ;
  assign n5772 = ( n5499 & ~n5770 ) | ( n5499 & n5771 ) | ( ~n5770 & n5771 ) ;
  assign n5773 = ( ~n1523 & n5767 ) | ( ~n1523 & n5772 ) | ( n5767 & n5772 ) ;
  assign n5774 = ~n1523 & n5500 ;
  assign n5775 = ( ~n1523 & n5500 ) | ( ~n1523 & n5642 ) | ( n5500 & n5642 ) ;
  assign n5776 = ( n5505 & n5774 ) | ( n5505 & n5775 ) | ( n5774 & n5775 ) ;
  assign n5777 = ( ~n5505 & n5774 ) | ( ~n5505 & n5775 ) | ( n5774 & n5775 ) ;
  assign n5778 = ( n5505 & ~n5776 ) | ( n5505 & n5777 ) | ( ~n5776 & n5777 ) ;
  assign n5779 = ( ~n1393 & n5773 ) | ( ~n1393 & n5778 ) | ( n5773 & n5778 ) ;
  assign n5780 = n1393 & ~n5506 ;
  assign n5781 = ( n1393 & ~n5506 ) | ( n1393 & n5642 ) | ( ~n5506 & n5642 ) ;
  assign n5782 = ( n5511 & n5780 ) | ( n5511 & n5781 ) | ( n5780 & n5781 ) ;
  assign n5783 = ( ~n5511 & n5780 ) | ( ~n5511 & n5781 ) | ( n5780 & n5781 ) ;
  assign n5784 = ( n5511 & ~n5782 ) | ( n5511 & n5783 ) | ( ~n5782 & n5783 ) ;
  assign n5785 = ( ~n1266 & n5779 ) | ( ~n1266 & n5784 ) | ( n5779 & n5784 ) ;
  assign n5786 = ( n1266 & ~n5512 ) | ( n1266 & n5642 ) | ( ~n5512 & n5642 ) ;
  assign n5787 = n1266 & ~n5512 ;
  assign n5788 = ( n5517 & n5786 ) | ( n5517 & n5787 ) | ( n5786 & n5787 ) ;
  assign n5789 = ( ~n5517 & n5786 ) | ( ~n5517 & n5787 ) | ( n5786 & n5787 ) ;
  assign n5790 = ( n5517 & ~n5788 ) | ( n5517 & n5789 ) | ( ~n5788 & n5789 ) ;
  assign n5791 = ( ~n1150 & n5785 ) | ( ~n1150 & n5790 ) | ( n5785 & n5790 ) ;
  assign n5792 = ~n1150 & n5518 ;
  assign n5793 = ( ~n1150 & n5518 ) | ( ~n1150 & n5642 ) | ( n5518 & n5642 ) ;
  assign n5794 = ( ~n5523 & n5792 ) | ( ~n5523 & n5793 ) | ( n5792 & n5793 ) ;
  assign n5795 = ( n5523 & n5792 ) | ( n5523 & n5793 ) | ( n5792 & n5793 ) ;
  assign n5796 = ( n5523 & n5794 ) | ( n5523 & ~n5795 ) | ( n5794 & ~n5795 ) ;
  assign n5797 = ( ~n1038 & n5791 ) | ( ~n1038 & n5796 ) | ( n5791 & n5796 ) ;
  assign n5798 = ~n1038 & n5524 ;
  assign n5799 = ( ~n1038 & n5524 ) | ( ~n1038 & n5642 ) | ( n5524 & n5642 ) ;
  assign n5800 = ( ~n5529 & n5798 ) | ( ~n5529 & n5799 ) | ( n5798 & n5799 ) ;
  assign n5801 = ( n5529 & n5798 ) | ( n5529 & n5799 ) | ( n5798 & n5799 ) ;
  assign n5802 = ( n5529 & n5800 ) | ( n5529 & ~n5801 ) | ( n5800 & ~n5801 ) ;
  assign n5803 = ( ~n933 & n5797 ) | ( ~n933 & n5802 ) | ( n5797 & n5802 ) ;
  assign n5804 = ( n933 & ~n5530 ) | ( n933 & n5642 ) | ( ~n5530 & n5642 ) ;
  assign n5805 = n933 & ~n5530 ;
  assign n5806 = ( n5535 & n5804 ) | ( n5535 & n5805 ) | ( n5804 & n5805 ) ;
  assign n5807 = ( ~n5535 & n5804 ) | ( ~n5535 & n5805 ) | ( n5804 & n5805 ) ;
  assign n5808 = ( n5535 & ~n5806 ) | ( n5535 & n5807 ) | ( ~n5806 & n5807 ) ;
  assign n5809 = ( ~n839 & n5803 ) | ( ~n839 & n5808 ) | ( n5803 & n5808 ) ;
  assign n5810 = ~n839 & n5536 ;
  assign n5811 = ( ~n839 & n5536 ) | ( ~n839 & n5642 ) | ( n5536 & n5642 ) ;
  assign n5812 = ( ~n5541 & n5810 ) | ( ~n5541 & n5811 ) | ( n5810 & n5811 ) ;
  assign n5813 = ( n5541 & n5810 ) | ( n5541 & n5811 ) | ( n5810 & n5811 ) ;
  assign n5814 = ( n5541 & n5812 ) | ( n5541 & ~n5813 ) | ( n5812 & ~n5813 ) ;
  assign n5815 = ( ~n746 & n5809 ) | ( ~n746 & n5814 ) | ( n5809 & n5814 ) ;
  assign n5816 = ( n746 & ~n5542 ) | ( n746 & n5642 ) | ( ~n5542 & n5642 ) ;
  assign n5817 = n746 & ~n5542 ;
  assign n5818 = ( n5547 & n5816 ) | ( n5547 & n5817 ) | ( n5816 & n5817 ) ;
  assign n5819 = ( ~n5547 & n5816 ) | ( ~n5547 & n5817 ) | ( n5816 & n5817 ) ;
  assign n5820 = ( n5547 & ~n5818 ) | ( n5547 & n5819 ) | ( ~n5818 & n5819 ) ;
  assign n5821 = ( ~n664 & n5815 ) | ( ~n664 & n5820 ) | ( n5815 & n5820 ) ;
  assign n5822 = ( n664 & ~n5548 ) | ( n664 & n5642 ) | ( ~n5548 & n5642 ) ;
  assign n5823 = n664 & ~n5548 ;
  assign n5824 = ( n5553 & n5822 ) | ( n5553 & n5823 ) | ( n5822 & n5823 ) ;
  assign n5825 = ( ~n5553 & n5822 ) | ( ~n5553 & n5823 ) | ( n5822 & n5823 ) ;
  assign n5826 = ( n5553 & ~n5824 ) | ( n5553 & n5825 ) | ( ~n5824 & n5825 ) ;
  assign n5827 = ( ~n588 & n5821 ) | ( ~n588 & n5826 ) | ( n5821 & n5826 ) ;
  assign n5828 = ( n588 & ~n5554 ) | ( n588 & n5642 ) | ( ~n5554 & n5642 ) ;
  assign n5829 = n588 & ~n5554 ;
  assign n5830 = ( n5559 & n5828 ) | ( n5559 & n5829 ) | ( n5828 & n5829 ) ;
  assign n5831 = ( ~n5559 & n5828 ) | ( ~n5559 & n5829 ) | ( n5828 & n5829 ) ;
  assign n5832 = ( n5559 & ~n5830 ) | ( n5559 & n5831 ) | ( ~n5830 & n5831 ) ;
  assign n5833 = ( ~n518 & n5827 ) | ( ~n518 & n5832 ) | ( n5827 & n5832 ) ;
  assign n5834 = ( n518 & ~n5560 ) | ( n518 & n5642 ) | ( ~n5560 & n5642 ) ;
  assign n5835 = n518 & ~n5560 ;
  assign n5836 = ( n5565 & n5834 ) | ( n5565 & n5835 ) | ( n5834 & n5835 ) ;
  assign n5837 = ( ~n5565 & n5834 ) | ( ~n5565 & n5835 ) | ( n5834 & n5835 ) ;
  assign n5838 = ( n5565 & ~n5836 ) | ( n5565 & n5837 ) | ( ~n5836 & n5837 ) ;
  assign n5839 = ( ~n454 & n5833 ) | ( ~n454 & n5838 ) | ( n5833 & n5838 ) ;
  assign n5840 = n454 & ~n5566 ;
  assign n5841 = ( n454 & ~n5566 ) | ( n454 & n5642 ) | ( ~n5566 & n5642 ) ;
  assign n5842 = ( ~n5571 & n5840 ) | ( ~n5571 & n5841 ) | ( n5840 & n5841 ) ;
  assign n5843 = ( n5571 & n5840 ) | ( n5571 & n5841 ) | ( n5840 & n5841 ) ;
  assign n5844 = ( n5571 & n5842 ) | ( n5571 & ~n5843 ) | ( n5842 & ~n5843 ) ;
  assign n5845 = ( ~n396 & n5839 ) | ( ~n396 & n5844 ) | ( n5839 & n5844 ) ;
  assign n5846 = ( n396 & ~n5572 ) | ( n396 & n5642 ) | ( ~n5572 & n5642 ) ;
  assign n5847 = n396 & ~n5572 ;
  assign n5848 = ( n5577 & n5846 ) | ( n5577 & n5847 ) | ( n5846 & n5847 ) ;
  assign n5849 = ( ~n5577 & n5846 ) | ( ~n5577 & n5847 ) | ( n5846 & n5847 ) ;
  assign n5850 = ( n5577 & ~n5848 ) | ( n5577 & n5849 ) | ( ~n5848 & n5849 ) ;
  assign n5851 = ( ~n344 & n5845 ) | ( ~n344 & n5850 ) | ( n5845 & n5850 ) ;
  assign n5852 = n344 & ~n5578 ;
  assign n5853 = ( n344 & ~n5578 ) | ( n344 & n5642 ) | ( ~n5578 & n5642 ) ;
  assign n5854 = ( n5583 & n5852 ) | ( n5583 & n5853 ) | ( n5852 & n5853 ) ;
  assign n5855 = ( ~n5583 & n5852 ) | ( ~n5583 & n5853 ) | ( n5852 & n5853 ) ;
  assign n5856 = ( n5583 & ~n5854 ) | ( n5583 & n5855 ) | ( ~n5854 & n5855 ) ;
  assign n5857 = ( ~n298 & n5851 ) | ( ~n298 & n5856 ) | ( n5851 & n5856 ) ;
  assign n5858 = ( n298 & ~n5584 ) | ( n298 & n5642 ) | ( ~n5584 & n5642 ) ;
  assign n5859 = n298 & ~n5584 ;
  assign n5860 = ( n5589 & n5858 ) | ( n5589 & n5859 ) | ( n5858 & n5859 ) ;
  assign n5861 = ( ~n5589 & n5858 ) | ( ~n5589 & n5859 ) | ( n5858 & n5859 ) ;
  assign n5862 = ( n5589 & ~n5860 ) | ( n5589 & n5861 ) | ( ~n5860 & n5861 ) ;
  assign n5863 = ( ~n258 & n5857 ) | ( ~n258 & n5862 ) | ( n5857 & n5862 ) ;
  assign n5864 = ( n258 & ~n5590 ) | ( n258 & n5642 ) | ( ~n5590 & n5642 ) ;
  assign n5865 = n258 & ~n5590 ;
  assign n5866 = ( n5595 & n5864 ) | ( n5595 & n5865 ) | ( n5864 & n5865 ) ;
  assign n5867 = ( ~n5595 & n5864 ) | ( ~n5595 & n5865 ) | ( n5864 & n5865 ) ;
  assign n5868 = ( n5595 & ~n5866 ) | ( n5595 & n5867 ) | ( ~n5866 & n5867 ) ;
  assign n5869 = ( ~n225 & n5863 ) | ( ~n225 & n5868 ) | ( n5863 & n5868 ) ;
  assign n5870 = n225 & ~n5596 ;
  assign n5871 = ( n225 & ~n5596 ) | ( n225 & n5642 ) | ( ~n5596 & n5642 ) ;
  assign n5872 = ( n5601 & n5870 ) | ( n5601 & n5871 ) | ( n5870 & n5871 ) ;
  assign n5873 = ( ~n5601 & n5870 ) | ( ~n5601 & n5871 ) | ( n5870 & n5871 ) ;
  assign n5874 = ( n5601 & ~n5872 ) | ( n5601 & n5873 ) | ( ~n5872 & n5873 ) ;
  assign n5875 = ( ~n197 & n5869 ) | ( ~n197 & n5874 ) | ( n5869 & n5874 ) ;
  assign n5876 = ( n197 & ~n5602 ) | ( n197 & n5642 ) | ( ~n5602 & n5642 ) ;
  assign n5877 = n197 & ~n5602 ;
  assign n5878 = ( n5607 & n5876 ) | ( n5607 & n5877 ) | ( n5876 & n5877 ) ;
  assign n5879 = ( ~n5607 & n5876 ) | ( ~n5607 & n5877 ) | ( n5876 & n5877 ) ;
  assign n5880 = ( n5607 & ~n5878 ) | ( n5607 & n5879 ) | ( ~n5878 & n5879 ) ;
  assign n5881 = ( ~n170 & n5875 ) | ( ~n170 & n5880 ) | ( n5875 & n5880 ) ;
  assign n5882 = n170 & ~n5608 ;
  assign n5883 = ( n170 & ~n5608 ) | ( n170 & n5642 ) | ( ~n5608 & n5642 ) ;
  assign n5884 = ( ~n5613 & n5882 ) | ( ~n5613 & n5883 ) | ( n5882 & n5883 ) ;
  assign n5885 = ( n5613 & n5882 ) | ( n5613 & n5883 ) | ( n5882 & n5883 ) ;
  assign n5886 = ( n5613 & n5884 ) | ( n5613 & ~n5885 ) | ( n5884 & ~n5885 ) ;
  assign n5887 = ( ~n142 & n5881 ) | ( ~n142 & n5886 ) | ( n5881 & n5886 ) ;
  assign n5888 = ( n142 & ~n5614 ) | ( n142 & n5642 ) | ( ~n5614 & n5642 ) ;
  assign n5889 = n142 & ~n5614 ;
  assign n5890 = ( n5619 & n5888 ) | ( n5619 & n5889 ) | ( n5888 & n5889 ) ;
  assign n5891 = ( ~n5619 & n5888 ) | ( ~n5619 & n5889 ) | ( n5888 & n5889 ) ;
  assign n5892 = ( n5619 & ~n5890 ) | ( n5619 & n5891 ) | ( ~n5890 & n5891 ) ;
  assign n5893 = ( ~n132 & n5887 ) | ( ~n132 & n5892 ) | ( n5887 & n5892 ) ;
  assign n5894 = ( n132 & ~n5620 ) | ( n132 & n5642 ) | ( ~n5620 & n5642 ) ;
  assign n5895 = n132 & ~n5620 ;
  assign n5896 = ( n5625 & n5894 ) | ( n5625 & n5895 ) | ( n5894 & n5895 ) ;
  assign n5897 = ( ~n5625 & n5894 ) | ( ~n5625 & n5895 ) | ( n5894 & n5895 ) ;
  assign n5898 = ( n5625 & ~n5896 ) | ( n5625 & n5897 ) | ( ~n5896 & n5897 ) ;
  assign n5899 = ~n5626 & n5638 ;
  assign n5900 = n5631 | n5899 ;
  assign n5901 = ~n5626 & n5631 ;
  assign n5902 = ( n5898 & n5900 ) | ( n5898 & ~n5901 ) | ( n5900 & ~n5901 ) ;
  assign n5903 = n131 | n5902 ;
  assign n5904 = ( ~n5647 & n5898 ) | ( ~n5647 & n5903 ) | ( n5898 & n5903 ) ;
  assign n5905 = ( ~n5647 & n5893 ) | ( ~n5647 & n5904 ) | ( n5893 & n5904 ) ;
  assign n5906 = ( ~n131 & n5893 ) | ( ~n131 & n5898 ) | ( n5893 & n5898 ) ;
  assign n5907 = ( n131 & ~n5647 ) | ( n131 & n5898 ) | ( ~n5647 & n5898 ) ;
  assign n5908 = ( n131 & ~n5893 ) | ( n131 & n5898 ) | ( ~n5893 & n5898 ) ;
  assign n5909 = n5907 & ~n5908 ;
  assign n5910 = ( ~n131 & n5898 ) | ( ~n131 & n5902 ) | ( n5898 & n5902 ) ;
  assign n5911 = ( ~n5906 & n5909 ) | ( ~n5906 & n5910 ) | ( n5909 & n5910 ) ;
  assign n5912 = ( n132 & ~n5887 ) | ( n132 & n5905 ) | ( ~n5887 & n5905 ) ;
  assign n5913 = n132 & ~n5887 ;
  assign n5914 = ( n5892 & ~n5912 ) | ( n5892 & n5913 ) | ( ~n5912 & n5913 ) ;
  assign n5915 = ( n5892 & n5912 ) | ( n5892 & n5913 ) | ( n5912 & n5913 ) ;
  assign n5916 = ( n5912 & n5914 ) | ( n5912 & ~n5915 ) | ( n5914 & ~n5915 ) ;
  assign n5917 = ~x41 & n5905 ;
  assign n5918 = x40 & n5917 ;
  assign n5919 = x41 & ~n5905 ;
  assign n5920 = n5917 | n5919 ;
  assign n5921 = x38 | x39 ;
  assign n5922 = x40 | n5921 ;
  assign n5923 = ( ~n5642 & n5920 ) | ( ~n5642 & n5922 ) | ( n5920 & n5922 ) ;
  assign n5924 = ~n5918 & n5923 ;
  assign n5925 = ~n5654 & n5905 ;
  assign n5926 = n5642 & ~n5905 ;
  assign n5927 = ( ~x42 & n5925 ) | ( ~x42 & n5926 ) | ( n5925 & n5926 ) ;
  assign n5928 = ( x42 & n5925 ) | ( x42 & n5926 ) | ( n5925 & n5926 ) ;
  assign n5929 = ( x42 & n5927 ) | ( x42 & ~n5928 ) | ( n5927 & ~n5928 ) ;
  assign n5930 = ( ~n5386 & n5924 ) | ( ~n5386 & n5929 ) | ( n5924 & n5929 ) ;
  assign n5931 = ~n5386 & n5642 ;
  assign n5932 = ( n5660 & n5905 ) | ( n5660 & n5931 ) | ( n5905 & n5931 ) ;
  assign n5933 = ( x43 & n5927 ) | ( x43 & n5932 ) | ( n5927 & n5932 ) ;
  assign n5934 = ( ~x43 & n5927 ) | ( ~x43 & n5932 ) | ( n5927 & n5932 ) ;
  assign n5935 = ( x43 & ~n5933 ) | ( x43 & n5934 ) | ( ~n5933 & n5934 ) ;
  assign n5936 = ( ~n5139 & n5930 ) | ( ~n5139 & n5935 ) | ( n5930 & n5935 ) ;
  assign n5937 = n5139 & ~n5659 ;
  assign n5938 = ( n5139 & ~n5659 ) | ( n5139 & n5905 ) | ( ~n5659 & n5905 ) ;
  assign n5939 = ( n5663 & n5937 ) | ( n5663 & n5938 ) | ( n5937 & n5938 ) ;
  assign n5940 = ( ~n5663 & n5937 ) | ( ~n5663 & n5938 ) | ( n5937 & n5938 ) ;
  assign n5941 = ( n5663 & ~n5939 ) | ( n5663 & n5940 ) | ( ~n5939 & n5940 ) ;
  assign n5942 = ( ~n4898 & n5936 ) | ( ~n4898 & n5941 ) | ( n5936 & n5941 ) ;
  assign n5943 = ( n4898 & ~n5664 ) | ( n4898 & n5905 ) | ( ~n5664 & n5905 ) ;
  assign n5944 = n4898 & ~n5664 ;
  assign n5945 = ( n5669 & n5943 ) | ( n5669 & n5944 ) | ( n5943 & n5944 ) ;
  assign n5946 = ( ~n5669 & n5943 ) | ( ~n5669 & n5944 ) | ( n5943 & n5944 ) ;
  assign n5947 = ( n5669 & ~n5945 ) | ( n5669 & n5946 ) | ( ~n5945 & n5946 ) ;
  assign n5948 = ( ~n4661 & n5942 ) | ( ~n4661 & n5947 ) | ( n5942 & n5947 ) ;
  assign n5949 = ( n4661 & ~n5670 ) | ( n4661 & n5905 ) | ( ~n5670 & n5905 ) ;
  assign n5950 = n4661 & ~n5670 ;
  assign n5951 = ( n5675 & n5949 ) | ( n5675 & n5950 ) | ( n5949 & n5950 ) ;
  assign n5952 = ( ~n5675 & n5949 ) | ( ~n5675 & n5950 ) | ( n5949 & n5950 ) ;
  assign n5953 = ( n5675 & ~n5951 ) | ( n5675 & n5952 ) | ( ~n5951 & n5952 ) ;
  assign n5954 = ( ~n4432 & n5948 ) | ( ~n4432 & n5953 ) | ( n5948 & n5953 ) ;
  assign n5955 = ( n4432 & ~n5676 ) | ( n4432 & n5905 ) | ( ~n5676 & n5905 ) ;
  assign n5956 = n4432 & ~n5676 ;
  assign n5957 = ( n5681 & n5955 ) | ( n5681 & n5956 ) | ( n5955 & n5956 ) ;
  assign n5958 = ( ~n5681 & n5955 ) | ( ~n5681 & n5956 ) | ( n5955 & n5956 ) ;
  assign n5959 = ( n5681 & ~n5957 ) | ( n5681 & n5958 ) | ( ~n5957 & n5958 ) ;
  assign n5960 = ( ~n4203 & n5954 ) | ( ~n4203 & n5959 ) | ( n5954 & n5959 ) ;
  assign n5961 = ( n4203 & ~n5682 ) | ( n4203 & n5905 ) | ( ~n5682 & n5905 ) ;
  assign n5962 = n4203 & ~n5682 ;
  assign n5963 = ( n5687 & n5961 ) | ( n5687 & n5962 ) | ( n5961 & n5962 ) ;
  assign n5964 = ( ~n5687 & n5961 ) | ( ~n5687 & n5962 ) | ( n5961 & n5962 ) ;
  assign n5965 = ( n5687 & ~n5963 ) | ( n5687 & n5964 ) | ( ~n5963 & n5964 ) ;
  assign n5966 = ( ~n3985 & n5960 ) | ( ~n3985 & n5965 ) | ( n5960 & n5965 ) ;
  assign n5967 = ( n3985 & ~n5688 ) | ( n3985 & n5905 ) | ( ~n5688 & n5905 ) ;
  assign n5968 = n3985 & ~n5688 ;
  assign n5969 = ( n5693 & n5967 ) | ( n5693 & n5968 ) | ( n5967 & n5968 ) ;
  assign n5970 = ( ~n5693 & n5967 ) | ( ~n5693 & n5968 ) | ( n5967 & n5968 ) ;
  assign n5971 = ( n5693 & ~n5969 ) | ( n5693 & n5970 ) | ( ~n5969 & n5970 ) ;
  assign n5972 = ( ~n3772 & n5966 ) | ( ~n3772 & n5971 ) | ( n5966 & n5971 ) ;
  assign n5973 = ~n3772 & n5694 ;
  assign n5974 = ( ~n3772 & n5694 ) | ( ~n3772 & n5905 ) | ( n5694 & n5905 ) ;
  assign n5975 = ( ~n5699 & n5973 ) | ( ~n5699 & n5974 ) | ( n5973 & n5974 ) ;
  assign n5976 = ( n5699 & n5973 ) | ( n5699 & n5974 ) | ( n5973 & n5974 ) ;
  assign n5977 = ( n5699 & n5975 ) | ( n5699 & ~n5976 ) | ( n5975 & ~n5976 ) ;
  assign n5978 = ( ~n3567 & n5972 ) | ( ~n3567 & n5977 ) | ( n5972 & n5977 ) ;
  assign n5979 = n3567 & ~n5700 ;
  assign n5980 = ( n3567 & ~n5700 ) | ( n3567 & n5905 ) | ( ~n5700 & n5905 ) ;
  assign n5981 = ( n5705 & n5979 ) | ( n5705 & n5980 ) | ( n5979 & n5980 ) ;
  assign n5982 = ( ~n5705 & n5979 ) | ( ~n5705 & n5980 ) | ( n5979 & n5980 ) ;
  assign n5983 = ( n5705 & ~n5981 ) | ( n5705 & n5982 ) | ( ~n5981 & n5982 ) ;
  assign n5984 = ( ~n3362 & n5978 ) | ( ~n3362 & n5983 ) | ( n5978 & n5983 ) ;
  assign n5985 = ~n3362 & n5706 ;
  assign n5986 = ( ~n3362 & n5706 ) | ( ~n3362 & n5905 ) | ( n5706 & n5905 ) ;
  assign n5987 = ( ~n5711 & n5985 ) | ( ~n5711 & n5986 ) | ( n5985 & n5986 ) ;
  assign n5988 = ( n5711 & n5985 ) | ( n5711 & n5986 ) | ( n5985 & n5986 ) ;
  assign n5989 = ( n5711 & n5987 ) | ( n5711 & ~n5988 ) | ( n5987 & ~n5988 ) ;
  assign n5990 = ( ~n3169 & n5984 ) | ( ~n3169 & n5989 ) | ( n5984 & n5989 ) ;
  assign n5991 = n3169 & ~n5712 ;
  assign n5992 = ( n3169 & ~n5712 ) | ( n3169 & n5905 ) | ( ~n5712 & n5905 ) ;
  assign n5993 = ( n5717 & n5991 ) | ( n5717 & n5992 ) | ( n5991 & n5992 ) ;
  assign n5994 = ( ~n5717 & n5991 ) | ( ~n5717 & n5992 ) | ( n5991 & n5992 ) ;
  assign n5995 = ( n5717 & ~n5993 ) | ( n5717 & n5994 ) | ( ~n5993 & n5994 ) ;
  assign n5996 = ( ~n2979 & n5990 ) | ( ~n2979 & n5995 ) | ( n5990 & n5995 ) ;
  assign n5997 = ~n2979 & n5718 ;
  assign n5998 = ( ~n2979 & n5718 ) | ( ~n2979 & n5905 ) | ( n5718 & n5905 ) ;
  assign n5999 = ( n5723 & n5997 ) | ( n5723 & n5998 ) | ( n5997 & n5998 ) ;
  assign n6000 = ( ~n5723 & n5997 ) | ( ~n5723 & n5998 ) | ( n5997 & n5998 ) ;
  assign n6001 = ( n5723 & ~n5999 ) | ( n5723 & n6000 ) | ( ~n5999 & n6000 ) ;
  assign n6002 = ( ~n2791 & n5996 ) | ( ~n2791 & n6001 ) | ( n5996 & n6001 ) ;
  assign n6003 = ( n2791 & ~n5724 ) | ( n2791 & n5905 ) | ( ~n5724 & n5905 ) ;
  assign n6004 = n2791 & ~n5724 ;
  assign n6005 = ( n5729 & n6003 ) | ( n5729 & n6004 ) | ( n6003 & n6004 ) ;
  assign n6006 = ( ~n5729 & n6003 ) | ( ~n5729 & n6004 ) | ( n6003 & n6004 ) ;
  assign n6007 = ( n5729 & ~n6005 ) | ( n5729 & n6006 ) | ( ~n6005 & n6006 ) ;
  assign n6008 = ( ~n2615 & n6002 ) | ( ~n2615 & n6007 ) | ( n6002 & n6007 ) ;
  assign n6009 = ( n2615 & ~n5730 ) | ( n2615 & n5905 ) | ( ~n5730 & n5905 ) ;
  assign n6010 = n2615 & ~n5730 ;
  assign n6011 = ( n5735 & n6009 ) | ( n5735 & n6010 ) | ( n6009 & n6010 ) ;
  assign n6012 = ( ~n5735 & n6009 ) | ( ~n5735 & n6010 ) | ( n6009 & n6010 ) ;
  assign n6013 = ( n5735 & ~n6011 ) | ( n5735 & n6012 ) | ( ~n6011 & n6012 ) ;
  assign n6014 = ( ~n2443 & n6008 ) | ( ~n2443 & n6013 ) | ( n6008 & n6013 ) ;
  assign n6015 = ~n2443 & n5736 ;
  assign n6016 = ( ~n2443 & n5736 ) | ( ~n2443 & n5905 ) | ( n5736 & n5905 ) ;
  assign n6017 = ( n5741 & n6015 ) | ( n5741 & n6016 ) | ( n6015 & n6016 ) ;
  assign n6018 = ( ~n5741 & n6015 ) | ( ~n5741 & n6016 ) | ( n6015 & n6016 ) ;
  assign n6019 = ( n5741 & ~n6017 ) | ( n5741 & n6018 ) | ( ~n6017 & n6018 ) ;
  assign n6020 = ( ~n2277 & n6014 ) | ( ~n2277 & n6019 ) | ( n6014 & n6019 ) ;
  assign n6021 = ~n2277 & n5742 ;
  assign n6022 = ( ~n2277 & n5742 ) | ( ~n2277 & n5905 ) | ( n5742 & n5905 ) ;
  assign n6023 = ( ~n5747 & n6021 ) | ( ~n5747 & n6022 ) | ( n6021 & n6022 ) ;
  assign n6024 = ( n5747 & n6021 ) | ( n5747 & n6022 ) | ( n6021 & n6022 ) ;
  assign n6025 = ( n5747 & n6023 ) | ( n5747 & ~n6024 ) | ( n6023 & ~n6024 ) ;
  assign n6026 = ( ~n2111 & n6020 ) | ( ~n2111 & n6025 ) | ( n6020 & n6025 ) ;
  assign n6027 = ( n2111 & ~n5748 ) | ( n2111 & n5905 ) | ( ~n5748 & n5905 ) ;
  assign n6028 = n2111 & ~n5748 ;
  assign n6029 = ( n5753 & n6027 ) | ( n5753 & n6028 ) | ( n6027 & n6028 ) ;
  assign n6030 = ( ~n5753 & n6027 ) | ( ~n5753 & n6028 ) | ( n6027 & n6028 ) ;
  assign n6031 = ( n5753 & ~n6029 ) | ( n5753 & n6030 ) | ( ~n6029 & n6030 ) ;
  assign n6032 = ( ~n1949 & n6026 ) | ( ~n1949 & n6031 ) | ( n6026 & n6031 ) ;
  assign n6033 = ~n1949 & n5754 ;
  assign n6034 = ( ~n1949 & n5754 ) | ( ~n1949 & n5905 ) | ( n5754 & n5905 ) ;
  assign n6035 = ( ~n5759 & n6033 ) | ( ~n5759 & n6034 ) | ( n6033 & n6034 ) ;
  assign n6036 = ( n5759 & n6033 ) | ( n5759 & n6034 ) | ( n6033 & n6034 ) ;
  assign n6037 = ( n5759 & n6035 ) | ( n5759 & ~n6036 ) | ( n6035 & ~n6036 ) ;
  assign n6038 = ( ~n1802 & n6032 ) | ( ~n1802 & n6037 ) | ( n6032 & n6037 ) ;
  assign n6039 = ~n1802 & n5760 ;
  assign n6040 = ( ~n1802 & n5760 ) | ( ~n1802 & n5905 ) | ( n5760 & n5905 ) ;
  assign n6041 = ( ~n5765 & n6039 ) | ( ~n5765 & n6040 ) | ( n6039 & n6040 ) ;
  assign n6042 = ( n5765 & n6039 ) | ( n5765 & n6040 ) | ( n6039 & n6040 ) ;
  assign n6043 = ( n5765 & n6041 ) | ( n5765 & ~n6042 ) | ( n6041 & ~n6042 ) ;
  assign n6044 = ( ~n1661 & n6038 ) | ( ~n1661 & n6043 ) | ( n6038 & n6043 ) ;
  assign n6045 = n1661 & ~n5766 ;
  assign n6046 = ( n1661 & ~n5766 ) | ( n1661 & n5905 ) | ( ~n5766 & n5905 ) ;
  assign n6047 = ( ~n5652 & n6045 ) | ( ~n5652 & n6046 ) | ( n6045 & n6046 ) ;
  assign n6048 = ( n5652 & n6045 ) | ( n5652 & n6046 ) | ( n6045 & n6046 ) ;
  assign n6049 = ( n5652 & n6047 ) | ( n5652 & ~n6048 ) | ( n6047 & ~n6048 ) ;
  assign n6050 = ( ~n1523 & n6044 ) | ( ~n1523 & n6049 ) | ( n6044 & n6049 ) ;
  assign n6051 = ( n1523 & ~n5767 ) | ( n1523 & n5905 ) | ( ~n5767 & n5905 ) ;
  assign n6052 = n1523 & ~n5767 ;
  assign n6053 = ( n5772 & n6051 ) | ( n5772 & n6052 ) | ( n6051 & n6052 ) ;
  assign n6054 = ( ~n5772 & n6051 ) | ( ~n5772 & n6052 ) | ( n6051 & n6052 ) ;
  assign n6055 = ( n5772 & ~n6053 ) | ( n5772 & n6054 ) | ( ~n6053 & n6054 ) ;
  assign n6056 = ( ~n1393 & n6050 ) | ( ~n1393 & n6055 ) | ( n6050 & n6055 ) ;
  assign n6057 = n1393 & ~n5773 ;
  assign n6058 = ( n1393 & ~n5773 ) | ( n1393 & n5905 ) | ( ~n5773 & n5905 ) ;
  assign n6059 = ( n5778 & n6057 ) | ( n5778 & n6058 ) | ( n6057 & n6058 ) ;
  assign n6060 = ( ~n5778 & n6057 ) | ( ~n5778 & n6058 ) | ( n6057 & n6058 ) ;
  assign n6061 = ( n5778 & ~n6059 ) | ( n5778 & n6060 ) | ( ~n6059 & n6060 ) ;
  assign n6062 = ( ~n1266 & n6056 ) | ( ~n1266 & n6061 ) | ( n6056 & n6061 ) ;
  assign n6063 = ( n1266 & ~n5779 ) | ( n1266 & n5905 ) | ( ~n5779 & n5905 ) ;
  assign n6064 = n1266 & ~n5779 ;
  assign n6065 = ( n5784 & n6063 ) | ( n5784 & n6064 ) | ( n6063 & n6064 ) ;
  assign n6066 = ( ~n5784 & n6063 ) | ( ~n5784 & n6064 ) | ( n6063 & n6064 ) ;
  assign n6067 = ( n5784 & ~n6065 ) | ( n5784 & n6066 ) | ( ~n6065 & n6066 ) ;
  assign n6068 = ( ~n1150 & n6062 ) | ( ~n1150 & n6067 ) | ( n6062 & n6067 ) ;
  assign n6069 = ( n1150 & ~n5785 ) | ( n1150 & n5905 ) | ( ~n5785 & n5905 ) ;
  assign n6070 = n1150 & ~n5785 ;
  assign n6071 = ( n5790 & n6069 ) | ( n5790 & n6070 ) | ( n6069 & n6070 ) ;
  assign n6072 = ( ~n5790 & n6069 ) | ( ~n5790 & n6070 ) | ( n6069 & n6070 ) ;
  assign n6073 = ( n5790 & ~n6071 ) | ( n5790 & n6072 ) | ( ~n6071 & n6072 ) ;
  assign n6074 = ( ~n1038 & n6068 ) | ( ~n1038 & n6073 ) | ( n6068 & n6073 ) ;
  assign n6075 = ~n1038 & n5791 ;
  assign n6076 = ( ~n1038 & n5791 ) | ( ~n1038 & n5905 ) | ( n5791 & n5905 ) ;
  assign n6077 = ( ~n5796 & n6075 ) | ( ~n5796 & n6076 ) | ( n6075 & n6076 ) ;
  assign n6078 = ( n5796 & n6075 ) | ( n5796 & n6076 ) | ( n6075 & n6076 ) ;
  assign n6079 = ( n5796 & n6077 ) | ( n5796 & ~n6078 ) | ( n6077 & ~n6078 ) ;
  assign n6080 = ( ~n933 & n6074 ) | ( ~n933 & n6079 ) | ( n6074 & n6079 ) ;
  assign n6081 = ~n933 & n5797 ;
  assign n6082 = ( ~n933 & n5797 ) | ( ~n933 & n5905 ) | ( n5797 & n5905 ) ;
  assign n6083 = ( n5802 & n6081 ) | ( n5802 & n6082 ) | ( n6081 & n6082 ) ;
  assign n6084 = ( ~n5802 & n6081 ) | ( ~n5802 & n6082 ) | ( n6081 & n6082 ) ;
  assign n6085 = ( n5802 & ~n6083 ) | ( n5802 & n6084 ) | ( ~n6083 & n6084 ) ;
  assign n6086 = ( ~n839 & n6080 ) | ( ~n839 & n6085 ) | ( n6080 & n6085 ) ;
  assign n6087 = ~n839 & n5803 ;
  assign n6088 = ( ~n839 & n5803 ) | ( ~n839 & n5905 ) | ( n5803 & n5905 ) ;
  assign n6089 = ( ~n5808 & n6087 ) | ( ~n5808 & n6088 ) | ( n6087 & n6088 ) ;
  assign n6090 = ( n5808 & n6087 ) | ( n5808 & n6088 ) | ( n6087 & n6088 ) ;
  assign n6091 = ( n5808 & n6089 ) | ( n5808 & ~n6090 ) | ( n6089 & ~n6090 ) ;
  assign n6092 = ( ~n746 & n6086 ) | ( ~n746 & n6091 ) | ( n6086 & n6091 ) ;
  assign n6093 = ( n746 & ~n5809 ) | ( n746 & n5905 ) | ( ~n5809 & n5905 ) ;
  assign n6094 = n746 & ~n5809 ;
  assign n6095 = ( n5814 & n6093 ) | ( n5814 & n6094 ) | ( n6093 & n6094 ) ;
  assign n6096 = ( ~n5814 & n6093 ) | ( ~n5814 & n6094 ) | ( n6093 & n6094 ) ;
  assign n6097 = ( n5814 & ~n6095 ) | ( n5814 & n6096 ) | ( ~n6095 & n6096 ) ;
  assign n6098 = ( ~n664 & n6092 ) | ( ~n664 & n6097 ) | ( n6092 & n6097 ) ;
  assign n6099 = ( n664 & ~n5815 ) | ( n664 & n5905 ) | ( ~n5815 & n5905 ) ;
  assign n6100 = n664 & ~n5815 ;
  assign n6101 = ( n5820 & n6099 ) | ( n5820 & n6100 ) | ( n6099 & n6100 ) ;
  assign n6102 = ( ~n5820 & n6099 ) | ( ~n5820 & n6100 ) | ( n6099 & n6100 ) ;
  assign n6103 = ( n5820 & ~n6101 ) | ( n5820 & n6102 ) | ( ~n6101 & n6102 ) ;
  assign n6104 = ( ~n588 & n6098 ) | ( ~n588 & n6103 ) | ( n6098 & n6103 ) ;
  assign n6105 = ~n588 & n5821 ;
  assign n6106 = ( ~n588 & n5821 ) | ( ~n588 & n5905 ) | ( n5821 & n5905 ) ;
  assign n6107 = ( ~n5826 & n6105 ) | ( ~n5826 & n6106 ) | ( n6105 & n6106 ) ;
  assign n6108 = ( n5826 & n6105 ) | ( n5826 & n6106 ) | ( n6105 & n6106 ) ;
  assign n6109 = ( n5826 & n6107 ) | ( n5826 & ~n6108 ) | ( n6107 & ~n6108 ) ;
  assign n6110 = ( ~n518 & n6104 ) | ( ~n518 & n6109 ) | ( n6104 & n6109 ) ;
  assign n6111 = ~n518 & n5827 ;
  assign n6112 = ( ~n518 & n5827 ) | ( ~n518 & n5905 ) | ( n5827 & n5905 ) ;
  assign n6113 = ( ~n5832 & n6111 ) | ( ~n5832 & n6112 ) | ( n6111 & n6112 ) ;
  assign n6114 = ( n5832 & n6111 ) | ( n5832 & n6112 ) | ( n6111 & n6112 ) ;
  assign n6115 = ( n5832 & n6113 ) | ( n5832 & ~n6114 ) | ( n6113 & ~n6114 ) ;
  assign n6116 = ( ~n454 & n6110 ) | ( ~n454 & n6115 ) | ( n6110 & n6115 ) ;
  assign n6117 = ( n454 & ~n5833 ) | ( n454 & n5905 ) | ( ~n5833 & n5905 ) ;
  assign n6118 = n454 & ~n5833 ;
  assign n6119 = ( n5838 & n6117 ) | ( n5838 & n6118 ) | ( n6117 & n6118 ) ;
  assign n6120 = ( ~n5838 & n6117 ) | ( ~n5838 & n6118 ) | ( n6117 & n6118 ) ;
  assign n6121 = ( n5838 & ~n6119 ) | ( n5838 & n6120 ) | ( ~n6119 & n6120 ) ;
  assign n6122 = ( ~n396 & n6116 ) | ( ~n396 & n6121 ) | ( n6116 & n6121 ) ;
  assign n6123 = ( n396 & ~n5839 ) | ( n396 & n5905 ) | ( ~n5839 & n5905 ) ;
  assign n6124 = n396 & ~n5839 ;
  assign n6125 = ( n5844 & n6123 ) | ( n5844 & n6124 ) | ( n6123 & n6124 ) ;
  assign n6126 = ( ~n5844 & n6123 ) | ( ~n5844 & n6124 ) | ( n6123 & n6124 ) ;
  assign n6127 = ( n5844 & ~n6125 ) | ( n5844 & n6126 ) | ( ~n6125 & n6126 ) ;
  assign n6128 = ( ~n344 & n6122 ) | ( ~n344 & n6127 ) | ( n6122 & n6127 ) ;
  assign n6129 = ( n344 & ~n5845 ) | ( n344 & n5905 ) | ( ~n5845 & n5905 ) ;
  assign n6130 = n344 & ~n5845 ;
  assign n6131 = ( n5850 & n6129 ) | ( n5850 & n6130 ) | ( n6129 & n6130 ) ;
  assign n6132 = ( ~n5850 & n6129 ) | ( ~n5850 & n6130 ) | ( n6129 & n6130 ) ;
  assign n6133 = ( n5850 & ~n6131 ) | ( n5850 & n6132 ) | ( ~n6131 & n6132 ) ;
  assign n6134 = ( ~n298 & n6128 ) | ( ~n298 & n6133 ) | ( n6128 & n6133 ) ;
  assign n6135 = ( n298 & ~n5851 ) | ( n298 & n5905 ) | ( ~n5851 & n5905 ) ;
  assign n6136 = n298 & ~n5851 ;
  assign n6137 = ( n5856 & n6135 ) | ( n5856 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6138 = ( ~n5856 & n6135 ) | ( ~n5856 & n6136 ) | ( n6135 & n6136 ) ;
  assign n6139 = ( n5856 & ~n6137 ) | ( n5856 & n6138 ) | ( ~n6137 & n6138 ) ;
  assign n6140 = ( ~n258 & n6134 ) | ( ~n258 & n6139 ) | ( n6134 & n6139 ) ;
  assign n6141 = ~n258 & n5857 ;
  assign n6142 = ( ~n258 & n5857 ) | ( ~n258 & n5905 ) | ( n5857 & n5905 ) ;
  assign n6143 = ( n5862 & n6141 ) | ( n5862 & n6142 ) | ( n6141 & n6142 ) ;
  assign n6144 = ( ~n5862 & n6141 ) | ( ~n5862 & n6142 ) | ( n6141 & n6142 ) ;
  assign n6145 = ( n5862 & ~n6143 ) | ( n5862 & n6144 ) | ( ~n6143 & n6144 ) ;
  assign n6146 = ( ~n225 & n6140 ) | ( ~n225 & n6145 ) | ( n6140 & n6145 ) ;
  assign n6147 = n225 & ~n5863 ;
  assign n6148 = ( n225 & ~n5863 ) | ( n225 & n5905 ) | ( ~n5863 & n5905 ) ;
  assign n6149 = ( ~n5868 & n6147 ) | ( ~n5868 & n6148 ) | ( n6147 & n6148 ) ;
  assign n6150 = ( n5868 & n6147 ) | ( n5868 & n6148 ) | ( n6147 & n6148 ) ;
  assign n6151 = ( n5868 & n6149 ) | ( n5868 & ~n6150 ) | ( n6149 & ~n6150 ) ;
  assign n6152 = ( ~n197 & n6146 ) | ( ~n197 & n6151 ) | ( n6146 & n6151 ) ;
  assign n6153 = ~n197 & n5869 ;
  assign n6154 = ( ~n197 & n5869 ) | ( ~n197 & n5905 ) | ( n5869 & n5905 ) ;
  assign n6155 = ( n5874 & n6153 ) | ( n5874 & n6154 ) | ( n6153 & n6154 ) ;
  assign n6156 = ( ~n5874 & n6153 ) | ( ~n5874 & n6154 ) | ( n6153 & n6154 ) ;
  assign n6157 = ( n5874 & ~n6155 ) | ( n5874 & n6156 ) | ( ~n6155 & n6156 ) ;
  assign n6158 = ( ~n170 & n6152 ) | ( ~n170 & n6157 ) | ( n6152 & n6157 ) ;
  assign n6159 = ~n170 & n5875 ;
  assign n6160 = ( ~n170 & n5875 ) | ( ~n170 & n5905 ) | ( n5875 & n5905 ) ;
  assign n6161 = ( ~n5880 & n6159 ) | ( ~n5880 & n6160 ) | ( n6159 & n6160 ) ;
  assign n6162 = ( n5880 & n6159 ) | ( n5880 & n6160 ) | ( n6159 & n6160 ) ;
  assign n6163 = ( n5880 & n6161 ) | ( n5880 & ~n6162 ) | ( n6161 & ~n6162 ) ;
  assign n6164 = ( ~n142 & n6158 ) | ( ~n142 & n6163 ) | ( n6158 & n6163 ) ;
  assign n6165 = ( n142 & ~n5881 ) | ( n142 & n5905 ) | ( ~n5881 & n5905 ) ;
  assign n6166 = n142 & ~n5881 ;
  assign n6167 = ( n5886 & n6165 ) | ( n5886 & n6166 ) | ( n6165 & n6166 ) ;
  assign n6168 = ( ~n5886 & n6165 ) | ( ~n5886 & n6166 ) | ( n6165 & n6166 ) ;
  assign n6169 = ( n5886 & ~n6167 ) | ( n5886 & n6168 ) | ( ~n6167 & n6168 ) ;
  assign n6170 = ( ~n132 & n6164 ) | ( ~n132 & n6169 ) | ( n6164 & n6169 ) ;
  assign n6171 = ( ~n131 & n5916 ) | ( ~n131 & n6170 ) | ( n5916 & n6170 ) ;
  assign n6172 = n5911 | n6171 ;
  assign n6173 = n5911 & ~n5916 ;
  assign n6174 = ( ~n131 & n6170 ) | ( ~n131 & n6173 ) | ( n6170 & n6173 ) ;
  assign n6175 = ( n5916 & ~n6171 ) | ( n5916 & n6174 ) | ( ~n6171 & n6174 ) ;
  assign n6176 = x36 | x37 ;
  assign n6177 = x38 | n6176 ;
  assign n6178 = ( x39 & n6172 ) | ( x39 & ~n6177 ) | ( n6172 & ~n6177 ) ;
  assign n6179 = n5921 & n6172 ;
  assign n6180 = ( n6177 & n6178 ) | ( n6177 & ~n6179 ) | ( n6178 & ~n6179 ) ;
  assign n6181 = x39 | n6172 ;
  assign n6182 = ( n5905 & n6178 ) | ( n5905 & ~n6181 ) | ( n6178 & ~n6181 ) ;
  assign n6183 = n6180 & ~n6182 ;
  assign n6184 = n5905 | n6172 ;
  assign n6185 = ( ~x40 & n6179 ) | ( ~x40 & n6184 ) | ( n6179 & n6184 ) ;
  assign n6186 = ( x40 & n6179 ) | ( x40 & n6184 ) | ( n6179 & n6184 ) ;
  assign n6187 = ( x40 & n6185 ) | ( x40 & ~n6186 ) | ( n6185 & ~n6186 ) ;
  assign n6188 = ( ~n5642 & n6183 ) | ( ~n5642 & n6187 ) | ( n6183 & n6187 ) ;
  assign n6189 = ~n6179 & n6185 ;
  assign n6190 = ~n5642 & n6172 ;
  assign n6191 = n6184 & ~n6190 ;
  assign n6192 = ( ~n5920 & n6189 ) | ( ~n5920 & n6191 ) | ( n6189 & n6191 ) ;
  assign n6193 = ( n5920 & n6189 ) | ( n5920 & n6191 ) | ( n6189 & n6191 ) ;
  assign n6194 = ( n5920 & n6192 ) | ( n5920 & ~n6193 ) | ( n6192 & ~n6193 ) ;
  assign n6195 = ( ~n5386 & n6188 ) | ( ~n5386 & n6194 ) | ( n6188 & n6194 ) ;
  assign n6196 = ( n5386 & n5918 ) | ( n5386 & ~n5923 ) | ( n5918 & ~n5923 ) ;
  assign n6197 = ( n5386 & ~n5924 ) | ( n5386 & n6172 ) | ( ~n5924 & n6172 ) ;
  assign n6198 = ( n5929 & n6196 ) | ( n5929 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6199 = ( ~n5929 & n6196 ) | ( ~n5929 & n6197 ) | ( n6196 & n6197 ) ;
  assign n6200 = ( n5929 & ~n6198 ) | ( n5929 & n6199 ) | ( ~n6198 & n6199 ) ;
  assign n6201 = ( ~n5139 & n6195 ) | ( ~n5139 & n6200 ) | ( n6195 & n6200 ) ;
  assign n6202 = n5139 & ~n5930 ;
  assign n6203 = ( n5139 & ~n5930 ) | ( n5139 & n6172 ) | ( ~n5930 & n6172 ) ;
  assign n6204 = ( ~n5935 & n6202 ) | ( ~n5935 & n6203 ) | ( n6202 & n6203 ) ;
  assign n6205 = ( n5935 & n6202 ) | ( n5935 & n6203 ) | ( n6202 & n6203 ) ;
  assign n6206 = ( n5935 & n6204 ) | ( n5935 & ~n6205 ) | ( n6204 & ~n6205 ) ;
  assign n6207 = ( ~n4898 & n6201 ) | ( ~n4898 & n6206 ) | ( n6201 & n6206 ) ;
  assign n6208 = n4898 & ~n5936 ;
  assign n6209 = ( n4898 & ~n5936 ) | ( n4898 & n6172 ) | ( ~n5936 & n6172 ) ;
  assign n6210 = ( n5941 & n6208 ) | ( n5941 & n6209 ) | ( n6208 & n6209 ) ;
  assign n6211 = ( ~n5941 & n6208 ) | ( ~n5941 & n6209 ) | ( n6208 & n6209 ) ;
  assign n6212 = ( n5941 & ~n6210 ) | ( n5941 & n6211 ) | ( ~n6210 & n6211 ) ;
  assign n6213 = ( ~n4661 & n6207 ) | ( ~n4661 & n6212 ) | ( n6207 & n6212 ) ;
  assign n6214 = ~n4661 & n5942 ;
  assign n6215 = ( ~n4661 & n5942 ) | ( ~n4661 & n6172 ) | ( n5942 & n6172 ) ;
  assign n6216 = ( ~n5947 & n6214 ) | ( ~n5947 & n6215 ) | ( n6214 & n6215 ) ;
  assign n6217 = ( n5947 & n6214 ) | ( n5947 & n6215 ) | ( n6214 & n6215 ) ;
  assign n6218 = ( n5947 & n6216 ) | ( n5947 & ~n6217 ) | ( n6216 & ~n6217 ) ;
  assign n6219 = ( ~n4432 & n6213 ) | ( ~n4432 & n6218 ) | ( n6213 & n6218 ) ;
  assign n6220 = n4432 & ~n5948 ;
  assign n6221 = ( n4432 & ~n5948 ) | ( n4432 & n6172 ) | ( ~n5948 & n6172 ) ;
  assign n6222 = ( n5953 & n6220 ) | ( n5953 & n6221 ) | ( n6220 & n6221 ) ;
  assign n6223 = ( ~n5953 & n6220 ) | ( ~n5953 & n6221 ) | ( n6220 & n6221 ) ;
  assign n6224 = ( n5953 & ~n6222 ) | ( n5953 & n6223 ) | ( ~n6222 & n6223 ) ;
  assign n6225 = ( ~n4203 & n6219 ) | ( ~n4203 & n6224 ) | ( n6219 & n6224 ) ;
  assign n6226 = ~n4203 & n5954 ;
  assign n6227 = ( ~n4203 & n5954 ) | ( ~n4203 & n6172 ) | ( n5954 & n6172 ) ;
  assign n6228 = ( n5959 & n6226 ) | ( n5959 & n6227 ) | ( n6226 & n6227 ) ;
  assign n6229 = ( ~n5959 & n6226 ) | ( ~n5959 & n6227 ) | ( n6226 & n6227 ) ;
  assign n6230 = ( n5959 & ~n6228 ) | ( n5959 & n6229 ) | ( ~n6228 & n6229 ) ;
  assign n6231 = ( ~n3985 & n6225 ) | ( ~n3985 & n6230 ) | ( n6225 & n6230 ) ;
  assign n6232 = ( n3985 & ~n5960 ) | ( n3985 & n6172 ) | ( ~n5960 & n6172 ) ;
  assign n6233 = n3985 & ~n5960 ;
  assign n6234 = ( n5965 & n6232 ) | ( n5965 & n6233 ) | ( n6232 & n6233 ) ;
  assign n6235 = ( ~n5965 & n6232 ) | ( ~n5965 & n6233 ) | ( n6232 & n6233 ) ;
  assign n6236 = ( n5965 & ~n6234 ) | ( n5965 & n6235 ) | ( ~n6234 & n6235 ) ;
  assign n6237 = ( ~n3772 & n6231 ) | ( ~n3772 & n6236 ) | ( n6231 & n6236 ) ;
  assign n6238 = ~n3772 & n5966 ;
  assign n6239 = ( ~n3772 & n5966 ) | ( ~n3772 & n6172 ) | ( n5966 & n6172 ) ;
  assign n6240 = ( ~n5971 & n6238 ) | ( ~n5971 & n6239 ) | ( n6238 & n6239 ) ;
  assign n6241 = ( n5971 & n6238 ) | ( n5971 & n6239 ) | ( n6238 & n6239 ) ;
  assign n6242 = ( n5971 & n6240 ) | ( n5971 & ~n6241 ) | ( n6240 & ~n6241 ) ;
  assign n6243 = ( ~n3567 & n6237 ) | ( ~n3567 & n6242 ) | ( n6237 & n6242 ) ;
  assign n6244 = ( n3567 & ~n5972 ) | ( n3567 & n6172 ) | ( ~n5972 & n6172 ) ;
  assign n6245 = n3567 & ~n5972 ;
  assign n6246 = ( n5977 & n6244 ) | ( n5977 & n6245 ) | ( n6244 & n6245 ) ;
  assign n6247 = ( ~n5977 & n6244 ) | ( ~n5977 & n6245 ) | ( n6244 & n6245 ) ;
  assign n6248 = ( n5977 & ~n6246 ) | ( n5977 & n6247 ) | ( ~n6246 & n6247 ) ;
  assign n6249 = ( ~n3362 & n6243 ) | ( ~n3362 & n6248 ) | ( n6243 & n6248 ) ;
  assign n6250 = ~n3362 & n5978 ;
  assign n6251 = ( ~n3362 & n5978 ) | ( ~n3362 & n6172 ) | ( n5978 & n6172 ) ;
  assign n6252 = ( ~n5983 & n6250 ) | ( ~n5983 & n6251 ) | ( n6250 & n6251 ) ;
  assign n6253 = ( n5983 & n6250 ) | ( n5983 & n6251 ) | ( n6250 & n6251 ) ;
  assign n6254 = ( n5983 & n6252 ) | ( n5983 & ~n6253 ) | ( n6252 & ~n6253 ) ;
  assign n6255 = ( ~n3169 & n6249 ) | ( ~n3169 & n6254 ) | ( n6249 & n6254 ) ;
  assign n6256 = ( n3169 & ~n5984 ) | ( n3169 & n6172 ) | ( ~n5984 & n6172 ) ;
  assign n6257 = n3169 & ~n5984 ;
  assign n6258 = ( n5989 & n6256 ) | ( n5989 & n6257 ) | ( n6256 & n6257 ) ;
  assign n6259 = ( ~n5989 & n6256 ) | ( ~n5989 & n6257 ) | ( n6256 & n6257 ) ;
  assign n6260 = ( n5989 & ~n6258 ) | ( n5989 & n6259 ) | ( ~n6258 & n6259 ) ;
  assign n6261 = ( ~n2979 & n6255 ) | ( ~n2979 & n6260 ) | ( n6255 & n6260 ) ;
  assign n6262 = n2979 & ~n5990 ;
  assign n6263 = ( n2979 & ~n5990 ) | ( n2979 & n6172 ) | ( ~n5990 & n6172 ) ;
  assign n6264 = ( n5995 & n6262 ) | ( n5995 & n6263 ) | ( n6262 & n6263 ) ;
  assign n6265 = ( ~n5995 & n6262 ) | ( ~n5995 & n6263 ) | ( n6262 & n6263 ) ;
  assign n6266 = ( n5995 & ~n6264 ) | ( n5995 & n6265 ) | ( ~n6264 & n6265 ) ;
  assign n6267 = ( ~n2791 & n6261 ) | ( ~n2791 & n6266 ) | ( n6261 & n6266 ) ;
  assign n6268 = ( n2791 & ~n5996 ) | ( n2791 & n6172 ) | ( ~n5996 & n6172 ) ;
  assign n6269 = n2791 & ~n5996 ;
  assign n6270 = ( n6001 & n6268 ) | ( n6001 & n6269 ) | ( n6268 & n6269 ) ;
  assign n6271 = ( ~n6001 & n6268 ) | ( ~n6001 & n6269 ) | ( n6268 & n6269 ) ;
  assign n6272 = ( n6001 & ~n6270 ) | ( n6001 & n6271 ) | ( ~n6270 & n6271 ) ;
  assign n6273 = ( ~n2615 & n6267 ) | ( ~n2615 & n6272 ) | ( n6267 & n6272 ) ;
  assign n6274 = ~n2615 & n6002 ;
  assign n6275 = ( ~n2615 & n6002 ) | ( ~n2615 & n6172 ) | ( n6002 & n6172 ) ;
  assign n6276 = ( ~n6007 & n6274 ) | ( ~n6007 & n6275 ) | ( n6274 & n6275 ) ;
  assign n6277 = ( n6007 & n6274 ) | ( n6007 & n6275 ) | ( n6274 & n6275 ) ;
  assign n6278 = ( n6007 & n6276 ) | ( n6007 & ~n6277 ) | ( n6276 & ~n6277 ) ;
  assign n6279 = ( ~n2443 & n6273 ) | ( ~n2443 & n6278 ) | ( n6273 & n6278 ) ;
  assign n6280 = n2443 & ~n6008 ;
  assign n6281 = ( n2443 & ~n6008 ) | ( n2443 & n6172 ) | ( ~n6008 & n6172 ) ;
  assign n6282 = ( ~n6013 & n6280 ) | ( ~n6013 & n6281 ) | ( n6280 & n6281 ) ;
  assign n6283 = ( n6013 & n6280 ) | ( n6013 & n6281 ) | ( n6280 & n6281 ) ;
  assign n6284 = ( n6013 & n6282 ) | ( n6013 & ~n6283 ) | ( n6282 & ~n6283 ) ;
  assign n6285 = ( ~n2277 & n6279 ) | ( ~n2277 & n6284 ) | ( n6279 & n6284 ) ;
  assign n6286 = ~n2277 & n6014 ;
  assign n6287 = ( ~n2277 & n6014 ) | ( ~n2277 & n6172 ) | ( n6014 & n6172 ) ;
  assign n6288 = ( ~n6019 & n6286 ) | ( ~n6019 & n6287 ) | ( n6286 & n6287 ) ;
  assign n6289 = ( n6019 & n6286 ) | ( n6019 & n6287 ) | ( n6286 & n6287 ) ;
  assign n6290 = ( n6019 & n6288 ) | ( n6019 & ~n6289 ) | ( n6288 & ~n6289 ) ;
  assign n6291 = ( ~n2111 & n6285 ) | ( ~n2111 & n6290 ) | ( n6285 & n6290 ) ;
  assign n6292 = ( n2111 & ~n6020 ) | ( n2111 & n6172 ) | ( ~n6020 & n6172 ) ;
  assign n6293 = n2111 & ~n6020 ;
  assign n6294 = ( n6025 & n6292 ) | ( n6025 & n6293 ) | ( n6292 & n6293 ) ;
  assign n6295 = ( ~n6025 & n6292 ) | ( ~n6025 & n6293 ) | ( n6292 & n6293 ) ;
  assign n6296 = ( n6025 & ~n6294 ) | ( n6025 & n6295 ) | ( ~n6294 & n6295 ) ;
  assign n6297 = ( ~n1949 & n6291 ) | ( ~n1949 & n6296 ) | ( n6291 & n6296 ) ;
  assign n6298 = ~n1949 & n6026 ;
  assign n6299 = ( ~n1949 & n6026 ) | ( ~n1949 & n6172 ) | ( n6026 & n6172 ) ;
  assign n6300 = ( ~n6031 & n6298 ) | ( ~n6031 & n6299 ) | ( n6298 & n6299 ) ;
  assign n6301 = ( n6031 & n6298 ) | ( n6031 & n6299 ) | ( n6298 & n6299 ) ;
  assign n6302 = ( n6031 & n6300 ) | ( n6031 & ~n6301 ) | ( n6300 & ~n6301 ) ;
  assign n6303 = ( ~n1802 & n6297 ) | ( ~n1802 & n6302 ) | ( n6297 & n6302 ) ;
  assign n6304 = n1802 & ~n6032 ;
  assign n6305 = ( n1802 & ~n6032 ) | ( n1802 & n6172 ) | ( ~n6032 & n6172 ) ;
  assign n6306 = ( n6037 & n6304 ) | ( n6037 & n6305 ) | ( n6304 & n6305 ) ;
  assign n6307 = ( ~n6037 & n6304 ) | ( ~n6037 & n6305 ) | ( n6304 & n6305 ) ;
  assign n6308 = ( n6037 & ~n6306 ) | ( n6037 & n6307 ) | ( ~n6306 & n6307 ) ;
  assign n6309 = ( ~n1661 & n6303 ) | ( ~n1661 & n6308 ) | ( n6303 & n6308 ) ;
  assign n6310 = n1661 & ~n6038 ;
  assign n6311 = ( n1661 & ~n6038 ) | ( n1661 & n6172 ) | ( ~n6038 & n6172 ) ;
  assign n6312 = ( n6043 & n6310 ) | ( n6043 & n6311 ) | ( n6310 & n6311 ) ;
  assign n6313 = ( ~n6043 & n6310 ) | ( ~n6043 & n6311 ) | ( n6310 & n6311 ) ;
  assign n6314 = ( n6043 & ~n6312 ) | ( n6043 & n6313 ) | ( ~n6312 & n6313 ) ;
  assign n6315 = ( ~n1523 & n6309 ) | ( ~n1523 & n6314 ) | ( n6309 & n6314 ) ;
  assign n6316 = ~n1523 & n6044 ;
  assign n6317 = ( ~n1523 & n6044 ) | ( ~n1523 & n6172 ) | ( n6044 & n6172 ) ;
  assign n6318 = ( ~n6049 & n6316 ) | ( ~n6049 & n6317 ) | ( n6316 & n6317 ) ;
  assign n6319 = ( n6049 & n6316 ) | ( n6049 & n6317 ) | ( n6316 & n6317 ) ;
  assign n6320 = ( n6049 & n6318 ) | ( n6049 & ~n6319 ) | ( n6318 & ~n6319 ) ;
  assign n6321 = ( ~n1393 & n6315 ) | ( ~n1393 & n6320 ) | ( n6315 & n6320 ) ;
  assign n6322 = ( n1393 & ~n6050 ) | ( n1393 & n6172 ) | ( ~n6050 & n6172 ) ;
  assign n6323 = n1393 & ~n6050 ;
  assign n6324 = ( n6055 & n6322 ) | ( n6055 & n6323 ) | ( n6322 & n6323 ) ;
  assign n6325 = ( ~n6055 & n6322 ) | ( ~n6055 & n6323 ) | ( n6322 & n6323 ) ;
  assign n6326 = ( n6055 & ~n6324 ) | ( n6055 & n6325 ) | ( ~n6324 & n6325 ) ;
  assign n6327 = ( ~n1266 & n6321 ) | ( ~n1266 & n6326 ) | ( n6321 & n6326 ) ;
  assign n6328 = ~n1266 & n6056 ;
  assign n6329 = ( ~n1266 & n6056 ) | ( ~n1266 & n6172 ) | ( n6056 & n6172 ) ;
  assign n6330 = ( ~n6061 & n6328 ) | ( ~n6061 & n6329 ) | ( n6328 & n6329 ) ;
  assign n6331 = ( n6061 & n6328 ) | ( n6061 & n6329 ) | ( n6328 & n6329 ) ;
  assign n6332 = ( n6061 & n6330 ) | ( n6061 & ~n6331 ) | ( n6330 & ~n6331 ) ;
  assign n6333 = ( ~n1150 & n6327 ) | ( ~n1150 & n6332 ) | ( n6327 & n6332 ) ;
  assign n6334 = ~n1150 & n6062 ;
  assign n6335 = ( ~n1150 & n6062 ) | ( ~n1150 & n6172 ) | ( n6062 & n6172 ) ;
  assign n6336 = ( ~n6067 & n6334 ) | ( ~n6067 & n6335 ) | ( n6334 & n6335 ) ;
  assign n6337 = ( n6067 & n6334 ) | ( n6067 & n6335 ) | ( n6334 & n6335 ) ;
  assign n6338 = ( n6067 & n6336 ) | ( n6067 & ~n6337 ) | ( n6336 & ~n6337 ) ;
  assign n6339 = ( ~n1038 & n6333 ) | ( ~n1038 & n6338 ) | ( n6333 & n6338 ) ;
  assign n6340 = ( n1038 & ~n6068 ) | ( n1038 & n6172 ) | ( ~n6068 & n6172 ) ;
  assign n6341 = n1038 & ~n6068 ;
  assign n6342 = ( n6073 & n6340 ) | ( n6073 & n6341 ) | ( n6340 & n6341 ) ;
  assign n6343 = ( ~n6073 & n6340 ) | ( ~n6073 & n6341 ) | ( n6340 & n6341 ) ;
  assign n6344 = ( n6073 & ~n6342 ) | ( n6073 & n6343 ) | ( ~n6342 & n6343 ) ;
  assign n6345 = ( ~n933 & n6339 ) | ( ~n933 & n6344 ) | ( n6339 & n6344 ) ;
  assign n6346 = ( n933 & ~n6074 ) | ( n933 & n6172 ) | ( ~n6074 & n6172 ) ;
  assign n6347 = n933 & ~n6074 ;
  assign n6348 = ( n6079 & n6346 ) | ( n6079 & n6347 ) | ( n6346 & n6347 ) ;
  assign n6349 = ( ~n6079 & n6346 ) | ( ~n6079 & n6347 ) | ( n6346 & n6347 ) ;
  assign n6350 = ( n6079 & ~n6348 ) | ( n6079 & n6349 ) | ( ~n6348 & n6349 ) ;
  assign n6351 = ( ~n839 & n6345 ) | ( ~n839 & n6350 ) | ( n6345 & n6350 ) ;
  assign n6352 = n839 & ~n6080 ;
  assign n6353 = ( n839 & ~n6080 ) | ( n839 & n6172 ) | ( ~n6080 & n6172 ) ;
  assign n6354 = ( ~n6085 & n6352 ) | ( ~n6085 & n6353 ) | ( n6352 & n6353 ) ;
  assign n6355 = ( n6085 & n6352 ) | ( n6085 & n6353 ) | ( n6352 & n6353 ) ;
  assign n6356 = ( n6085 & n6354 ) | ( n6085 & ~n6355 ) | ( n6354 & ~n6355 ) ;
  assign n6357 = ( ~n746 & n6351 ) | ( ~n746 & n6356 ) | ( n6351 & n6356 ) ;
  assign n6358 = ( n746 & ~n6086 ) | ( n746 & n6172 ) | ( ~n6086 & n6172 ) ;
  assign n6359 = n746 & ~n6086 ;
  assign n6360 = ( n6091 & n6358 ) | ( n6091 & n6359 ) | ( n6358 & n6359 ) ;
  assign n6361 = ( ~n6091 & n6358 ) | ( ~n6091 & n6359 ) | ( n6358 & n6359 ) ;
  assign n6362 = ( n6091 & ~n6360 ) | ( n6091 & n6361 ) | ( ~n6360 & n6361 ) ;
  assign n6363 = ( ~n664 & n6357 ) | ( ~n664 & n6362 ) | ( n6357 & n6362 ) ;
  assign n6364 = ~n664 & n6092 ;
  assign n6365 = ( ~n664 & n6092 ) | ( ~n664 & n6172 ) | ( n6092 & n6172 ) ;
  assign n6366 = ( ~n6097 & n6364 ) | ( ~n6097 & n6365 ) | ( n6364 & n6365 ) ;
  assign n6367 = ( n6097 & n6364 ) | ( n6097 & n6365 ) | ( n6364 & n6365 ) ;
  assign n6368 = ( n6097 & n6366 ) | ( n6097 & ~n6367 ) | ( n6366 & ~n6367 ) ;
  assign n6369 = ( ~n588 & n6363 ) | ( ~n588 & n6368 ) | ( n6363 & n6368 ) ;
  assign n6370 = ( n588 & ~n6098 ) | ( n588 & n6172 ) | ( ~n6098 & n6172 ) ;
  assign n6371 = n588 & ~n6098 ;
  assign n6372 = ( n6103 & n6370 ) | ( n6103 & n6371 ) | ( n6370 & n6371 ) ;
  assign n6373 = ( ~n6103 & n6370 ) | ( ~n6103 & n6371 ) | ( n6370 & n6371 ) ;
  assign n6374 = ( n6103 & ~n6372 ) | ( n6103 & n6373 ) | ( ~n6372 & n6373 ) ;
  assign n6375 = ( ~n518 & n6369 ) | ( ~n518 & n6374 ) | ( n6369 & n6374 ) ;
  assign n6376 = ~n518 & n6104 ;
  assign n6377 = ( ~n518 & n6104 ) | ( ~n518 & n6172 ) | ( n6104 & n6172 ) ;
  assign n6378 = ( ~n6109 & n6376 ) | ( ~n6109 & n6377 ) | ( n6376 & n6377 ) ;
  assign n6379 = ( n6109 & n6376 ) | ( n6109 & n6377 ) | ( n6376 & n6377 ) ;
  assign n6380 = ( n6109 & n6378 ) | ( n6109 & ~n6379 ) | ( n6378 & ~n6379 ) ;
  assign n6381 = ( ~n454 & n6375 ) | ( ~n454 & n6380 ) | ( n6375 & n6380 ) ;
  assign n6382 = ( n454 & ~n6110 ) | ( n454 & n6172 ) | ( ~n6110 & n6172 ) ;
  assign n6383 = n454 & ~n6110 ;
  assign n6384 = ( n6115 & n6382 ) | ( n6115 & n6383 ) | ( n6382 & n6383 ) ;
  assign n6385 = ( ~n6115 & n6382 ) | ( ~n6115 & n6383 ) | ( n6382 & n6383 ) ;
  assign n6386 = ( n6115 & ~n6384 ) | ( n6115 & n6385 ) | ( ~n6384 & n6385 ) ;
  assign n6387 = ( ~n396 & n6381 ) | ( ~n396 & n6386 ) | ( n6381 & n6386 ) ;
  assign n6388 = ( n396 & ~n6116 ) | ( n396 & n6172 ) | ( ~n6116 & n6172 ) ;
  assign n6389 = n396 & ~n6116 ;
  assign n6390 = ( n6121 & n6388 ) | ( n6121 & n6389 ) | ( n6388 & n6389 ) ;
  assign n6391 = ( ~n6121 & n6388 ) | ( ~n6121 & n6389 ) | ( n6388 & n6389 ) ;
  assign n6392 = ( n6121 & ~n6390 ) | ( n6121 & n6391 ) | ( ~n6390 & n6391 ) ;
  assign n6393 = ( ~n344 & n6387 ) | ( ~n344 & n6392 ) | ( n6387 & n6392 ) ;
  assign n6394 = ( n344 & ~n6122 ) | ( n344 & n6172 ) | ( ~n6122 & n6172 ) ;
  assign n6395 = n344 & ~n6122 ;
  assign n6396 = ( n6127 & n6394 ) | ( n6127 & n6395 ) | ( n6394 & n6395 ) ;
  assign n6397 = ( ~n6127 & n6394 ) | ( ~n6127 & n6395 ) | ( n6394 & n6395 ) ;
  assign n6398 = ( n6127 & ~n6396 ) | ( n6127 & n6397 ) | ( ~n6396 & n6397 ) ;
  assign n6399 = ( ~n298 & n6393 ) | ( ~n298 & n6398 ) | ( n6393 & n6398 ) ;
  assign n6400 = ( n298 & ~n6128 ) | ( n298 & n6172 ) | ( ~n6128 & n6172 ) ;
  assign n6401 = n298 & ~n6128 ;
  assign n6402 = ( n6133 & n6400 ) | ( n6133 & n6401 ) | ( n6400 & n6401 ) ;
  assign n6403 = ( ~n6133 & n6400 ) | ( ~n6133 & n6401 ) | ( n6400 & n6401 ) ;
  assign n6404 = ( n6133 & ~n6402 ) | ( n6133 & n6403 ) | ( ~n6402 & n6403 ) ;
  assign n6405 = ( ~n258 & n6399 ) | ( ~n258 & n6404 ) | ( n6399 & n6404 ) ;
  assign n6406 = ( n258 & ~n6134 ) | ( n258 & n6172 ) | ( ~n6134 & n6172 ) ;
  assign n6407 = n258 & ~n6134 ;
  assign n6408 = ( n6139 & n6406 ) | ( n6139 & n6407 ) | ( n6406 & n6407 ) ;
  assign n6409 = ( ~n6139 & n6406 ) | ( ~n6139 & n6407 ) | ( n6406 & n6407 ) ;
  assign n6410 = ( n6139 & ~n6408 ) | ( n6139 & n6409 ) | ( ~n6408 & n6409 ) ;
  assign n6411 = ( ~n225 & n6405 ) | ( ~n225 & n6410 ) | ( n6405 & n6410 ) ;
  assign n6412 = ~n225 & n6140 ;
  assign n6413 = ( ~n225 & n6140 ) | ( ~n225 & n6172 ) | ( n6140 & n6172 ) ;
  assign n6414 = ( ~n6145 & n6412 ) | ( ~n6145 & n6413 ) | ( n6412 & n6413 ) ;
  assign n6415 = ( n6145 & n6412 ) | ( n6145 & n6413 ) | ( n6412 & n6413 ) ;
  assign n6416 = ( n6145 & n6414 ) | ( n6145 & ~n6415 ) | ( n6414 & ~n6415 ) ;
  assign n6417 = ( ~n197 & n6411 ) | ( ~n197 & n6416 ) | ( n6411 & n6416 ) ;
  assign n6418 = n197 & ~n6146 ;
  assign n6419 = ( n197 & ~n6146 ) | ( n197 & n6172 ) | ( ~n6146 & n6172 ) ;
  assign n6420 = ( ~n6151 & n6418 ) | ( ~n6151 & n6419 ) | ( n6418 & n6419 ) ;
  assign n6421 = ( n6151 & n6418 ) | ( n6151 & n6419 ) | ( n6418 & n6419 ) ;
  assign n6422 = ( n6151 & n6420 ) | ( n6151 & ~n6421 ) | ( n6420 & ~n6421 ) ;
  assign n6423 = ( ~n170 & n6417 ) | ( ~n170 & n6422 ) | ( n6417 & n6422 ) ;
  assign n6424 = ( n170 & ~n6152 ) | ( n170 & n6172 ) | ( ~n6152 & n6172 ) ;
  assign n6425 = n170 & ~n6152 ;
  assign n6426 = ( n6157 & n6424 ) | ( n6157 & n6425 ) | ( n6424 & n6425 ) ;
  assign n6427 = ( ~n6157 & n6424 ) | ( ~n6157 & n6425 ) | ( n6424 & n6425 ) ;
  assign n6428 = ( n6157 & ~n6426 ) | ( n6157 & n6427 ) | ( ~n6426 & n6427 ) ;
  assign n6429 = ( ~n142 & n6423 ) | ( ~n142 & n6428 ) | ( n6423 & n6428 ) ;
  assign n6430 = ~n142 & n6158 ;
  assign n6431 = ( ~n142 & n6158 ) | ( ~n142 & n6172 ) | ( n6158 & n6172 ) ;
  assign n6432 = ( ~n6163 & n6430 ) | ( ~n6163 & n6431 ) | ( n6430 & n6431 ) ;
  assign n6433 = ( n6163 & n6430 ) | ( n6163 & n6431 ) | ( n6430 & n6431 ) ;
  assign n6434 = ( n6163 & n6432 ) | ( n6163 & ~n6433 ) | ( n6432 & ~n6433 ) ;
  assign n6435 = ( ~n132 & n6429 ) | ( ~n132 & n6434 ) | ( n6429 & n6434 ) ;
  assign n6436 = ( n132 & ~n6164 ) | ( n132 & n6172 ) | ( ~n6164 & n6172 ) ;
  assign n6437 = n132 & ~n6164 ;
  assign n6438 = ( n6169 & n6436 ) | ( n6169 & n6437 ) | ( n6436 & n6437 ) ;
  assign n6439 = ( ~n6169 & n6436 ) | ( ~n6169 & n6437 ) | ( n6436 & n6437 ) ;
  assign n6440 = ( n6169 & ~n6438 ) | ( n6169 & n6439 ) | ( ~n6438 & n6439 ) ;
  assign n6441 = ( ~n131 & n6435 ) | ( ~n131 & n6440 ) | ( n6435 & n6440 ) ;
  assign n6442 = n6175 | n6441 ;
  assign n6443 = n6435 & ~n6440 ;
  assign n6444 = n6175 | n6440 ;
  assign n6445 = ~n6435 & n6440 ;
  assign n6446 = ( n6443 & n6444 ) | ( n6443 & n6445 ) | ( n6444 & n6445 ) ;
  assign n6447 = n131 & n6446 ;
  assign n6448 = n132 & ~n6429 ;
  assign n6449 = ( n132 & ~n6429 ) | ( n132 & n6442 ) | ( ~n6429 & n6442 ) ;
  assign n6450 = ( n6434 & n6448 ) | ( n6434 & n6449 ) | ( n6448 & n6449 ) ;
  assign n6451 = ( ~n6434 & n6448 ) | ( ~n6434 & n6449 ) | ( n6448 & n6449 ) ;
  assign n6452 = ( n6434 & ~n6450 ) | ( n6434 & n6451 ) | ( ~n6450 & n6451 ) ;
  assign n6453 = x34 | x35 ;
  assign n6454 = x36 | n6453 ;
  assign n6455 = ~n6172 & n6454 ;
  assign n6456 = ( x37 & ~n6442 ) | ( x37 & n6455 ) | ( ~n6442 & n6455 ) ;
  assign n6457 = n6172 & ~n6454 ;
  assign n6458 = ~n6176 & n6442 ;
  assign n6459 = ( n6456 & ~n6457 ) | ( n6456 & n6458 ) | ( ~n6457 & n6458 ) ;
  assign n6460 = n6172 & ~n6442 ;
  assign n6461 = ( x38 & n6458 ) | ( x38 & n6460 ) | ( n6458 & n6460 ) ;
  assign n6462 = ( ~x38 & n6458 ) | ( ~x38 & n6460 ) | ( n6458 & n6460 ) ;
  assign n6463 = ( x38 & ~n6461 ) | ( x38 & n6462 ) | ( ~n6461 & n6462 ) ;
  assign n6464 = ( ~n5905 & n6459 ) | ( ~n5905 & n6463 ) | ( n6459 & n6463 ) ;
  assign n6465 = ( n5905 & n6172 ) | ( n5905 & ~n6442 ) | ( n6172 & ~n6442 ) ;
  assign n6466 = n6184 & ~n6465 ;
  assign n6467 = ( ~x39 & n6462 ) | ( ~x39 & n6466 ) | ( n6462 & n6466 ) ;
  assign n6468 = ( x39 & n6462 ) | ( x39 & n6466 ) | ( n6462 & n6466 ) ;
  assign n6469 = ( x39 & n6467 ) | ( x39 & ~n6468 ) | ( n6467 & ~n6468 ) ;
  assign n6470 = ( ~n5642 & n6464 ) | ( ~n5642 & n6469 ) | ( n6464 & n6469 ) ;
  assign n6471 = ( n5642 & ~n6183 ) | ( n5642 & n6442 ) | ( ~n6183 & n6442 ) ;
  assign n6472 = n5642 & ~n6183 ;
  assign n6473 = ( n6187 & n6471 ) | ( n6187 & n6472 ) | ( n6471 & n6472 ) ;
  assign n6474 = ( ~n6187 & n6471 ) | ( ~n6187 & n6472 ) | ( n6471 & n6472 ) ;
  assign n6475 = ( n6187 & ~n6473 ) | ( n6187 & n6474 ) | ( ~n6473 & n6474 ) ;
  assign n6476 = ( ~n5386 & n6470 ) | ( ~n5386 & n6475 ) | ( n6470 & n6475 ) ;
  assign n6477 = n5386 & ~n6188 ;
  assign n6478 = ( n5386 & ~n6188 ) | ( n5386 & n6442 ) | ( ~n6188 & n6442 ) ;
  assign n6479 = ( ~n6194 & n6477 ) | ( ~n6194 & n6478 ) | ( n6477 & n6478 ) ;
  assign n6480 = ( n6194 & n6477 ) | ( n6194 & n6478 ) | ( n6477 & n6478 ) ;
  assign n6481 = ( n6194 & n6479 ) | ( n6194 & ~n6480 ) | ( n6479 & ~n6480 ) ;
  assign n6482 = ( ~n5139 & n6476 ) | ( ~n5139 & n6481 ) | ( n6476 & n6481 ) ;
  assign n6483 = ( n5139 & ~n6195 ) | ( n5139 & n6442 ) | ( ~n6195 & n6442 ) ;
  assign n6484 = n5139 & ~n6195 ;
  assign n6485 = ( n6200 & n6483 ) | ( n6200 & n6484 ) | ( n6483 & n6484 ) ;
  assign n6486 = ( ~n6200 & n6483 ) | ( ~n6200 & n6484 ) | ( n6483 & n6484 ) ;
  assign n6487 = ( n6200 & ~n6485 ) | ( n6200 & n6486 ) | ( ~n6485 & n6486 ) ;
  assign n6488 = ( ~n4898 & n6482 ) | ( ~n4898 & n6487 ) | ( n6482 & n6487 ) ;
  assign n6489 = ( n4898 & ~n6201 ) | ( n4898 & n6442 ) | ( ~n6201 & n6442 ) ;
  assign n6490 = n4898 & ~n6201 ;
  assign n6491 = ( n6206 & n6489 ) | ( n6206 & n6490 ) | ( n6489 & n6490 ) ;
  assign n6492 = ( ~n6206 & n6489 ) | ( ~n6206 & n6490 ) | ( n6489 & n6490 ) ;
  assign n6493 = ( n6206 & ~n6491 ) | ( n6206 & n6492 ) | ( ~n6491 & n6492 ) ;
  assign n6494 = ( ~n4661 & n6488 ) | ( ~n4661 & n6493 ) | ( n6488 & n6493 ) ;
  assign n6495 = ( n4661 & ~n6207 ) | ( n4661 & n6442 ) | ( ~n6207 & n6442 ) ;
  assign n6496 = n4661 & ~n6207 ;
  assign n6497 = ( n6212 & n6495 ) | ( n6212 & n6496 ) | ( n6495 & n6496 ) ;
  assign n6498 = ( ~n6212 & n6495 ) | ( ~n6212 & n6496 ) | ( n6495 & n6496 ) ;
  assign n6499 = ( n6212 & ~n6497 ) | ( n6212 & n6498 ) | ( ~n6497 & n6498 ) ;
  assign n6500 = ( ~n4432 & n6494 ) | ( ~n4432 & n6499 ) | ( n6494 & n6499 ) ;
  assign n6501 = ( n4432 & ~n6213 ) | ( n4432 & n6442 ) | ( ~n6213 & n6442 ) ;
  assign n6502 = n4432 & ~n6213 ;
  assign n6503 = ( n6218 & n6501 ) | ( n6218 & n6502 ) | ( n6501 & n6502 ) ;
  assign n6504 = ( ~n6218 & n6501 ) | ( ~n6218 & n6502 ) | ( n6501 & n6502 ) ;
  assign n6505 = ( n6218 & ~n6503 ) | ( n6218 & n6504 ) | ( ~n6503 & n6504 ) ;
  assign n6506 = ( ~n4203 & n6500 ) | ( ~n4203 & n6505 ) | ( n6500 & n6505 ) ;
  assign n6507 = ~n4203 & n6219 ;
  assign n6508 = ( ~n4203 & n6219 ) | ( ~n4203 & n6442 ) | ( n6219 & n6442 ) ;
  assign n6509 = ( n6224 & n6507 ) | ( n6224 & n6508 ) | ( n6507 & n6508 ) ;
  assign n6510 = ( ~n6224 & n6507 ) | ( ~n6224 & n6508 ) | ( n6507 & n6508 ) ;
  assign n6511 = ( n6224 & ~n6509 ) | ( n6224 & n6510 ) | ( ~n6509 & n6510 ) ;
  assign n6512 = ( ~n3985 & n6506 ) | ( ~n3985 & n6511 ) | ( n6506 & n6511 ) ;
  assign n6513 = ~n3985 & n6225 ;
  assign n6514 = ( ~n3985 & n6225 ) | ( ~n3985 & n6442 ) | ( n6225 & n6442 ) ;
  assign n6515 = ( ~n6230 & n6513 ) | ( ~n6230 & n6514 ) | ( n6513 & n6514 ) ;
  assign n6516 = ( n6230 & n6513 ) | ( n6230 & n6514 ) | ( n6513 & n6514 ) ;
  assign n6517 = ( n6230 & n6515 ) | ( n6230 & ~n6516 ) | ( n6515 & ~n6516 ) ;
  assign n6518 = ( ~n3772 & n6512 ) | ( ~n3772 & n6517 ) | ( n6512 & n6517 ) ;
  assign n6519 = ~n3772 & n6231 ;
  assign n6520 = ( ~n3772 & n6231 ) | ( ~n3772 & n6442 ) | ( n6231 & n6442 ) ;
  assign n6521 = ( n6236 & n6519 ) | ( n6236 & n6520 ) | ( n6519 & n6520 ) ;
  assign n6522 = ( ~n6236 & n6519 ) | ( ~n6236 & n6520 ) | ( n6519 & n6520 ) ;
  assign n6523 = ( n6236 & ~n6521 ) | ( n6236 & n6522 ) | ( ~n6521 & n6522 ) ;
  assign n6524 = ( ~n3567 & n6518 ) | ( ~n3567 & n6523 ) | ( n6518 & n6523 ) ;
  assign n6525 = ( n3567 & ~n6237 ) | ( n3567 & n6442 ) | ( ~n6237 & n6442 ) ;
  assign n6526 = n3567 & ~n6237 ;
  assign n6527 = ( n6242 & n6525 ) | ( n6242 & n6526 ) | ( n6525 & n6526 ) ;
  assign n6528 = ( ~n6242 & n6525 ) | ( ~n6242 & n6526 ) | ( n6525 & n6526 ) ;
  assign n6529 = ( n6242 & ~n6527 ) | ( n6242 & n6528 ) | ( ~n6527 & n6528 ) ;
  assign n6530 = ( ~n3362 & n6524 ) | ( ~n3362 & n6529 ) | ( n6524 & n6529 ) ;
  assign n6531 = ~n3362 & n6243 ;
  assign n6532 = ( ~n3362 & n6243 ) | ( ~n3362 & n6442 ) | ( n6243 & n6442 ) ;
  assign n6533 = ( ~n6248 & n6531 ) | ( ~n6248 & n6532 ) | ( n6531 & n6532 ) ;
  assign n6534 = ( n6248 & n6531 ) | ( n6248 & n6532 ) | ( n6531 & n6532 ) ;
  assign n6535 = ( n6248 & n6533 ) | ( n6248 & ~n6534 ) | ( n6533 & ~n6534 ) ;
  assign n6536 = ( ~n3169 & n6530 ) | ( ~n3169 & n6535 ) | ( n6530 & n6535 ) ;
  assign n6537 = ( n3169 & ~n6249 ) | ( n3169 & n6442 ) | ( ~n6249 & n6442 ) ;
  assign n6538 = n3169 & ~n6249 ;
  assign n6539 = ( n6254 & n6537 ) | ( n6254 & n6538 ) | ( n6537 & n6538 ) ;
  assign n6540 = ( ~n6254 & n6537 ) | ( ~n6254 & n6538 ) | ( n6537 & n6538 ) ;
  assign n6541 = ( n6254 & ~n6539 ) | ( n6254 & n6540 ) | ( ~n6539 & n6540 ) ;
  assign n6542 = ( ~n2979 & n6536 ) | ( ~n2979 & n6541 ) | ( n6536 & n6541 ) ;
  assign n6543 = ( n2979 & ~n6255 ) | ( n2979 & n6442 ) | ( ~n6255 & n6442 ) ;
  assign n6544 = n2979 & ~n6255 ;
  assign n6545 = ( n6260 & n6543 ) | ( n6260 & n6544 ) | ( n6543 & n6544 ) ;
  assign n6546 = ( ~n6260 & n6543 ) | ( ~n6260 & n6544 ) | ( n6543 & n6544 ) ;
  assign n6547 = ( n6260 & ~n6545 ) | ( n6260 & n6546 ) | ( ~n6545 & n6546 ) ;
  assign n6548 = ( ~n2791 & n6542 ) | ( ~n2791 & n6547 ) | ( n6542 & n6547 ) ;
  assign n6549 = n2791 & ~n6261 ;
  assign n6550 = ( n2791 & ~n6261 ) | ( n2791 & n6442 ) | ( ~n6261 & n6442 ) ;
  assign n6551 = ( n6266 & n6549 ) | ( n6266 & n6550 ) | ( n6549 & n6550 ) ;
  assign n6552 = ( ~n6266 & n6549 ) | ( ~n6266 & n6550 ) | ( n6549 & n6550 ) ;
  assign n6553 = ( n6266 & ~n6551 ) | ( n6266 & n6552 ) | ( ~n6551 & n6552 ) ;
  assign n6554 = ( ~n2615 & n6548 ) | ( ~n2615 & n6553 ) | ( n6548 & n6553 ) ;
  assign n6555 = ~n2615 & n6267 ;
  assign n6556 = ( ~n2615 & n6267 ) | ( ~n2615 & n6442 ) | ( n6267 & n6442 ) ;
  assign n6557 = ( ~n6272 & n6555 ) | ( ~n6272 & n6556 ) | ( n6555 & n6556 ) ;
  assign n6558 = ( n6272 & n6555 ) | ( n6272 & n6556 ) | ( n6555 & n6556 ) ;
  assign n6559 = ( n6272 & n6557 ) | ( n6272 & ~n6558 ) | ( n6557 & ~n6558 ) ;
  assign n6560 = ( ~n2443 & n6554 ) | ( ~n2443 & n6559 ) | ( n6554 & n6559 ) ;
  assign n6561 = ( n2443 & ~n6273 ) | ( n2443 & n6442 ) | ( ~n6273 & n6442 ) ;
  assign n6562 = n2443 & ~n6273 ;
  assign n6563 = ( n6278 & n6561 ) | ( n6278 & n6562 ) | ( n6561 & n6562 ) ;
  assign n6564 = ( ~n6278 & n6561 ) | ( ~n6278 & n6562 ) | ( n6561 & n6562 ) ;
  assign n6565 = ( n6278 & ~n6563 ) | ( n6278 & n6564 ) | ( ~n6563 & n6564 ) ;
  assign n6566 = ( ~n2277 & n6560 ) | ( ~n2277 & n6565 ) | ( n6560 & n6565 ) ;
  assign n6567 = ( n2277 & ~n6279 ) | ( n2277 & n6442 ) | ( ~n6279 & n6442 ) ;
  assign n6568 = n2277 & ~n6279 ;
  assign n6569 = ( n6284 & n6567 ) | ( n6284 & n6568 ) | ( n6567 & n6568 ) ;
  assign n6570 = ( ~n6284 & n6567 ) | ( ~n6284 & n6568 ) | ( n6567 & n6568 ) ;
  assign n6571 = ( n6284 & ~n6569 ) | ( n6284 & n6570 ) | ( ~n6569 & n6570 ) ;
  assign n6572 = ( ~n2111 & n6566 ) | ( ~n2111 & n6571 ) | ( n6566 & n6571 ) ;
  assign n6573 = ~n2111 & n6285 ;
  assign n6574 = ( ~n2111 & n6285 ) | ( ~n2111 & n6442 ) | ( n6285 & n6442 ) ;
  assign n6575 = ( n6290 & n6573 ) | ( n6290 & n6574 ) | ( n6573 & n6574 ) ;
  assign n6576 = ( ~n6290 & n6573 ) | ( ~n6290 & n6574 ) | ( n6573 & n6574 ) ;
  assign n6577 = ( n6290 & ~n6575 ) | ( n6290 & n6576 ) | ( ~n6575 & n6576 ) ;
  assign n6578 = ( ~n1949 & n6572 ) | ( ~n1949 & n6577 ) | ( n6572 & n6577 ) ;
  assign n6579 = ~n1949 & n6291 ;
  assign n6580 = ( ~n1949 & n6291 ) | ( ~n1949 & n6442 ) | ( n6291 & n6442 ) ;
  assign n6581 = ( ~n6296 & n6579 ) | ( ~n6296 & n6580 ) | ( n6579 & n6580 ) ;
  assign n6582 = ( n6296 & n6579 ) | ( n6296 & n6580 ) | ( n6579 & n6580 ) ;
  assign n6583 = ( n6296 & n6581 ) | ( n6296 & ~n6582 ) | ( n6581 & ~n6582 ) ;
  assign n6584 = ( ~n1802 & n6578 ) | ( ~n1802 & n6583 ) | ( n6578 & n6583 ) ;
  assign n6585 = ( n1802 & ~n6297 ) | ( n1802 & n6442 ) | ( ~n6297 & n6442 ) ;
  assign n6586 = n1802 & ~n6297 ;
  assign n6587 = ( n6302 & n6585 ) | ( n6302 & n6586 ) | ( n6585 & n6586 ) ;
  assign n6588 = ( ~n6302 & n6585 ) | ( ~n6302 & n6586 ) | ( n6585 & n6586 ) ;
  assign n6589 = ( n6302 & ~n6587 ) | ( n6302 & n6588 ) | ( ~n6587 & n6588 ) ;
  assign n6590 = ( ~n1661 & n6584 ) | ( ~n1661 & n6589 ) | ( n6584 & n6589 ) ;
  assign n6591 = n1661 & ~n6303 ;
  assign n6592 = ( n1661 & ~n6303 ) | ( n1661 & n6442 ) | ( ~n6303 & n6442 ) ;
  assign n6593 = ( n6308 & n6591 ) | ( n6308 & n6592 ) | ( n6591 & n6592 ) ;
  assign n6594 = ( ~n6308 & n6591 ) | ( ~n6308 & n6592 ) | ( n6591 & n6592 ) ;
  assign n6595 = ( n6308 & ~n6593 ) | ( n6308 & n6594 ) | ( ~n6593 & n6594 ) ;
  assign n6596 = ( ~n1523 & n6590 ) | ( ~n1523 & n6595 ) | ( n6590 & n6595 ) ;
  assign n6597 = ( n1523 & ~n6309 ) | ( n1523 & n6442 ) | ( ~n6309 & n6442 ) ;
  assign n6598 = n1523 & ~n6309 ;
  assign n6599 = ( n6314 & n6597 ) | ( n6314 & n6598 ) | ( n6597 & n6598 ) ;
  assign n6600 = ( ~n6314 & n6597 ) | ( ~n6314 & n6598 ) | ( n6597 & n6598 ) ;
  assign n6601 = ( n6314 & ~n6599 ) | ( n6314 & n6600 ) | ( ~n6599 & n6600 ) ;
  assign n6602 = ( ~n1393 & n6596 ) | ( ~n1393 & n6601 ) | ( n6596 & n6601 ) ;
  assign n6603 = ~n1393 & n6315 ;
  assign n6604 = ( ~n1393 & n6315 ) | ( ~n1393 & n6442 ) | ( n6315 & n6442 ) ;
  assign n6605 = ( ~n6320 & n6603 ) | ( ~n6320 & n6604 ) | ( n6603 & n6604 ) ;
  assign n6606 = ( n6320 & n6603 ) | ( n6320 & n6604 ) | ( n6603 & n6604 ) ;
  assign n6607 = ( n6320 & n6605 ) | ( n6320 & ~n6606 ) | ( n6605 & ~n6606 ) ;
  assign n6608 = ( ~n1266 & n6602 ) | ( ~n1266 & n6607 ) | ( n6602 & n6607 ) ;
  assign n6609 = ~n1266 & n6321 ;
  assign n6610 = ( ~n1266 & n6321 ) | ( ~n1266 & n6442 ) | ( n6321 & n6442 ) ;
  assign n6611 = ( ~n6326 & n6609 ) | ( ~n6326 & n6610 ) | ( n6609 & n6610 ) ;
  assign n6612 = ( n6326 & n6609 ) | ( n6326 & n6610 ) | ( n6609 & n6610 ) ;
  assign n6613 = ( n6326 & n6611 ) | ( n6326 & ~n6612 ) | ( n6611 & ~n6612 ) ;
  assign n6614 = ( ~n1150 & n6608 ) | ( ~n1150 & n6613 ) | ( n6608 & n6613 ) ;
  assign n6615 = ( n1150 & ~n6327 ) | ( n1150 & n6442 ) | ( ~n6327 & n6442 ) ;
  assign n6616 = n1150 & ~n6327 ;
  assign n6617 = ( n6332 & n6615 ) | ( n6332 & n6616 ) | ( n6615 & n6616 ) ;
  assign n6618 = ( ~n6332 & n6615 ) | ( ~n6332 & n6616 ) | ( n6615 & n6616 ) ;
  assign n6619 = ( n6332 & ~n6617 ) | ( n6332 & n6618 ) | ( ~n6617 & n6618 ) ;
  assign n6620 = ( ~n1038 & n6614 ) | ( ~n1038 & n6619 ) | ( n6614 & n6619 ) ;
  assign n6621 = n1038 & ~n6333 ;
  assign n6622 = ( n1038 & ~n6333 ) | ( n1038 & n6442 ) | ( ~n6333 & n6442 ) ;
  assign n6623 = ( n6338 & n6621 ) | ( n6338 & n6622 ) | ( n6621 & n6622 ) ;
  assign n6624 = ( ~n6338 & n6621 ) | ( ~n6338 & n6622 ) | ( n6621 & n6622 ) ;
  assign n6625 = ( n6338 & ~n6623 ) | ( n6338 & n6624 ) | ( ~n6623 & n6624 ) ;
  assign n6626 = ( ~n933 & n6620 ) | ( ~n933 & n6625 ) | ( n6620 & n6625 ) ;
  assign n6627 = ( n933 & ~n6339 ) | ( n933 & n6442 ) | ( ~n6339 & n6442 ) ;
  assign n6628 = n933 & ~n6339 ;
  assign n6629 = ( n6344 & n6627 ) | ( n6344 & n6628 ) | ( n6627 & n6628 ) ;
  assign n6630 = ( ~n6344 & n6627 ) | ( ~n6344 & n6628 ) | ( n6627 & n6628 ) ;
  assign n6631 = ( n6344 & ~n6629 ) | ( n6344 & n6630 ) | ( ~n6629 & n6630 ) ;
  assign n6632 = ( ~n839 & n6626 ) | ( ~n839 & n6631 ) | ( n6626 & n6631 ) ;
  assign n6633 = ( n839 & ~n6345 ) | ( n839 & n6442 ) | ( ~n6345 & n6442 ) ;
  assign n6634 = n839 & ~n6345 ;
  assign n6635 = ( n6350 & n6633 ) | ( n6350 & n6634 ) | ( n6633 & n6634 ) ;
  assign n6636 = ( ~n6350 & n6633 ) | ( ~n6350 & n6634 ) | ( n6633 & n6634 ) ;
  assign n6637 = ( n6350 & ~n6635 ) | ( n6350 & n6636 ) | ( ~n6635 & n6636 ) ;
  assign n6638 = ( ~n746 & n6632 ) | ( ~n746 & n6637 ) | ( n6632 & n6637 ) ;
  assign n6639 = ~n746 & n6351 ;
  assign n6640 = ( ~n746 & n6351 ) | ( ~n746 & n6442 ) | ( n6351 & n6442 ) ;
  assign n6641 = ( ~n6356 & n6639 ) | ( ~n6356 & n6640 ) | ( n6639 & n6640 ) ;
  assign n6642 = ( n6356 & n6639 ) | ( n6356 & n6640 ) | ( n6639 & n6640 ) ;
  assign n6643 = ( n6356 & n6641 ) | ( n6356 & ~n6642 ) | ( n6641 & ~n6642 ) ;
  assign n6644 = ( ~n664 & n6638 ) | ( ~n664 & n6643 ) | ( n6638 & n6643 ) ;
  assign n6645 = ( n664 & ~n6357 ) | ( n664 & n6442 ) | ( ~n6357 & n6442 ) ;
  assign n6646 = n664 & ~n6357 ;
  assign n6647 = ( n6362 & n6645 ) | ( n6362 & n6646 ) | ( n6645 & n6646 ) ;
  assign n6648 = ( ~n6362 & n6645 ) | ( ~n6362 & n6646 ) | ( n6645 & n6646 ) ;
  assign n6649 = ( n6362 & ~n6647 ) | ( n6362 & n6648 ) | ( ~n6647 & n6648 ) ;
  assign n6650 = ( ~n588 & n6644 ) | ( ~n588 & n6649 ) | ( n6644 & n6649 ) ;
  assign n6651 = ( n588 & ~n6363 ) | ( n588 & n6442 ) | ( ~n6363 & n6442 ) ;
  assign n6652 = n588 & ~n6363 ;
  assign n6653 = ( n6368 & n6651 ) | ( n6368 & n6652 ) | ( n6651 & n6652 ) ;
  assign n6654 = ( ~n6368 & n6651 ) | ( ~n6368 & n6652 ) | ( n6651 & n6652 ) ;
  assign n6655 = ( n6368 & ~n6653 ) | ( n6368 & n6654 ) | ( ~n6653 & n6654 ) ;
  assign n6656 = ( ~n518 & n6650 ) | ( ~n518 & n6655 ) | ( n6650 & n6655 ) ;
  assign n6657 = ( n518 & ~n6369 ) | ( n518 & n6442 ) | ( ~n6369 & n6442 ) ;
  assign n6658 = n518 & ~n6369 ;
  assign n6659 = ( n6374 & n6657 ) | ( n6374 & n6658 ) | ( n6657 & n6658 ) ;
  assign n6660 = ( ~n6374 & n6657 ) | ( ~n6374 & n6658 ) | ( n6657 & n6658 ) ;
  assign n6661 = ( n6374 & ~n6659 ) | ( n6374 & n6660 ) | ( ~n6659 & n6660 ) ;
  assign n6662 = ( ~n454 & n6656 ) | ( ~n454 & n6661 ) | ( n6656 & n6661 ) ;
  assign n6663 = ( n454 & ~n6375 ) | ( n454 & n6442 ) | ( ~n6375 & n6442 ) ;
  assign n6664 = n454 & ~n6375 ;
  assign n6665 = ( n6380 & n6663 ) | ( n6380 & n6664 ) | ( n6663 & n6664 ) ;
  assign n6666 = ( ~n6380 & n6663 ) | ( ~n6380 & n6664 ) | ( n6663 & n6664 ) ;
  assign n6667 = ( n6380 & ~n6665 ) | ( n6380 & n6666 ) | ( ~n6665 & n6666 ) ;
  assign n6668 = ( ~n396 & n6662 ) | ( ~n396 & n6667 ) | ( n6662 & n6667 ) ;
  assign n6669 = ( n396 & ~n6381 ) | ( n396 & n6442 ) | ( ~n6381 & n6442 ) ;
  assign n6670 = n396 & ~n6381 ;
  assign n6671 = ( n6386 & n6669 ) | ( n6386 & n6670 ) | ( n6669 & n6670 ) ;
  assign n6672 = ( ~n6386 & n6669 ) | ( ~n6386 & n6670 ) | ( n6669 & n6670 ) ;
  assign n6673 = ( n6386 & ~n6671 ) | ( n6386 & n6672 ) | ( ~n6671 & n6672 ) ;
  assign n6674 = ( ~n344 & n6668 ) | ( ~n344 & n6673 ) | ( n6668 & n6673 ) ;
  assign n6675 = ~n344 & n6387 ;
  assign n6676 = ( ~n344 & n6387 ) | ( ~n344 & n6442 ) | ( n6387 & n6442 ) ;
  assign n6677 = ( n6392 & n6675 ) | ( n6392 & n6676 ) | ( n6675 & n6676 ) ;
  assign n6678 = ( ~n6392 & n6675 ) | ( ~n6392 & n6676 ) | ( n6675 & n6676 ) ;
  assign n6679 = ( n6392 & ~n6677 ) | ( n6392 & n6678 ) | ( ~n6677 & n6678 ) ;
  assign n6680 = ( ~n298 & n6674 ) | ( ~n298 & n6679 ) | ( n6674 & n6679 ) ;
  assign n6681 = ( n298 & ~n6393 ) | ( n298 & n6442 ) | ( ~n6393 & n6442 ) ;
  assign n6682 = n298 & ~n6393 ;
  assign n6683 = ( n6398 & n6681 ) | ( n6398 & n6682 ) | ( n6681 & n6682 ) ;
  assign n6684 = ( ~n6398 & n6681 ) | ( ~n6398 & n6682 ) | ( n6681 & n6682 ) ;
  assign n6685 = ( n6398 & ~n6683 ) | ( n6398 & n6684 ) | ( ~n6683 & n6684 ) ;
  assign n6686 = ( ~n258 & n6680 ) | ( ~n258 & n6685 ) | ( n6680 & n6685 ) ;
  assign n6687 = ~n258 & n6399 ;
  assign n6688 = ( ~n258 & n6399 ) | ( ~n258 & n6442 ) | ( n6399 & n6442 ) ;
  assign n6689 = ( n6404 & n6687 ) | ( n6404 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6690 = ( ~n6404 & n6687 ) | ( ~n6404 & n6688 ) | ( n6687 & n6688 ) ;
  assign n6691 = ( n6404 & ~n6689 ) | ( n6404 & n6690 ) | ( ~n6689 & n6690 ) ;
  assign n6692 = ( ~n225 & n6686 ) | ( ~n225 & n6691 ) | ( n6686 & n6691 ) ;
  assign n6693 = ~n225 & n6405 ;
  assign n6694 = ( ~n225 & n6405 ) | ( ~n225 & n6442 ) | ( n6405 & n6442 ) ;
  assign n6695 = ( ~n6410 & n6693 ) | ( ~n6410 & n6694 ) | ( n6693 & n6694 ) ;
  assign n6696 = ( n6410 & n6693 ) | ( n6410 & n6694 ) | ( n6693 & n6694 ) ;
  assign n6697 = ( n6410 & n6695 ) | ( n6410 & ~n6696 ) | ( n6695 & ~n6696 ) ;
  assign n6698 = ( ~n197 & n6692 ) | ( ~n197 & n6697 ) | ( n6692 & n6697 ) ;
  assign n6699 = ~n197 & n6411 ;
  assign n6700 = ( ~n197 & n6411 ) | ( ~n197 & n6442 ) | ( n6411 & n6442 ) ;
  assign n6701 = ( ~n6416 & n6699 ) | ( ~n6416 & n6700 ) | ( n6699 & n6700 ) ;
  assign n6702 = ( n6416 & n6699 ) | ( n6416 & n6700 ) | ( n6699 & n6700 ) ;
  assign n6703 = ( n6416 & n6701 ) | ( n6416 & ~n6702 ) | ( n6701 & ~n6702 ) ;
  assign n6704 = ( ~n170 & n6698 ) | ( ~n170 & n6703 ) | ( n6698 & n6703 ) ;
  assign n6705 = ( n170 & ~n6417 ) | ( n170 & n6442 ) | ( ~n6417 & n6442 ) ;
  assign n6706 = n170 & ~n6417 ;
  assign n6707 = ( n6422 & n6705 ) | ( n6422 & n6706 ) | ( n6705 & n6706 ) ;
  assign n6708 = ( ~n6422 & n6705 ) | ( ~n6422 & n6706 ) | ( n6705 & n6706 ) ;
  assign n6709 = ( n6422 & ~n6707 ) | ( n6422 & n6708 ) | ( ~n6707 & n6708 ) ;
  assign n6710 = ( ~n142 & n6704 ) | ( ~n142 & n6709 ) | ( n6704 & n6709 ) ;
  assign n6711 = ~n142 & n6423 ;
  assign n6712 = ( ~n142 & n6423 ) | ( ~n142 & n6442 ) | ( n6423 & n6442 ) ;
  assign n6713 = ( ~n6428 & n6711 ) | ( ~n6428 & n6712 ) | ( n6711 & n6712 ) ;
  assign n6714 = ( n6428 & n6711 ) | ( n6428 & n6712 ) | ( n6711 & n6712 ) ;
  assign n6715 = ( n6428 & n6713 ) | ( n6428 & ~n6714 ) | ( n6713 & ~n6714 ) ;
  assign n6716 = ( ~n132 & n6710 ) | ( ~n132 & n6715 ) | ( n6710 & n6715 ) ;
  assign n6717 = n6452 & n6716 ;
  assign n6718 = ( ~n131 & n6452 ) | ( ~n131 & n6717 ) | ( n6452 & n6717 ) ;
  assign n6719 = n6447 | n6718 ;
  assign n6720 = ( ~n131 & n6444 ) | ( ~n131 & n6446 ) | ( n6444 & n6446 ) ;
  assign n6721 = ~n6446 & n6720 ;
  assign n6722 = ( ~n131 & n6716 ) | ( ~n131 & n6721 ) | ( n6716 & n6721 ) ;
  assign n6723 = n6719 | n6722 ;
  assign n6724 = x32 | x33 ;
  assign n6725 = x34 | n6724 ;
  assign n6726 = ~n6442 & n6725 ;
  assign n6727 = ( x35 & ~n6723 ) | ( x35 & n6726 ) | ( ~n6723 & n6726 ) ;
  assign n6728 = n6442 & ~n6725 ;
  assign n6729 = ~n6453 & n6723 ;
  assign n6730 = ( n6727 & ~n6728 ) | ( n6727 & n6729 ) | ( ~n6728 & n6729 ) ;
  assign n6731 = n6442 & ~n6723 ;
  assign n6732 = ( x36 & n6729 ) | ( x36 & n6731 ) | ( n6729 & n6731 ) ;
  assign n6733 = ( ~x36 & n6729 ) | ( ~x36 & n6731 ) | ( n6729 & n6731 ) ;
  assign n6734 = ( x36 & ~n6732 ) | ( x36 & n6733 ) | ( ~n6732 & n6733 ) ;
  assign n6735 = ( ~n6172 & n6730 ) | ( ~n6172 & n6734 ) | ( n6730 & n6734 ) ;
  assign n6736 = ~n6172 & n6442 ;
  assign n6737 = ( n6460 & n6723 ) | ( n6460 & n6736 ) | ( n6723 & n6736 ) ;
  assign n6738 = ( x37 & n6733 ) | ( x37 & n6737 ) | ( n6733 & n6737 ) ;
  assign n6739 = ( ~x37 & n6733 ) | ( ~x37 & n6737 ) | ( n6733 & n6737 ) ;
  assign n6740 = ( x37 & ~n6738 ) | ( x37 & n6739 ) | ( ~n6738 & n6739 ) ;
  assign n6741 = ( ~n5905 & n6735 ) | ( ~n5905 & n6740 ) | ( n6735 & n6740 ) ;
  assign n6742 = n5905 & ~n6459 ;
  assign n6743 = ( n5905 & ~n6459 ) | ( n5905 & n6723 ) | ( ~n6459 & n6723 ) ;
  assign n6744 = ( ~n6463 & n6742 ) | ( ~n6463 & n6743 ) | ( n6742 & n6743 ) ;
  assign n6745 = ( n6463 & n6742 ) | ( n6463 & n6743 ) | ( n6742 & n6743 ) ;
  assign n6746 = ( n6463 & n6744 ) | ( n6463 & ~n6745 ) | ( n6744 & ~n6745 ) ;
  assign n6747 = ( ~n5642 & n6741 ) | ( ~n5642 & n6746 ) | ( n6741 & n6746 ) ;
  assign n6748 = n5642 & ~n6464 ;
  assign n6749 = ( n5642 & ~n6464 ) | ( n5642 & n6723 ) | ( ~n6464 & n6723 ) ;
  assign n6750 = ( n6469 & n6748 ) | ( n6469 & n6749 ) | ( n6748 & n6749 ) ;
  assign n6751 = ( ~n6469 & n6748 ) | ( ~n6469 & n6749 ) | ( n6748 & n6749 ) ;
  assign n6752 = ( n6469 & ~n6750 ) | ( n6469 & n6751 ) | ( ~n6750 & n6751 ) ;
  assign n6753 = ( ~n5386 & n6747 ) | ( ~n5386 & n6752 ) | ( n6747 & n6752 ) ;
  assign n6754 = ( n5386 & ~n6470 ) | ( n5386 & n6723 ) | ( ~n6470 & n6723 ) ;
  assign n6755 = n5386 & ~n6470 ;
  assign n6756 = ( n6475 & n6754 ) | ( n6475 & n6755 ) | ( n6754 & n6755 ) ;
  assign n6757 = ( ~n6475 & n6754 ) | ( ~n6475 & n6755 ) | ( n6754 & n6755 ) ;
  assign n6758 = ( n6475 & ~n6756 ) | ( n6475 & n6757 ) | ( ~n6756 & n6757 ) ;
  assign n6759 = ( ~n5139 & n6753 ) | ( ~n5139 & n6758 ) | ( n6753 & n6758 ) ;
  assign n6760 = ( n5139 & ~n6476 ) | ( n5139 & n6723 ) | ( ~n6476 & n6723 ) ;
  assign n6761 = n5139 & ~n6476 ;
  assign n6762 = ( n6481 & n6760 ) | ( n6481 & n6761 ) | ( n6760 & n6761 ) ;
  assign n6763 = ( ~n6481 & n6760 ) | ( ~n6481 & n6761 ) | ( n6760 & n6761 ) ;
  assign n6764 = ( n6481 & ~n6762 ) | ( n6481 & n6763 ) | ( ~n6762 & n6763 ) ;
  assign n6765 = ( ~n4898 & n6759 ) | ( ~n4898 & n6764 ) | ( n6759 & n6764 ) ;
  assign n6766 = ~n4898 & n6482 ;
  assign n6767 = ( ~n4898 & n6482 ) | ( ~n4898 & n6723 ) | ( n6482 & n6723 ) ;
  assign n6768 = ( ~n6487 & n6766 ) | ( ~n6487 & n6767 ) | ( n6766 & n6767 ) ;
  assign n6769 = ( n6487 & n6766 ) | ( n6487 & n6767 ) | ( n6766 & n6767 ) ;
  assign n6770 = ( n6487 & n6768 ) | ( n6487 & ~n6769 ) | ( n6768 & ~n6769 ) ;
  assign n6771 = ( ~n4661 & n6765 ) | ( ~n4661 & n6770 ) | ( n6765 & n6770 ) ;
  assign n6772 = ~n4661 & n6488 ;
  assign n6773 = ( ~n4661 & n6488 ) | ( ~n4661 & n6723 ) | ( n6488 & n6723 ) ;
  assign n6774 = ( ~n6493 & n6772 ) | ( ~n6493 & n6773 ) | ( n6772 & n6773 ) ;
  assign n6775 = ( n6493 & n6772 ) | ( n6493 & n6773 ) | ( n6772 & n6773 ) ;
  assign n6776 = ( n6493 & n6774 ) | ( n6493 & ~n6775 ) | ( n6774 & ~n6775 ) ;
  assign n6777 = ( ~n4432 & n6771 ) | ( ~n4432 & n6776 ) | ( n6771 & n6776 ) ;
  assign n6778 = ( n4432 & ~n6494 ) | ( n4432 & n6723 ) | ( ~n6494 & n6723 ) ;
  assign n6779 = n4432 & ~n6494 ;
  assign n6780 = ( n6499 & n6778 ) | ( n6499 & n6779 ) | ( n6778 & n6779 ) ;
  assign n6781 = ( ~n6499 & n6778 ) | ( ~n6499 & n6779 ) | ( n6778 & n6779 ) ;
  assign n6782 = ( n6499 & ~n6780 ) | ( n6499 & n6781 ) | ( ~n6780 & n6781 ) ;
  assign n6783 = ( ~n4203 & n6777 ) | ( ~n4203 & n6782 ) | ( n6777 & n6782 ) ;
  assign n6784 = ( n4203 & ~n6500 ) | ( n4203 & n6723 ) | ( ~n6500 & n6723 ) ;
  assign n6785 = n4203 & ~n6500 ;
  assign n6786 = ( n6505 & n6784 ) | ( n6505 & n6785 ) | ( n6784 & n6785 ) ;
  assign n6787 = ( ~n6505 & n6784 ) | ( ~n6505 & n6785 ) | ( n6784 & n6785 ) ;
  assign n6788 = ( n6505 & ~n6786 ) | ( n6505 & n6787 ) | ( ~n6786 & n6787 ) ;
  assign n6789 = ( ~n3985 & n6783 ) | ( ~n3985 & n6788 ) | ( n6783 & n6788 ) ;
  assign n6790 = n3985 & ~n6506 ;
  assign n6791 = ( n3985 & ~n6506 ) | ( n3985 & n6723 ) | ( ~n6506 & n6723 ) ;
  assign n6792 = ( n6511 & n6790 ) | ( n6511 & n6791 ) | ( n6790 & n6791 ) ;
  assign n6793 = ( ~n6511 & n6790 ) | ( ~n6511 & n6791 ) | ( n6790 & n6791 ) ;
  assign n6794 = ( n6511 & ~n6792 ) | ( n6511 & n6793 ) | ( ~n6792 & n6793 ) ;
  assign n6795 = ( ~n3772 & n6789 ) | ( ~n3772 & n6794 ) | ( n6789 & n6794 ) ;
  assign n6796 = ( n3772 & ~n6512 ) | ( n3772 & n6723 ) | ( ~n6512 & n6723 ) ;
  assign n6797 = n3772 & ~n6512 ;
  assign n6798 = ( n6517 & n6796 ) | ( n6517 & n6797 ) | ( n6796 & n6797 ) ;
  assign n6799 = ( ~n6517 & n6796 ) | ( ~n6517 & n6797 ) | ( n6796 & n6797 ) ;
  assign n6800 = ( n6517 & ~n6798 ) | ( n6517 & n6799 ) | ( ~n6798 & n6799 ) ;
  assign n6801 = ( ~n3567 & n6795 ) | ( ~n3567 & n6800 ) | ( n6795 & n6800 ) ;
  assign n6802 = ( n3567 & ~n6518 ) | ( n3567 & n6723 ) | ( ~n6518 & n6723 ) ;
  assign n6803 = n3567 & ~n6518 ;
  assign n6804 = ( n6523 & n6802 ) | ( n6523 & n6803 ) | ( n6802 & n6803 ) ;
  assign n6805 = ( ~n6523 & n6802 ) | ( ~n6523 & n6803 ) | ( n6802 & n6803 ) ;
  assign n6806 = ( n6523 & ~n6804 ) | ( n6523 & n6805 ) | ( ~n6804 & n6805 ) ;
  assign n6807 = ( ~n3362 & n6801 ) | ( ~n3362 & n6806 ) | ( n6801 & n6806 ) ;
  assign n6808 = ~n3362 & n6524 ;
  assign n6809 = ( ~n3362 & n6524 ) | ( ~n3362 & n6723 ) | ( n6524 & n6723 ) ;
  assign n6810 = ( n6529 & n6808 ) | ( n6529 & n6809 ) | ( n6808 & n6809 ) ;
  assign n6811 = ( ~n6529 & n6808 ) | ( ~n6529 & n6809 ) | ( n6808 & n6809 ) ;
  assign n6812 = ( n6529 & ~n6810 ) | ( n6529 & n6811 ) | ( ~n6810 & n6811 ) ;
  assign n6813 = ( ~n3169 & n6807 ) | ( ~n3169 & n6812 ) | ( n6807 & n6812 ) ;
  assign n6814 = ~n3169 & n6530 ;
  assign n6815 = ( ~n3169 & n6530 ) | ( ~n3169 & n6723 ) | ( n6530 & n6723 ) ;
  assign n6816 = ( n6535 & n6814 ) | ( n6535 & n6815 ) | ( n6814 & n6815 ) ;
  assign n6817 = ( ~n6535 & n6814 ) | ( ~n6535 & n6815 ) | ( n6814 & n6815 ) ;
  assign n6818 = ( n6535 & ~n6816 ) | ( n6535 & n6817 ) | ( ~n6816 & n6817 ) ;
  assign n6819 = ( ~n2979 & n6813 ) | ( ~n2979 & n6818 ) | ( n6813 & n6818 ) ;
  assign n6820 = n2979 & ~n6536 ;
  assign n6821 = ( n2979 & ~n6536 ) | ( n2979 & n6723 ) | ( ~n6536 & n6723 ) ;
  assign n6822 = ( ~n6541 & n6820 ) | ( ~n6541 & n6821 ) | ( n6820 & n6821 ) ;
  assign n6823 = ( n6541 & n6820 ) | ( n6541 & n6821 ) | ( n6820 & n6821 ) ;
  assign n6824 = ( n6541 & n6822 ) | ( n6541 & ~n6823 ) | ( n6822 & ~n6823 ) ;
  assign n6825 = ( ~n2791 & n6819 ) | ( ~n2791 & n6824 ) | ( n6819 & n6824 ) ;
  assign n6826 = ~n2791 & n6542 ;
  assign n6827 = ( ~n2791 & n6542 ) | ( ~n2791 & n6723 ) | ( n6542 & n6723 ) ;
  assign n6828 = ( n6547 & n6826 ) | ( n6547 & n6827 ) | ( n6826 & n6827 ) ;
  assign n6829 = ( ~n6547 & n6826 ) | ( ~n6547 & n6827 ) | ( n6826 & n6827 ) ;
  assign n6830 = ( n6547 & ~n6828 ) | ( n6547 & n6829 ) | ( ~n6828 & n6829 ) ;
  assign n6831 = ( ~n2615 & n6825 ) | ( ~n2615 & n6830 ) | ( n6825 & n6830 ) ;
  assign n6832 = ( n2615 & ~n6548 ) | ( n2615 & n6723 ) | ( ~n6548 & n6723 ) ;
  assign n6833 = n2615 & ~n6548 ;
  assign n6834 = ( n6553 & n6832 ) | ( n6553 & n6833 ) | ( n6832 & n6833 ) ;
  assign n6835 = ( ~n6553 & n6832 ) | ( ~n6553 & n6833 ) | ( n6832 & n6833 ) ;
  assign n6836 = ( n6553 & ~n6834 ) | ( n6553 & n6835 ) | ( ~n6834 & n6835 ) ;
  assign n6837 = ( ~n2443 & n6831 ) | ( ~n2443 & n6836 ) | ( n6831 & n6836 ) ;
  assign n6838 = ~n2443 & n6554 ;
  assign n6839 = ( ~n2443 & n6554 ) | ( ~n2443 & n6723 ) | ( n6554 & n6723 ) ;
  assign n6840 = ( ~n6559 & n6838 ) | ( ~n6559 & n6839 ) | ( n6838 & n6839 ) ;
  assign n6841 = ( n6559 & n6838 ) | ( n6559 & n6839 ) | ( n6838 & n6839 ) ;
  assign n6842 = ( n6559 & n6840 ) | ( n6559 & ~n6841 ) | ( n6840 & ~n6841 ) ;
  assign n6843 = ( ~n2277 & n6837 ) | ( ~n2277 & n6842 ) | ( n6837 & n6842 ) ;
  assign n6844 = ~n2277 & n6560 ;
  assign n6845 = ( ~n2277 & n6560 ) | ( ~n2277 & n6723 ) | ( n6560 & n6723 ) ;
  assign n6846 = ( n6565 & n6844 ) | ( n6565 & n6845 ) | ( n6844 & n6845 ) ;
  assign n6847 = ( ~n6565 & n6844 ) | ( ~n6565 & n6845 ) | ( n6844 & n6845 ) ;
  assign n6848 = ( n6565 & ~n6846 ) | ( n6565 & n6847 ) | ( ~n6846 & n6847 ) ;
  assign n6849 = ( ~n2111 & n6843 ) | ( ~n2111 & n6848 ) | ( n6843 & n6848 ) ;
  assign n6850 = ~n2111 & n6566 ;
  assign n6851 = ( ~n2111 & n6566 ) | ( ~n2111 & n6723 ) | ( n6566 & n6723 ) ;
  assign n6852 = ( n6571 & n6850 ) | ( n6571 & n6851 ) | ( n6850 & n6851 ) ;
  assign n6853 = ( ~n6571 & n6850 ) | ( ~n6571 & n6851 ) | ( n6850 & n6851 ) ;
  assign n6854 = ( n6571 & ~n6852 ) | ( n6571 & n6853 ) | ( ~n6852 & n6853 ) ;
  assign n6855 = ( ~n1949 & n6849 ) | ( ~n1949 & n6854 ) | ( n6849 & n6854 ) ;
  assign n6856 = ( n1949 & ~n6572 ) | ( n1949 & n6723 ) | ( ~n6572 & n6723 ) ;
  assign n6857 = n1949 & ~n6572 ;
  assign n6858 = ( n6577 & n6856 ) | ( n6577 & n6857 ) | ( n6856 & n6857 ) ;
  assign n6859 = ( ~n6577 & n6856 ) | ( ~n6577 & n6857 ) | ( n6856 & n6857 ) ;
  assign n6860 = ( n6577 & ~n6858 ) | ( n6577 & n6859 ) | ( ~n6858 & n6859 ) ;
  assign n6861 = ( ~n1802 & n6855 ) | ( ~n1802 & n6860 ) | ( n6855 & n6860 ) ;
  assign n6862 = ( n1802 & ~n6578 ) | ( n1802 & n6723 ) | ( ~n6578 & n6723 ) ;
  assign n6863 = n1802 & ~n6578 ;
  assign n6864 = ( n6583 & n6862 ) | ( n6583 & n6863 ) | ( n6862 & n6863 ) ;
  assign n6865 = ( ~n6583 & n6862 ) | ( ~n6583 & n6863 ) | ( n6862 & n6863 ) ;
  assign n6866 = ( n6583 & ~n6864 ) | ( n6583 & n6865 ) | ( ~n6864 & n6865 ) ;
  assign n6867 = ( ~n1661 & n6861 ) | ( ~n1661 & n6866 ) | ( n6861 & n6866 ) ;
  assign n6868 = ~n1661 & n6584 ;
  assign n6869 = ( ~n1661 & n6584 ) | ( ~n1661 & n6723 ) | ( n6584 & n6723 ) ;
  assign n6870 = ( n6589 & n6868 ) | ( n6589 & n6869 ) | ( n6868 & n6869 ) ;
  assign n6871 = ( ~n6589 & n6868 ) | ( ~n6589 & n6869 ) | ( n6868 & n6869 ) ;
  assign n6872 = ( n6589 & ~n6870 ) | ( n6589 & n6871 ) | ( ~n6870 & n6871 ) ;
  assign n6873 = ( ~n1523 & n6867 ) | ( ~n1523 & n6872 ) | ( n6867 & n6872 ) ;
  assign n6874 = ~n1523 & n6590 ;
  assign n6875 = ( ~n1523 & n6590 ) | ( ~n1523 & n6723 ) | ( n6590 & n6723 ) ;
  assign n6876 = ( ~n6595 & n6874 ) | ( ~n6595 & n6875 ) | ( n6874 & n6875 ) ;
  assign n6877 = ( n6595 & n6874 ) | ( n6595 & n6875 ) | ( n6874 & n6875 ) ;
  assign n6878 = ( n6595 & n6876 ) | ( n6595 & ~n6877 ) | ( n6876 & ~n6877 ) ;
  assign n6879 = ( ~n1393 & n6873 ) | ( ~n1393 & n6878 ) | ( n6873 & n6878 ) ;
  assign n6880 = ~n1393 & n6596 ;
  assign n6881 = ( ~n1393 & n6596 ) | ( ~n1393 & n6723 ) | ( n6596 & n6723 ) ;
  assign n6882 = ( ~n6601 & n6880 ) | ( ~n6601 & n6881 ) | ( n6880 & n6881 ) ;
  assign n6883 = ( n6601 & n6880 ) | ( n6601 & n6881 ) | ( n6880 & n6881 ) ;
  assign n6884 = ( n6601 & n6882 ) | ( n6601 & ~n6883 ) | ( n6882 & ~n6883 ) ;
  assign n6885 = ( ~n1266 & n6879 ) | ( ~n1266 & n6884 ) | ( n6879 & n6884 ) ;
  assign n6886 = ( n1266 & ~n6602 ) | ( n1266 & n6723 ) | ( ~n6602 & n6723 ) ;
  assign n6887 = n1266 & ~n6602 ;
  assign n6888 = ( n6607 & n6886 ) | ( n6607 & n6887 ) | ( n6886 & n6887 ) ;
  assign n6889 = ( ~n6607 & n6886 ) | ( ~n6607 & n6887 ) | ( n6886 & n6887 ) ;
  assign n6890 = ( n6607 & ~n6888 ) | ( n6607 & n6889 ) | ( ~n6888 & n6889 ) ;
  assign n6891 = ( ~n1150 & n6885 ) | ( ~n1150 & n6890 ) | ( n6885 & n6890 ) ;
  assign n6892 = ( n1150 & ~n6608 ) | ( n1150 & n6723 ) | ( ~n6608 & n6723 ) ;
  assign n6893 = n1150 & ~n6608 ;
  assign n6894 = ( n6613 & n6892 ) | ( n6613 & n6893 ) | ( n6892 & n6893 ) ;
  assign n6895 = ( ~n6613 & n6892 ) | ( ~n6613 & n6893 ) | ( n6892 & n6893 ) ;
  assign n6896 = ( n6613 & ~n6894 ) | ( n6613 & n6895 ) | ( ~n6894 & n6895 ) ;
  assign n6897 = ( ~n1038 & n6891 ) | ( ~n1038 & n6896 ) | ( n6891 & n6896 ) ;
  assign n6898 = ( n1038 & ~n6614 ) | ( n1038 & n6723 ) | ( ~n6614 & n6723 ) ;
  assign n6899 = n1038 & ~n6614 ;
  assign n6900 = ( n6619 & n6898 ) | ( n6619 & n6899 ) | ( n6898 & n6899 ) ;
  assign n6901 = ( ~n6619 & n6898 ) | ( ~n6619 & n6899 ) | ( n6898 & n6899 ) ;
  assign n6902 = ( n6619 & ~n6900 ) | ( n6619 & n6901 ) | ( ~n6900 & n6901 ) ;
  assign n6903 = ( ~n933 & n6897 ) | ( ~n933 & n6902 ) | ( n6897 & n6902 ) ;
  assign n6904 = ~n933 & n6620 ;
  assign n6905 = ( ~n933 & n6620 ) | ( ~n933 & n6723 ) | ( n6620 & n6723 ) ;
  assign n6906 = ( n6625 & n6904 ) | ( n6625 & n6905 ) | ( n6904 & n6905 ) ;
  assign n6907 = ( ~n6625 & n6904 ) | ( ~n6625 & n6905 ) | ( n6904 & n6905 ) ;
  assign n6908 = ( n6625 & ~n6906 ) | ( n6625 & n6907 ) | ( ~n6906 & n6907 ) ;
  assign n6909 = ( ~n839 & n6903 ) | ( ~n839 & n6908 ) | ( n6903 & n6908 ) ;
  assign n6910 = ( n839 & ~n6626 ) | ( n839 & n6723 ) | ( ~n6626 & n6723 ) ;
  assign n6911 = n839 & ~n6626 ;
  assign n6912 = ( n6631 & n6910 ) | ( n6631 & n6911 ) | ( n6910 & n6911 ) ;
  assign n6913 = ( ~n6631 & n6910 ) | ( ~n6631 & n6911 ) | ( n6910 & n6911 ) ;
  assign n6914 = ( n6631 & ~n6912 ) | ( n6631 & n6913 ) | ( ~n6912 & n6913 ) ;
  assign n6915 = ( ~n746 & n6909 ) | ( ~n746 & n6914 ) | ( n6909 & n6914 ) ;
  assign n6916 = ~n746 & n6632 ;
  assign n6917 = ( ~n746 & n6632 ) | ( ~n746 & n6723 ) | ( n6632 & n6723 ) ;
  assign n6918 = ( n6637 & n6916 ) | ( n6637 & n6917 ) | ( n6916 & n6917 ) ;
  assign n6919 = ( ~n6637 & n6916 ) | ( ~n6637 & n6917 ) | ( n6916 & n6917 ) ;
  assign n6920 = ( n6637 & ~n6918 ) | ( n6637 & n6919 ) | ( ~n6918 & n6919 ) ;
  assign n6921 = ( ~n664 & n6915 ) | ( ~n664 & n6920 ) | ( n6915 & n6920 ) ;
  assign n6922 = ( n664 & ~n6638 ) | ( n664 & n6723 ) | ( ~n6638 & n6723 ) ;
  assign n6923 = n664 & ~n6638 ;
  assign n6924 = ( n6643 & n6922 ) | ( n6643 & n6923 ) | ( n6922 & n6923 ) ;
  assign n6925 = ( ~n6643 & n6922 ) | ( ~n6643 & n6923 ) | ( n6922 & n6923 ) ;
  assign n6926 = ( n6643 & ~n6924 ) | ( n6643 & n6925 ) | ( ~n6924 & n6925 ) ;
  assign n6927 = ( ~n588 & n6921 ) | ( ~n588 & n6926 ) | ( n6921 & n6926 ) ;
  assign n6928 = ~n588 & n6644 ;
  assign n6929 = ( ~n588 & n6644 ) | ( ~n588 & n6723 ) | ( n6644 & n6723 ) ;
  assign n6930 = ( n6649 & n6928 ) | ( n6649 & n6929 ) | ( n6928 & n6929 ) ;
  assign n6931 = ( ~n6649 & n6928 ) | ( ~n6649 & n6929 ) | ( n6928 & n6929 ) ;
  assign n6932 = ( n6649 & ~n6930 ) | ( n6649 & n6931 ) | ( ~n6930 & n6931 ) ;
  assign n6933 = ( ~n518 & n6927 ) | ( ~n518 & n6932 ) | ( n6927 & n6932 ) ;
  assign n6934 = ( n518 & ~n6650 ) | ( n518 & n6723 ) | ( ~n6650 & n6723 ) ;
  assign n6935 = n518 & ~n6650 ;
  assign n6936 = ( n6655 & n6934 ) | ( n6655 & n6935 ) | ( n6934 & n6935 ) ;
  assign n6937 = ( ~n6655 & n6934 ) | ( ~n6655 & n6935 ) | ( n6934 & n6935 ) ;
  assign n6938 = ( n6655 & ~n6936 ) | ( n6655 & n6937 ) | ( ~n6936 & n6937 ) ;
  assign n6939 = ( ~n454 & n6933 ) | ( ~n454 & n6938 ) | ( n6933 & n6938 ) ;
  assign n6940 = n454 & ~n6656 ;
  assign n6941 = ( n454 & ~n6656 ) | ( n454 & n6723 ) | ( ~n6656 & n6723 ) ;
  assign n6942 = ( ~n6661 & n6940 ) | ( ~n6661 & n6941 ) | ( n6940 & n6941 ) ;
  assign n6943 = ( n6661 & n6940 ) | ( n6661 & n6941 ) | ( n6940 & n6941 ) ;
  assign n6944 = ( n6661 & n6942 ) | ( n6661 & ~n6943 ) | ( n6942 & ~n6943 ) ;
  assign n6945 = ( ~n396 & n6939 ) | ( ~n396 & n6944 ) | ( n6939 & n6944 ) ;
  assign n6946 = ( n396 & ~n6662 ) | ( n396 & n6723 ) | ( ~n6662 & n6723 ) ;
  assign n6947 = n396 & ~n6662 ;
  assign n6948 = ( n6667 & n6946 ) | ( n6667 & n6947 ) | ( n6946 & n6947 ) ;
  assign n6949 = ( ~n6667 & n6946 ) | ( ~n6667 & n6947 ) | ( n6946 & n6947 ) ;
  assign n6950 = ( n6667 & ~n6948 ) | ( n6667 & n6949 ) | ( ~n6948 & n6949 ) ;
  assign n6951 = ( ~n344 & n6945 ) | ( ~n344 & n6950 ) | ( n6945 & n6950 ) ;
  assign n6952 = ~n344 & n6668 ;
  assign n6953 = ( ~n344 & n6668 ) | ( ~n344 & n6723 ) | ( n6668 & n6723 ) ;
  assign n6954 = ( n6673 & n6952 ) | ( n6673 & n6953 ) | ( n6952 & n6953 ) ;
  assign n6955 = ( ~n6673 & n6952 ) | ( ~n6673 & n6953 ) | ( n6952 & n6953 ) ;
  assign n6956 = ( n6673 & ~n6954 ) | ( n6673 & n6955 ) | ( ~n6954 & n6955 ) ;
  assign n6957 = ( ~n298 & n6951 ) | ( ~n298 & n6956 ) | ( n6951 & n6956 ) ;
  assign n6958 = ( n298 & ~n6674 ) | ( n298 & n6723 ) | ( ~n6674 & n6723 ) ;
  assign n6959 = n298 & ~n6674 ;
  assign n6960 = ( n6679 & n6958 ) | ( n6679 & n6959 ) | ( n6958 & n6959 ) ;
  assign n6961 = ( ~n6679 & n6958 ) | ( ~n6679 & n6959 ) | ( n6958 & n6959 ) ;
  assign n6962 = ( n6679 & ~n6960 ) | ( n6679 & n6961 ) | ( ~n6960 & n6961 ) ;
  assign n6963 = ( ~n258 & n6957 ) | ( ~n258 & n6962 ) | ( n6957 & n6962 ) ;
  assign n6964 = n258 & ~n6680 ;
  assign n6965 = ( n258 & ~n6680 ) | ( n258 & n6723 ) | ( ~n6680 & n6723 ) ;
  assign n6966 = ( ~n6685 & n6964 ) | ( ~n6685 & n6965 ) | ( n6964 & n6965 ) ;
  assign n6967 = ( n6685 & n6964 ) | ( n6685 & n6965 ) | ( n6964 & n6965 ) ;
  assign n6968 = ( n6685 & n6966 ) | ( n6685 & ~n6967 ) | ( n6966 & ~n6967 ) ;
  assign n6969 = ( ~n225 & n6963 ) | ( ~n225 & n6968 ) | ( n6963 & n6968 ) ;
  assign n6970 = ( n225 & ~n6686 ) | ( n225 & n6723 ) | ( ~n6686 & n6723 ) ;
  assign n6971 = n225 & ~n6686 ;
  assign n6972 = ( n6691 & n6970 ) | ( n6691 & n6971 ) | ( n6970 & n6971 ) ;
  assign n6973 = ( ~n6691 & n6970 ) | ( ~n6691 & n6971 ) | ( n6970 & n6971 ) ;
  assign n6974 = ( n6691 & ~n6972 ) | ( n6691 & n6973 ) | ( ~n6972 & n6973 ) ;
  assign n6975 = ( ~n197 & n6969 ) | ( ~n197 & n6974 ) | ( n6969 & n6974 ) ;
  assign n6976 = ( n197 & ~n6692 ) | ( n197 & n6723 ) | ( ~n6692 & n6723 ) ;
  assign n6977 = n197 & ~n6692 ;
  assign n6978 = ( n6697 & n6976 ) | ( n6697 & n6977 ) | ( n6976 & n6977 ) ;
  assign n6979 = ( ~n6697 & n6976 ) | ( ~n6697 & n6977 ) | ( n6976 & n6977 ) ;
  assign n6980 = ( n6697 & ~n6978 ) | ( n6697 & n6979 ) | ( ~n6978 & n6979 ) ;
  assign n6981 = ( ~n170 & n6975 ) | ( ~n170 & n6980 ) | ( n6975 & n6980 ) ;
  assign n6982 = ~n170 & n6698 ;
  assign n6983 = ( ~n170 & n6698 ) | ( ~n170 & n6723 ) | ( n6698 & n6723 ) ;
  assign n6984 = ( ~n6703 & n6982 ) | ( ~n6703 & n6983 ) | ( n6982 & n6983 ) ;
  assign n6985 = ( n6703 & n6982 ) | ( n6703 & n6983 ) | ( n6982 & n6983 ) ;
  assign n6986 = ( n6703 & n6984 ) | ( n6703 & ~n6985 ) | ( n6984 & ~n6985 ) ;
  assign n6987 = ( ~n142 & n6981 ) | ( ~n142 & n6986 ) | ( n6981 & n6986 ) ;
  assign n6988 = ~n142 & n6704 ;
  assign n6989 = ( ~n142 & n6704 ) | ( ~n142 & n6723 ) | ( n6704 & n6723 ) ;
  assign n6990 = ( ~n6709 & n6988 ) | ( ~n6709 & n6989 ) | ( n6988 & n6989 ) ;
  assign n6991 = ( n6709 & n6988 ) | ( n6709 & n6989 ) | ( n6988 & n6989 ) ;
  assign n6992 = ( n6709 & n6990 ) | ( n6709 & ~n6991 ) | ( n6990 & ~n6991 ) ;
  assign n6993 = ( ~n132 & n6987 ) | ( ~n132 & n6992 ) | ( n6987 & n6992 ) ;
  assign n6994 = ( n132 & ~n6710 ) | ( n132 & n6723 ) | ( ~n6710 & n6723 ) ;
  assign n6995 = n132 & ~n6710 ;
  assign n6996 = ( n6715 & n6994 ) | ( n6715 & n6995 ) | ( n6994 & n6995 ) ;
  assign n6997 = ( ~n6715 & n6994 ) | ( ~n6715 & n6995 ) | ( n6994 & n6995 ) ;
  assign n6998 = ( n6715 & ~n6996 ) | ( n6715 & n6997 ) | ( ~n6996 & n6997 ) ;
  assign n6999 = ( ~n131 & n6993 ) | ( ~n131 & n6998 ) | ( n6993 & n6998 ) ;
  assign n7000 = n6452 | n6716 ;
  assign n7001 = ( n6717 & n6722 ) | ( n6717 & ~n7000 ) | ( n6722 & ~n7000 ) ;
  assign n7002 = ( n131 & n6452 ) | ( n131 & n6716 ) | ( n6452 & n6716 ) ;
  assign n7003 = n6446 & ~n6452 ;
  assign n7004 = n6716 & ~n7003 ;
  assign n7005 = ( n7001 & n7002 ) | ( n7001 & ~n7004 ) | ( n7002 & ~n7004 ) ;
  assign n7006 = n6999 | n7005 ;
  assign n7007 = ~n131 & n6998 ;
  assign n7008 = n6998 | n7001 ;
  assign n7009 = ( ~n6993 & n7007 ) | ( ~n6993 & n7008 ) | ( n7007 & n7008 ) ;
  assign n7010 = ( ~n6998 & n7002 ) | ( ~n6998 & n7004 ) | ( n7002 & n7004 ) ;
  assign n7011 = ~n7004 & n7010 ;
  assign n7012 = ( n6993 & ~n7007 ) | ( n6993 & n7008 ) | ( ~n7007 & n7008 ) ;
  assign n7013 = ( n7009 & n7011 ) | ( n7009 & n7012 ) | ( n7011 & n7012 ) ;
  assign n7014 = ( n132 & ~n6987 ) | ( n132 & n7006 ) | ( ~n6987 & n7006 ) ;
  assign n7015 = n132 & ~n6987 ;
  assign n7016 = ( n6992 & ~n7014 ) | ( n6992 & n7015 ) | ( ~n7014 & n7015 ) ;
  assign n7017 = ( n6992 & n7014 ) | ( n6992 & n7015 ) | ( n7014 & n7015 ) ;
  assign n7018 = ( n7014 & n7016 ) | ( n7014 & ~n7017 ) | ( n7016 & ~n7017 ) ;
  assign n7019 = n6723 & ~n7006 ;
  assign n7020 = ~n6724 & n7006 ;
  assign n7021 = ( x34 & n7019 ) | ( x34 & n7020 ) | ( n7019 & n7020 ) ;
  assign n7022 = ( ~x34 & n7019 ) | ( ~x34 & n7020 ) | ( n7019 & n7020 ) ;
  assign n7023 = ( x34 & ~n7021 ) | ( x34 & n7022 ) | ( ~n7021 & n7022 ) ;
  assign n7024 = x30 | x31 ;
  assign n7025 = x32 | n7024 ;
  assign n7026 = ~n6723 & n7025 ;
  assign n7027 = ( x33 & ~n7006 ) | ( x33 & n7026 ) | ( ~n7006 & n7026 ) ;
  assign n7028 = n6723 & ~n7025 ;
  assign n7029 = ( n7020 & n7027 ) | ( n7020 & ~n7028 ) | ( n7027 & ~n7028 ) ;
  assign n7030 = ( ~n6442 & n7023 ) | ( ~n6442 & n7029 ) | ( n7023 & n7029 ) ;
  assign n7031 = ~n6442 & n6723 ;
  assign n7032 = ( n6731 & n7006 ) | ( n6731 & n7031 ) | ( n7006 & n7031 ) ;
  assign n7033 = ( x35 & n7022 ) | ( x35 & n7032 ) | ( n7022 & n7032 ) ;
  assign n7034 = ( ~x35 & n7022 ) | ( ~x35 & n7032 ) | ( n7022 & n7032 ) ;
  assign n7035 = ( x35 & ~n7033 ) | ( x35 & n7034 ) | ( ~n7033 & n7034 ) ;
  assign n7036 = ( ~n6172 & n7030 ) | ( ~n6172 & n7035 ) | ( n7030 & n7035 ) ;
  assign n7037 = ( n6172 & ~n6730 ) | ( n6172 & n7006 ) | ( ~n6730 & n7006 ) ;
  assign n7038 = n6172 & ~n6730 ;
  assign n7039 = ( n6734 & n7037 ) | ( n6734 & n7038 ) | ( n7037 & n7038 ) ;
  assign n7040 = ( ~n6734 & n7037 ) | ( ~n6734 & n7038 ) | ( n7037 & n7038 ) ;
  assign n7041 = ( n6734 & ~n7039 ) | ( n6734 & n7040 ) | ( ~n7039 & n7040 ) ;
  assign n7042 = ( ~n5905 & n7036 ) | ( ~n5905 & n7041 ) | ( n7036 & n7041 ) ;
  assign n7043 = ( n5905 & ~n6735 ) | ( n5905 & n7006 ) | ( ~n6735 & n7006 ) ;
  assign n7044 = n5905 & ~n6735 ;
  assign n7045 = ( n6740 & n7043 ) | ( n6740 & n7044 ) | ( n7043 & n7044 ) ;
  assign n7046 = ( ~n6740 & n7043 ) | ( ~n6740 & n7044 ) | ( n7043 & n7044 ) ;
  assign n7047 = ( n6740 & ~n7045 ) | ( n6740 & n7046 ) | ( ~n7045 & n7046 ) ;
  assign n7048 = ( ~n5642 & n7042 ) | ( ~n5642 & n7047 ) | ( n7042 & n7047 ) ;
  assign n7049 = n5642 & ~n6741 ;
  assign n7050 = ( n5642 & ~n6741 ) | ( n5642 & n7006 ) | ( ~n6741 & n7006 ) ;
  assign n7051 = ( n6746 & n7049 ) | ( n6746 & n7050 ) | ( n7049 & n7050 ) ;
  assign n7052 = ( ~n6746 & n7049 ) | ( ~n6746 & n7050 ) | ( n7049 & n7050 ) ;
  assign n7053 = ( n6746 & ~n7051 ) | ( n6746 & n7052 ) | ( ~n7051 & n7052 ) ;
  assign n7054 = ( ~n5386 & n7048 ) | ( ~n5386 & n7053 ) | ( n7048 & n7053 ) ;
  assign n7055 = ~n5386 & n6747 ;
  assign n7056 = ( ~n5386 & n6747 ) | ( ~n5386 & n7006 ) | ( n6747 & n7006 ) ;
  assign n7057 = ( ~n6752 & n7055 ) | ( ~n6752 & n7056 ) | ( n7055 & n7056 ) ;
  assign n7058 = ( n6752 & n7055 ) | ( n6752 & n7056 ) | ( n7055 & n7056 ) ;
  assign n7059 = ( n6752 & n7057 ) | ( n6752 & ~n7058 ) | ( n7057 & ~n7058 ) ;
  assign n7060 = ( ~n5139 & n7054 ) | ( ~n5139 & n7059 ) | ( n7054 & n7059 ) ;
  assign n7061 = n5139 & ~n6753 ;
  assign n7062 = ( n5139 & ~n6753 ) | ( n5139 & n7006 ) | ( ~n6753 & n7006 ) ;
  assign n7063 = ( n6758 & n7061 ) | ( n6758 & n7062 ) | ( n7061 & n7062 ) ;
  assign n7064 = ( ~n6758 & n7061 ) | ( ~n6758 & n7062 ) | ( n7061 & n7062 ) ;
  assign n7065 = ( n6758 & ~n7063 ) | ( n6758 & n7064 ) | ( ~n7063 & n7064 ) ;
  assign n7066 = ( ~n4898 & n7060 ) | ( ~n4898 & n7065 ) | ( n7060 & n7065 ) ;
  assign n7067 = ~n4898 & n6759 ;
  assign n7068 = ( ~n4898 & n6759 ) | ( ~n4898 & n7006 ) | ( n6759 & n7006 ) ;
  assign n7069 = ( ~n6764 & n7067 ) | ( ~n6764 & n7068 ) | ( n7067 & n7068 ) ;
  assign n7070 = ( n6764 & n7067 ) | ( n6764 & n7068 ) | ( n7067 & n7068 ) ;
  assign n7071 = ( n6764 & n7069 ) | ( n6764 & ~n7070 ) | ( n7069 & ~n7070 ) ;
  assign n7072 = ( ~n4661 & n7066 ) | ( ~n4661 & n7071 ) | ( n7066 & n7071 ) ;
  assign n7073 = ( n4661 & ~n6765 ) | ( n4661 & n7006 ) | ( ~n6765 & n7006 ) ;
  assign n7074 = n4661 & ~n6765 ;
  assign n7075 = ( n6770 & n7073 ) | ( n6770 & n7074 ) | ( n7073 & n7074 ) ;
  assign n7076 = ( ~n6770 & n7073 ) | ( ~n6770 & n7074 ) | ( n7073 & n7074 ) ;
  assign n7077 = ( n6770 & ~n7075 ) | ( n6770 & n7076 ) | ( ~n7075 & n7076 ) ;
  assign n7078 = ( ~n4432 & n7072 ) | ( ~n4432 & n7077 ) | ( n7072 & n7077 ) ;
  assign n7079 = ( n4432 & ~n6771 ) | ( n4432 & n7006 ) | ( ~n6771 & n7006 ) ;
  assign n7080 = n4432 & ~n6771 ;
  assign n7081 = ( n6776 & n7079 ) | ( n6776 & n7080 ) | ( n7079 & n7080 ) ;
  assign n7082 = ( ~n6776 & n7079 ) | ( ~n6776 & n7080 ) | ( n7079 & n7080 ) ;
  assign n7083 = ( n6776 & ~n7081 ) | ( n6776 & n7082 ) | ( ~n7081 & n7082 ) ;
  assign n7084 = ( ~n4203 & n7078 ) | ( ~n4203 & n7083 ) | ( n7078 & n7083 ) ;
  assign n7085 = ( n4203 & ~n6777 ) | ( n4203 & n7006 ) | ( ~n6777 & n7006 ) ;
  assign n7086 = n4203 & ~n6777 ;
  assign n7087 = ( n6782 & n7085 ) | ( n6782 & n7086 ) | ( n7085 & n7086 ) ;
  assign n7088 = ( ~n6782 & n7085 ) | ( ~n6782 & n7086 ) | ( n7085 & n7086 ) ;
  assign n7089 = ( n6782 & ~n7087 ) | ( n6782 & n7088 ) | ( ~n7087 & n7088 ) ;
  assign n7090 = ( ~n3985 & n7084 ) | ( ~n3985 & n7089 ) | ( n7084 & n7089 ) ;
  assign n7091 = ~n3985 & n6783 ;
  assign n7092 = ( ~n3985 & n6783 ) | ( ~n3985 & n7006 ) | ( n6783 & n7006 ) ;
  assign n7093 = ( n6788 & n7091 ) | ( n6788 & n7092 ) | ( n7091 & n7092 ) ;
  assign n7094 = ( ~n6788 & n7091 ) | ( ~n6788 & n7092 ) | ( n7091 & n7092 ) ;
  assign n7095 = ( n6788 & ~n7093 ) | ( n6788 & n7094 ) | ( ~n7093 & n7094 ) ;
  assign n7096 = ( ~n3772 & n7090 ) | ( ~n3772 & n7095 ) | ( n7090 & n7095 ) ;
  assign n7097 = ( n3772 & ~n6789 ) | ( n3772 & n7006 ) | ( ~n6789 & n7006 ) ;
  assign n7098 = n3772 & ~n6789 ;
  assign n7099 = ( n6794 & n7097 ) | ( n6794 & n7098 ) | ( n7097 & n7098 ) ;
  assign n7100 = ( ~n6794 & n7097 ) | ( ~n6794 & n7098 ) | ( n7097 & n7098 ) ;
  assign n7101 = ( n6794 & ~n7099 ) | ( n6794 & n7100 ) | ( ~n7099 & n7100 ) ;
  assign n7102 = ( ~n3567 & n7096 ) | ( ~n3567 & n7101 ) | ( n7096 & n7101 ) ;
  assign n7103 = ~n3567 & n6795 ;
  assign n7104 = ( ~n3567 & n6795 ) | ( ~n3567 & n7006 ) | ( n6795 & n7006 ) ;
  assign n7105 = ( ~n6800 & n7103 ) | ( ~n6800 & n7104 ) | ( n7103 & n7104 ) ;
  assign n7106 = ( n6800 & n7103 ) | ( n6800 & n7104 ) | ( n7103 & n7104 ) ;
  assign n7107 = ( n6800 & n7105 ) | ( n6800 & ~n7106 ) | ( n7105 & ~n7106 ) ;
  assign n7108 = ( ~n3362 & n7102 ) | ( ~n3362 & n7107 ) | ( n7102 & n7107 ) ;
  assign n7109 = ~n3362 & n6801 ;
  assign n7110 = ( ~n3362 & n6801 ) | ( ~n3362 & n7006 ) | ( n6801 & n7006 ) ;
  assign n7111 = ( n6806 & n7109 ) | ( n6806 & n7110 ) | ( n7109 & n7110 ) ;
  assign n7112 = ( ~n6806 & n7109 ) | ( ~n6806 & n7110 ) | ( n7109 & n7110 ) ;
  assign n7113 = ( n6806 & ~n7111 ) | ( n6806 & n7112 ) | ( ~n7111 & n7112 ) ;
  assign n7114 = ( ~n3169 & n7108 ) | ( ~n3169 & n7113 ) | ( n7108 & n7113 ) ;
  assign n7115 = ~n3169 & n6807 ;
  assign n7116 = ( ~n3169 & n6807 ) | ( ~n3169 & n7006 ) | ( n6807 & n7006 ) ;
  assign n7117 = ( ~n6812 & n7115 ) | ( ~n6812 & n7116 ) | ( n7115 & n7116 ) ;
  assign n7118 = ( n6812 & n7115 ) | ( n6812 & n7116 ) | ( n7115 & n7116 ) ;
  assign n7119 = ( n6812 & n7117 ) | ( n6812 & ~n7118 ) | ( n7117 & ~n7118 ) ;
  assign n7120 = ( ~n2979 & n7114 ) | ( ~n2979 & n7119 ) | ( n7114 & n7119 ) ;
  assign n7121 = ( n2979 & ~n6813 ) | ( n2979 & n7006 ) | ( ~n6813 & n7006 ) ;
  assign n7122 = n2979 & ~n6813 ;
  assign n7123 = ( n6818 & n7121 ) | ( n6818 & n7122 ) | ( n7121 & n7122 ) ;
  assign n7124 = ( ~n6818 & n7121 ) | ( ~n6818 & n7122 ) | ( n7121 & n7122 ) ;
  assign n7125 = ( n6818 & ~n7123 ) | ( n6818 & n7124 ) | ( ~n7123 & n7124 ) ;
  assign n7126 = ( ~n2791 & n7120 ) | ( ~n2791 & n7125 ) | ( n7120 & n7125 ) ;
  assign n7127 = ( n2791 & ~n6819 ) | ( n2791 & n7006 ) | ( ~n6819 & n7006 ) ;
  assign n7128 = n2791 & ~n6819 ;
  assign n7129 = ( n6824 & n7127 ) | ( n6824 & n7128 ) | ( n7127 & n7128 ) ;
  assign n7130 = ( ~n6824 & n7127 ) | ( ~n6824 & n7128 ) | ( n7127 & n7128 ) ;
  assign n7131 = ( n6824 & ~n7129 ) | ( n6824 & n7130 ) | ( ~n7129 & n7130 ) ;
  assign n7132 = ( ~n2615 & n7126 ) | ( ~n2615 & n7131 ) | ( n7126 & n7131 ) ;
  assign n7133 = ~n2615 & n6825 ;
  assign n7134 = ( ~n2615 & n6825 ) | ( ~n2615 & n7006 ) | ( n6825 & n7006 ) ;
  assign n7135 = ( n6830 & n7133 ) | ( n6830 & n7134 ) | ( n7133 & n7134 ) ;
  assign n7136 = ( ~n6830 & n7133 ) | ( ~n6830 & n7134 ) | ( n7133 & n7134 ) ;
  assign n7137 = ( n6830 & ~n7135 ) | ( n6830 & n7136 ) | ( ~n7135 & n7136 ) ;
  assign n7138 = ( ~n2443 & n7132 ) | ( ~n2443 & n7137 ) | ( n7132 & n7137 ) ;
  assign n7139 = ~n2443 & n6831 ;
  assign n7140 = ( ~n2443 & n6831 ) | ( ~n2443 & n7006 ) | ( n6831 & n7006 ) ;
  assign n7141 = ( n6836 & n7139 ) | ( n6836 & n7140 ) | ( n7139 & n7140 ) ;
  assign n7142 = ( ~n6836 & n7139 ) | ( ~n6836 & n7140 ) | ( n7139 & n7140 ) ;
  assign n7143 = ( n6836 & ~n7141 ) | ( n6836 & n7142 ) | ( ~n7141 & n7142 ) ;
  assign n7144 = ( ~n2277 & n7138 ) | ( ~n2277 & n7143 ) | ( n7138 & n7143 ) ;
  assign n7145 = ~n2277 & n6837 ;
  assign n7146 = ( ~n2277 & n6837 ) | ( ~n2277 & n7006 ) | ( n6837 & n7006 ) ;
  assign n7147 = ( ~n6842 & n7145 ) | ( ~n6842 & n7146 ) | ( n7145 & n7146 ) ;
  assign n7148 = ( n6842 & n7145 ) | ( n6842 & n7146 ) | ( n7145 & n7146 ) ;
  assign n7149 = ( n6842 & n7147 ) | ( n6842 & ~n7148 ) | ( n7147 & ~n7148 ) ;
  assign n7150 = ( ~n2111 & n7144 ) | ( ~n2111 & n7149 ) | ( n7144 & n7149 ) ;
  assign n7151 = n2111 & ~n6843 ;
  assign n7152 = ( n2111 & ~n6843 ) | ( n2111 & n7006 ) | ( ~n6843 & n7006 ) ;
  assign n7153 = ( n6848 & n7151 ) | ( n6848 & n7152 ) | ( n7151 & n7152 ) ;
  assign n7154 = ( ~n6848 & n7151 ) | ( ~n6848 & n7152 ) | ( n7151 & n7152 ) ;
  assign n7155 = ( n6848 & ~n7153 ) | ( n6848 & n7154 ) | ( ~n7153 & n7154 ) ;
  assign n7156 = ( ~n1949 & n7150 ) | ( ~n1949 & n7155 ) | ( n7150 & n7155 ) ;
  assign n7157 = ( n1949 & ~n6849 ) | ( n1949 & n7006 ) | ( ~n6849 & n7006 ) ;
  assign n7158 = n1949 & ~n6849 ;
  assign n7159 = ( n6854 & n7157 ) | ( n6854 & n7158 ) | ( n7157 & n7158 ) ;
  assign n7160 = ( ~n6854 & n7157 ) | ( ~n6854 & n7158 ) | ( n7157 & n7158 ) ;
  assign n7161 = ( n6854 & ~n7159 ) | ( n6854 & n7160 ) | ( ~n7159 & n7160 ) ;
  assign n7162 = ( ~n1802 & n7156 ) | ( ~n1802 & n7161 ) | ( n7156 & n7161 ) ;
  assign n7163 = ~n1802 & n6855 ;
  assign n7164 = ( ~n1802 & n6855 ) | ( ~n1802 & n7006 ) | ( n6855 & n7006 ) ;
  assign n7165 = ( ~n6860 & n7163 ) | ( ~n6860 & n7164 ) | ( n7163 & n7164 ) ;
  assign n7166 = ( n6860 & n7163 ) | ( n6860 & n7164 ) | ( n7163 & n7164 ) ;
  assign n7167 = ( n6860 & n7165 ) | ( n6860 & ~n7166 ) | ( n7165 & ~n7166 ) ;
  assign n7168 = ( ~n1661 & n7162 ) | ( ~n1661 & n7167 ) | ( n7162 & n7167 ) ;
  assign n7169 = ~n1661 & n6861 ;
  assign n7170 = ( ~n1661 & n6861 ) | ( ~n1661 & n7006 ) | ( n6861 & n7006 ) ;
  assign n7171 = ( ~n6866 & n7169 ) | ( ~n6866 & n7170 ) | ( n7169 & n7170 ) ;
  assign n7172 = ( n6866 & n7169 ) | ( n6866 & n7170 ) | ( n7169 & n7170 ) ;
  assign n7173 = ( n6866 & n7171 ) | ( n6866 & ~n7172 ) | ( n7171 & ~n7172 ) ;
  assign n7174 = ( ~n1523 & n7168 ) | ( ~n1523 & n7173 ) | ( n7168 & n7173 ) ;
  assign n7175 = ~n1523 & n6867 ;
  assign n7176 = ( ~n1523 & n6867 ) | ( ~n1523 & n7006 ) | ( n6867 & n7006 ) ;
  assign n7177 = ( ~n6872 & n7175 ) | ( ~n6872 & n7176 ) | ( n7175 & n7176 ) ;
  assign n7178 = ( n6872 & n7175 ) | ( n6872 & n7176 ) | ( n7175 & n7176 ) ;
  assign n7179 = ( n6872 & n7177 ) | ( n6872 & ~n7178 ) | ( n7177 & ~n7178 ) ;
  assign n7180 = ( ~n1393 & n7174 ) | ( ~n1393 & n7179 ) | ( n7174 & n7179 ) ;
  assign n7181 = n1393 & ~n6873 ;
  assign n7182 = ( n1393 & ~n6873 ) | ( n1393 & n7006 ) | ( ~n6873 & n7006 ) ;
  assign n7183 = ( n6878 & n7181 ) | ( n6878 & n7182 ) | ( n7181 & n7182 ) ;
  assign n7184 = ( ~n6878 & n7181 ) | ( ~n6878 & n7182 ) | ( n7181 & n7182 ) ;
  assign n7185 = ( n6878 & ~n7183 ) | ( n6878 & n7184 ) | ( ~n7183 & n7184 ) ;
  assign n7186 = ( ~n1266 & n7180 ) | ( ~n1266 & n7185 ) | ( n7180 & n7185 ) ;
  assign n7187 = ( n1266 & ~n6879 ) | ( n1266 & n7006 ) | ( ~n6879 & n7006 ) ;
  assign n7188 = n1266 & ~n6879 ;
  assign n7189 = ( n6884 & n7187 ) | ( n6884 & n7188 ) | ( n7187 & n7188 ) ;
  assign n7190 = ( ~n6884 & n7187 ) | ( ~n6884 & n7188 ) | ( n7187 & n7188 ) ;
  assign n7191 = ( n6884 & ~n7189 ) | ( n6884 & n7190 ) | ( ~n7189 & n7190 ) ;
  assign n7192 = ( ~n1150 & n7186 ) | ( ~n1150 & n7191 ) | ( n7186 & n7191 ) ;
  assign n7193 = ~n1150 & n6885 ;
  assign n7194 = ( ~n1150 & n6885 ) | ( ~n1150 & n7006 ) | ( n6885 & n7006 ) ;
  assign n7195 = ( ~n6890 & n7193 ) | ( ~n6890 & n7194 ) | ( n7193 & n7194 ) ;
  assign n7196 = ( n6890 & n7193 ) | ( n6890 & n7194 ) | ( n7193 & n7194 ) ;
  assign n7197 = ( n6890 & n7195 ) | ( n6890 & ~n7196 ) | ( n7195 & ~n7196 ) ;
  assign n7198 = ( ~n1038 & n7192 ) | ( ~n1038 & n7197 ) | ( n7192 & n7197 ) ;
  assign n7199 = ( n1038 & ~n6891 ) | ( n1038 & n7006 ) | ( ~n6891 & n7006 ) ;
  assign n7200 = n1038 & ~n6891 ;
  assign n7201 = ( n6896 & n7199 ) | ( n6896 & n7200 ) | ( n7199 & n7200 ) ;
  assign n7202 = ( ~n6896 & n7199 ) | ( ~n6896 & n7200 ) | ( n7199 & n7200 ) ;
  assign n7203 = ( n6896 & ~n7201 ) | ( n6896 & n7202 ) | ( ~n7201 & n7202 ) ;
  assign n7204 = ( ~n933 & n7198 ) | ( ~n933 & n7203 ) | ( n7198 & n7203 ) ;
  assign n7205 = ~n933 & n6897 ;
  assign n7206 = ( ~n933 & n6897 ) | ( ~n933 & n7006 ) | ( n6897 & n7006 ) ;
  assign n7207 = ( n6902 & n7205 ) | ( n6902 & n7206 ) | ( n7205 & n7206 ) ;
  assign n7208 = ( ~n6902 & n7205 ) | ( ~n6902 & n7206 ) | ( n7205 & n7206 ) ;
  assign n7209 = ( n6902 & ~n7207 ) | ( n6902 & n7208 ) | ( ~n7207 & n7208 ) ;
  assign n7210 = ( ~n839 & n7204 ) | ( ~n839 & n7209 ) | ( n7204 & n7209 ) ;
  assign n7211 = ( n839 & ~n6903 ) | ( n839 & n7006 ) | ( ~n6903 & n7006 ) ;
  assign n7212 = n839 & ~n6903 ;
  assign n7213 = ( n6908 & n7211 ) | ( n6908 & n7212 ) | ( n7211 & n7212 ) ;
  assign n7214 = ( ~n6908 & n7211 ) | ( ~n6908 & n7212 ) | ( n7211 & n7212 ) ;
  assign n7215 = ( n6908 & ~n7213 ) | ( n6908 & n7214 ) | ( ~n7213 & n7214 ) ;
  assign n7216 = ( ~n746 & n7210 ) | ( ~n746 & n7215 ) | ( n7210 & n7215 ) ;
  assign n7217 = ( n746 & ~n6909 ) | ( n746 & n7006 ) | ( ~n6909 & n7006 ) ;
  assign n7218 = n746 & ~n6909 ;
  assign n7219 = ( n6914 & n7217 ) | ( n6914 & n7218 ) | ( n7217 & n7218 ) ;
  assign n7220 = ( ~n6914 & n7217 ) | ( ~n6914 & n7218 ) | ( n7217 & n7218 ) ;
  assign n7221 = ( n6914 & ~n7219 ) | ( n6914 & n7220 ) | ( ~n7219 & n7220 ) ;
  assign n7222 = ( ~n664 & n7216 ) | ( ~n664 & n7221 ) | ( n7216 & n7221 ) ;
  assign n7223 = ( n664 & ~n6915 ) | ( n664 & n7006 ) | ( ~n6915 & n7006 ) ;
  assign n7224 = n664 & ~n6915 ;
  assign n7225 = ( n6920 & n7223 ) | ( n6920 & n7224 ) | ( n7223 & n7224 ) ;
  assign n7226 = ( ~n6920 & n7223 ) | ( ~n6920 & n7224 ) | ( n7223 & n7224 ) ;
  assign n7227 = ( n6920 & ~n7225 ) | ( n6920 & n7226 ) | ( ~n7225 & n7226 ) ;
  assign n7228 = ( ~n588 & n7222 ) | ( ~n588 & n7227 ) | ( n7222 & n7227 ) ;
  assign n7229 = ( n588 & ~n6921 ) | ( n588 & n7006 ) | ( ~n6921 & n7006 ) ;
  assign n7230 = n588 & ~n6921 ;
  assign n7231 = ( n6926 & n7229 ) | ( n6926 & n7230 ) | ( n7229 & n7230 ) ;
  assign n7232 = ( ~n6926 & n7229 ) | ( ~n6926 & n7230 ) | ( n7229 & n7230 ) ;
  assign n7233 = ( n6926 & ~n7231 ) | ( n6926 & n7232 ) | ( ~n7231 & n7232 ) ;
  assign n7234 = ( ~n518 & n7228 ) | ( ~n518 & n7233 ) | ( n7228 & n7233 ) ;
  assign n7235 = ( n518 & ~n6927 ) | ( n518 & n7006 ) | ( ~n6927 & n7006 ) ;
  assign n7236 = n518 & ~n6927 ;
  assign n7237 = ( n6932 & n7235 ) | ( n6932 & n7236 ) | ( n7235 & n7236 ) ;
  assign n7238 = ( ~n6932 & n7235 ) | ( ~n6932 & n7236 ) | ( n7235 & n7236 ) ;
  assign n7239 = ( n6932 & ~n7237 ) | ( n6932 & n7238 ) | ( ~n7237 & n7238 ) ;
  assign n7240 = ( ~n454 & n7234 ) | ( ~n454 & n7239 ) | ( n7234 & n7239 ) ;
  assign n7241 = ( n454 & ~n6933 ) | ( n454 & n7006 ) | ( ~n6933 & n7006 ) ;
  assign n7242 = n454 & ~n6933 ;
  assign n7243 = ( n6938 & n7241 ) | ( n6938 & n7242 ) | ( n7241 & n7242 ) ;
  assign n7244 = ( ~n6938 & n7241 ) | ( ~n6938 & n7242 ) | ( n7241 & n7242 ) ;
  assign n7245 = ( n6938 & ~n7243 ) | ( n6938 & n7244 ) | ( ~n7243 & n7244 ) ;
  assign n7246 = ( ~n396 & n7240 ) | ( ~n396 & n7245 ) | ( n7240 & n7245 ) ;
  assign n7247 = ( n396 & ~n6939 ) | ( n396 & n7006 ) | ( ~n6939 & n7006 ) ;
  assign n7248 = n396 & ~n6939 ;
  assign n7249 = ( n6944 & n7247 ) | ( n6944 & n7248 ) | ( n7247 & n7248 ) ;
  assign n7250 = ( ~n6944 & n7247 ) | ( ~n6944 & n7248 ) | ( n7247 & n7248 ) ;
  assign n7251 = ( n6944 & ~n7249 ) | ( n6944 & n7250 ) | ( ~n7249 & n7250 ) ;
  assign n7252 = ( ~n344 & n7246 ) | ( ~n344 & n7251 ) | ( n7246 & n7251 ) ;
  assign n7253 = ( n344 & ~n6945 ) | ( n344 & n7006 ) | ( ~n6945 & n7006 ) ;
  assign n7254 = n344 & ~n6945 ;
  assign n7255 = ( n6950 & n7253 ) | ( n6950 & n7254 ) | ( n7253 & n7254 ) ;
  assign n7256 = ( ~n6950 & n7253 ) | ( ~n6950 & n7254 ) | ( n7253 & n7254 ) ;
  assign n7257 = ( n6950 & ~n7255 ) | ( n6950 & n7256 ) | ( ~n7255 & n7256 ) ;
  assign n7258 = ( ~n298 & n7252 ) | ( ~n298 & n7257 ) | ( n7252 & n7257 ) ;
  assign n7259 = n298 & ~n6951 ;
  assign n7260 = ( n298 & ~n6951 ) | ( n298 & n7006 ) | ( ~n6951 & n7006 ) ;
  assign n7261 = ( n6956 & n7259 ) | ( n6956 & n7260 ) | ( n7259 & n7260 ) ;
  assign n7262 = ( ~n6956 & n7259 ) | ( ~n6956 & n7260 ) | ( n7259 & n7260 ) ;
  assign n7263 = ( n6956 & ~n7261 ) | ( n6956 & n7262 ) | ( ~n7261 & n7262 ) ;
  assign n7264 = ( ~n258 & n7258 ) | ( ~n258 & n7263 ) | ( n7258 & n7263 ) ;
  assign n7265 = ( n258 & ~n6957 ) | ( n258 & n7006 ) | ( ~n6957 & n7006 ) ;
  assign n7266 = n258 & ~n6957 ;
  assign n7267 = ( n6962 & n7265 ) | ( n6962 & n7266 ) | ( n7265 & n7266 ) ;
  assign n7268 = ( ~n6962 & n7265 ) | ( ~n6962 & n7266 ) | ( n7265 & n7266 ) ;
  assign n7269 = ( n6962 & ~n7267 ) | ( n6962 & n7268 ) | ( ~n7267 & n7268 ) ;
  assign n7270 = ( ~n225 & n7264 ) | ( ~n225 & n7269 ) | ( n7264 & n7269 ) ;
  assign n7271 = ( n225 & ~n6963 ) | ( n225 & n7006 ) | ( ~n6963 & n7006 ) ;
  assign n7272 = n225 & ~n6963 ;
  assign n7273 = ( n6968 & n7271 ) | ( n6968 & n7272 ) | ( n7271 & n7272 ) ;
  assign n7274 = ( ~n6968 & n7271 ) | ( ~n6968 & n7272 ) | ( n7271 & n7272 ) ;
  assign n7275 = ( n6968 & ~n7273 ) | ( n6968 & n7274 ) | ( ~n7273 & n7274 ) ;
  assign n7276 = ( ~n197 & n7270 ) | ( ~n197 & n7275 ) | ( n7270 & n7275 ) ;
  assign n7277 = ( n197 & ~n6969 ) | ( n197 & n7006 ) | ( ~n6969 & n7006 ) ;
  assign n7278 = n197 & ~n6969 ;
  assign n7279 = ( n6974 & n7277 ) | ( n6974 & n7278 ) | ( n7277 & n7278 ) ;
  assign n7280 = ( ~n6974 & n7277 ) | ( ~n6974 & n7278 ) | ( n7277 & n7278 ) ;
  assign n7281 = ( n6974 & ~n7279 ) | ( n6974 & n7280 ) | ( ~n7279 & n7280 ) ;
  assign n7282 = ( ~n170 & n7276 ) | ( ~n170 & n7281 ) | ( n7276 & n7281 ) ;
  assign n7283 = ~n170 & n6975 ;
  assign n7284 = ( ~n170 & n6975 ) | ( ~n170 & n7006 ) | ( n6975 & n7006 ) ;
  assign n7285 = ( ~n6980 & n7283 ) | ( ~n6980 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7286 = ( n6980 & n7283 ) | ( n6980 & n7284 ) | ( n7283 & n7284 ) ;
  assign n7287 = ( n6980 & n7285 ) | ( n6980 & ~n7286 ) | ( n7285 & ~n7286 ) ;
  assign n7288 = ( ~n142 & n7282 ) | ( ~n142 & n7287 ) | ( n7282 & n7287 ) ;
  assign n7289 = ~n142 & n6981 ;
  assign n7290 = ( ~n142 & n6981 ) | ( ~n142 & n7006 ) | ( n6981 & n7006 ) ;
  assign n7291 = ( ~n6986 & n7289 ) | ( ~n6986 & n7290 ) | ( n7289 & n7290 ) ;
  assign n7292 = ( n6986 & n7289 ) | ( n6986 & n7290 ) | ( n7289 & n7290 ) ;
  assign n7293 = ( n6986 & n7291 ) | ( n6986 & ~n7292 ) | ( n7291 & ~n7292 ) ;
  assign n7294 = ( ~n132 & n7288 ) | ( ~n132 & n7293 ) | ( n7288 & n7293 ) ;
  assign n7295 = ( ~n131 & n7018 ) | ( ~n131 & n7294 ) | ( n7018 & n7294 ) ;
  assign n7296 = n7013 | n7295 ;
  assign n7297 = n6993 & ~n7011 ;
  assign n7298 = n6993 | n6998 ;
  assign n7299 = ( n7018 & ~n7297 ) | ( n7018 & n7298 ) | ( ~n7297 & n7298 ) ;
  assign n7300 = ( n7018 & n7294 ) | ( n7018 & n7299 ) | ( n7294 & n7299 ) ;
  assign n7301 = ~n7295 & n7300 ;
  assign n7302 = ( ~n7018 & n7294 ) | ( ~n7018 & n7296 ) | ( n7294 & n7296 ) ;
  assign n7303 = ( n131 & ~n7018 ) | ( n131 & n7294 ) | ( ~n7018 & n7294 ) ;
  assign n7304 = n7302 & ~n7303 ;
  assign n7305 = n7301 | n7304 ;
  assign n7306 = ( n132 & ~n7288 ) | ( n132 & n7296 ) | ( ~n7288 & n7296 ) ;
  assign n7307 = n132 & ~n7288 ;
  assign n7308 = ( n7293 & n7306 ) | ( n7293 & n7307 ) | ( n7306 & n7307 ) ;
  assign n7309 = ( n7293 & ~n7306 ) | ( n7293 & n7307 ) | ( ~n7306 & n7307 ) ;
  assign n7310 = ( n7306 & ~n7308 ) | ( n7306 & n7309 ) | ( ~n7308 & n7309 ) ;
  assign n7311 = ~n7024 & n7296 ;
  assign n7312 = x28 | x29 ;
  assign n7313 = x30 | n7312 ;
  assign n7314 = n7006 & ~n7313 ;
  assign n7315 = ~n7006 & n7313 ;
  assign n7316 = ( x31 & ~n7296 ) | ( x31 & n7315 ) | ( ~n7296 & n7315 ) ;
  assign n7317 = ( n7311 & ~n7314 ) | ( n7311 & n7316 ) | ( ~n7314 & n7316 ) ;
  assign n7318 = n7006 & ~n7296 ;
  assign n7319 = ( ~x32 & n7311 ) | ( ~x32 & n7318 ) | ( n7311 & n7318 ) ;
  assign n7320 = ( x32 & n7311 ) | ( x32 & n7318 ) | ( n7311 & n7318 ) ;
  assign n7321 = ( x32 & n7319 ) | ( x32 & ~n7320 ) | ( n7319 & ~n7320 ) ;
  assign n7322 = ( ~n6723 & n7317 ) | ( ~n6723 & n7321 ) | ( n7317 & n7321 ) ;
  assign n7323 = ~n6723 & n7006 ;
  assign n7324 = ( n7019 & n7296 ) | ( n7019 & n7323 ) | ( n7296 & n7323 ) ;
  assign n7325 = ( x33 & n7319 ) | ( x33 & n7324 ) | ( n7319 & n7324 ) ;
  assign n7326 = ( ~x33 & n7319 ) | ( ~x33 & n7324 ) | ( n7319 & n7324 ) ;
  assign n7327 = ( x33 & ~n7325 ) | ( x33 & n7326 ) | ( ~n7325 & n7326 ) ;
  assign n7328 = ( ~n6442 & n7322 ) | ( ~n6442 & n7327 ) | ( n7322 & n7327 ) ;
  assign n7329 = ( ~n6442 & n7029 ) | ( ~n6442 & n7296 ) | ( n7029 & n7296 ) ;
  assign n7330 = ~n6442 & n7029 ;
  assign n7331 = ( ~n7023 & n7329 ) | ( ~n7023 & n7330 ) | ( n7329 & n7330 ) ;
  assign n7332 = ( n7023 & n7329 ) | ( n7023 & n7330 ) | ( n7329 & n7330 ) ;
  assign n7333 = ( n7023 & n7331 ) | ( n7023 & ~n7332 ) | ( n7331 & ~n7332 ) ;
  assign n7334 = ( ~n6172 & n7328 ) | ( ~n6172 & n7333 ) | ( n7328 & n7333 ) ;
  assign n7335 = n6172 & ~n7030 ;
  assign n7336 = ( n6172 & ~n7030 ) | ( n6172 & n7296 ) | ( ~n7030 & n7296 ) ;
  assign n7337 = ( n7035 & n7335 ) | ( n7035 & n7336 ) | ( n7335 & n7336 ) ;
  assign n7338 = ( ~n7035 & n7335 ) | ( ~n7035 & n7336 ) | ( n7335 & n7336 ) ;
  assign n7339 = ( n7035 & ~n7337 ) | ( n7035 & n7338 ) | ( ~n7337 & n7338 ) ;
  assign n7340 = ( ~n5905 & n7334 ) | ( ~n5905 & n7339 ) | ( n7334 & n7339 ) ;
  assign n7341 = n5905 & ~n7036 ;
  assign n7342 = ( n5905 & ~n7036 ) | ( n5905 & n7296 ) | ( ~n7036 & n7296 ) ;
  assign n7343 = ( ~n7041 & n7341 ) | ( ~n7041 & n7342 ) | ( n7341 & n7342 ) ;
  assign n7344 = ( n7041 & n7341 ) | ( n7041 & n7342 ) | ( n7341 & n7342 ) ;
  assign n7345 = ( n7041 & n7343 ) | ( n7041 & ~n7344 ) | ( n7343 & ~n7344 ) ;
  assign n7346 = ( ~n5642 & n7340 ) | ( ~n5642 & n7345 ) | ( n7340 & n7345 ) ;
  assign n7347 = ( n5642 & ~n7042 ) | ( n5642 & n7296 ) | ( ~n7042 & n7296 ) ;
  assign n7348 = n5642 & ~n7042 ;
  assign n7349 = ( n7047 & n7347 ) | ( n7047 & n7348 ) | ( n7347 & n7348 ) ;
  assign n7350 = ( ~n7047 & n7347 ) | ( ~n7047 & n7348 ) | ( n7347 & n7348 ) ;
  assign n7351 = ( n7047 & ~n7349 ) | ( n7047 & n7350 ) | ( ~n7349 & n7350 ) ;
  assign n7352 = ( ~n5386 & n7346 ) | ( ~n5386 & n7351 ) | ( n7346 & n7351 ) ;
  assign n7353 = ~n5386 & n7048 ;
  assign n7354 = ( ~n5386 & n7048 ) | ( ~n5386 & n7296 ) | ( n7048 & n7296 ) ;
  assign n7355 = ( ~n7053 & n7353 ) | ( ~n7053 & n7354 ) | ( n7353 & n7354 ) ;
  assign n7356 = ( n7053 & n7353 ) | ( n7053 & n7354 ) | ( n7353 & n7354 ) ;
  assign n7357 = ( n7053 & n7355 ) | ( n7053 & ~n7356 ) | ( n7355 & ~n7356 ) ;
  assign n7358 = ( ~n5139 & n7352 ) | ( ~n5139 & n7357 ) | ( n7352 & n7357 ) ;
  assign n7359 = ~n5139 & n7054 ;
  assign n7360 = ( ~n5139 & n7054 ) | ( ~n5139 & n7296 ) | ( n7054 & n7296 ) ;
  assign n7361 = ( ~n7059 & n7359 ) | ( ~n7059 & n7360 ) | ( n7359 & n7360 ) ;
  assign n7362 = ( n7059 & n7359 ) | ( n7059 & n7360 ) | ( n7359 & n7360 ) ;
  assign n7363 = ( n7059 & n7361 ) | ( n7059 & ~n7362 ) | ( n7361 & ~n7362 ) ;
  assign n7364 = ( ~n4898 & n7358 ) | ( ~n4898 & n7363 ) | ( n7358 & n7363 ) ;
  assign n7365 = ~n4898 & n7060 ;
  assign n7366 = ( ~n4898 & n7060 ) | ( ~n4898 & n7296 ) | ( n7060 & n7296 ) ;
  assign n7367 = ( ~n7065 & n7365 ) | ( ~n7065 & n7366 ) | ( n7365 & n7366 ) ;
  assign n7368 = ( n7065 & n7365 ) | ( n7065 & n7366 ) | ( n7365 & n7366 ) ;
  assign n7369 = ( n7065 & n7367 ) | ( n7065 & ~n7368 ) | ( n7367 & ~n7368 ) ;
  assign n7370 = ( ~n4661 & n7364 ) | ( ~n4661 & n7369 ) | ( n7364 & n7369 ) ;
  assign n7371 = ( n4661 & ~n7066 ) | ( n4661 & n7296 ) | ( ~n7066 & n7296 ) ;
  assign n7372 = n4661 & ~n7066 ;
  assign n7373 = ( n7071 & n7371 ) | ( n7071 & n7372 ) | ( n7371 & n7372 ) ;
  assign n7374 = ( ~n7071 & n7371 ) | ( ~n7071 & n7372 ) | ( n7371 & n7372 ) ;
  assign n7375 = ( n7071 & ~n7373 ) | ( n7071 & n7374 ) | ( ~n7373 & n7374 ) ;
  assign n7376 = ( ~n4432 & n7370 ) | ( ~n4432 & n7375 ) | ( n7370 & n7375 ) ;
  assign n7377 = ( n4432 & ~n7072 ) | ( n4432 & n7296 ) | ( ~n7072 & n7296 ) ;
  assign n7378 = n4432 & ~n7072 ;
  assign n7379 = ( n7077 & n7377 ) | ( n7077 & n7378 ) | ( n7377 & n7378 ) ;
  assign n7380 = ( ~n7077 & n7377 ) | ( ~n7077 & n7378 ) | ( n7377 & n7378 ) ;
  assign n7381 = ( n7077 & ~n7379 ) | ( n7077 & n7380 ) | ( ~n7379 & n7380 ) ;
  assign n7382 = ( ~n4203 & n7376 ) | ( ~n4203 & n7381 ) | ( n7376 & n7381 ) ;
  assign n7383 = ( n4203 & ~n7078 ) | ( n4203 & n7296 ) | ( ~n7078 & n7296 ) ;
  assign n7384 = n4203 & ~n7078 ;
  assign n7385 = ( n7083 & n7383 ) | ( n7083 & n7384 ) | ( n7383 & n7384 ) ;
  assign n7386 = ( ~n7083 & n7383 ) | ( ~n7083 & n7384 ) | ( n7383 & n7384 ) ;
  assign n7387 = ( n7083 & ~n7385 ) | ( n7083 & n7386 ) | ( ~n7385 & n7386 ) ;
  assign n7388 = ( ~n3985 & n7382 ) | ( ~n3985 & n7387 ) | ( n7382 & n7387 ) ;
  assign n7389 = ~n3985 & n7084 ;
  assign n7390 = ( ~n3985 & n7084 ) | ( ~n3985 & n7296 ) | ( n7084 & n7296 ) ;
  assign n7391 = ( ~n7089 & n7389 ) | ( ~n7089 & n7390 ) | ( n7389 & n7390 ) ;
  assign n7392 = ( n7089 & n7389 ) | ( n7089 & n7390 ) | ( n7389 & n7390 ) ;
  assign n7393 = ( n7089 & n7391 ) | ( n7089 & ~n7392 ) | ( n7391 & ~n7392 ) ;
  assign n7394 = ( ~n3772 & n7388 ) | ( ~n3772 & n7393 ) | ( n7388 & n7393 ) ;
  assign n7395 = ~n3772 & n7090 ;
  assign n7396 = ( ~n3772 & n7090 ) | ( ~n3772 & n7296 ) | ( n7090 & n7296 ) ;
  assign n7397 = ( ~n7095 & n7395 ) | ( ~n7095 & n7396 ) | ( n7395 & n7396 ) ;
  assign n7398 = ( n7095 & n7395 ) | ( n7095 & n7396 ) | ( n7395 & n7396 ) ;
  assign n7399 = ( n7095 & n7397 ) | ( n7095 & ~n7398 ) | ( n7397 & ~n7398 ) ;
  assign n7400 = ( ~n3567 & n7394 ) | ( ~n3567 & n7399 ) | ( n7394 & n7399 ) ;
  assign n7401 = ~n3567 & n7096 ;
  assign n7402 = ( ~n3567 & n7096 ) | ( ~n3567 & n7296 ) | ( n7096 & n7296 ) ;
  assign n7403 = ( ~n7101 & n7401 ) | ( ~n7101 & n7402 ) | ( n7401 & n7402 ) ;
  assign n7404 = ( n7101 & n7401 ) | ( n7101 & n7402 ) | ( n7401 & n7402 ) ;
  assign n7405 = ( n7101 & n7403 ) | ( n7101 & ~n7404 ) | ( n7403 & ~n7404 ) ;
  assign n7406 = ( ~n3362 & n7400 ) | ( ~n3362 & n7405 ) | ( n7400 & n7405 ) ;
  assign n7407 = ~n3362 & n7102 ;
  assign n7408 = ( ~n3362 & n7102 ) | ( ~n3362 & n7296 ) | ( n7102 & n7296 ) ;
  assign n7409 = ( ~n7107 & n7407 ) | ( ~n7107 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7410 = ( n7107 & n7407 ) | ( n7107 & n7408 ) | ( n7407 & n7408 ) ;
  assign n7411 = ( n7107 & n7409 ) | ( n7107 & ~n7410 ) | ( n7409 & ~n7410 ) ;
  assign n7412 = ( ~n3169 & n7406 ) | ( ~n3169 & n7411 ) | ( n7406 & n7411 ) ;
  assign n7413 = ( n3169 & ~n7108 ) | ( n3169 & n7296 ) | ( ~n7108 & n7296 ) ;
  assign n7414 = n3169 & ~n7108 ;
  assign n7415 = ( n7113 & n7413 ) | ( n7113 & n7414 ) | ( n7413 & n7414 ) ;
  assign n7416 = ( ~n7113 & n7413 ) | ( ~n7113 & n7414 ) | ( n7413 & n7414 ) ;
  assign n7417 = ( n7113 & ~n7415 ) | ( n7113 & n7416 ) | ( ~n7415 & n7416 ) ;
  assign n7418 = ( ~n2979 & n7412 ) | ( ~n2979 & n7417 ) | ( n7412 & n7417 ) ;
  assign n7419 = ~n2979 & n7114 ;
  assign n7420 = ( ~n2979 & n7114 ) | ( ~n2979 & n7296 ) | ( n7114 & n7296 ) ;
  assign n7421 = ( ~n7119 & n7419 ) | ( ~n7119 & n7420 ) | ( n7419 & n7420 ) ;
  assign n7422 = ( n7119 & n7419 ) | ( n7119 & n7420 ) | ( n7419 & n7420 ) ;
  assign n7423 = ( n7119 & n7421 ) | ( n7119 & ~n7422 ) | ( n7421 & ~n7422 ) ;
  assign n7424 = ( ~n2791 & n7418 ) | ( ~n2791 & n7423 ) | ( n7418 & n7423 ) ;
  assign n7425 = n2791 & ~n7120 ;
  assign n7426 = ( n2791 & ~n7120 ) | ( n2791 & n7296 ) | ( ~n7120 & n7296 ) ;
  assign n7427 = ( n7125 & n7425 ) | ( n7125 & n7426 ) | ( n7425 & n7426 ) ;
  assign n7428 = ( ~n7125 & n7425 ) | ( ~n7125 & n7426 ) | ( n7425 & n7426 ) ;
  assign n7429 = ( n7125 & ~n7427 ) | ( n7125 & n7428 ) | ( ~n7427 & n7428 ) ;
  assign n7430 = ( ~n2615 & n7424 ) | ( ~n2615 & n7429 ) | ( n7424 & n7429 ) ;
  assign n7431 = ( n2615 & ~n7126 ) | ( n2615 & n7296 ) | ( ~n7126 & n7296 ) ;
  assign n7432 = n2615 & ~n7126 ;
  assign n7433 = ( n7131 & n7431 ) | ( n7131 & n7432 ) | ( n7431 & n7432 ) ;
  assign n7434 = ( ~n7131 & n7431 ) | ( ~n7131 & n7432 ) | ( n7431 & n7432 ) ;
  assign n7435 = ( n7131 & ~n7433 ) | ( n7131 & n7434 ) | ( ~n7433 & n7434 ) ;
  assign n7436 = ( ~n2443 & n7430 ) | ( ~n2443 & n7435 ) | ( n7430 & n7435 ) ;
  assign n7437 = ( n2443 & ~n7132 ) | ( n2443 & n7296 ) | ( ~n7132 & n7296 ) ;
  assign n7438 = n2443 & ~n7132 ;
  assign n7439 = ( n7137 & n7437 ) | ( n7137 & n7438 ) | ( n7437 & n7438 ) ;
  assign n7440 = ( ~n7137 & n7437 ) | ( ~n7137 & n7438 ) | ( n7437 & n7438 ) ;
  assign n7441 = ( n7137 & ~n7439 ) | ( n7137 & n7440 ) | ( ~n7439 & n7440 ) ;
  assign n7442 = ( ~n2277 & n7436 ) | ( ~n2277 & n7441 ) | ( n7436 & n7441 ) ;
  assign n7443 = n2277 & ~n7138 ;
  assign n7444 = ( n2277 & ~n7138 ) | ( n2277 & n7296 ) | ( ~n7138 & n7296 ) ;
  assign n7445 = ( n7143 & n7443 ) | ( n7143 & n7444 ) | ( n7443 & n7444 ) ;
  assign n7446 = ( ~n7143 & n7443 ) | ( ~n7143 & n7444 ) | ( n7443 & n7444 ) ;
  assign n7447 = ( n7143 & ~n7445 ) | ( n7143 & n7446 ) | ( ~n7445 & n7446 ) ;
  assign n7448 = ( ~n2111 & n7442 ) | ( ~n2111 & n7447 ) | ( n7442 & n7447 ) ;
  assign n7449 = ( n2111 & ~n7144 ) | ( n2111 & n7296 ) | ( ~n7144 & n7296 ) ;
  assign n7450 = n2111 & ~n7144 ;
  assign n7451 = ( n7149 & n7449 ) | ( n7149 & n7450 ) | ( n7449 & n7450 ) ;
  assign n7452 = ( ~n7149 & n7449 ) | ( ~n7149 & n7450 ) | ( n7449 & n7450 ) ;
  assign n7453 = ( n7149 & ~n7451 ) | ( n7149 & n7452 ) | ( ~n7451 & n7452 ) ;
  assign n7454 = ( ~n1949 & n7448 ) | ( ~n1949 & n7453 ) | ( n7448 & n7453 ) ;
  assign n7455 = ( n1949 & ~n7150 ) | ( n1949 & n7296 ) | ( ~n7150 & n7296 ) ;
  assign n7456 = n1949 & ~n7150 ;
  assign n7457 = ( n7155 & n7455 ) | ( n7155 & n7456 ) | ( n7455 & n7456 ) ;
  assign n7458 = ( ~n7155 & n7455 ) | ( ~n7155 & n7456 ) | ( n7455 & n7456 ) ;
  assign n7459 = ( n7155 & ~n7457 ) | ( n7155 & n7458 ) | ( ~n7457 & n7458 ) ;
  assign n7460 = ( ~n1802 & n7454 ) | ( ~n1802 & n7459 ) | ( n7454 & n7459 ) ;
  assign n7461 = ( n1802 & ~n7156 ) | ( n1802 & n7296 ) | ( ~n7156 & n7296 ) ;
  assign n7462 = n1802 & ~n7156 ;
  assign n7463 = ( n7161 & n7461 ) | ( n7161 & n7462 ) | ( n7461 & n7462 ) ;
  assign n7464 = ( ~n7161 & n7461 ) | ( ~n7161 & n7462 ) | ( n7461 & n7462 ) ;
  assign n7465 = ( n7161 & ~n7463 ) | ( n7161 & n7464 ) | ( ~n7463 & n7464 ) ;
  assign n7466 = ( ~n1661 & n7460 ) | ( ~n1661 & n7465 ) | ( n7460 & n7465 ) ;
  assign n7467 = ~n1661 & n7162 ;
  assign n7468 = ( ~n1661 & n7162 ) | ( ~n1661 & n7296 ) | ( n7162 & n7296 ) ;
  assign n7469 = ( n7167 & n7467 ) | ( n7167 & n7468 ) | ( n7467 & n7468 ) ;
  assign n7470 = ( ~n7167 & n7467 ) | ( ~n7167 & n7468 ) | ( n7467 & n7468 ) ;
  assign n7471 = ( n7167 & ~n7469 ) | ( n7167 & n7470 ) | ( ~n7469 & n7470 ) ;
  assign n7472 = ( ~n1523 & n7466 ) | ( ~n1523 & n7471 ) | ( n7466 & n7471 ) ;
  assign n7473 = ( n1523 & ~n7168 ) | ( n1523 & n7296 ) | ( ~n7168 & n7296 ) ;
  assign n7474 = n1523 & ~n7168 ;
  assign n7475 = ( n7173 & n7473 ) | ( n7173 & n7474 ) | ( n7473 & n7474 ) ;
  assign n7476 = ( ~n7173 & n7473 ) | ( ~n7173 & n7474 ) | ( n7473 & n7474 ) ;
  assign n7477 = ( n7173 & ~n7475 ) | ( n7173 & n7476 ) | ( ~n7475 & n7476 ) ;
  assign n7478 = ( ~n1393 & n7472 ) | ( ~n1393 & n7477 ) | ( n7472 & n7477 ) ;
  assign n7479 = ~n1393 & n7174 ;
  assign n7480 = ( ~n1393 & n7174 ) | ( ~n1393 & n7296 ) | ( n7174 & n7296 ) ;
  assign n7481 = ( n7179 & n7479 ) | ( n7179 & n7480 ) | ( n7479 & n7480 ) ;
  assign n7482 = ( ~n7179 & n7479 ) | ( ~n7179 & n7480 ) | ( n7479 & n7480 ) ;
  assign n7483 = ( n7179 & ~n7481 ) | ( n7179 & n7482 ) | ( ~n7481 & n7482 ) ;
  assign n7484 = ( ~n1266 & n7478 ) | ( ~n1266 & n7483 ) | ( n7478 & n7483 ) ;
  assign n7485 = ( n1266 & ~n7180 ) | ( n1266 & n7296 ) | ( ~n7180 & n7296 ) ;
  assign n7486 = n1266 & ~n7180 ;
  assign n7487 = ( n7185 & n7485 ) | ( n7185 & n7486 ) | ( n7485 & n7486 ) ;
  assign n7488 = ( ~n7185 & n7485 ) | ( ~n7185 & n7486 ) | ( n7485 & n7486 ) ;
  assign n7489 = ( n7185 & ~n7487 ) | ( n7185 & n7488 ) | ( ~n7487 & n7488 ) ;
  assign n7490 = ( ~n1150 & n7484 ) | ( ~n1150 & n7489 ) | ( n7484 & n7489 ) ;
  assign n7491 = ( n1150 & ~n7186 ) | ( n1150 & n7296 ) | ( ~n7186 & n7296 ) ;
  assign n7492 = n1150 & ~n7186 ;
  assign n7493 = ( n7191 & n7491 ) | ( n7191 & n7492 ) | ( n7491 & n7492 ) ;
  assign n7494 = ( ~n7191 & n7491 ) | ( ~n7191 & n7492 ) | ( n7491 & n7492 ) ;
  assign n7495 = ( n7191 & ~n7493 ) | ( n7191 & n7494 ) | ( ~n7493 & n7494 ) ;
  assign n7496 = ( ~n1038 & n7490 ) | ( ~n1038 & n7495 ) | ( n7490 & n7495 ) ;
  assign n7497 = ~n1038 & n7192 ;
  assign n7498 = ( ~n1038 & n7192 ) | ( ~n1038 & n7296 ) | ( n7192 & n7296 ) ;
  assign n7499 = ( ~n7197 & n7497 ) | ( ~n7197 & n7498 ) | ( n7497 & n7498 ) ;
  assign n7500 = ( n7197 & n7497 ) | ( n7197 & n7498 ) | ( n7497 & n7498 ) ;
  assign n7501 = ( n7197 & n7499 ) | ( n7197 & ~n7500 ) | ( n7499 & ~n7500 ) ;
  assign n7502 = ( ~n933 & n7496 ) | ( ~n933 & n7501 ) | ( n7496 & n7501 ) ;
  assign n7503 = ( n933 & ~n7198 ) | ( n933 & n7296 ) | ( ~n7198 & n7296 ) ;
  assign n7504 = n933 & ~n7198 ;
  assign n7505 = ( n7203 & n7503 ) | ( n7203 & n7504 ) | ( n7503 & n7504 ) ;
  assign n7506 = ( ~n7203 & n7503 ) | ( ~n7203 & n7504 ) | ( n7503 & n7504 ) ;
  assign n7507 = ( n7203 & ~n7505 ) | ( n7203 & n7506 ) | ( ~n7505 & n7506 ) ;
  assign n7508 = ( ~n839 & n7502 ) | ( ~n839 & n7507 ) | ( n7502 & n7507 ) ;
  assign n7509 = ( n839 & ~n7204 ) | ( n839 & n7296 ) | ( ~n7204 & n7296 ) ;
  assign n7510 = n839 & ~n7204 ;
  assign n7511 = ( n7209 & n7509 ) | ( n7209 & n7510 ) | ( n7509 & n7510 ) ;
  assign n7512 = ( ~n7209 & n7509 ) | ( ~n7209 & n7510 ) | ( n7509 & n7510 ) ;
  assign n7513 = ( n7209 & ~n7511 ) | ( n7209 & n7512 ) | ( ~n7511 & n7512 ) ;
  assign n7514 = ( ~n746 & n7508 ) | ( ~n746 & n7513 ) | ( n7508 & n7513 ) ;
  assign n7515 = ( n746 & ~n7210 ) | ( n746 & n7296 ) | ( ~n7210 & n7296 ) ;
  assign n7516 = n746 & ~n7210 ;
  assign n7517 = ( n7215 & n7515 ) | ( n7215 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7518 = ( ~n7215 & n7515 ) | ( ~n7215 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7519 = ( n7215 & ~n7517 ) | ( n7215 & n7518 ) | ( ~n7517 & n7518 ) ;
  assign n7520 = ( ~n664 & n7514 ) | ( ~n664 & n7519 ) | ( n7514 & n7519 ) ;
  assign n7521 = ~n664 & n7216 ;
  assign n7522 = ( ~n664 & n7216 ) | ( ~n664 & n7296 ) | ( n7216 & n7296 ) ;
  assign n7523 = ( ~n7221 & n7521 ) | ( ~n7221 & n7522 ) | ( n7521 & n7522 ) ;
  assign n7524 = ( n7221 & n7521 ) | ( n7221 & n7522 ) | ( n7521 & n7522 ) ;
  assign n7525 = ( n7221 & n7523 ) | ( n7221 & ~n7524 ) | ( n7523 & ~n7524 ) ;
  assign n7526 = ( ~n588 & n7520 ) | ( ~n588 & n7525 ) | ( n7520 & n7525 ) ;
  assign n7527 = ~n588 & n7222 ;
  assign n7528 = ( ~n588 & n7222 ) | ( ~n588 & n7296 ) | ( n7222 & n7296 ) ;
  assign n7529 = ( ~n7227 & n7527 ) | ( ~n7227 & n7528 ) | ( n7527 & n7528 ) ;
  assign n7530 = ( n7227 & n7527 ) | ( n7227 & n7528 ) | ( n7527 & n7528 ) ;
  assign n7531 = ( n7227 & n7529 ) | ( n7227 & ~n7530 ) | ( n7529 & ~n7530 ) ;
  assign n7532 = ( ~n518 & n7526 ) | ( ~n518 & n7531 ) | ( n7526 & n7531 ) ;
  assign n7533 = ( n518 & ~n7228 ) | ( n518 & n7296 ) | ( ~n7228 & n7296 ) ;
  assign n7534 = n518 & ~n7228 ;
  assign n7535 = ( n7233 & n7533 ) | ( n7233 & n7534 ) | ( n7533 & n7534 ) ;
  assign n7536 = ( ~n7233 & n7533 ) | ( ~n7233 & n7534 ) | ( n7533 & n7534 ) ;
  assign n7537 = ( n7233 & ~n7535 ) | ( n7233 & n7536 ) | ( ~n7535 & n7536 ) ;
  assign n7538 = ( ~n454 & n7532 ) | ( ~n454 & n7537 ) | ( n7532 & n7537 ) ;
  assign n7539 = ~n454 & n7234 ;
  assign n7540 = ( ~n454 & n7234 ) | ( ~n454 & n7296 ) | ( n7234 & n7296 ) ;
  assign n7541 = ( ~n7239 & n7539 ) | ( ~n7239 & n7540 ) | ( n7539 & n7540 ) ;
  assign n7542 = ( n7239 & n7539 ) | ( n7239 & n7540 ) | ( n7539 & n7540 ) ;
  assign n7543 = ( n7239 & n7541 ) | ( n7239 & ~n7542 ) | ( n7541 & ~n7542 ) ;
  assign n7544 = ( ~n396 & n7538 ) | ( ~n396 & n7543 ) | ( n7538 & n7543 ) ;
  assign n7545 = ~n396 & n7240 ;
  assign n7546 = ( ~n396 & n7240 ) | ( ~n396 & n7296 ) | ( n7240 & n7296 ) ;
  assign n7547 = ( ~n7245 & n7545 ) | ( ~n7245 & n7546 ) | ( n7545 & n7546 ) ;
  assign n7548 = ( n7245 & n7545 ) | ( n7245 & n7546 ) | ( n7545 & n7546 ) ;
  assign n7549 = ( n7245 & n7547 ) | ( n7245 & ~n7548 ) | ( n7547 & ~n7548 ) ;
  assign n7550 = ( ~n344 & n7544 ) | ( ~n344 & n7549 ) | ( n7544 & n7549 ) ;
  assign n7551 = ( n344 & ~n7246 ) | ( n344 & n7296 ) | ( ~n7246 & n7296 ) ;
  assign n7552 = n344 & ~n7246 ;
  assign n7553 = ( n7251 & n7551 ) | ( n7251 & n7552 ) | ( n7551 & n7552 ) ;
  assign n7554 = ( ~n7251 & n7551 ) | ( ~n7251 & n7552 ) | ( n7551 & n7552 ) ;
  assign n7555 = ( n7251 & ~n7553 ) | ( n7251 & n7554 ) | ( ~n7553 & n7554 ) ;
  assign n7556 = ( ~n298 & n7550 ) | ( ~n298 & n7555 ) | ( n7550 & n7555 ) ;
  assign n7557 = ~n298 & n7252 ;
  assign n7558 = ( ~n298 & n7252 ) | ( ~n298 & n7296 ) | ( n7252 & n7296 ) ;
  assign n7559 = ( n7257 & n7557 ) | ( n7257 & n7558 ) | ( n7557 & n7558 ) ;
  assign n7560 = ( ~n7257 & n7557 ) | ( ~n7257 & n7558 ) | ( n7557 & n7558 ) ;
  assign n7561 = ( n7257 & ~n7559 ) | ( n7257 & n7560 ) | ( ~n7559 & n7560 ) ;
  assign n7562 = ( ~n258 & n7556 ) | ( ~n258 & n7561 ) | ( n7556 & n7561 ) ;
  assign n7563 = ( n258 & ~n7258 ) | ( n258 & n7296 ) | ( ~n7258 & n7296 ) ;
  assign n7564 = n258 & ~n7258 ;
  assign n7565 = ( n7263 & n7563 ) | ( n7263 & n7564 ) | ( n7563 & n7564 ) ;
  assign n7566 = ( ~n7263 & n7563 ) | ( ~n7263 & n7564 ) | ( n7563 & n7564 ) ;
  assign n7567 = ( n7263 & ~n7565 ) | ( n7263 & n7566 ) | ( ~n7565 & n7566 ) ;
  assign n7568 = ( ~n225 & n7562 ) | ( ~n225 & n7567 ) | ( n7562 & n7567 ) ;
  assign n7569 = ~n225 & n7264 ;
  assign n7570 = ( ~n225 & n7264 ) | ( ~n225 & n7296 ) | ( n7264 & n7296 ) ;
  assign n7571 = ( ~n7269 & n7569 ) | ( ~n7269 & n7570 ) | ( n7569 & n7570 ) ;
  assign n7572 = ( n7269 & n7569 ) | ( n7269 & n7570 ) | ( n7569 & n7570 ) ;
  assign n7573 = ( n7269 & n7571 ) | ( n7269 & ~n7572 ) | ( n7571 & ~n7572 ) ;
  assign n7574 = ( ~n197 & n7568 ) | ( ~n197 & n7573 ) | ( n7568 & n7573 ) ;
  assign n7575 = ( n197 & ~n7270 ) | ( n197 & n7296 ) | ( ~n7270 & n7296 ) ;
  assign n7576 = n197 & ~n7270 ;
  assign n7577 = ( n7275 & n7575 ) | ( n7275 & n7576 ) | ( n7575 & n7576 ) ;
  assign n7578 = ( ~n7275 & n7575 ) | ( ~n7275 & n7576 ) | ( n7575 & n7576 ) ;
  assign n7579 = ( n7275 & ~n7577 ) | ( n7275 & n7578 ) | ( ~n7577 & n7578 ) ;
  assign n7580 = ( ~n170 & n7574 ) | ( ~n170 & n7579 ) | ( n7574 & n7579 ) ;
  assign n7581 = ( n170 & ~n7276 ) | ( n170 & n7296 ) | ( ~n7276 & n7296 ) ;
  assign n7582 = n170 & ~n7276 ;
  assign n7583 = ( n7281 & n7581 ) | ( n7281 & n7582 ) | ( n7581 & n7582 ) ;
  assign n7584 = ( ~n7281 & n7581 ) | ( ~n7281 & n7582 ) | ( n7581 & n7582 ) ;
  assign n7585 = ( n7281 & ~n7583 ) | ( n7281 & n7584 ) | ( ~n7583 & n7584 ) ;
  assign n7586 = ( ~n142 & n7580 ) | ( ~n142 & n7585 ) | ( n7580 & n7585 ) ;
  assign n7587 = ( n142 & ~n7282 ) | ( n142 & n7296 ) | ( ~n7282 & n7296 ) ;
  assign n7588 = n142 & ~n7282 ;
  assign n7589 = ( n7287 & n7587 ) | ( n7287 & n7588 ) | ( n7587 & n7588 ) ;
  assign n7590 = ( ~n7287 & n7587 ) | ( ~n7287 & n7588 ) | ( n7587 & n7588 ) ;
  assign n7591 = ( n7287 & ~n7589 ) | ( n7287 & n7590 ) | ( ~n7589 & n7590 ) ;
  assign n7592 = ( ~n132 & n7586 ) | ( ~n132 & n7591 ) | ( n7586 & n7591 ) ;
  assign n7593 = ( ~n131 & n7310 ) | ( ~n131 & n7592 ) | ( n7310 & n7592 ) ;
  assign n7594 = n7305 | n7593 ;
  assign n7595 = ( n132 & ~n7586 ) | ( n132 & n7594 ) | ( ~n7586 & n7594 ) ;
  assign n7596 = n132 & ~n7586 ;
  assign n7597 = ( n7591 & ~n7595 ) | ( n7591 & n7596 ) | ( ~n7595 & n7596 ) ;
  assign n7598 = ( n7591 & n7595 ) | ( n7591 & n7596 ) | ( n7595 & n7596 ) ;
  assign n7599 = ( n7595 & n7597 ) | ( n7595 & ~n7598 ) | ( n7597 & ~n7598 ) ;
  assign n7600 = n7310 & ~n7592 ;
  assign n7601 = ( n7304 & ~n7592 ) | ( n7304 & n7600 ) | ( ~n7592 & n7600 ) ;
  assign n7602 = ( ~n131 & n7310 ) | ( ~n131 & n7601 ) | ( n7310 & n7601 ) ;
  assign n7603 = ~n7600 & n7602 ;
  assign n7604 = ( ~n131 & n7599 ) | ( ~n131 & n7603 ) | ( n7599 & n7603 ) ;
  assign n7605 = n7301 & n7592 ;
  assign n7606 = ( ~n7593 & n7600 ) | ( ~n7593 & n7605 ) | ( n7600 & n7605 ) ;
  assign n7607 = n7604 | n7606 ;
  assign n7608 = ~n7312 & n7594 ;
  assign n7609 = x26 | x27 ;
  assign n7610 = x28 | n7609 ;
  assign n7611 = n7296 & ~n7610 ;
  assign n7612 = ~n7296 & n7610 ;
  assign n7613 = ( x29 & ~n7594 ) | ( x29 & n7612 ) | ( ~n7594 & n7612 ) ;
  assign n7614 = ( n7608 & ~n7611 ) | ( n7608 & n7613 ) | ( ~n7611 & n7613 ) ;
  assign n7615 = n7296 & ~n7594 ;
  assign n7616 = ( x30 & n7608 ) | ( x30 & n7615 ) | ( n7608 & n7615 ) ;
  assign n7617 = ( ~x30 & n7608 ) | ( ~x30 & n7615 ) | ( n7608 & n7615 ) ;
  assign n7618 = ( x30 & ~n7616 ) | ( x30 & n7617 ) | ( ~n7616 & n7617 ) ;
  assign n7619 = ( ~n7006 & n7614 ) | ( ~n7006 & n7618 ) | ( n7614 & n7618 ) ;
  assign n7620 = ~n7006 & n7296 ;
  assign n7621 = ( n7318 & n7594 ) | ( n7318 & n7620 ) | ( n7594 & n7620 ) ;
  assign n7622 = ( ~x31 & n7617 ) | ( ~x31 & n7621 ) | ( n7617 & n7621 ) ;
  assign n7623 = ( x31 & n7617 ) | ( x31 & n7621 ) | ( n7617 & n7621 ) ;
  assign n7624 = ( x31 & n7622 ) | ( x31 & ~n7623 ) | ( n7622 & ~n7623 ) ;
  assign n7625 = ( ~n6723 & n7619 ) | ( ~n6723 & n7624 ) | ( n7619 & n7624 ) ;
  assign n7626 = n6723 & ~n7317 ;
  assign n7627 = ( n6723 & ~n7317 ) | ( n6723 & n7594 ) | ( ~n7317 & n7594 ) ;
  assign n7628 = ( n7321 & n7626 ) | ( n7321 & n7627 ) | ( n7626 & n7627 ) ;
  assign n7629 = ( ~n7321 & n7626 ) | ( ~n7321 & n7627 ) | ( n7626 & n7627 ) ;
  assign n7630 = ( n7321 & ~n7628 ) | ( n7321 & n7629 ) | ( ~n7628 & n7629 ) ;
  assign n7631 = ( ~n6442 & n7625 ) | ( ~n6442 & n7630 ) | ( n7625 & n7630 ) ;
  assign n7632 = ( n6442 & ~n7322 ) | ( n6442 & n7594 ) | ( ~n7322 & n7594 ) ;
  assign n7633 = n6442 & ~n7322 ;
  assign n7634 = ( n7327 & n7632 ) | ( n7327 & n7633 ) | ( n7632 & n7633 ) ;
  assign n7635 = ( ~n7327 & n7632 ) | ( ~n7327 & n7633 ) | ( n7632 & n7633 ) ;
  assign n7636 = ( n7327 & ~n7634 ) | ( n7327 & n7635 ) | ( ~n7634 & n7635 ) ;
  assign n7637 = ( ~n6172 & n7631 ) | ( ~n6172 & n7636 ) | ( n7631 & n7636 ) ;
  assign n7638 = ( n6172 & ~n7328 ) | ( n6172 & n7594 ) | ( ~n7328 & n7594 ) ;
  assign n7639 = n6172 & ~n7328 ;
  assign n7640 = ( n7333 & n7638 ) | ( n7333 & n7639 ) | ( n7638 & n7639 ) ;
  assign n7641 = ( ~n7333 & n7638 ) | ( ~n7333 & n7639 ) | ( n7638 & n7639 ) ;
  assign n7642 = ( n7333 & ~n7640 ) | ( n7333 & n7641 ) | ( ~n7640 & n7641 ) ;
  assign n7643 = ( ~n5905 & n7637 ) | ( ~n5905 & n7642 ) | ( n7637 & n7642 ) ;
  assign n7644 = n5905 & ~n7334 ;
  assign n7645 = ( n5905 & ~n7334 ) | ( n5905 & n7594 ) | ( ~n7334 & n7594 ) ;
  assign n7646 = ( ~n7339 & n7644 ) | ( ~n7339 & n7645 ) | ( n7644 & n7645 ) ;
  assign n7647 = ( n7339 & n7644 ) | ( n7339 & n7645 ) | ( n7644 & n7645 ) ;
  assign n7648 = ( n7339 & n7646 ) | ( n7339 & ~n7647 ) | ( n7646 & ~n7647 ) ;
  assign n7649 = ( ~n5642 & n7643 ) | ( ~n5642 & n7648 ) | ( n7643 & n7648 ) ;
  assign n7650 = ~n5642 & n7340 ;
  assign n7651 = ( ~n5642 & n7340 ) | ( ~n5642 & n7594 ) | ( n7340 & n7594 ) ;
  assign n7652 = ( n7345 & n7650 ) | ( n7345 & n7651 ) | ( n7650 & n7651 ) ;
  assign n7653 = ( ~n7345 & n7650 ) | ( ~n7345 & n7651 ) | ( n7650 & n7651 ) ;
  assign n7654 = ( n7345 & ~n7652 ) | ( n7345 & n7653 ) | ( ~n7652 & n7653 ) ;
  assign n7655 = ( ~n5386 & n7649 ) | ( ~n5386 & n7654 ) | ( n7649 & n7654 ) ;
  assign n7656 = ( n5386 & ~n7346 ) | ( n5386 & n7594 ) | ( ~n7346 & n7594 ) ;
  assign n7657 = n5386 & ~n7346 ;
  assign n7658 = ( n7351 & n7656 ) | ( n7351 & n7657 ) | ( n7656 & n7657 ) ;
  assign n7659 = ( ~n7351 & n7656 ) | ( ~n7351 & n7657 ) | ( n7656 & n7657 ) ;
  assign n7660 = ( n7351 & ~n7658 ) | ( n7351 & n7659 ) | ( ~n7658 & n7659 ) ;
  assign n7661 = ( ~n5139 & n7655 ) | ( ~n5139 & n7660 ) | ( n7655 & n7660 ) ;
  assign n7662 = ( n5139 & ~n7352 ) | ( n5139 & n7594 ) | ( ~n7352 & n7594 ) ;
  assign n7663 = n5139 & ~n7352 ;
  assign n7664 = ( n7357 & n7662 ) | ( n7357 & n7663 ) | ( n7662 & n7663 ) ;
  assign n7665 = ( ~n7357 & n7662 ) | ( ~n7357 & n7663 ) | ( n7662 & n7663 ) ;
  assign n7666 = ( n7357 & ~n7664 ) | ( n7357 & n7665 ) | ( ~n7664 & n7665 ) ;
  assign n7667 = ( ~n4898 & n7661 ) | ( ~n4898 & n7666 ) | ( n7661 & n7666 ) ;
  assign n7668 = ~n4898 & n7358 ;
  assign n7669 = ( ~n4898 & n7358 ) | ( ~n4898 & n7594 ) | ( n7358 & n7594 ) ;
  assign n7670 = ( ~n7363 & n7668 ) | ( ~n7363 & n7669 ) | ( n7668 & n7669 ) ;
  assign n7671 = ( n7363 & n7668 ) | ( n7363 & n7669 ) | ( n7668 & n7669 ) ;
  assign n7672 = ( n7363 & n7670 ) | ( n7363 & ~n7671 ) | ( n7670 & ~n7671 ) ;
  assign n7673 = ( ~n4661 & n7667 ) | ( ~n4661 & n7672 ) | ( n7667 & n7672 ) ;
  assign n7674 = ( n4661 & ~n7364 ) | ( n4661 & n7594 ) | ( ~n7364 & n7594 ) ;
  assign n7675 = n4661 & ~n7364 ;
  assign n7676 = ( n7369 & n7674 ) | ( n7369 & n7675 ) | ( n7674 & n7675 ) ;
  assign n7677 = ( ~n7369 & n7674 ) | ( ~n7369 & n7675 ) | ( n7674 & n7675 ) ;
  assign n7678 = ( n7369 & ~n7676 ) | ( n7369 & n7677 ) | ( ~n7676 & n7677 ) ;
  assign n7679 = ( ~n4432 & n7673 ) | ( ~n4432 & n7678 ) | ( n7673 & n7678 ) ;
  assign n7680 = n4432 & ~n7370 ;
  assign n7681 = ( n4432 & ~n7370 ) | ( n4432 & n7594 ) | ( ~n7370 & n7594 ) ;
  assign n7682 = ( n7375 & n7680 ) | ( n7375 & n7681 ) | ( n7680 & n7681 ) ;
  assign n7683 = ( ~n7375 & n7680 ) | ( ~n7375 & n7681 ) | ( n7680 & n7681 ) ;
  assign n7684 = ( n7375 & ~n7682 ) | ( n7375 & n7683 ) | ( ~n7682 & n7683 ) ;
  assign n7685 = ( ~n4203 & n7679 ) | ( ~n4203 & n7684 ) | ( n7679 & n7684 ) ;
  assign n7686 = ~n4203 & n7376 ;
  assign n7687 = ( ~n4203 & n7376 ) | ( ~n4203 & n7594 ) | ( n7376 & n7594 ) ;
  assign n7688 = ( ~n7381 & n7686 ) | ( ~n7381 & n7687 ) | ( n7686 & n7687 ) ;
  assign n7689 = ( n7381 & n7686 ) | ( n7381 & n7687 ) | ( n7686 & n7687 ) ;
  assign n7690 = ( n7381 & n7688 ) | ( n7381 & ~n7689 ) | ( n7688 & ~n7689 ) ;
  assign n7691 = ( ~n3985 & n7685 ) | ( ~n3985 & n7690 ) | ( n7685 & n7690 ) ;
  assign n7692 = ~n3985 & n7382 ;
  assign n7693 = ( ~n3985 & n7382 ) | ( ~n3985 & n7594 ) | ( n7382 & n7594 ) ;
  assign n7694 = ( ~n7387 & n7692 ) | ( ~n7387 & n7693 ) | ( n7692 & n7693 ) ;
  assign n7695 = ( n7387 & n7692 ) | ( n7387 & n7693 ) | ( n7692 & n7693 ) ;
  assign n7696 = ( n7387 & n7694 ) | ( n7387 & ~n7695 ) | ( n7694 & ~n7695 ) ;
  assign n7697 = ( ~n3772 & n7691 ) | ( ~n3772 & n7696 ) | ( n7691 & n7696 ) ;
  assign n7698 = ( n3772 & ~n7388 ) | ( n3772 & n7594 ) | ( ~n7388 & n7594 ) ;
  assign n7699 = n3772 & ~n7388 ;
  assign n7700 = ( n7393 & n7698 ) | ( n7393 & n7699 ) | ( n7698 & n7699 ) ;
  assign n7701 = ( ~n7393 & n7698 ) | ( ~n7393 & n7699 ) | ( n7698 & n7699 ) ;
  assign n7702 = ( n7393 & ~n7700 ) | ( n7393 & n7701 ) | ( ~n7700 & n7701 ) ;
  assign n7703 = ( ~n3567 & n7697 ) | ( ~n3567 & n7702 ) | ( n7697 & n7702 ) ;
  assign n7704 = ( n3567 & ~n7394 ) | ( n3567 & n7594 ) | ( ~n7394 & n7594 ) ;
  assign n7705 = n3567 & ~n7394 ;
  assign n7706 = ( n7399 & n7704 ) | ( n7399 & n7705 ) | ( n7704 & n7705 ) ;
  assign n7707 = ( ~n7399 & n7704 ) | ( ~n7399 & n7705 ) | ( n7704 & n7705 ) ;
  assign n7708 = ( n7399 & ~n7706 ) | ( n7399 & n7707 ) | ( ~n7706 & n7707 ) ;
  assign n7709 = ( ~n3362 & n7703 ) | ( ~n3362 & n7708 ) | ( n7703 & n7708 ) ;
  assign n7710 = ~n3362 & n7400 ;
  assign n7711 = ( ~n3362 & n7400 ) | ( ~n3362 & n7594 ) | ( n7400 & n7594 ) ;
  assign n7712 = ( n7405 & n7710 ) | ( n7405 & n7711 ) | ( n7710 & n7711 ) ;
  assign n7713 = ( ~n7405 & n7710 ) | ( ~n7405 & n7711 ) | ( n7710 & n7711 ) ;
  assign n7714 = ( n7405 & ~n7712 ) | ( n7405 & n7713 ) | ( ~n7712 & n7713 ) ;
  assign n7715 = ( ~n3169 & n7709 ) | ( ~n3169 & n7714 ) | ( n7709 & n7714 ) ;
  assign n7716 = ~n3169 & n7406 ;
  assign n7717 = ( ~n3169 & n7406 ) | ( ~n3169 & n7594 ) | ( n7406 & n7594 ) ;
  assign n7718 = ( n7411 & n7716 ) | ( n7411 & n7717 ) | ( n7716 & n7717 ) ;
  assign n7719 = ( ~n7411 & n7716 ) | ( ~n7411 & n7717 ) | ( n7716 & n7717 ) ;
  assign n7720 = ( n7411 & ~n7718 ) | ( n7411 & n7719 ) | ( ~n7718 & n7719 ) ;
  assign n7721 = ( ~n2979 & n7715 ) | ( ~n2979 & n7720 ) | ( n7715 & n7720 ) ;
  assign n7722 = ~n2979 & n7412 ;
  assign n7723 = ( ~n2979 & n7412 ) | ( ~n2979 & n7594 ) | ( n7412 & n7594 ) ;
  assign n7724 = ( ~n7417 & n7722 ) | ( ~n7417 & n7723 ) | ( n7722 & n7723 ) ;
  assign n7725 = ( n7417 & n7722 ) | ( n7417 & n7723 ) | ( n7722 & n7723 ) ;
  assign n7726 = ( n7417 & n7724 ) | ( n7417 & ~n7725 ) | ( n7724 & ~n7725 ) ;
  assign n7727 = ( ~n2791 & n7721 ) | ( ~n2791 & n7726 ) | ( n7721 & n7726 ) ;
  assign n7728 = ~n2791 & n7418 ;
  assign n7729 = ( ~n2791 & n7418 ) | ( ~n2791 & n7594 ) | ( n7418 & n7594 ) ;
  assign n7730 = ( ~n7423 & n7728 ) | ( ~n7423 & n7729 ) | ( n7728 & n7729 ) ;
  assign n7731 = ( n7423 & n7728 ) | ( n7423 & n7729 ) | ( n7728 & n7729 ) ;
  assign n7732 = ( n7423 & n7730 ) | ( n7423 & ~n7731 ) | ( n7730 & ~n7731 ) ;
  assign n7733 = ( ~n2615 & n7727 ) | ( ~n2615 & n7732 ) | ( n7727 & n7732 ) ;
  assign n7734 = ( n2615 & ~n7424 ) | ( n2615 & n7594 ) | ( ~n7424 & n7594 ) ;
  assign n7735 = n2615 & ~n7424 ;
  assign n7736 = ( n7429 & n7734 ) | ( n7429 & n7735 ) | ( n7734 & n7735 ) ;
  assign n7737 = ( ~n7429 & n7734 ) | ( ~n7429 & n7735 ) | ( n7734 & n7735 ) ;
  assign n7738 = ( n7429 & ~n7736 ) | ( n7429 & n7737 ) | ( ~n7736 & n7737 ) ;
  assign n7739 = ( ~n2443 & n7733 ) | ( ~n2443 & n7738 ) | ( n7733 & n7738 ) ;
  assign n7740 = ( n2443 & ~n7430 ) | ( n2443 & n7594 ) | ( ~n7430 & n7594 ) ;
  assign n7741 = n2443 & ~n7430 ;
  assign n7742 = ( n7435 & n7740 ) | ( n7435 & n7741 ) | ( n7740 & n7741 ) ;
  assign n7743 = ( ~n7435 & n7740 ) | ( ~n7435 & n7741 ) | ( n7740 & n7741 ) ;
  assign n7744 = ( n7435 & ~n7742 ) | ( n7435 & n7743 ) | ( ~n7742 & n7743 ) ;
  assign n7745 = ( ~n2277 & n7739 ) | ( ~n2277 & n7744 ) | ( n7739 & n7744 ) ;
  assign n7746 = ~n2277 & n7436 ;
  assign n7747 = ( ~n2277 & n7436 ) | ( ~n2277 & n7594 ) | ( n7436 & n7594 ) ;
  assign n7748 = ( ~n7441 & n7746 ) | ( ~n7441 & n7747 ) | ( n7746 & n7747 ) ;
  assign n7749 = ( n7441 & n7746 ) | ( n7441 & n7747 ) | ( n7746 & n7747 ) ;
  assign n7750 = ( n7441 & n7748 ) | ( n7441 & ~n7749 ) | ( n7748 & ~n7749 ) ;
  assign n7751 = ( ~n2111 & n7745 ) | ( ~n2111 & n7750 ) | ( n7745 & n7750 ) ;
  assign n7752 = ( n2111 & ~n7442 ) | ( n2111 & n7594 ) | ( ~n7442 & n7594 ) ;
  assign n7753 = n2111 & ~n7442 ;
  assign n7754 = ( n7447 & n7752 ) | ( n7447 & n7753 ) | ( n7752 & n7753 ) ;
  assign n7755 = ( ~n7447 & n7752 ) | ( ~n7447 & n7753 ) | ( n7752 & n7753 ) ;
  assign n7756 = ( n7447 & ~n7754 ) | ( n7447 & n7755 ) | ( ~n7754 & n7755 ) ;
  assign n7757 = ( ~n1949 & n7751 ) | ( ~n1949 & n7756 ) | ( n7751 & n7756 ) ;
  assign n7758 = ~n1949 & n7448 ;
  assign n7759 = ( ~n1949 & n7448 ) | ( ~n1949 & n7594 ) | ( n7448 & n7594 ) ;
  assign n7760 = ( ~n7453 & n7758 ) | ( ~n7453 & n7759 ) | ( n7758 & n7759 ) ;
  assign n7761 = ( n7453 & n7758 ) | ( n7453 & n7759 ) | ( n7758 & n7759 ) ;
  assign n7762 = ( n7453 & n7760 ) | ( n7453 & ~n7761 ) | ( n7760 & ~n7761 ) ;
  assign n7763 = ( ~n1802 & n7757 ) | ( ~n1802 & n7762 ) | ( n7757 & n7762 ) ;
  assign n7764 = n1802 & ~n7454 ;
  assign n7765 = ( n1802 & ~n7454 ) | ( n1802 & n7594 ) | ( ~n7454 & n7594 ) ;
  assign n7766 = ( n7459 & n7764 ) | ( n7459 & n7765 ) | ( n7764 & n7765 ) ;
  assign n7767 = ( ~n7459 & n7764 ) | ( ~n7459 & n7765 ) | ( n7764 & n7765 ) ;
  assign n7768 = ( n7459 & ~n7766 ) | ( n7459 & n7767 ) | ( ~n7766 & n7767 ) ;
  assign n7769 = ( ~n1661 & n7763 ) | ( ~n1661 & n7768 ) | ( n7763 & n7768 ) ;
  assign n7770 = ~n1661 & n7460 ;
  assign n7771 = ( ~n1661 & n7460 ) | ( ~n1661 & n7594 ) | ( n7460 & n7594 ) ;
  assign n7772 = ( ~n7465 & n7770 ) | ( ~n7465 & n7771 ) | ( n7770 & n7771 ) ;
  assign n7773 = ( n7465 & n7770 ) | ( n7465 & n7771 ) | ( n7770 & n7771 ) ;
  assign n7774 = ( n7465 & n7772 ) | ( n7465 & ~n7773 ) | ( n7772 & ~n7773 ) ;
  assign n7775 = ( ~n1523 & n7769 ) | ( ~n1523 & n7774 ) | ( n7769 & n7774 ) ;
  assign n7776 = n1523 & ~n7466 ;
  assign n7777 = ( n1523 & ~n7466 ) | ( n1523 & n7594 ) | ( ~n7466 & n7594 ) ;
  assign n7778 = ( n7471 & n7776 ) | ( n7471 & n7777 ) | ( n7776 & n7777 ) ;
  assign n7779 = ( ~n7471 & n7776 ) | ( ~n7471 & n7777 ) | ( n7776 & n7777 ) ;
  assign n7780 = ( n7471 & ~n7778 ) | ( n7471 & n7779 ) | ( ~n7778 & n7779 ) ;
  assign n7781 = ( ~n1393 & n7775 ) | ( ~n1393 & n7780 ) | ( n7775 & n7780 ) ;
  assign n7782 = ( n1393 & ~n7472 ) | ( n1393 & n7594 ) | ( ~n7472 & n7594 ) ;
  assign n7783 = n1393 & ~n7472 ;
  assign n7784 = ( n7477 & n7782 ) | ( n7477 & n7783 ) | ( n7782 & n7783 ) ;
  assign n7785 = ( ~n7477 & n7782 ) | ( ~n7477 & n7783 ) | ( n7782 & n7783 ) ;
  assign n7786 = ( n7477 & ~n7784 ) | ( n7477 & n7785 ) | ( ~n7784 & n7785 ) ;
  assign n7787 = ( ~n1266 & n7781 ) | ( ~n1266 & n7786 ) | ( n7781 & n7786 ) ;
  assign n7788 = ( n1266 & ~n7478 ) | ( n1266 & n7594 ) | ( ~n7478 & n7594 ) ;
  assign n7789 = n1266 & ~n7478 ;
  assign n7790 = ( n7483 & n7788 ) | ( n7483 & n7789 ) | ( n7788 & n7789 ) ;
  assign n7791 = ( ~n7483 & n7788 ) | ( ~n7483 & n7789 ) | ( n7788 & n7789 ) ;
  assign n7792 = ( n7483 & ~n7790 ) | ( n7483 & n7791 ) | ( ~n7790 & n7791 ) ;
  assign n7793 = ( ~n1150 & n7787 ) | ( ~n1150 & n7792 ) | ( n7787 & n7792 ) ;
  assign n7794 = ( n1150 & ~n7484 ) | ( n1150 & n7594 ) | ( ~n7484 & n7594 ) ;
  assign n7795 = n1150 & ~n7484 ;
  assign n7796 = ( n7489 & n7794 ) | ( n7489 & n7795 ) | ( n7794 & n7795 ) ;
  assign n7797 = ( ~n7489 & n7794 ) | ( ~n7489 & n7795 ) | ( n7794 & n7795 ) ;
  assign n7798 = ( n7489 & ~n7796 ) | ( n7489 & n7797 ) | ( ~n7796 & n7797 ) ;
  assign n7799 = ( ~n1038 & n7793 ) | ( ~n1038 & n7798 ) | ( n7793 & n7798 ) ;
  assign n7800 = ~n1038 & n7490 ;
  assign n7801 = ( ~n1038 & n7490 ) | ( ~n1038 & n7594 ) | ( n7490 & n7594 ) ;
  assign n7802 = ( ~n7495 & n7800 ) | ( ~n7495 & n7801 ) | ( n7800 & n7801 ) ;
  assign n7803 = ( n7495 & n7800 ) | ( n7495 & n7801 ) | ( n7800 & n7801 ) ;
  assign n7804 = ( n7495 & n7802 ) | ( n7495 & ~n7803 ) | ( n7802 & ~n7803 ) ;
  assign n7805 = ( ~n933 & n7799 ) | ( ~n933 & n7804 ) | ( n7799 & n7804 ) ;
  assign n7806 = ( n933 & ~n7496 ) | ( n933 & n7594 ) | ( ~n7496 & n7594 ) ;
  assign n7807 = n933 & ~n7496 ;
  assign n7808 = ( n7501 & n7806 ) | ( n7501 & n7807 ) | ( n7806 & n7807 ) ;
  assign n7809 = ( ~n7501 & n7806 ) | ( ~n7501 & n7807 ) | ( n7806 & n7807 ) ;
  assign n7810 = ( n7501 & ~n7808 ) | ( n7501 & n7809 ) | ( ~n7808 & n7809 ) ;
  assign n7811 = ( ~n839 & n7805 ) | ( ~n839 & n7810 ) | ( n7805 & n7810 ) ;
  assign n7812 = ~n839 & n7502 ;
  assign n7813 = ( ~n839 & n7502 ) | ( ~n839 & n7594 ) | ( n7502 & n7594 ) ;
  assign n7814 = ( ~n7507 & n7812 ) | ( ~n7507 & n7813 ) | ( n7812 & n7813 ) ;
  assign n7815 = ( n7507 & n7812 ) | ( n7507 & n7813 ) | ( n7812 & n7813 ) ;
  assign n7816 = ( n7507 & n7814 ) | ( n7507 & ~n7815 ) | ( n7814 & ~n7815 ) ;
  assign n7817 = ( ~n746 & n7811 ) | ( ~n746 & n7816 ) | ( n7811 & n7816 ) ;
  assign n7818 = ~n746 & n7508 ;
  assign n7819 = ( ~n746 & n7508 ) | ( ~n746 & n7594 ) | ( n7508 & n7594 ) ;
  assign n7820 = ( ~n7513 & n7818 ) | ( ~n7513 & n7819 ) | ( n7818 & n7819 ) ;
  assign n7821 = ( n7513 & n7818 ) | ( n7513 & n7819 ) | ( n7818 & n7819 ) ;
  assign n7822 = ( n7513 & n7820 ) | ( n7513 & ~n7821 ) | ( n7820 & ~n7821 ) ;
  assign n7823 = ( ~n664 & n7817 ) | ( ~n664 & n7822 ) | ( n7817 & n7822 ) ;
  assign n7824 = ( n664 & ~n7514 ) | ( n664 & n7594 ) | ( ~n7514 & n7594 ) ;
  assign n7825 = n664 & ~n7514 ;
  assign n7826 = ( n7519 & n7824 ) | ( n7519 & n7825 ) | ( n7824 & n7825 ) ;
  assign n7827 = ( ~n7519 & n7824 ) | ( ~n7519 & n7825 ) | ( n7824 & n7825 ) ;
  assign n7828 = ( n7519 & ~n7826 ) | ( n7519 & n7827 ) | ( ~n7826 & n7827 ) ;
  assign n7829 = ( ~n588 & n7823 ) | ( ~n588 & n7828 ) | ( n7823 & n7828 ) ;
  assign n7830 = ( n588 & ~n7520 ) | ( n588 & n7594 ) | ( ~n7520 & n7594 ) ;
  assign n7831 = n588 & ~n7520 ;
  assign n7832 = ( n7525 & n7830 ) | ( n7525 & n7831 ) | ( n7830 & n7831 ) ;
  assign n7833 = ( ~n7525 & n7830 ) | ( ~n7525 & n7831 ) | ( n7830 & n7831 ) ;
  assign n7834 = ( n7525 & ~n7832 ) | ( n7525 & n7833 ) | ( ~n7832 & n7833 ) ;
  assign n7835 = ( ~n518 & n7829 ) | ( ~n518 & n7834 ) | ( n7829 & n7834 ) ;
  assign n7836 = n518 & ~n7526 ;
  assign n7837 = ( n518 & ~n7526 ) | ( n518 & n7594 ) | ( ~n7526 & n7594 ) ;
  assign n7838 = ( n7531 & n7836 ) | ( n7531 & n7837 ) | ( n7836 & n7837 ) ;
  assign n7839 = ( ~n7531 & n7836 ) | ( ~n7531 & n7837 ) | ( n7836 & n7837 ) ;
  assign n7840 = ( n7531 & ~n7838 ) | ( n7531 & n7839 ) | ( ~n7838 & n7839 ) ;
  assign n7841 = ( ~n454 & n7835 ) | ( ~n454 & n7840 ) | ( n7835 & n7840 ) ;
  assign n7842 = ( n454 & ~n7532 ) | ( n454 & n7594 ) | ( ~n7532 & n7594 ) ;
  assign n7843 = n454 & ~n7532 ;
  assign n7844 = ( n7537 & n7842 ) | ( n7537 & n7843 ) | ( n7842 & n7843 ) ;
  assign n7845 = ( ~n7537 & n7842 ) | ( ~n7537 & n7843 ) | ( n7842 & n7843 ) ;
  assign n7846 = ( n7537 & ~n7844 ) | ( n7537 & n7845 ) | ( ~n7844 & n7845 ) ;
  assign n7847 = ( ~n396 & n7841 ) | ( ~n396 & n7846 ) | ( n7841 & n7846 ) ;
  assign n7848 = ( n396 & ~n7538 ) | ( n396 & n7594 ) | ( ~n7538 & n7594 ) ;
  assign n7849 = n396 & ~n7538 ;
  assign n7850 = ( n7543 & n7848 ) | ( n7543 & n7849 ) | ( n7848 & n7849 ) ;
  assign n7851 = ( ~n7543 & n7848 ) | ( ~n7543 & n7849 ) | ( n7848 & n7849 ) ;
  assign n7852 = ( n7543 & ~n7850 ) | ( n7543 & n7851 ) | ( ~n7850 & n7851 ) ;
  assign n7853 = ( ~n344 & n7847 ) | ( ~n344 & n7852 ) | ( n7847 & n7852 ) ;
  assign n7854 = ( n344 & ~n7544 ) | ( n344 & n7594 ) | ( ~n7544 & n7594 ) ;
  assign n7855 = n344 & ~n7544 ;
  assign n7856 = ( n7549 & n7854 ) | ( n7549 & n7855 ) | ( n7854 & n7855 ) ;
  assign n7857 = ( ~n7549 & n7854 ) | ( ~n7549 & n7855 ) | ( n7854 & n7855 ) ;
  assign n7858 = ( n7549 & ~n7856 ) | ( n7549 & n7857 ) | ( ~n7856 & n7857 ) ;
  assign n7859 = ( ~n298 & n7853 ) | ( ~n298 & n7858 ) | ( n7853 & n7858 ) ;
  assign n7860 = ~n298 & n7550 ;
  assign n7861 = ( ~n298 & n7550 ) | ( ~n298 & n7594 ) | ( n7550 & n7594 ) ;
  assign n7862 = ( ~n7555 & n7860 ) | ( ~n7555 & n7861 ) | ( n7860 & n7861 ) ;
  assign n7863 = ( n7555 & n7860 ) | ( n7555 & n7861 ) | ( n7860 & n7861 ) ;
  assign n7864 = ( n7555 & n7862 ) | ( n7555 & ~n7863 ) | ( n7862 & ~n7863 ) ;
  assign n7865 = ( ~n258 & n7859 ) | ( ~n258 & n7864 ) | ( n7859 & n7864 ) ;
  assign n7866 = ~n258 & n7556 ;
  assign n7867 = ( ~n258 & n7556 ) | ( ~n258 & n7594 ) | ( n7556 & n7594 ) ;
  assign n7868 = ( n7561 & n7866 ) | ( n7561 & n7867 ) | ( n7866 & n7867 ) ;
  assign n7869 = ( ~n7561 & n7866 ) | ( ~n7561 & n7867 ) | ( n7866 & n7867 ) ;
  assign n7870 = ( n7561 & ~n7868 ) | ( n7561 & n7869 ) | ( ~n7868 & n7869 ) ;
  assign n7871 = ( ~n225 & n7865 ) | ( ~n225 & n7870 ) | ( n7865 & n7870 ) ;
  assign n7872 = ( n225 & ~n7562 ) | ( n225 & n7594 ) | ( ~n7562 & n7594 ) ;
  assign n7873 = n225 & ~n7562 ;
  assign n7874 = ( n7567 & n7872 ) | ( n7567 & n7873 ) | ( n7872 & n7873 ) ;
  assign n7875 = ( ~n7567 & n7872 ) | ( ~n7567 & n7873 ) | ( n7872 & n7873 ) ;
  assign n7876 = ( n7567 & ~n7874 ) | ( n7567 & n7875 ) | ( ~n7874 & n7875 ) ;
  assign n7877 = ( ~n197 & n7871 ) | ( ~n197 & n7876 ) | ( n7871 & n7876 ) ;
  assign n7878 = ~n197 & n7568 ;
  assign n7879 = ( ~n197 & n7568 ) | ( ~n197 & n7594 ) | ( n7568 & n7594 ) ;
  assign n7880 = ( n7573 & n7878 ) | ( n7573 & n7879 ) | ( n7878 & n7879 ) ;
  assign n7881 = ( ~n7573 & n7878 ) | ( ~n7573 & n7879 ) | ( n7878 & n7879 ) ;
  assign n7882 = ( n7573 & ~n7880 ) | ( n7573 & n7881 ) | ( ~n7880 & n7881 ) ;
  assign n7883 = ( ~n170 & n7877 ) | ( ~n170 & n7882 ) | ( n7877 & n7882 ) ;
  assign n7884 = ~n170 & n7574 ;
  assign n7885 = ( ~n170 & n7574 ) | ( ~n170 & n7594 ) | ( n7574 & n7594 ) ;
  assign n7886 = ( n7579 & n7884 ) | ( n7579 & n7885 ) | ( n7884 & n7885 ) ;
  assign n7887 = ( ~n7579 & n7884 ) | ( ~n7579 & n7885 ) | ( n7884 & n7885 ) ;
  assign n7888 = ( n7579 & ~n7886 ) | ( n7579 & n7887 ) | ( ~n7886 & n7887 ) ;
  assign n7889 = ( ~n142 & n7883 ) | ( ~n142 & n7888 ) | ( n7883 & n7888 ) ;
  assign n7890 = ~n142 & n7580 ;
  assign n7891 = ( ~n142 & n7580 ) | ( ~n142 & n7594 ) | ( n7580 & n7594 ) ;
  assign n7892 = ( n7585 & n7890 ) | ( n7585 & n7891 ) | ( n7890 & n7891 ) ;
  assign n7893 = ( ~n7585 & n7890 ) | ( ~n7585 & n7891 ) | ( n7890 & n7891 ) ;
  assign n7894 = ( n7585 & ~n7892 ) | ( n7585 & n7893 ) | ( ~n7892 & n7893 ) ;
  assign n7895 = ( ~n132 & n7889 ) | ( ~n132 & n7894 ) | ( n7889 & n7894 ) ;
  assign n7896 = ( ~n131 & n7599 ) | ( ~n131 & n7895 ) | ( n7599 & n7895 ) ;
  assign n7897 = n7607 | n7896 ;
  assign n7898 = ( n132 & ~n7889 ) | ( n132 & n7897 ) | ( ~n7889 & n7897 ) ;
  assign n7899 = n132 & ~n7889 ;
  assign n7900 = ( n7894 & ~n7898 ) | ( n7894 & n7899 ) | ( ~n7898 & n7899 ) ;
  assign n7901 = ( n7894 & n7898 ) | ( n7894 & n7899 ) | ( n7898 & n7899 ) ;
  assign n7902 = ( n7898 & n7900 ) | ( n7898 & ~n7901 ) | ( n7900 & ~n7901 ) ;
  assign n7903 = ~n7609 & n7897 ;
  assign n7904 = x24 | x25 ;
  assign n7905 = x26 | n7904 ;
  assign n7906 = n7594 & ~n7905 ;
  assign n7907 = ~n7594 & n7905 ;
  assign n7908 = ( x27 & ~n7897 ) | ( x27 & n7907 ) | ( ~n7897 & n7907 ) ;
  assign n7909 = ( n7903 & ~n7906 ) | ( n7903 & n7908 ) | ( ~n7906 & n7908 ) ;
  assign n7910 = n7594 & ~n7897 ;
  assign n7911 = ( x28 & n7903 ) | ( x28 & n7910 ) | ( n7903 & n7910 ) ;
  assign n7912 = ( ~x28 & n7903 ) | ( ~x28 & n7910 ) | ( n7903 & n7910 ) ;
  assign n7913 = ( x28 & ~n7911 ) | ( x28 & n7912 ) | ( ~n7911 & n7912 ) ;
  assign n7914 = ( ~n7296 & n7909 ) | ( ~n7296 & n7913 ) | ( n7909 & n7913 ) ;
  assign n7915 = ~n7296 & n7594 ;
  assign n7916 = ( n7615 & n7897 ) | ( n7615 & n7915 ) | ( n7897 & n7915 ) ;
  assign n7917 = ( ~x29 & n7912 ) | ( ~x29 & n7916 ) | ( n7912 & n7916 ) ;
  assign n7918 = ( x29 & n7912 ) | ( x29 & n7916 ) | ( n7912 & n7916 ) ;
  assign n7919 = ( x29 & n7917 ) | ( x29 & ~n7918 ) | ( n7917 & ~n7918 ) ;
  assign n7920 = ( ~n7006 & n7914 ) | ( ~n7006 & n7919 ) | ( n7914 & n7919 ) ;
  assign n7921 = ( n7006 & ~n7614 ) | ( n7006 & n7897 ) | ( ~n7614 & n7897 ) ;
  assign n7922 = n7006 & ~n7614 ;
  assign n7923 = ( n7618 & n7921 ) | ( n7618 & n7922 ) | ( n7921 & n7922 ) ;
  assign n7924 = ( ~n7618 & n7921 ) | ( ~n7618 & n7922 ) | ( n7921 & n7922 ) ;
  assign n7925 = ( n7618 & ~n7923 ) | ( n7618 & n7924 ) | ( ~n7923 & n7924 ) ;
  assign n7926 = ( ~n6723 & n7920 ) | ( ~n6723 & n7925 ) | ( n7920 & n7925 ) ;
  assign n7927 = n6723 & ~n7619 ;
  assign n7928 = ( n6723 & ~n7619 ) | ( n6723 & n7897 ) | ( ~n7619 & n7897 ) ;
  assign n7929 = ( n7624 & n7927 ) | ( n7624 & n7928 ) | ( n7927 & n7928 ) ;
  assign n7930 = ( ~n7624 & n7927 ) | ( ~n7624 & n7928 ) | ( n7927 & n7928 ) ;
  assign n7931 = ( n7624 & ~n7929 ) | ( n7624 & n7930 ) | ( ~n7929 & n7930 ) ;
  assign n7932 = ( ~n6442 & n7926 ) | ( ~n6442 & n7931 ) | ( n7926 & n7931 ) ;
  assign n7933 = n6442 & ~n7625 ;
  assign n7934 = ( n6442 & ~n7625 ) | ( n6442 & n7897 ) | ( ~n7625 & n7897 ) ;
  assign n7935 = ( ~n7630 & n7933 ) | ( ~n7630 & n7934 ) | ( n7933 & n7934 ) ;
  assign n7936 = ( n7630 & n7933 ) | ( n7630 & n7934 ) | ( n7933 & n7934 ) ;
  assign n7937 = ( n7630 & n7935 ) | ( n7630 & ~n7936 ) | ( n7935 & ~n7936 ) ;
  assign n7938 = ( ~n6172 & n7932 ) | ( ~n6172 & n7937 ) | ( n7932 & n7937 ) ;
  assign n7939 = ( n6172 & ~n7631 ) | ( n6172 & n7897 ) | ( ~n7631 & n7897 ) ;
  assign n7940 = n6172 & ~n7631 ;
  assign n7941 = ( n7636 & n7939 ) | ( n7636 & n7940 ) | ( n7939 & n7940 ) ;
  assign n7942 = ( ~n7636 & n7939 ) | ( ~n7636 & n7940 ) | ( n7939 & n7940 ) ;
  assign n7943 = ( n7636 & ~n7941 ) | ( n7636 & n7942 ) | ( ~n7941 & n7942 ) ;
  assign n7944 = ( ~n5905 & n7938 ) | ( ~n5905 & n7943 ) | ( n7938 & n7943 ) ;
  assign n7945 = ~n5905 & n7637 ;
  assign n7946 = ( ~n5905 & n7637 ) | ( ~n5905 & n7897 ) | ( n7637 & n7897 ) ;
  assign n7947 = ( ~n7642 & n7945 ) | ( ~n7642 & n7946 ) | ( n7945 & n7946 ) ;
  assign n7948 = ( n7642 & n7945 ) | ( n7642 & n7946 ) | ( n7945 & n7946 ) ;
  assign n7949 = ( n7642 & n7947 ) | ( n7642 & ~n7948 ) | ( n7947 & ~n7948 ) ;
  assign n7950 = ( ~n5642 & n7944 ) | ( ~n5642 & n7949 ) | ( n7944 & n7949 ) ;
  assign n7951 = ~n5642 & n7643 ;
  assign n7952 = ( ~n5642 & n7643 ) | ( ~n5642 & n7897 ) | ( n7643 & n7897 ) ;
  assign n7953 = ( n7648 & n7951 ) | ( n7648 & n7952 ) | ( n7951 & n7952 ) ;
  assign n7954 = ( ~n7648 & n7951 ) | ( ~n7648 & n7952 ) | ( n7951 & n7952 ) ;
  assign n7955 = ( n7648 & ~n7953 ) | ( n7648 & n7954 ) | ( ~n7953 & n7954 ) ;
  assign n7956 = ( ~n5386 & n7950 ) | ( ~n5386 & n7955 ) | ( n7950 & n7955 ) ;
  assign n7957 = ~n5386 & n7649 ;
  assign n7958 = ( ~n5386 & n7649 ) | ( ~n5386 & n7897 ) | ( n7649 & n7897 ) ;
  assign n7959 = ( ~n7654 & n7957 ) | ( ~n7654 & n7958 ) | ( n7957 & n7958 ) ;
  assign n7960 = ( n7654 & n7957 ) | ( n7654 & n7958 ) | ( n7957 & n7958 ) ;
  assign n7961 = ( n7654 & n7959 ) | ( n7654 & ~n7960 ) | ( n7959 & ~n7960 ) ;
  assign n7962 = ( ~n5139 & n7956 ) | ( ~n5139 & n7961 ) | ( n7956 & n7961 ) ;
  assign n7963 = ( n5139 & ~n7655 ) | ( n5139 & n7897 ) | ( ~n7655 & n7897 ) ;
  assign n7964 = n5139 & ~n7655 ;
  assign n7965 = ( n7660 & n7963 ) | ( n7660 & n7964 ) | ( n7963 & n7964 ) ;
  assign n7966 = ( ~n7660 & n7963 ) | ( ~n7660 & n7964 ) | ( n7963 & n7964 ) ;
  assign n7967 = ( n7660 & ~n7965 ) | ( n7660 & n7966 ) | ( ~n7965 & n7966 ) ;
  assign n7968 = ( ~n4898 & n7962 ) | ( ~n4898 & n7967 ) | ( n7962 & n7967 ) ;
  assign n7969 = ( n4898 & ~n7661 ) | ( n4898 & n7897 ) | ( ~n7661 & n7897 ) ;
  assign n7970 = n4898 & ~n7661 ;
  assign n7971 = ( n7666 & n7969 ) | ( n7666 & n7970 ) | ( n7969 & n7970 ) ;
  assign n7972 = ( ~n7666 & n7969 ) | ( ~n7666 & n7970 ) | ( n7969 & n7970 ) ;
  assign n7973 = ( n7666 & ~n7971 ) | ( n7666 & n7972 ) | ( ~n7971 & n7972 ) ;
  assign n7974 = ( ~n4661 & n7968 ) | ( ~n4661 & n7973 ) | ( n7968 & n7973 ) ;
  assign n7975 = ( n4661 & ~n7667 ) | ( n4661 & n7897 ) | ( ~n7667 & n7897 ) ;
  assign n7976 = n4661 & ~n7667 ;
  assign n7977 = ( n7672 & n7975 ) | ( n7672 & n7976 ) | ( n7975 & n7976 ) ;
  assign n7978 = ( ~n7672 & n7975 ) | ( ~n7672 & n7976 ) | ( n7975 & n7976 ) ;
  assign n7979 = ( n7672 & ~n7977 ) | ( n7672 & n7978 ) | ( ~n7977 & n7978 ) ;
  assign n7980 = ( ~n4432 & n7974 ) | ( ~n4432 & n7979 ) | ( n7974 & n7979 ) ;
  assign n7981 = ~n4432 & n7673 ;
  assign n7982 = ( ~n4432 & n7673 ) | ( ~n4432 & n7897 ) | ( n7673 & n7897 ) ;
  assign n7983 = ( ~n7678 & n7981 ) | ( ~n7678 & n7982 ) | ( n7981 & n7982 ) ;
  assign n7984 = ( n7678 & n7981 ) | ( n7678 & n7982 ) | ( n7981 & n7982 ) ;
  assign n7985 = ( n7678 & n7983 ) | ( n7678 & ~n7984 ) | ( n7983 & ~n7984 ) ;
  assign n7986 = ( ~n4203 & n7980 ) | ( ~n4203 & n7985 ) | ( n7980 & n7985 ) ;
  assign n7987 = ( n4203 & ~n7679 ) | ( n4203 & n7897 ) | ( ~n7679 & n7897 ) ;
  assign n7988 = n4203 & ~n7679 ;
  assign n7989 = ( n7684 & n7987 ) | ( n7684 & n7988 ) | ( n7987 & n7988 ) ;
  assign n7990 = ( ~n7684 & n7987 ) | ( ~n7684 & n7988 ) | ( n7987 & n7988 ) ;
  assign n7991 = ( n7684 & ~n7989 ) | ( n7684 & n7990 ) | ( ~n7989 & n7990 ) ;
  assign n7992 = ( ~n3985 & n7986 ) | ( ~n3985 & n7991 ) | ( n7986 & n7991 ) ;
  assign n7993 = ( n3985 & ~n7685 ) | ( n3985 & n7897 ) | ( ~n7685 & n7897 ) ;
  assign n7994 = n3985 & ~n7685 ;
  assign n7995 = ( n7690 & n7993 ) | ( n7690 & n7994 ) | ( n7993 & n7994 ) ;
  assign n7996 = ( ~n7690 & n7993 ) | ( ~n7690 & n7994 ) | ( n7993 & n7994 ) ;
  assign n7997 = ( n7690 & ~n7995 ) | ( n7690 & n7996 ) | ( ~n7995 & n7996 ) ;
  assign n7998 = ( ~n3772 & n7992 ) | ( ~n3772 & n7997 ) | ( n7992 & n7997 ) ;
  assign n7999 = ( n3772 & ~n7691 ) | ( n3772 & n7897 ) | ( ~n7691 & n7897 ) ;
  assign n8000 = n3772 & ~n7691 ;
  assign n8001 = ( n7696 & n7999 ) | ( n7696 & n8000 ) | ( n7999 & n8000 ) ;
  assign n8002 = ( ~n7696 & n7999 ) | ( ~n7696 & n8000 ) | ( n7999 & n8000 ) ;
  assign n8003 = ( n7696 & ~n8001 ) | ( n7696 & n8002 ) | ( ~n8001 & n8002 ) ;
  assign n8004 = ( ~n3567 & n7998 ) | ( ~n3567 & n8003 ) | ( n7998 & n8003 ) ;
  assign n8005 = ( n3567 & ~n7697 ) | ( n3567 & n7897 ) | ( ~n7697 & n7897 ) ;
  assign n8006 = n3567 & ~n7697 ;
  assign n8007 = ( ~n7702 & n8005 ) | ( ~n7702 & n8006 ) | ( n8005 & n8006 ) ;
  assign n8008 = ( n7702 & n8005 ) | ( n7702 & n8006 ) | ( n8005 & n8006 ) ;
  assign n8009 = ( n7702 & n8007 ) | ( n7702 & ~n8008 ) | ( n8007 & ~n8008 ) ;
  assign n8010 = ( ~n3362 & n8004 ) | ( ~n3362 & n8009 ) | ( n8004 & n8009 ) ;
  assign n8011 = ~n3362 & n7703 ;
  assign n8012 = ( ~n3362 & n7703 ) | ( ~n3362 & n7897 ) | ( n7703 & n7897 ) ;
  assign n8013 = ( ~n7708 & n8011 ) | ( ~n7708 & n8012 ) | ( n8011 & n8012 ) ;
  assign n8014 = ( n7708 & n8011 ) | ( n7708 & n8012 ) | ( n8011 & n8012 ) ;
  assign n8015 = ( n7708 & n8013 ) | ( n7708 & ~n8014 ) | ( n8013 & ~n8014 ) ;
  assign n8016 = ( ~n3169 & n8010 ) | ( ~n3169 & n8015 ) | ( n8010 & n8015 ) ;
  assign n8017 = ~n3169 & n7709 ;
  assign n8018 = ( ~n3169 & n7709 ) | ( ~n3169 & n7897 ) | ( n7709 & n7897 ) ;
  assign n8019 = ( n7714 & n8017 ) | ( n7714 & n8018 ) | ( n8017 & n8018 ) ;
  assign n8020 = ( ~n7714 & n8017 ) | ( ~n7714 & n8018 ) | ( n8017 & n8018 ) ;
  assign n8021 = ( n7714 & ~n8019 ) | ( n7714 & n8020 ) | ( ~n8019 & n8020 ) ;
  assign n8022 = ( ~n2979 & n8016 ) | ( ~n2979 & n8021 ) | ( n8016 & n8021 ) ;
  assign n8023 = ( n2979 & ~n7715 ) | ( n2979 & n7897 ) | ( ~n7715 & n7897 ) ;
  assign n8024 = n2979 & ~n7715 ;
  assign n8025 = ( n7720 & n8023 ) | ( n7720 & n8024 ) | ( n8023 & n8024 ) ;
  assign n8026 = ( ~n7720 & n8023 ) | ( ~n7720 & n8024 ) | ( n8023 & n8024 ) ;
  assign n8027 = ( n7720 & ~n8025 ) | ( n7720 & n8026 ) | ( ~n8025 & n8026 ) ;
  assign n8028 = ( ~n2791 & n8022 ) | ( ~n2791 & n8027 ) | ( n8022 & n8027 ) ;
  assign n8029 = ( n2791 & ~n7721 ) | ( n2791 & n7897 ) | ( ~n7721 & n7897 ) ;
  assign n8030 = n2791 & ~n7721 ;
  assign n8031 = ( n7726 & n8029 ) | ( n7726 & n8030 ) | ( n8029 & n8030 ) ;
  assign n8032 = ( ~n7726 & n8029 ) | ( ~n7726 & n8030 ) | ( n8029 & n8030 ) ;
  assign n8033 = ( n7726 & ~n8031 ) | ( n7726 & n8032 ) | ( ~n8031 & n8032 ) ;
  assign n8034 = ( ~n2615 & n8028 ) | ( ~n2615 & n8033 ) | ( n8028 & n8033 ) ;
  assign n8035 = ( n2615 & ~n7727 ) | ( n2615 & n7897 ) | ( ~n7727 & n7897 ) ;
  assign n8036 = n2615 & ~n7727 ;
  assign n8037 = ( n7732 & n8035 ) | ( n7732 & n8036 ) | ( n8035 & n8036 ) ;
  assign n8038 = ( ~n7732 & n8035 ) | ( ~n7732 & n8036 ) | ( n8035 & n8036 ) ;
  assign n8039 = ( n7732 & ~n8037 ) | ( n7732 & n8038 ) | ( ~n8037 & n8038 ) ;
  assign n8040 = ( ~n2443 & n8034 ) | ( ~n2443 & n8039 ) | ( n8034 & n8039 ) ;
  assign n8041 = ( n2443 & ~n7733 ) | ( n2443 & n7897 ) | ( ~n7733 & n7897 ) ;
  assign n8042 = n2443 & ~n7733 ;
  assign n8043 = ( n7738 & n8041 ) | ( n7738 & n8042 ) | ( n8041 & n8042 ) ;
  assign n8044 = ( ~n7738 & n8041 ) | ( ~n7738 & n8042 ) | ( n8041 & n8042 ) ;
  assign n8045 = ( n7738 & ~n8043 ) | ( n7738 & n8044 ) | ( ~n8043 & n8044 ) ;
  assign n8046 = ( ~n2277 & n8040 ) | ( ~n2277 & n8045 ) | ( n8040 & n8045 ) ;
  assign n8047 = ( n2277 & ~n7739 ) | ( n2277 & n7897 ) | ( ~n7739 & n7897 ) ;
  assign n8048 = n2277 & ~n7739 ;
  assign n8049 = ( n7744 & n8047 ) | ( n7744 & n8048 ) | ( n8047 & n8048 ) ;
  assign n8050 = ( ~n7744 & n8047 ) | ( ~n7744 & n8048 ) | ( n8047 & n8048 ) ;
  assign n8051 = ( n7744 & ~n8049 ) | ( n7744 & n8050 ) | ( ~n8049 & n8050 ) ;
  assign n8052 = ( ~n2111 & n8046 ) | ( ~n2111 & n8051 ) | ( n8046 & n8051 ) ;
  assign n8053 = ( n2111 & ~n7745 ) | ( n2111 & n7897 ) | ( ~n7745 & n7897 ) ;
  assign n8054 = n2111 & ~n7745 ;
  assign n8055 = ( n7750 & n8053 ) | ( n7750 & n8054 ) | ( n8053 & n8054 ) ;
  assign n8056 = ( ~n7750 & n8053 ) | ( ~n7750 & n8054 ) | ( n8053 & n8054 ) ;
  assign n8057 = ( n7750 & ~n8055 ) | ( n7750 & n8056 ) | ( ~n8055 & n8056 ) ;
  assign n8058 = ( ~n1949 & n8052 ) | ( ~n1949 & n8057 ) | ( n8052 & n8057 ) ;
  assign n8059 = ( n1949 & ~n7751 ) | ( n1949 & n7897 ) | ( ~n7751 & n7897 ) ;
  assign n8060 = n1949 & ~n7751 ;
  assign n8061 = ( n7756 & n8059 ) | ( n7756 & n8060 ) | ( n8059 & n8060 ) ;
  assign n8062 = ( ~n7756 & n8059 ) | ( ~n7756 & n8060 ) | ( n8059 & n8060 ) ;
  assign n8063 = ( n7756 & ~n8061 ) | ( n7756 & n8062 ) | ( ~n8061 & n8062 ) ;
  assign n8064 = ( ~n1802 & n8058 ) | ( ~n1802 & n8063 ) | ( n8058 & n8063 ) ;
  assign n8065 = ( n1802 & ~n7757 ) | ( n1802 & n7897 ) | ( ~n7757 & n7897 ) ;
  assign n8066 = n1802 & ~n7757 ;
  assign n8067 = ( n7762 & n8065 ) | ( n7762 & n8066 ) | ( n8065 & n8066 ) ;
  assign n8068 = ( ~n7762 & n8065 ) | ( ~n7762 & n8066 ) | ( n8065 & n8066 ) ;
  assign n8069 = ( n7762 & ~n8067 ) | ( n7762 & n8068 ) | ( ~n8067 & n8068 ) ;
  assign n8070 = ( ~n1661 & n8064 ) | ( ~n1661 & n8069 ) | ( n8064 & n8069 ) ;
  assign n8071 = ~n1661 & n7763 ;
  assign n8072 = ( ~n1661 & n7763 ) | ( ~n1661 & n7897 ) | ( n7763 & n7897 ) ;
  assign n8073 = ( ~n7768 & n8071 ) | ( ~n7768 & n8072 ) | ( n8071 & n8072 ) ;
  assign n8074 = ( n7768 & n8071 ) | ( n7768 & n8072 ) | ( n8071 & n8072 ) ;
  assign n8075 = ( n7768 & n8073 ) | ( n7768 & ~n8074 ) | ( n8073 & ~n8074 ) ;
  assign n8076 = ( ~n1523 & n8070 ) | ( ~n1523 & n8075 ) | ( n8070 & n8075 ) ;
  assign n8077 = n1523 & ~n7769 ;
  assign n8078 = ( n1523 & ~n7769 ) | ( n1523 & n7897 ) | ( ~n7769 & n7897 ) ;
  assign n8079 = ( ~n7774 & n8077 ) | ( ~n7774 & n8078 ) | ( n8077 & n8078 ) ;
  assign n8080 = ( n7774 & n8077 ) | ( n7774 & n8078 ) | ( n8077 & n8078 ) ;
  assign n8081 = ( n7774 & n8079 ) | ( n7774 & ~n8080 ) | ( n8079 & ~n8080 ) ;
  assign n8082 = ( ~n1393 & n8076 ) | ( ~n1393 & n8081 ) | ( n8076 & n8081 ) ;
  assign n8083 = ( n1393 & ~n7775 ) | ( n1393 & n7897 ) | ( ~n7775 & n7897 ) ;
  assign n8084 = n1393 & ~n7775 ;
  assign n8085 = ( n7780 & n8083 ) | ( n7780 & n8084 ) | ( n8083 & n8084 ) ;
  assign n8086 = ( ~n7780 & n8083 ) | ( ~n7780 & n8084 ) | ( n8083 & n8084 ) ;
  assign n8087 = ( n7780 & ~n8085 ) | ( n7780 & n8086 ) | ( ~n8085 & n8086 ) ;
  assign n8088 = ( ~n1266 & n8082 ) | ( ~n1266 & n8087 ) | ( n8082 & n8087 ) ;
  assign n8089 = ~n1266 & n7781 ;
  assign n8090 = ( ~n1266 & n7781 ) | ( ~n1266 & n7897 ) | ( n7781 & n7897 ) ;
  assign n8091 = ( ~n7786 & n8089 ) | ( ~n7786 & n8090 ) | ( n8089 & n8090 ) ;
  assign n8092 = ( n7786 & n8089 ) | ( n7786 & n8090 ) | ( n8089 & n8090 ) ;
  assign n8093 = ( n7786 & n8091 ) | ( n7786 & ~n8092 ) | ( n8091 & ~n8092 ) ;
  assign n8094 = ( ~n1150 & n8088 ) | ( ~n1150 & n8093 ) | ( n8088 & n8093 ) ;
  assign n8095 = n1150 & ~n7787 ;
  assign n8096 = ( n1150 & ~n7787 ) | ( n1150 & n7897 ) | ( ~n7787 & n7897 ) ;
  assign n8097 = ( n7792 & n8095 ) | ( n7792 & n8096 ) | ( n8095 & n8096 ) ;
  assign n8098 = ( ~n7792 & n8095 ) | ( ~n7792 & n8096 ) | ( n8095 & n8096 ) ;
  assign n8099 = ( n7792 & ~n8097 ) | ( n7792 & n8098 ) | ( ~n8097 & n8098 ) ;
  assign n8100 = ( ~n1038 & n8094 ) | ( ~n1038 & n8099 ) | ( n8094 & n8099 ) ;
  assign n8101 = n1038 & ~n7793 ;
  assign n8102 = ( n1038 & ~n7793 ) | ( n1038 & n7897 ) | ( ~n7793 & n7897 ) ;
  assign n8103 = ( n7798 & n8101 ) | ( n7798 & n8102 ) | ( n8101 & n8102 ) ;
  assign n8104 = ( ~n7798 & n8101 ) | ( ~n7798 & n8102 ) | ( n8101 & n8102 ) ;
  assign n8105 = ( n7798 & ~n8103 ) | ( n7798 & n8104 ) | ( ~n8103 & n8104 ) ;
  assign n8106 = ( ~n933 & n8100 ) | ( ~n933 & n8105 ) | ( n8100 & n8105 ) ;
  assign n8107 = n933 & ~n7799 ;
  assign n8108 = ( n933 & ~n7799 ) | ( n933 & n7897 ) | ( ~n7799 & n7897 ) ;
  assign n8109 = ( n7804 & n8107 ) | ( n7804 & n8108 ) | ( n8107 & n8108 ) ;
  assign n8110 = ( ~n7804 & n8107 ) | ( ~n7804 & n8108 ) | ( n8107 & n8108 ) ;
  assign n8111 = ( n7804 & ~n8109 ) | ( n7804 & n8110 ) | ( ~n8109 & n8110 ) ;
  assign n8112 = ( ~n839 & n8106 ) | ( ~n839 & n8111 ) | ( n8106 & n8111 ) ;
  assign n8113 = ~n839 & n7805 ;
  assign n8114 = ( ~n839 & n7805 ) | ( ~n839 & n7897 ) | ( n7805 & n7897 ) ;
  assign n8115 = ( ~n7810 & n8113 ) | ( ~n7810 & n8114 ) | ( n8113 & n8114 ) ;
  assign n8116 = ( n7810 & n8113 ) | ( n7810 & n8114 ) | ( n8113 & n8114 ) ;
  assign n8117 = ( n7810 & n8115 ) | ( n7810 & ~n8116 ) | ( n8115 & ~n8116 ) ;
  assign n8118 = ( ~n746 & n8112 ) | ( ~n746 & n8117 ) | ( n8112 & n8117 ) ;
  assign n8119 = ~n746 & n7811 ;
  assign n8120 = ( ~n746 & n7811 ) | ( ~n746 & n7897 ) | ( n7811 & n7897 ) ;
  assign n8121 = ( ~n7816 & n8119 ) | ( ~n7816 & n8120 ) | ( n8119 & n8120 ) ;
  assign n8122 = ( n7816 & n8119 ) | ( n7816 & n8120 ) | ( n8119 & n8120 ) ;
  assign n8123 = ( n7816 & n8121 ) | ( n7816 & ~n8122 ) | ( n8121 & ~n8122 ) ;
  assign n8124 = ( ~n664 & n8118 ) | ( ~n664 & n8123 ) | ( n8118 & n8123 ) ;
  assign n8125 = ~n664 & n7817 ;
  assign n8126 = ( ~n664 & n7817 ) | ( ~n664 & n7897 ) | ( n7817 & n7897 ) ;
  assign n8127 = ( ~n7822 & n8125 ) | ( ~n7822 & n8126 ) | ( n8125 & n8126 ) ;
  assign n8128 = ( n7822 & n8125 ) | ( n7822 & n8126 ) | ( n8125 & n8126 ) ;
  assign n8129 = ( n7822 & n8127 ) | ( n7822 & ~n8128 ) | ( n8127 & ~n8128 ) ;
  assign n8130 = ( ~n588 & n8124 ) | ( ~n588 & n8129 ) | ( n8124 & n8129 ) ;
  assign n8131 = ( n588 & ~n7823 ) | ( n588 & n7897 ) | ( ~n7823 & n7897 ) ;
  assign n8132 = n588 & ~n7823 ;
  assign n8133 = ( n7828 & n8131 ) | ( n7828 & n8132 ) | ( n8131 & n8132 ) ;
  assign n8134 = ( ~n7828 & n8131 ) | ( ~n7828 & n8132 ) | ( n8131 & n8132 ) ;
  assign n8135 = ( n7828 & ~n8133 ) | ( n7828 & n8134 ) | ( ~n8133 & n8134 ) ;
  assign n8136 = ( ~n518 & n8130 ) | ( ~n518 & n8135 ) | ( n8130 & n8135 ) ;
  assign n8137 = ~n518 & n7829 ;
  assign n8138 = ( ~n518 & n7829 ) | ( ~n518 & n7897 ) | ( n7829 & n7897 ) ;
  assign n8139 = ( ~n7834 & n8137 ) | ( ~n7834 & n8138 ) | ( n8137 & n8138 ) ;
  assign n8140 = ( n7834 & n8137 ) | ( n7834 & n8138 ) | ( n8137 & n8138 ) ;
  assign n8141 = ( n7834 & n8139 ) | ( n7834 & ~n8140 ) | ( n8139 & ~n8140 ) ;
  assign n8142 = ( ~n454 & n8136 ) | ( ~n454 & n8141 ) | ( n8136 & n8141 ) ;
  assign n8143 = ( n454 & ~n7835 ) | ( n454 & n7897 ) | ( ~n7835 & n7897 ) ;
  assign n8144 = n454 & ~n7835 ;
  assign n8145 = ( n7840 & n8143 ) | ( n7840 & n8144 ) | ( n8143 & n8144 ) ;
  assign n8146 = ( ~n7840 & n8143 ) | ( ~n7840 & n8144 ) | ( n8143 & n8144 ) ;
  assign n8147 = ( n7840 & ~n8145 ) | ( n7840 & n8146 ) | ( ~n8145 & n8146 ) ;
  assign n8148 = ( ~n396 & n8142 ) | ( ~n396 & n8147 ) | ( n8142 & n8147 ) ;
  assign n8149 = ~n396 & n7841 ;
  assign n8150 = ( ~n396 & n7841 ) | ( ~n396 & n7897 ) | ( n7841 & n7897 ) ;
  assign n8151 = ( ~n7846 & n8149 ) | ( ~n7846 & n8150 ) | ( n8149 & n8150 ) ;
  assign n8152 = ( n7846 & n8149 ) | ( n7846 & n8150 ) | ( n8149 & n8150 ) ;
  assign n8153 = ( n7846 & n8151 ) | ( n7846 & ~n8152 ) | ( n8151 & ~n8152 ) ;
  assign n8154 = ( ~n344 & n8148 ) | ( ~n344 & n8153 ) | ( n8148 & n8153 ) ;
  assign n8155 = ~n344 & n7847 ;
  assign n8156 = ( ~n344 & n7847 ) | ( ~n344 & n7897 ) | ( n7847 & n7897 ) ;
  assign n8157 = ( ~n7852 & n8155 ) | ( ~n7852 & n8156 ) | ( n8155 & n8156 ) ;
  assign n8158 = ( n7852 & n8155 ) | ( n7852 & n8156 ) | ( n8155 & n8156 ) ;
  assign n8159 = ( n7852 & n8157 ) | ( n7852 & ~n8158 ) | ( n8157 & ~n8158 ) ;
  assign n8160 = ( ~n298 & n8154 ) | ( ~n298 & n8159 ) | ( n8154 & n8159 ) ;
  assign n8161 = ( n298 & ~n7853 ) | ( n298 & n7897 ) | ( ~n7853 & n7897 ) ;
  assign n8162 = n298 & ~n7853 ;
  assign n8163 = ( n7858 & n8161 ) | ( n7858 & n8162 ) | ( n8161 & n8162 ) ;
  assign n8164 = ( ~n7858 & n8161 ) | ( ~n7858 & n8162 ) | ( n8161 & n8162 ) ;
  assign n8165 = ( n7858 & ~n8163 ) | ( n7858 & n8164 ) | ( ~n8163 & n8164 ) ;
  assign n8166 = ( ~n258 & n8160 ) | ( ~n258 & n8165 ) | ( n8160 & n8165 ) ;
  assign n8167 = ( n258 & ~n7859 ) | ( n258 & n7897 ) | ( ~n7859 & n7897 ) ;
  assign n8168 = n258 & ~n7859 ;
  assign n8169 = ( n7864 & n8167 ) | ( n7864 & n8168 ) | ( n8167 & n8168 ) ;
  assign n8170 = ( ~n7864 & n8167 ) | ( ~n7864 & n8168 ) | ( n8167 & n8168 ) ;
  assign n8171 = ( n7864 & ~n8169 ) | ( n7864 & n8170 ) | ( ~n8169 & n8170 ) ;
  assign n8172 = ( ~n225 & n8166 ) | ( ~n225 & n8171 ) | ( n8166 & n8171 ) ;
  assign n8173 = ~n225 & n7865 ;
  assign n8174 = ( ~n225 & n7865 ) | ( ~n225 & n7897 ) | ( n7865 & n7897 ) ;
  assign n8175 = ( n7870 & n8173 ) | ( n7870 & n8174 ) | ( n8173 & n8174 ) ;
  assign n8176 = ( ~n7870 & n8173 ) | ( ~n7870 & n8174 ) | ( n8173 & n8174 ) ;
  assign n8177 = ( n7870 & ~n8175 ) | ( n7870 & n8176 ) | ( ~n8175 & n8176 ) ;
  assign n8178 = ( ~n197 & n8172 ) | ( ~n197 & n8177 ) | ( n8172 & n8177 ) ;
  assign n8179 = n197 & ~n7871 ;
  assign n8180 = ( n197 & ~n7871 ) | ( n197 & n7897 ) | ( ~n7871 & n7897 ) ;
  assign n8181 = ( n7876 & n8179 ) | ( n7876 & n8180 ) | ( n8179 & n8180 ) ;
  assign n8182 = ( ~n7876 & n8179 ) | ( ~n7876 & n8180 ) | ( n8179 & n8180 ) ;
  assign n8183 = ( n7876 & ~n8181 ) | ( n7876 & n8182 ) | ( ~n8181 & n8182 ) ;
  assign n8184 = ( ~n170 & n8178 ) | ( ~n170 & n8183 ) | ( n8178 & n8183 ) ;
  assign n8185 = ( n170 & ~n7877 ) | ( n170 & n7897 ) | ( ~n7877 & n7897 ) ;
  assign n8186 = n170 & ~n7877 ;
  assign n8187 = ( n7882 & n8185 ) | ( n7882 & n8186 ) | ( n8185 & n8186 ) ;
  assign n8188 = ( ~n7882 & n8185 ) | ( ~n7882 & n8186 ) | ( n8185 & n8186 ) ;
  assign n8189 = ( n7882 & ~n8187 ) | ( n7882 & n8188 ) | ( ~n8187 & n8188 ) ;
  assign n8190 = ( ~n142 & n8184 ) | ( ~n142 & n8189 ) | ( n8184 & n8189 ) ;
  assign n8191 = ( n142 & ~n7883 ) | ( n142 & n7897 ) | ( ~n7883 & n7897 ) ;
  assign n8192 = n142 & ~n7883 ;
  assign n8193 = ( n7888 & n8191 ) | ( n7888 & n8192 ) | ( n8191 & n8192 ) ;
  assign n8194 = ( ~n7888 & n8191 ) | ( ~n7888 & n8192 ) | ( n8191 & n8192 ) ;
  assign n8195 = ( n7888 & ~n8193 ) | ( n7888 & n8194 ) | ( ~n8193 & n8194 ) ;
  assign n8196 = ( ~n132 & n8190 ) | ( ~n132 & n8195 ) | ( n8190 & n8195 ) ;
  assign n8197 = ( ~n131 & n7902 ) | ( ~n131 & n8196 ) | ( n7902 & n8196 ) ;
  assign n8198 = ( n7599 & n7606 ) | ( n7599 & n7895 ) | ( n7606 & n7895 ) ;
  assign n8199 = ( n7599 & n7604 ) | ( n7599 & ~n7895 ) | ( n7604 & ~n7895 ) ;
  assign n8200 = ( ~n7896 & n8198 ) | ( ~n7896 & n8199 ) | ( n8198 & n8199 ) ;
  assign n8201 = n8197 | n8200 ;
  assign n8202 = n131 & n7902 ;
  assign n8203 = n7599 & ~n7895 ;
  assign n8204 = ( ~n7896 & n8198 ) | ( ~n7896 & n8203 ) | ( n8198 & n8203 ) ;
  assign n8205 = n7902 | n8204 ;
  assign n8206 = ( n8196 & n8202 ) | ( n8196 & ~n8205 ) | ( n8202 & ~n8205 ) ;
  assign n8207 = ( n7902 & n8199 ) | ( n7902 & n8203 ) | ( n8199 & n8203 ) ;
  assign n8208 = n8199 & ~n8207 ;
  assign n8209 = ( n131 & n7902 ) | ( n131 & n8196 ) | ( n7902 & n8196 ) ;
  assign n8210 = ( ~n8206 & n8208 ) | ( ~n8206 & n8209 ) | ( n8208 & n8209 ) ;
  assign n8211 = ( n132 & ~n8190 ) | ( n132 & n8201 ) | ( ~n8190 & n8201 ) ;
  assign n8212 = n132 & ~n8190 ;
  assign n8213 = ( n8195 & n8211 ) | ( n8195 & n8212 ) | ( n8211 & n8212 ) ;
  assign n8214 = ( n8195 & ~n8211 ) | ( n8195 & n8212 ) | ( ~n8211 & n8212 ) ;
  assign n8215 = ( n8211 & ~n8213 ) | ( n8211 & n8214 ) | ( ~n8213 & n8214 ) ;
  assign n8216 = ~n746 & n8112 ;
  assign n8217 = ( ~n746 & n8112 ) | ( ~n746 & n8201 ) | ( n8112 & n8201 ) ;
  assign n8218 = ( n8117 & n8216 ) | ( n8117 & n8217 ) | ( n8216 & n8217 ) ;
  assign n8219 = ( ~n8117 & n8216 ) | ( ~n8117 & n8217 ) | ( n8216 & n8217 ) ;
  assign n8220 = ( n8117 & ~n8218 ) | ( n8117 & n8219 ) | ( ~n8218 & n8219 ) ;
  assign n8221 = x22 | x23 ;
  assign n8222 = x24 | n8221 ;
  assign n8223 = n7897 & ~n8222 ;
  assign n8224 = ~n7904 & n8201 ;
  assign n8225 = ~n7897 & n8222 ;
  assign n8226 = ( x25 & ~n8201 ) | ( x25 & n8225 ) | ( ~n8201 & n8225 ) ;
  assign n8227 = ( ~n8223 & n8224 ) | ( ~n8223 & n8226 ) | ( n8224 & n8226 ) ;
  assign n8228 = n7897 & ~n8201 ;
  assign n8229 = ( x26 & n8224 ) | ( x26 & n8228 ) | ( n8224 & n8228 ) ;
  assign n8230 = ( ~x26 & n8224 ) | ( ~x26 & n8228 ) | ( n8224 & n8228 ) ;
  assign n8231 = ( x26 & ~n8229 ) | ( x26 & n8230 ) | ( ~n8229 & n8230 ) ;
  assign n8232 = ( ~n7594 & n8227 ) | ( ~n7594 & n8231 ) | ( n8227 & n8231 ) ;
  assign n8233 = ~n7594 & n7897 ;
  assign n8234 = ( n7910 & n8201 ) | ( n7910 & n8233 ) | ( n8201 & n8233 ) ;
  assign n8235 = ( x27 & n8230 ) | ( x27 & n8234 ) | ( n8230 & n8234 ) ;
  assign n8236 = ( ~x27 & n8230 ) | ( ~x27 & n8234 ) | ( n8230 & n8234 ) ;
  assign n8237 = ( x27 & ~n8235 ) | ( x27 & n8236 ) | ( ~n8235 & n8236 ) ;
  assign n8238 = ( ~n7296 & n8232 ) | ( ~n7296 & n8237 ) | ( n8232 & n8237 ) ;
  assign n8239 = ( n7296 & ~n7909 ) | ( n7296 & n8201 ) | ( ~n7909 & n8201 ) ;
  assign n8240 = n7296 & ~n7909 ;
  assign n8241 = ( n7913 & n8239 ) | ( n7913 & n8240 ) | ( n8239 & n8240 ) ;
  assign n8242 = ( ~n7913 & n8239 ) | ( ~n7913 & n8240 ) | ( n8239 & n8240 ) ;
  assign n8243 = ( n7913 & ~n8241 ) | ( n7913 & n8242 ) | ( ~n8241 & n8242 ) ;
  assign n8244 = ( ~n7006 & n8238 ) | ( ~n7006 & n8243 ) | ( n8238 & n8243 ) ;
  assign n8245 = ( n7006 & ~n7914 ) | ( n7006 & n8201 ) | ( ~n7914 & n8201 ) ;
  assign n8246 = n7006 & ~n7914 ;
  assign n8247 = ( n7919 & n8245 ) | ( n7919 & n8246 ) | ( n8245 & n8246 ) ;
  assign n8248 = ( ~n7919 & n8245 ) | ( ~n7919 & n8246 ) | ( n8245 & n8246 ) ;
  assign n8249 = ( n7919 & ~n8247 ) | ( n7919 & n8248 ) | ( ~n8247 & n8248 ) ;
  assign n8250 = ( ~n6723 & n8244 ) | ( ~n6723 & n8249 ) | ( n8244 & n8249 ) ;
  assign n8251 = ( n6723 & ~n7920 ) | ( n6723 & n8201 ) | ( ~n7920 & n8201 ) ;
  assign n8252 = n6723 & ~n7920 ;
  assign n8253 = ( n7925 & n8251 ) | ( n7925 & n8252 ) | ( n8251 & n8252 ) ;
  assign n8254 = ( ~n7925 & n8251 ) | ( ~n7925 & n8252 ) | ( n8251 & n8252 ) ;
  assign n8255 = ( n7925 & ~n8253 ) | ( n7925 & n8254 ) | ( ~n8253 & n8254 ) ;
  assign n8256 = ( ~n6442 & n8250 ) | ( ~n6442 & n8255 ) | ( n8250 & n8255 ) ;
  assign n8257 = ( n6442 & ~n7926 ) | ( n6442 & n8201 ) | ( ~n7926 & n8201 ) ;
  assign n8258 = n6442 & ~n7926 ;
  assign n8259 = ( n7931 & n8257 ) | ( n7931 & n8258 ) | ( n8257 & n8258 ) ;
  assign n8260 = ( ~n7931 & n8257 ) | ( ~n7931 & n8258 ) | ( n8257 & n8258 ) ;
  assign n8261 = ( n7931 & ~n8259 ) | ( n7931 & n8260 ) | ( ~n8259 & n8260 ) ;
  assign n8262 = ( ~n6172 & n8256 ) | ( ~n6172 & n8261 ) | ( n8256 & n8261 ) ;
  assign n8263 = ~n6172 & n7932 ;
  assign n8264 = ( ~n6172 & n7932 ) | ( ~n6172 & n8201 ) | ( n7932 & n8201 ) ;
  assign n8265 = ( n7937 & n8263 ) | ( n7937 & n8264 ) | ( n8263 & n8264 ) ;
  assign n8266 = ( ~n7937 & n8263 ) | ( ~n7937 & n8264 ) | ( n8263 & n8264 ) ;
  assign n8267 = ( n7937 & ~n8265 ) | ( n7937 & n8266 ) | ( ~n8265 & n8266 ) ;
  assign n8268 = ( ~n5905 & n8262 ) | ( ~n5905 & n8267 ) | ( n8262 & n8267 ) ;
  assign n8269 = ( n5905 & ~n7938 ) | ( n5905 & n8201 ) | ( ~n7938 & n8201 ) ;
  assign n8270 = n5905 & ~n7938 ;
  assign n8271 = ( n7943 & n8269 ) | ( n7943 & n8270 ) | ( n8269 & n8270 ) ;
  assign n8272 = ( ~n7943 & n8269 ) | ( ~n7943 & n8270 ) | ( n8269 & n8270 ) ;
  assign n8273 = ( n7943 & ~n8271 ) | ( n7943 & n8272 ) | ( ~n8271 & n8272 ) ;
  assign n8274 = ( ~n5642 & n8268 ) | ( ~n5642 & n8273 ) | ( n8268 & n8273 ) ;
  assign n8275 = ( n5642 & ~n7944 ) | ( n5642 & n8201 ) | ( ~n7944 & n8201 ) ;
  assign n8276 = n5642 & ~n7944 ;
  assign n8277 = ( n7949 & n8275 ) | ( n7949 & n8276 ) | ( n8275 & n8276 ) ;
  assign n8278 = ( ~n7949 & n8275 ) | ( ~n7949 & n8276 ) | ( n8275 & n8276 ) ;
  assign n8279 = ( n7949 & ~n8277 ) | ( n7949 & n8278 ) | ( ~n8277 & n8278 ) ;
  assign n8280 = ( ~n5386 & n8274 ) | ( ~n5386 & n8279 ) | ( n8274 & n8279 ) ;
  assign n8281 = ( n5386 & ~n7950 ) | ( n5386 & n8201 ) | ( ~n7950 & n8201 ) ;
  assign n8282 = n5386 & ~n7950 ;
  assign n8283 = ( n7955 & n8281 ) | ( n7955 & n8282 ) | ( n8281 & n8282 ) ;
  assign n8284 = ( ~n7955 & n8281 ) | ( ~n7955 & n8282 ) | ( n8281 & n8282 ) ;
  assign n8285 = ( n7955 & ~n8283 ) | ( n7955 & n8284 ) | ( ~n8283 & n8284 ) ;
  assign n8286 = ( ~n5139 & n8280 ) | ( ~n5139 & n8285 ) | ( n8280 & n8285 ) ;
  assign n8287 = ( n5139 & ~n7956 ) | ( n5139 & n8201 ) | ( ~n7956 & n8201 ) ;
  assign n8288 = n5139 & ~n7956 ;
  assign n8289 = ( n7961 & n8287 ) | ( n7961 & n8288 ) | ( n8287 & n8288 ) ;
  assign n8290 = ( ~n7961 & n8287 ) | ( ~n7961 & n8288 ) | ( n8287 & n8288 ) ;
  assign n8291 = ( n7961 & ~n8289 ) | ( n7961 & n8290 ) | ( ~n8289 & n8290 ) ;
  assign n8292 = ( ~n4898 & n8286 ) | ( ~n4898 & n8291 ) | ( n8286 & n8291 ) ;
  assign n8293 = ( n4898 & ~n7962 ) | ( n4898 & n8201 ) | ( ~n7962 & n8201 ) ;
  assign n8294 = n4898 & ~n7962 ;
  assign n8295 = ( n7967 & n8293 ) | ( n7967 & n8294 ) | ( n8293 & n8294 ) ;
  assign n8296 = ( ~n7967 & n8293 ) | ( ~n7967 & n8294 ) | ( n8293 & n8294 ) ;
  assign n8297 = ( n7967 & ~n8295 ) | ( n7967 & n8296 ) | ( ~n8295 & n8296 ) ;
  assign n8298 = ( ~n4661 & n8292 ) | ( ~n4661 & n8297 ) | ( n8292 & n8297 ) ;
  assign n8299 = ( n4661 & ~n7968 ) | ( n4661 & n8201 ) | ( ~n7968 & n8201 ) ;
  assign n8300 = n4661 & ~n7968 ;
  assign n8301 = ( n7973 & n8299 ) | ( n7973 & n8300 ) | ( n8299 & n8300 ) ;
  assign n8302 = ( ~n7973 & n8299 ) | ( ~n7973 & n8300 ) | ( n8299 & n8300 ) ;
  assign n8303 = ( n7973 & ~n8301 ) | ( n7973 & n8302 ) | ( ~n8301 & n8302 ) ;
  assign n8304 = ( ~n4432 & n8298 ) | ( ~n4432 & n8303 ) | ( n8298 & n8303 ) ;
  assign n8305 = n4432 & ~n7974 ;
  assign n8306 = ( n4432 & ~n7974 ) | ( n4432 & n8201 ) | ( ~n7974 & n8201 ) ;
  assign n8307 = ( ~n7979 & n8305 ) | ( ~n7979 & n8306 ) | ( n8305 & n8306 ) ;
  assign n8308 = ( n7979 & n8305 ) | ( n7979 & n8306 ) | ( n8305 & n8306 ) ;
  assign n8309 = ( n7979 & n8307 ) | ( n7979 & ~n8308 ) | ( n8307 & ~n8308 ) ;
  assign n8310 = ( ~n4203 & n8304 ) | ( ~n4203 & n8309 ) | ( n8304 & n8309 ) ;
  assign n8311 = ~n4203 & n7980 ;
  assign n8312 = ( ~n4203 & n7980 ) | ( ~n4203 & n8201 ) | ( n7980 & n8201 ) ;
  assign n8313 = ( ~n7985 & n8311 ) | ( ~n7985 & n8312 ) | ( n8311 & n8312 ) ;
  assign n8314 = ( n7985 & n8311 ) | ( n7985 & n8312 ) | ( n8311 & n8312 ) ;
  assign n8315 = ( n7985 & n8313 ) | ( n7985 & ~n8314 ) | ( n8313 & ~n8314 ) ;
  assign n8316 = ( ~n3985 & n8310 ) | ( ~n3985 & n8315 ) | ( n8310 & n8315 ) ;
  assign n8317 = ( n3985 & ~n7986 ) | ( n3985 & n8201 ) | ( ~n7986 & n8201 ) ;
  assign n8318 = n3985 & ~n7986 ;
  assign n8319 = ( n7991 & n8317 ) | ( n7991 & n8318 ) | ( n8317 & n8318 ) ;
  assign n8320 = ( ~n7991 & n8317 ) | ( ~n7991 & n8318 ) | ( n8317 & n8318 ) ;
  assign n8321 = ( n7991 & ~n8319 ) | ( n7991 & n8320 ) | ( ~n8319 & n8320 ) ;
  assign n8322 = ( ~n3772 & n8316 ) | ( ~n3772 & n8321 ) | ( n8316 & n8321 ) ;
  assign n8323 = ( n3772 & ~n7992 ) | ( n3772 & n8201 ) | ( ~n7992 & n8201 ) ;
  assign n8324 = n3772 & ~n7992 ;
  assign n8325 = ( n7997 & n8323 ) | ( n7997 & n8324 ) | ( n8323 & n8324 ) ;
  assign n8326 = ( ~n7997 & n8323 ) | ( ~n7997 & n8324 ) | ( n8323 & n8324 ) ;
  assign n8327 = ( n7997 & ~n8325 ) | ( n7997 & n8326 ) | ( ~n8325 & n8326 ) ;
  assign n8328 = ( ~n3567 & n8322 ) | ( ~n3567 & n8327 ) | ( n8322 & n8327 ) ;
  assign n8329 = ( n3567 & ~n7998 ) | ( n3567 & n8201 ) | ( ~n7998 & n8201 ) ;
  assign n8330 = n3567 & ~n7998 ;
  assign n8331 = ( n8003 & n8329 ) | ( n8003 & n8330 ) | ( n8329 & n8330 ) ;
  assign n8332 = ( ~n8003 & n8329 ) | ( ~n8003 & n8330 ) | ( n8329 & n8330 ) ;
  assign n8333 = ( n8003 & ~n8331 ) | ( n8003 & n8332 ) | ( ~n8331 & n8332 ) ;
  assign n8334 = ( ~n3362 & n8328 ) | ( ~n3362 & n8333 ) | ( n8328 & n8333 ) ;
  assign n8335 = ( n3362 & ~n8004 ) | ( n3362 & n8201 ) | ( ~n8004 & n8201 ) ;
  assign n8336 = n3362 & ~n8004 ;
  assign n8337 = ( n8009 & n8335 ) | ( n8009 & n8336 ) | ( n8335 & n8336 ) ;
  assign n8338 = ( ~n8009 & n8335 ) | ( ~n8009 & n8336 ) | ( n8335 & n8336 ) ;
  assign n8339 = ( n8009 & ~n8337 ) | ( n8009 & n8338 ) | ( ~n8337 & n8338 ) ;
  assign n8340 = ( ~n3169 & n8334 ) | ( ~n3169 & n8339 ) | ( n8334 & n8339 ) ;
  assign n8341 = ~n3169 & n8010 ;
  assign n8342 = ( ~n3169 & n8010 ) | ( ~n3169 & n8201 ) | ( n8010 & n8201 ) ;
  assign n8343 = ( ~n8015 & n8341 ) | ( ~n8015 & n8342 ) | ( n8341 & n8342 ) ;
  assign n8344 = ( n8015 & n8341 ) | ( n8015 & n8342 ) | ( n8341 & n8342 ) ;
  assign n8345 = ( n8015 & n8343 ) | ( n8015 & ~n8344 ) | ( n8343 & ~n8344 ) ;
  assign n8346 = ( ~n2979 & n8340 ) | ( ~n2979 & n8345 ) | ( n8340 & n8345 ) ;
  assign n8347 = n2979 & ~n8016 ;
  assign n8348 = ( n2979 & ~n8016 ) | ( n2979 & n8201 ) | ( ~n8016 & n8201 ) ;
  assign n8349 = ( n8021 & n8347 ) | ( n8021 & n8348 ) | ( n8347 & n8348 ) ;
  assign n8350 = ( ~n8021 & n8347 ) | ( ~n8021 & n8348 ) | ( n8347 & n8348 ) ;
  assign n8351 = ( n8021 & ~n8349 ) | ( n8021 & n8350 ) | ( ~n8349 & n8350 ) ;
  assign n8352 = ( ~n2791 & n8346 ) | ( ~n2791 & n8351 ) | ( n8346 & n8351 ) ;
  assign n8353 = ~n2791 & n8022 ;
  assign n8354 = ( ~n2791 & n8022 ) | ( ~n2791 & n8201 ) | ( n8022 & n8201 ) ;
  assign n8355 = ( ~n8027 & n8353 ) | ( ~n8027 & n8354 ) | ( n8353 & n8354 ) ;
  assign n8356 = ( n8027 & n8353 ) | ( n8027 & n8354 ) | ( n8353 & n8354 ) ;
  assign n8357 = ( n8027 & n8355 ) | ( n8027 & ~n8356 ) | ( n8355 & ~n8356 ) ;
  assign n8358 = ( ~n2615 & n8352 ) | ( ~n2615 & n8357 ) | ( n8352 & n8357 ) ;
  assign n8359 = ~n2615 & n8028 ;
  assign n8360 = ( ~n2615 & n8028 ) | ( ~n2615 & n8201 ) | ( n8028 & n8201 ) ;
  assign n8361 = ( ~n8033 & n8359 ) | ( ~n8033 & n8360 ) | ( n8359 & n8360 ) ;
  assign n8362 = ( n8033 & n8359 ) | ( n8033 & n8360 ) | ( n8359 & n8360 ) ;
  assign n8363 = ( n8033 & n8361 ) | ( n8033 & ~n8362 ) | ( n8361 & ~n8362 ) ;
  assign n8364 = ( ~n2443 & n8358 ) | ( ~n2443 & n8363 ) | ( n8358 & n8363 ) ;
  assign n8365 = ( n2443 & ~n8034 ) | ( n2443 & n8201 ) | ( ~n8034 & n8201 ) ;
  assign n8366 = n2443 & ~n8034 ;
  assign n8367 = ( n8039 & n8365 ) | ( n8039 & n8366 ) | ( n8365 & n8366 ) ;
  assign n8368 = ( ~n8039 & n8365 ) | ( ~n8039 & n8366 ) | ( n8365 & n8366 ) ;
  assign n8369 = ( n8039 & ~n8367 ) | ( n8039 & n8368 ) | ( ~n8367 & n8368 ) ;
  assign n8370 = ( ~n2277 & n8364 ) | ( ~n2277 & n8369 ) | ( n8364 & n8369 ) ;
  assign n8371 = ~n2277 & n8040 ;
  assign n8372 = ( ~n2277 & n8040 ) | ( ~n2277 & n8201 ) | ( n8040 & n8201 ) ;
  assign n8373 = ( n8045 & n8371 ) | ( n8045 & n8372 ) | ( n8371 & n8372 ) ;
  assign n8374 = ( ~n8045 & n8371 ) | ( ~n8045 & n8372 ) | ( n8371 & n8372 ) ;
  assign n8375 = ( n8045 & ~n8373 ) | ( n8045 & n8374 ) | ( ~n8373 & n8374 ) ;
  assign n8376 = ( ~n2111 & n8370 ) | ( ~n2111 & n8375 ) | ( n8370 & n8375 ) ;
  assign n8377 = ( n2111 & ~n8046 ) | ( n2111 & n8201 ) | ( ~n8046 & n8201 ) ;
  assign n8378 = n2111 & ~n8046 ;
  assign n8379 = ( n8051 & n8377 ) | ( n8051 & n8378 ) | ( n8377 & n8378 ) ;
  assign n8380 = ( ~n8051 & n8377 ) | ( ~n8051 & n8378 ) | ( n8377 & n8378 ) ;
  assign n8381 = ( n8051 & ~n8379 ) | ( n8051 & n8380 ) | ( ~n8379 & n8380 ) ;
  assign n8382 = ( ~n1949 & n8376 ) | ( ~n1949 & n8381 ) | ( n8376 & n8381 ) ;
  assign n8383 = ( n1949 & ~n8052 ) | ( n1949 & n8201 ) | ( ~n8052 & n8201 ) ;
  assign n8384 = n1949 & ~n8052 ;
  assign n8385 = ( n8057 & n8383 ) | ( n8057 & n8384 ) | ( n8383 & n8384 ) ;
  assign n8386 = ( ~n8057 & n8383 ) | ( ~n8057 & n8384 ) | ( n8383 & n8384 ) ;
  assign n8387 = ( n8057 & ~n8385 ) | ( n8057 & n8386 ) | ( ~n8385 & n8386 ) ;
  assign n8388 = ( ~n1802 & n8382 ) | ( ~n1802 & n8387 ) | ( n8382 & n8387 ) ;
  assign n8389 = n1802 & ~n8058 ;
  assign n8390 = ( n1802 & ~n8058 ) | ( n1802 & n8201 ) | ( ~n8058 & n8201 ) ;
  assign n8391 = ( n8063 & n8389 ) | ( n8063 & n8390 ) | ( n8389 & n8390 ) ;
  assign n8392 = ( ~n8063 & n8389 ) | ( ~n8063 & n8390 ) | ( n8389 & n8390 ) ;
  assign n8393 = ( n8063 & ~n8391 ) | ( n8063 & n8392 ) | ( ~n8391 & n8392 ) ;
  assign n8394 = ( ~n1661 & n8388 ) | ( ~n1661 & n8393 ) | ( n8388 & n8393 ) ;
  assign n8395 = n1661 & ~n8064 ;
  assign n8396 = ( n1661 & ~n8064 ) | ( n1661 & n8201 ) | ( ~n8064 & n8201 ) ;
  assign n8397 = ( n8069 & n8395 ) | ( n8069 & n8396 ) | ( n8395 & n8396 ) ;
  assign n8398 = ( ~n8069 & n8395 ) | ( ~n8069 & n8396 ) | ( n8395 & n8396 ) ;
  assign n8399 = ( n8069 & ~n8397 ) | ( n8069 & n8398 ) | ( ~n8397 & n8398 ) ;
  assign n8400 = ( ~n1523 & n8394 ) | ( ~n1523 & n8399 ) | ( n8394 & n8399 ) ;
  assign n8401 = ~n1523 & n8070 ;
  assign n8402 = ( ~n1523 & n8070 ) | ( ~n1523 & n8201 ) | ( n8070 & n8201 ) ;
  assign n8403 = ( n8075 & n8401 ) | ( n8075 & n8402 ) | ( n8401 & n8402 ) ;
  assign n8404 = ( ~n8075 & n8401 ) | ( ~n8075 & n8402 ) | ( n8401 & n8402 ) ;
  assign n8405 = ( n8075 & ~n8403 ) | ( n8075 & n8404 ) | ( ~n8403 & n8404 ) ;
  assign n8406 = ( ~n1393 & n8400 ) | ( ~n1393 & n8405 ) | ( n8400 & n8405 ) ;
  assign n8407 = ~n1393 & n8076 ;
  assign n8408 = ( ~n1393 & n8076 ) | ( ~n1393 & n8201 ) | ( n8076 & n8201 ) ;
  assign n8409 = ( ~n8081 & n8407 ) | ( ~n8081 & n8408 ) | ( n8407 & n8408 ) ;
  assign n8410 = ( n8081 & n8407 ) | ( n8081 & n8408 ) | ( n8407 & n8408 ) ;
  assign n8411 = ( n8081 & n8409 ) | ( n8081 & ~n8410 ) | ( n8409 & ~n8410 ) ;
  assign n8412 = ( ~n1266 & n8406 ) | ( ~n1266 & n8411 ) | ( n8406 & n8411 ) ;
  assign n8413 = ~n1266 & n8082 ;
  assign n8414 = ( ~n1266 & n8082 ) | ( ~n1266 & n8201 ) | ( n8082 & n8201 ) ;
  assign n8415 = ( n8087 & n8413 ) | ( n8087 & n8414 ) | ( n8413 & n8414 ) ;
  assign n8416 = ( ~n8087 & n8413 ) | ( ~n8087 & n8414 ) | ( n8413 & n8414 ) ;
  assign n8417 = ( n8087 & ~n8415 ) | ( n8087 & n8416 ) | ( ~n8415 & n8416 ) ;
  assign n8418 = ( ~n1150 & n8412 ) | ( ~n1150 & n8417 ) | ( n8412 & n8417 ) ;
  assign n8419 = ~n1150 & n8088 ;
  assign n8420 = ( ~n1150 & n8088 ) | ( ~n1150 & n8201 ) | ( n8088 & n8201 ) ;
  assign n8421 = ( ~n8093 & n8419 ) | ( ~n8093 & n8420 ) | ( n8419 & n8420 ) ;
  assign n8422 = ( n8093 & n8419 ) | ( n8093 & n8420 ) | ( n8419 & n8420 ) ;
  assign n8423 = ( n8093 & n8421 ) | ( n8093 & ~n8422 ) | ( n8421 & ~n8422 ) ;
  assign n8424 = ( ~n1038 & n8418 ) | ( ~n1038 & n8423 ) | ( n8418 & n8423 ) ;
  assign n8425 = ~n1038 & n8094 ;
  assign n8426 = ( ~n1038 & n8094 ) | ( ~n1038 & n8201 ) | ( n8094 & n8201 ) ;
  assign n8427 = ( n8099 & n8425 ) | ( n8099 & n8426 ) | ( n8425 & n8426 ) ;
  assign n8428 = ( ~n8099 & n8425 ) | ( ~n8099 & n8426 ) | ( n8425 & n8426 ) ;
  assign n8429 = ( n8099 & ~n8427 ) | ( n8099 & n8428 ) | ( ~n8427 & n8428 ) ;
  assign n8430 = ( ~n933 & n8424 ) | ( ~n933 & n8429 ) | ( n8424 & n8429 ) ;
  assign n8431 = ~n933 & n8100 ;
  assign n8432 = ( ~n933 & n8100 ) | ( ~n933 & n8201 ) | ( n8100 & n8201 ) ;
  assign n8433 = ( ~n8105 & n8431 ) | ( ~n8105 & n8432 ) | ( n8431 & n8432 ) ;
  assign n8434 = ( n8105 & n8431 ) | ( n8105 & n8432 ) | ( n8431 & n8432 ) ;
  assign n8435 = ( n8105 & n8433 ) | ( n8105 & ~n8434 ) | ( n8433 & ~n8434 ) ;
  assign n8436 = ( ~n839 & n8430 ) | ( ~n839 & n8435 ) | ( n8430 & n8435 ) ;
  assign n8437 = ( n839 & ~n8106 ) | ( n839 & n8201 ) | ( ~n8106 & n8201 ) ;
  assign n8438 = n839 & ~n8106 ;
  assign n8439 = ( n8111 & n8437 ) | ( n8111 & n8438 ) | ( n8437 & n8438 ) ;
  assign n8440 = ( ~n8111 & n8437 ) | ( ~n8111 & n8438 ) | ( n8437 & n8438 ) ;
  assign n8441 = ( n8111 & ~n8439 ) | ( n8111 & n8440 ) | ( ~n8439 & n8440 ) ;
  assign n8442 = ( ~n746 & n8436 ) | ( ~n746 & n8441 ) | ( n8436 & n8441 ) ;
  assign n8443 = ( ~n664 & n8220 ) | ( ~n664 & n8442 ) | ( n8220 & n8442 ) ;
  assign n8444 = ( n664 & ~n8118 ) | ( n664 & n8201 ) | ( ~n8118 & n8201 ) ;
  assign n8445 = n664 & ~n8118 ;
  assign n8446 = ( n8123 & n8444 ) | ( n8123 & n8445 ) | ( n8444 & n8445 ) ;
  assign n8447 = ( ~n8123 & n8444 ) | ( ~n8123 & n8445 ) | ( n8444 & n8445 ) ;
  assign n8448 = ( n8123 & ~n8446 ) | ( n8123 & n8447 ) | ( ~n8446 & n8447 ) ;
  assign n8449 = ( ~n588 & n8443 ) | ( ~n588 & n8448 ) | ( n8443 & n8448 ) ;
  assign n8450 = ~n588 & n8124 ;
  assign n8451 = ( ~n588 & n8124 ) | ( ~n588 & n8201 ) | ( n8124 & n8201 ) ;
  assign n8452 = ( ~n8129 & n8450 ) | ( ~n8129 & n8451 ) | ( n8450 & n8451 ) ;
  assign n8453 = ( n8129 & n8450 ) | ( n8129 & n8451 ) | ( n8450 & n8451 ) ;
  assign n8454 = ( n8129 & n8452 ) | ( n8129 & ~n8453 ) | ( n8452 & ~n8453 ) ;
  assign n8455 = ( ~n518 & n8449 ) | ( ~n518 & n8454 ) | ( n8449 & n8454 ) ;
  assign n8456 = ( n518 & ~n8130 ) | ( n518 & n8201 ) | ( ~n8130 & n8201 ) ;
  assign n8457 = n518 & ~n8130 ;
  assign n8458 = ( n8135 & n8456 ) | ( n8135 & n8457 ) | ( n8456 & n8457 ) ;
  assign n8459 = ( ~n8135 & n8456 ) | ( ~n8135 & n8457 ) | ( n8456 & n8457 ) ;
  assign n8460 = ( n8135 & ~n8458 ) | ( n8135 & n8459 ) | ( ~n8458 & n8459 ) ;
  assign n8461 = ( ~n454 & n8455 ) | ( ~n454 & n8460 ) | ( n8455 & n8460 ) ;
  assign n8462 = n454 & ~n8136 ;
  assign n8463 = ( n454 & ~n8136 ) | ( n454 & n8201 ) | ( ~n8136 & n8201 ) ;
  assign n8464 = ( n8141 & n8462 ) | ( n8141 & n8463 ) | ( n8462 & n8463 ) ;
  assign n8465 = ( ~n8141 & n8462 ) | ( ~n8141 & n8463 ) | ( n8462 & n8463 ) ;
  assign n8466 = ( n8141 & ~n8464 ) | ( n8141 & n8465 ) | ( ~n8464 & n8465 ) ;
  assign n8467 = ( ~n396 & n8461 ) | ( ~n396 & n8466 ) | ( n8461 & n8466 ) ;
  assign n8468 = ( n396 & ~n8142 ) | ( n396 & n8201 ) | ( ~n8142 & n8201 ) ;
  assign n8469 = n396 & ~n8142 ;
  assign n8470 = ( n8147 & n8468 ) | ( n8147 & n8469 ) | ( n8468 & n8469 ) ;
  assign n8471 = ( ~n8147 & n8468 ) | ( ~n8147 & n8469 ) | ( n8468 & n8469 ) ;
  assign n8472 = ( n8147 & ~n8470 ) | ( n8147 & n8471 ) | ( ~n8470 & n8471 ) ;
  assign n8473 = ( ~n344 & n8467 ) | ( ~n344 & n8472 ) | ( n8467 & n8472 ) ;
  assign n8474 = ~n344 & n8148 ;
  assign n8475 = ( ~n344 & n8148 ) | ( ~n344 & n8201 ) | ( n8148 & n8201 ) ;
  assign n8476 = ( ~n8153 & n8474 ) | ( ~n8153 & n8475 ) | ( n8474 & n8475 ) ;
  assign n8477 = ( n8153 & n8474 ) | ( n8153 & n8475 ) | ( n8474 & n8475 ) ;
  assign n8478 = ( n8153 & n8476 ) | ( n8153 & ~n8477 ) | ( n8476 & ~n8477 ) ;
  assign n8479 = ( ~n298 & n8473 ) | ( ~n298 & n8478 ) | ( n8473 & n8478 ) ;
  assign n8480 = ( n298 & ~n8154 ) | ( n298 & n8201 ) | ( ~n8154 & n8201 ) ;
  assign n8481 = n298 & ~n8154 ;
  assign n8482 = ( n8159 & n8480 ) | ( n8159 & n8481 ) | ( n8480 & n8481 ) ;
  assign n8483 = ( ~n8159 & n8480 ) | ( ~n8159 & n8481 ) | ( n8480 & n8481 ) ;
  assign n8484 = ( n8159 & ~n8482 ) | ( n8159 & n8483 ) | ( ~n8482 & n8483 ) ;
  assign n8485 = ( ~n258 & n8479 ) | ( ~n258 & n8484 ) | ( n8479 & n8484 ) ;
  assign n8486 = n258 & ~n8160 ;
  assign n8487 = ( n258 & ~n8160 ) | ( n258 & n8201 ) | ( ~n8160 & n8201 ) ;
  assign n8488 = ( n8165 & n8486 ) | ( n8165 & n8487 ) | ( n8486 & n8487 ) ;
  assign n8489 = ( ~n8165 & n8486 ) | ( ~n8165 & n8487 ) | ( n8486 & n8487 ) ;
  assign n8490 = ( n8165 & ~n8488 ) | ( n8165 & n8489 ) | ( ~n8488 & n8489 ) ;
  assign n8491 = ( ~n225 & n8485 ) | ( ~n225 & n8490 ) | ( n8485 & n8490 ) ;
  assign n8492 = ( n225 & ~n8166 ) | ( n225 & n8201 ) | ( ~n8166 & n8201 ) ;
  assign n8493 = n225 & ~n8166 ;
  assign n8494 = ( n8171 & n8492 ) | ( n8171 & n8493 ) | ( n8492 & n8493 ) ;
  assign n8495 = ( ~n8171 & n8492 ) | ( ~n8171 & n8493 ) | ( n8492 & n8493 ) ;
  assign n8496 = ( n8171 & ~n8494 ) | ( n8171 & n8495 ) | ( ~n8494 & n8495 ) ;
  assign n8497 = ( ~n197 & n8491 ) | ( ~n197 & n8496 ) | ( n8491 & n8496 ) ;
  assign n8498 = ( n197 & ~n8172 ) | ( n197 & n8201 ) | ( ~n8172 & n8201 ) ;
  assign n8499 = n197 & ~n8172 ;
  assign n8500 = ( n8177 & n8498 ) | ( n8177 & n8499 ) | ( n8498 & n8499 ) ;
  assign n8501 = ( ~n8177 & n8498 ) | ( ~n8177 & n8499 ) | ( n8498 & n8499 ) ;
  assign n8502 = ( n8177 & ~n8500 ) | ( n8177 & n8501 ) | ( ~n8500 & n8501 ) ;
  assign n8503 = ( ~n170 & n8497 ) | ( ~n170 & n8502 ) | ( n8497 & n8502 ) ;
  assign n8504 = ~n170 & n8178 ;
  assign n8505 = ( ~n170 & n8178 ) | ( ~n170 & n8201 ) | ( n8178 & n8201 ) ;
  assign n8506 = ( ~n8183 & n8504 ) | ( ~n8183 & n8505 ) | ( n8504 & n8505 ) ;
  assign n8507 = ( n8183 & n8504 ) | ( n8183 & n8505 ) | ( n8504 & n8505 ) ;
  assign n8508 = ( n8183 & n8506 ) | ( n8183 & ~n8507 ) | ( n8506 & ~n8507 ) ;
  assign n8509 = ( ~n142 & n8503 ) | ( ~n142 & n8508 ) | ( n8503 & n8508 ) ;
  assign n8510 = ( n142 & ~n8184 ) | ( n142 & n8201 ) | ( ~n8184 & n8201 ) ;
  assign n8511 = n142 & ~n8184 ;
  assign n8512 = ( n8189 & n8510 ) | ( n8189 & n8511 ) | ( n8510 & n8511 ) ;
  assign n8513 = ( ~n8189 & n8510 ) | ( ~n8189 & n8511 ) | ( n8510 & n8511 ) ;
  assign n8514 = ( n8189 & ~n8512 ) | ( n8189 & n8513 ) | ( ~n8512 & n8513 ) ;
  assign n8515 = ( ~n132 & n8509 ) | ( ~n132 & n8514 ) | ( n8509 & n8514 ) ;
  assign n8516 = ( ~n131 & n8215 ) | ( ~n131 & n8515 ) | ( n8215 & n8515 ) ;
  assign n8517 = n8210 | n8516 ;
  assign n8518 = ~n8221 & n8517 ;
  assign n8519 = x20 | x21 ;
  assign n8520 = x22 | n8519 ;
  assign n8521 = n8201 & ~n8520 ;
  assign n8522 = ~n8201 & n8520 ;
  assign n8523 = ( x23 & ~n8517 ) | ( x23 & n8522 ) | ( ~n8517 & n8522 ) ;
  assign n8524 = ( n8518 & ~n8521 ) | ( n8518 & n8523 ) | ( ~n8521 & n8523 ) ;
  assign n8525 = n8201 & ~n8517 ;
  assign n8526 = ( x24 & n8518 ) | ( x24 & n8525 ) | ( n8518 & n8525 ) ;
  assign n8527 = ( ~x24 & n8518 ) | ( ~x24 & n8525 ) | ( n8518 & n8525 ) ;
  assign n8528 = ( x24 & ~n8526 ) | ( x24 & n8527 ) | ( ~n8526 & n8527 ) ;
  assign n8529 = ( ~n7897 & n8524 ) | ( ~n7897 & n8528 ) | ( n8524 & n8528 ) ;
  assign n8530 = ~n7897 & n8201 ;
  assign n8531 = ( n8228 & n8517 ) | ( n8228 & n8530 ) | ( n8517 & n8530 ) ;
  assign n8532 = ( ~x25 & n8527 ) | ( ~x25 & n8531 ) | ( n8527 & n8531 ) ;
  assign n8533 = ( x25 & n8527 ) | ( x25 & n8531 ) | ( n8527 & n8531 ) ;
  assign n8534 = ( x25 & n8532 ) | ( x25 & ~n8533 ) | ( n8532 & ~n8533 ) ;
  assign n8535 = ( ~n7594 & n8529 ) | ( ~n7594 & n8534 ) | ( n8529 & n8534 ) ;
  assign n8536 = n7594 & ~n8227 ;
  assign n8537 = ( n7594 & ~n8227 ) | ( n7594 & n8517 ) | ( ~n8227 & n8517 ) ;
  assign n8538 = ( n8231 & n8536 ) | ( n8231 & n8537 ) | ( n8536 & n8537 ) ;
  assign n8539 = ( ~n8231 & n8536 ) | ( ~n8231 & n8537 ) | ( n8536 & n8537 ) ;
  assign n8540 = ( n8231 & ~n8538 ) | ( n8231 & n8539 ) | ( ~n8538 & n8539 ) ;
  assign n8541 = ( ~n7296 & n8535 ) | ( ~n7296 & n8540 ) | ( n8535 & n8540 ) ;
  assign n8542 = ( n7296 & ~n8232 ) | ( n7296 & n8517 ) | ( ~n8232 & n8517 ) ;
  assign n8543 = n7296 & ~n8232 ;
  assign n8544 = ( n8237 & n8542 ) | ( n8237 & n8543 ) | ( n8542 & n8543 ) ;
  assign n8545 = ( ~n8237 & n8542 ) | ( ~n8237 & n8543 ) | ( n8542 & n8543 ) ;
  assign n8546 = ( n8237 & ~n8544 ) | ( n8237 & n8545 ) | ( ~n8544 & n8545 ) ;
  assign n8547 = ( ~n7006 & n8541 ) | ( ~n7006 & n8546 ) | ( n8541 & n8546 ) ;
  assign n8548 = n7006 & ~n8238 ;
  assign n8549 = ( n7006 & ~n8238 ) | ( n7006 & n8517 ) | ( ~n8238 & n8517 ) ;
  assign n8550 = ( ~n8243 & n8548 ) | ( ~n8243 & n8549 ) | ( n8548 & n8549 ) ;
  assign n8551 = ( n8243 & n8548 ) | ( n8243 & n8549 ) | ( n8548 & n8549 ) ;
  assign n8552 = ( n8243 & n8550 ) | ( n8243 & ~n8551 ) | ( n8550 & ~n8551 ) ;
  assign n8553 = ( ~n6723 & n8547 ) | ( ~n6723 & n8552 ) | ( n8547 & n8552 ) ;
  assign n8554 = ~n6723 & n8244 ;
  assign n8555 = ( ~n6723 & n8244 ) | ( ~n6723 & n8517 ) | ( n8244 & n8517 ) ;
  assign n8556 = ( ~n8249 & n8554 ) | ( ~n8249 & n8555 ) | ( n8554 & n8555 ) ;
  assign n8557 = ( n8249 & n8554 ) | ( n8249 & n8555 ) | ( n8554 & n8555 ) ;
  assign n8558 = ( n8249 & n8556 ) | ( n8249 & ~n8557 ) | ( n8556 & ~n8557 ) ;
  assign n8559 = ( ~n6442 & n8553 ) | ( ~n6442 & n8558 ) | ( n8553 & n8558 ) ;
  assign n8560 = ( n6442 & ~n8250 ) | ( n6442 & n8517 ) | ( ~n8250 & n8517 ) ;
  assign n8561 = n6442 & ~n8250 ;
  assign n8562 = ( n8255 & n8560 ) | ( n8255 & n8561 ) | ( n8560 & n8561 ) ;
  assign n8563 = ( ~n8255 & n8560 ) | ( ~n8255 & n8561 ) | ( n8560 & n8561 ) ;
  assign n8564 = ( n8255 & ~n8562 ) | ( n8255 & n8563 ) | ( ~n8562 & n8563 ) ;
  assign n8565 = ( ~n6172 & n8559 ) | ( ~n6172 & n8564 ) | ( n8559 & n8564 ) ;
  assign n8566 = n6172 & ~n8256 ;
  assign n8567 = ( n6172 & ~n8256 ) | ( n6172 & n8517 ) | ( ~n8256 & n8517 ) ;
  assign n8568 = ( n8261 & n8566 ) | ( n8261 & n8567 ) | ( n8566 & n8567 ) ;
  assign n8569 = ( ~n8261 & n8566 ) | ( ~n8261 & n8567 ) | ( n8566 & n8567 ) ;
  assign n8570 = ( n8261 & ~n8568 ) | ( n8261 & n8569 ) | ( ~n8568 & n8569 ) ;
  assign n8571 = ( ~n5905 & n8565 ) | ( ~n5905 & n8570 ) | ( n8565 & n8570 ) ;
  assign n8572 = n5905 & ~n8262 ;
  assign n8573 = ( n5905 & ~n8262 ) | ( n5905 & n8517 ) | ( ~n8262 & n8517 ) ;
  assign n8574 = ( ~n8267 & n8572 ) | ( ~n8267 & n8573 ) | ( n8572 & n8573 ) ;
  assign n8575 = ( n8267 & n8572 ) | ( n8267 & n8573 ) | ( n8572 & n8573 ) ;
  assign n8576 = ( n8267 & n8574 ) | ( n8267 & ~n8575 ) | ( n8574 & ~n8575 ) ;
  assign n8577 = ( ~n5642 & n8571 ) | ( ~n5642 & n8576 ) | ( n8571 & n8576 ) ;
  assign n8578 = ~n5642 & n8268 ;
  assign n8579 = ( ~n5642 & n8268 ) | ( ~n5642 & n8517 ) | ( n8268 & n8517 ) ;
  assign n8580 = ( ~n8273 & n8578 ) | ( ~n8273 & n8579 ) | ( n8578 & n8579 ) ;
  assign n8581 = ( n8273 & n8578 ) | ( n8273 & n8579 ) | ( n8578 & n8579 ) ;
  assign n8582 = ( n8273 & n8580 ) | ( n8273 & ~n8581 ) | ( n8580 & ~n8581 ) ;
  assign n8583 = ( ~n5386 & n8577 ) | ( ~n5386 & n8582 ) | ( n8577 & n8582 ) ;
  assign n8584 = ~n5386 & n8274 ;
  assign n8585 = ( ~n5386 & n8274 ) | ( ~n5386 & n8517 ) | ( n8274 & n8517 ) ;
  assign n8586 = ( ~n8279 & n8584 ) | ( ~n8279 & n8585 ) | ( n8584 & n8585 ) ;
  assign n8587 = ( n8279 & n8584 ) | ( n8279 & n8585 ) | ( n8584 & n8585 ) ;
  assign n8588 = ( n8279 & n8586 ) | ( n8279 & ~n8587 ) | ( n8586 & ~n8587 ) ;
  assign n8589 = ( ~n5139 & n8583 ) | ( ~n5139 & n8588 ) | ( n8583 & n8588 ) ;
  assign n8590 = ( n5139 & ~n8280 ) | ( n5139 & n8517 ) | ( ~n8280 & n8517 ) ;
  assign n8591 = n5139 & ~n8280 ;
  assign n8592 = ( n8285 & n8590 ) | ( n8285 & n8591 ) | ( n8590 & n8591 ) ;
  assign n8593 = ( ~n8285 & n8590 ) | ( ~n8285 & n8591 ) | ( n8590 & n8591 ) ;
  assign n8594 = ( n8285 & ~n8592 ) | ( n8285 & n8593 ) | ( ~n8592 & n8593 ) ;
  assign n8595 = ( ~n4898 & n8589 ) | ( ~n4898 & n8594 ) | ( n8589 & n8594 ) ;
  assign n8596 = ~n4898 & n8286 ;
  assign n8597 = ( ~n4898 & n8286 ) | ( ~n4898 & n8517 ) | ( n8286 & n8517 ) ;
  assign n8598 = ( n8291 & n8596 ) | ( n8291 & n8597 ) | ( n8596 & n8597 ) ;
  assign n8599 = ( ~n8291 & n8596 ) | ( ~n8291 & n8597 ) | ( n8596 & n8597 ) ;
  assign n8600 = ( n8291 & ~n8598 ) | ( n8291 & n8599 ) | ( ~n8598 & n8599 ) ;
  assign n8601 = ( ~n4661 & n8595 ) | ( ~n4661 & n8600 ) | ( n8595 & n8600 ) ;
  assign n8602 = ( n4661 & ~n8292 ) | ( n4661 & n8517 ) | ( ~n8292 & n8517 ) ;
  assign n8603 = n4661 & ~n8292 ;
  assign n8604 = ( n8297 & n8602 ) | ( n8297 & n8603 ) | ( n8602 & n8603 ) ;
  assign n8605 = ( ~n8297 & n8602 ) | ( ~n8297 & n8603 ) | ( n8602 & n8603 ) ;
  assign n8606 = ( n8297 & ~n8604 ) | ( n8297 & n8605 ) | ( ~n8604 & n8605 ) ;
  assign n8607 = ( ~n4432 & n8601 ) | ( ~n4432 & n8606 ) | ( n8601 & n8606 ) ;
  assign n8608 = ( n4432 & ~n8298 ) | ( n4432 & n8517 ) | ( ~n8298 & n8517 ) ;
  assign n8609 = n4432 & ~n8298 ;
  assign n8610 = ( n8303 & n8608 ) | ( n8303 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8611 = ( ~n8303 & n8608 ) | ( ~n8303 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8612 = ( n8303 & ~n8610 ) | ( n8303 & n8611 ) | ( ~n8610 & n8611 ) ;
  assign n8613 = ( ~n4203 & n8607 ) | ( ~n4203 & n8612 ) | ( n8607 & n8612 ) ;
  assign n8614 = ( n4203 & ~n8304 ) | ( n4203 & n8517 ) | ( ~n8304 & n8517 ) ;
  assign n8615 = n4203 & ~n8304 ;
  assign n8616 = ( n8309 & n8614 ) | ( n8309 & n8615 ) | ( n8614 & n8615 ) ;
  assign n8617 = ( ~n8309 & n8614 ) | ( ~n8309 & n8615 ) | ( n8614 & n8615 ) ;
  assign n8618 = ( n8309 & ~n8616 ) | ( n8309 & n8617 ) | ( ~n8616 & n8617 ) ;
  assign n8619 = ( ~n3985 & n8613 ) | ( ~n3985 & n8618 ) | ( n8613 & n8618 ) ;
  assign n8620 = ( n3985 & ~n8310 ) | ( n3985 & n8517 ) | ( ~n8310 & n8517 ) ;
  assign n8621 = n3985 & ~n8310 ;
  assign n8622 = ( n8315 & n8620 ) | ( n8315 & n8621 ) | ( n8620 & n8621 ) ;
  assign n8623 = ( ~n8315 & n8620 ) | ( ~n8315 & n8621 ) | ( n8620 & n8621 ) ;
  assign n8624 = ( n8315 & ~n8622 ) | ( n8315 & n8623 ) | ( ~n8622 & n8623 ) ;
  assign n8625 = ( ~n3772 & n8619 ) | ( ~n3772 & n8624 ) | ( n8619 & n8624 ) ;
  assign n8626 = n3772 & ~n8316 ;
  assign n8627 = ( n3772 & ~n8316 ) | ( n3772 & n8517 ) | ( ~n8316 & n8517 ) ;
  assign n8628 = ( n8321 & n8626 ) | ( n8321 & n8627 ) | ( n8626 & n8627 ) ;
  assign n8629 = ( ~n8321 & n8626 ) | ( ~n8321 & n8627 ) | ( n8626 & n8627 ) ;
  assign n8630 = ( n8321 & ~n8628 ) | ( n8321 & n8629 ) | ( ~n8628 & n8629 ) ;
  assign n8631 = ( ~n3567 & n8625 ) | ( ~n3567 & n8630 ) | ( n8625 & n8630 ) ;
  assign n8632 = ( n3567 & ~n8322 ) | ( n3567 & n8517 ) | ( ~n8322 & n8517 ) ;
  assign n8633 = n3567 & ~n8322 ;
  assign n8634 = ( n8327 & n8632 ) | ( n8327 & n8633 ) | ( n8632 & n8633 ) ;
  assign n8635 = ( ~n8327 & n8632 ) | ( ~n8327 & n8633 ) | ( n8632 & n8633 ) ;
  assign n8636 = ( n8327 & ~n8634 ) | ( n8327 & n8635 ) | ( ~n8634 & n8635 ) ;
  assign n8637 = ( ~n3362 & n8631 ) | ( ~n3362 & n8636 ) | ( n8631 & n8636 ) ;
  assign n8638 = ~n3362 & n8328 ;
  assign n8639 = ( ~n3362 & n8328 ) | ( ~n3362 & n8517 ) | ( n8328 & n8517 ) ;
  assign n8640 = ( ~n8333 & n8638 ) | ( ~n8333 & n8639 ) | ( n8638 & n8639 ) ;
  assign n8641 = ( n8333 & n8638 ) | ( n8333 & n8639 ) | ( n8638 & n8639 ) ;
  assign n8642 = ( n8333 & n8640 ) | ( n8333 & ~n8641 ) | ( n8640 & ~n8641 ) ;
  assign n8643 = ( ~n3169 & n8637 ) | ( ~n3169 & n8642 ) | ( n8637 & n8642 ) ;
  assign n8644 = ( n3169 & ~n8334 ) | ( n3169 & n8517 ) | ( ~n8334 & n8517 ) ;
  assign n8645 = n3169 & ~n8334 ;
  assign n8646 = ( n8339 & n8644 ) | ( n8339 & n8645 ) | ( n8644 & n8645 ) ;
  assign n8647 = ( ~n8339 & n8644 ) | ( ~n8339 & n8645 ) | ( n8644 & n8645 ) ;
  assign n8648 = ( n8339 & ~n8646 ) | ( n8339 & n8647 ) | ( ~n8646 & n8647 ) ;
  assign n8649 = ( ~n2979 & n8643 ) | ( ~n2979 & n8648 ) | ( n8643 & n8648 ) ;
  assign n8650 = ( n2979 & ~n8340 ) | ( n2979 & n8517 ) | ( ~n8340 & n8517 ) ;
  assign n8651 = n2979 & ~n8340 ;
  assign n8652 = ( n8345 & n8650 ) | ( n8345 & n8651 ) | ( n8650 & n8651 ) ;
  assign n8653 = ( ~n8345 & n8650 ) | ( ~n8345 & n8651 ) | ( n8650 & n8651 ) ;
  assign n8654 = ( n8345 & ~n8652 ) | ( n8345 & n8653 ) | ( ~n8652 & n8653 ) ;
  assign n8655 = ( ~n2791 & n8649 ) | ( ~n2791 & n8654 ) | ( n8649 & n8654 ) ;
  assign n8656 = ( n2791 & ~n8346 ) | ( n2791 & n8517 ) | ( ~n8346 & n8517 ) ;
  assign n8657 = n2791 & ~n8346 ;
  assign n8658 = ( n8351 & n8656 ) | ( n8351 & n8657 ) | ( n8656 & n8657 ) ;
  assign n8659 = ( ~n8351 & n8656 ) | ( ~n8351 & n8657 ) | ( n8656 & n8657 ) ;
  assign n8660 = ( n8351 & ~n8658 ) | ( n8351 & n8659 ) | ( ~n8658 & n8659 ) ;
  assign n8661 = ( ~n2615 & n8655 ) | ( ~n2615 & n8660 ) | ( n8655 & n8660 ) ;
  assign n8662 = ( n2615 & ~n8352 ) | ( n2615 & n8517 ) | ( ~n8352 & n8517 ) ;
  assign n8663 = n2615 & ~n8352 ;
  assign n8664 = ( n8357 & n8662 ) | ( n8357 & n8663 ) | ( n8662 & n8663 ) ;
  assign n8665 = ( ~n8357 & n8662 ) | ( ~n8357 & n8663 ) | ( n8662 & n8663 ) ;
  assign n8666 = ( n8357 & ~n8664 ) | ( n8357 & n8665 ) | ( ~n8664 & n8665 ) ;
  assign n8667 = ( ~n2443 & n8661 ) | ( ~n2443 & n8666 ) | ( n8661 & n8666 ) ;
  assign n8668 = n2443 & ~n8358 ;
  assign n8669 = ( n2443 & ~n8358 ) | ( n2443 & n8517 ) | ( ~n8358 & n8517 ) ;
  assign n8670 = ( n8363 & n8668 ) | ( n8363 & n8669 ) | ( n8668 & n8669 ) ;
  assign n8671 = ( ~n8363 & n8668 ) | ( ~n8363 & n8669 ) | ( n8668 & n8669 ) ;
  assign n8672 = ( n8363 & ~n8670 ) | ( n8363 & n8671 ) | ( ~n8670 & n8671 ) ;
  assign n8673 = ( ~n2277 & n8667 ) | ( ~n2277 & n8672 ) | ( n8667 & n8672 ) ;
  assign n8674 = ( n2277 & ~n8364 ) | ( n2277 & n8517 ) | ( ~n8364 & n8517 ) ;
  assign n8675 = n2277 & ~n8364 ;
  assign n8676 = ( n8369 & n8674 ) | ( n8369 & n8675 ) | ( n8674 & n8675 ) ;
  assign n8677 = ( ~n8369 & n8674 ) | ( ~n8369 & n8675 ) | ( n8674 & n8675 ) ;
  assign n8678 = ( n8369 & ~n8676 ) | ( n8369 & n8677 ) | ( ~n8676 & n8677 ) ;
  assign n8679 = ( ~n2111 & n8673 ) | ( ~n2111 & n8678 ) | ( n8673 & n8678 ) ;
  assign n8680 = ( n2111 & ~n8370 ) | ( n2111 & n8517 ) | ( ~n8370 & n8517 ) ;
  assign n8681 = n2111 & ~n8370 ;
  assign n8682 = ( n8375 & n8680 ) | ( n8375 & n8681 ) | ( n8680 & n8681 ) ;
  assign n8683 = ( ~n8375 & n8680 ) | ( ~n8375 & n8681 ) | ( n8680 & n8681 ) ;
  assign n8684 = ( n8375 & ~n8682 ) | ( n8375 & n8683 ) | ( ~n8682 & n8683 ) ;
  assign n8685 = ( ~n1949 & n8679 ) | ( ~n1949 & n8684 ) | ( n8679 & n8684 ) ;
  assign n8686 = ( n1949 & ~n8376 ) | ( n1949 & n8517 ) | ( ~n8376 & n8517 ) ;
  assign n8687 = n1949 & ~n8376 ;
  assign n8688 = ( n8381 & n8686 ) | ( n8381 & n8687 ) | ( n8686 & n8687 ) ;
  assign n8689 = ( ~n8381 & n8686 ) | ( ~n8381 & n8687 ) | ( n8686 & n8687 ) ;
  assign n8690 = ( n8381 & ~n8688 ) | ( n8381 & n8689 ) | ( ~n8688 & n8689 ) ;
  assign n8691 = ( ~n1802 & n8685 ) | ( ~n1802 & n8690 ) | ( n8685 & n8690 ) ;
  assign n8692 = ( n1802 & ~n8382 ) | ( n1802 & n8517 ) | ( ~n8382 & n8517 ) ;
  assign n8693 = n1802 & ~n8382 ;
  assign n8694 = ( n8387 & n8692 ) | ( n8387 & n8693 ) | ( n8692 & n8693 ) ;
  assign n8695 = ( ~n8387 & n8692 ) | ( ~n8387 & n8693 ) | ( n8692 & n8693 ) ;
  assign n8696 = ( n8387 & ~n8694 ) | ( n8387 & n8695 ) | ( ~n8694 & n8695 ) ;
  assign n8697 = ( ~n1661 & n8691 ) | ( ~n1661 & n8696 ) | ( n8691 & n8696 ) ;
  assign n8698 = ( n1661 & ~n8388 ) | ( n1661 & n8517 ) | ( ~n8388 & n8517 ) ;
  assign n8699 = n1661 & ~n8388 ;
  assign n8700 = ( n8393 & n8698 ) | ( n8393 & n8699 ) | ( n8698 & n8699 ) ;
  assign n8701 = ( ~n8393 & n8698 ) | ( ~n8393 & n8699 ) | ( n8698 & n8699 ) ;
  assign n8702 = ( n8393 & ~n8700 ) | ( n8393 & n8701 ) | ( ~n8700 & n8701 ) ;
  assign n8703 = ( ~n1523 & n8697 ) | ( ~n1523 & n8702 ) | ( n8697 & n8702 ) ;
  assign n8704 = ~n1523 & n8394 ;
  assign n8705 = ( ~n1523 & n8394 ) | ( ~n1523 & n8517 ) | ( n8394 & n8517 ) ;
  assign n8706 = ( n8399 & n8704 ) | ( n8399 & n8705 ) | ( n8704 & n8705 ) ;
  assign n8707 = ( ~n8399 & n8704 ) | ( ~n8399 & n8705 ) | ( n8704 & n8705 ) ;
  assign n8708 = ( n8399 & ~n8706 ) | ( n8399 & n8707 ) | ( ~n8706 & n8707 ) ;
  assign n8709 = ( ~n1393 & n8703 ) | ( ~n1393 & n8708 ) | ( n8703 & n8708 ) ;
  assign n8710 = ( n1393 & ~n8400 ) | ( n1393 & n8517 ) | ( ~n8400 & n8517 ) ;
  assign n8711 = n1393 & ~n8400 ;
  assign n8712 = ( n8405 & n8710 ) | ( n8405 & n8711 ) | ( n8710 & n8711 ) ;
  assign n8713 = ( ~n8405 & n8710 ) | ( ~n8405 & n8711 ) | ( n8710 & n8711 ) ;
  assign n8714 = ( n8405 & ~n8712 ) | ( n8405 & n8713 ) | ( ~n8712 & n8713 ) ;
  assign n8715 = ( ~n1266 & n8709 ) | ( ~n1266 & n8714 ) | ( n8709 & n8714 ) ;
  assign n8716 = n1266 & ~n8406 ;
  assign n8717 = ( n1266 & ~n8406 ) | ( n1266 & n8517 ) | ( ~n8406 & n8517 ) ;
  assign n8718 = ( ~n8411 & n8716 ) | ( ~n8411 & n8717 ) | ( n8716 & n8717 ) ;
  assign n8719 = ( n8411 & n8716 ) | ( n8411 & n8717 ) | ( n8716 & n8717 ) ;
  assign n8720 = ( n8411 & n8718 ) | ( n8411 & ~n8719 ) | ( n8718 & ~n8719 ) ;
  assign n8721 = ( ~n1150 & n8715 ) | ( ~n1150 & n8720 ) | ( n8715 & n8720 ) ;
  assign n8722 = ( n1150 & ~n8412 ) | ( n1150 & n8517 ) | ( ~n8412 & n8517 ) ;
  assign n8723 = n1150 & ~n8412 ;
  assign n8724 = ( n8417 & n8722 ) | ( n8417 & n8723 ) | ( n8722 & n8723 ) ;
  assign n8725 = ( ~n8417 & n8722 ) | ( ~n8417 & n8723 ) | ( n8722 & n8723 ) ;
  assign n8726 = ( n8417 & ~n8724 ) | ( n8417 & n8725 ) | ( ~n8724 & n8725 ) ;
  assign n8727 = ( ~n1038 & n8721 ) | ( ~n1038 & n8726 ) | ( n8721 & n8726 ) ;
  assign n8728 = n1038 & ~n8418 ;
  assign n8729 = ( n1038 & ~n8418 ) | ( n1038 & n8517 ) | ( ~n8418 & n8517 ) ;
  assign n8730 = ( n8423 & n8728 ) | ( n8423 & n8729 ) | ( n8728 & n8729 ) ;
  assign n8731 = ( ~n8423 & n8728 ) | ( ~n8423 & n8729 ) | ( n8728 & n8729 ) ;
  assign n8732 = ( n8423 & ~n8730 ) | ( n8423 & n8731 ) | ( ~n8730 & n8731 ) ;
  assign n8733 = ( ~n933 & n8727 ) | ( ~n933 & n8732 ) | ( n8727 & n8732 ) ;
  assign n8734 = ~n933 & n8424 ;
  assign n8735 = ( ~n933 & n8424 ) | ( ~n933 & n8517 ) | ( n8424 & n8517 ) ;
  assign n8736 = ( ~n8429 & n8734 ) | ( ~n8429 & n8735 ) | ( n8734 & n8735 ) ;
  assign n8737 = ( n8429 & n8734 ) | ( n8429 & n8735 ) | ( n8734 & n8735 ) ;
  assign n8738 = ( n8429 & n8736 ) | ( n8429 & ~n8737 ) | ( n8736 & ~n8737 ) ;
  assign n8739 = ( ~n839 & n8733 ) | ( ~n839 & n8738 ) | ( n8733 & n8738 ) ;
  assign n8740 = ( n839 & ~n8430 ) | ( n839 & n8517 ) | ( ~n8430 & n8517 ) ;
  assign n8741 = n839 & ~n8430 ;
  assign n8742 = ( n8435 & n8740 ) | ( n8435 & n8741 ) | ( n8740 & n8741 ) ;
  assign n8743 = ( ~n8435 & n8740 ) | ( ~n8435 & n8741 ) | ( n8740 & n8741 ) ;
  assign n8744 = ( n8435 & ~n8742 ) | ( n8435 & n8743 ) | ( ~n8742 & n8743 ) ;
  assign n8745 = ( ~n746 & n8739 ) | ( ~n746 & n8744 ) | ( n8739 & n8744 ) ;
  assign n8746 = n746 & ~n8436 ;
  assign n8747 = ( n746 & ~n8436 ) | ( n746 & n8517 ) | ( ~n8436 & n8517 ) ;
  assign n8748 = ( n8441 & n8746 ) | ( n8441 & n8747 ) | ( n8746 & n8747 ) ;
  assign n8749 = ( ~n8441 & n8746 ) | ( ~n8441 & n8747 ) | ( n8746 & n8747 ) ;
  assign n8750 = ( n8441 & ~n8748 ) | ( n8441 & n8749 ) | ( ~n8748 & n8749 ) ;
  assign n8751 = ( ~n664 & n8745 ) | ( ~n664 & n8750 ) | ( n8745 & n8750 ) ;
  assign n8752 = ~n664 & n8442 ;
  assign n8753 = ( ~n664 & n8442 ) | ( ~n664 & n8517 ) | ( n8442 & n8517 ) ;
  assign n8754 = ( ~n8220 & n8752 ) | ( ~n8220 & n8753 ) | ( n8752 & n8753 ) ;
  assign n8755 = ( n8220 & n8752 ) | ( n8220 & n8753 ) | ( n8752 & n8753 ) ;
  assign n8756 = ( n8220 & n8754 ) | ( n8220 & ~n8755 ) | ( n8754 & ~n8755 ) ;
  assign n8757 = ( ~n588 & n8751 ) | ( ~n588 & n8756 ) | ( n8751 & n8756 ) ;
  assign n8758 = ( n588 & ~n8443 ) | ( n588 & n8517 ) | ( ~n8443 & n8517 ) ;
  assign n8759 = n588 & ~n8443 ;
  assign n8760 = ( n8448 & n8758 ) | ( n8448 & n8759 ) | ( n8758 & n8759 ) ;
  assign n8761 = ( ~n8448 & n8758 ) | ( ~n8448 & n8759 ) | ( n8758 & n8759 ) ;
  assign n8762 = ( n8448 & ~n8760 ) | ( n8448 & n8761 ) | ( ~n8760 & n8761 ) ;
  assign n8763 = ( ~n518 & n8757 ) | ( ~n518 & n8762 ) | ( n8757 & n8762 ) ;
  assign n8764 = ( n518 & ~n8449 ) | ( n518 & n8517 ) | ( ~n8449 & n8517 ) ;
  assign n8765 = n518 & ~n8449 ;
  assign n8766 = ( n8454 & n8764 ) | ( n8454 & n8765 ) | ( n8764 & n8765 ) ;
  assign n8767 = ( ~n8454 & n8764 ) | ( ~n8454 & n8765 ) | ( n8764 & n8765 ) ;
  assign n8768 = ( n8454 & ~n8766 ) | ( n8454 & n8767 ) | ( ~n8766 & n8767 ) ;
  assign n8769 = ( ~n454 & n8763 ) | ( ~n454 & n8768 ) | ( n8763 & n8768 ) ;
  assign n8770 = ( n454 & ~n8455 ) | ( n454 & n8517 ) | ( ~n8455 & n8517 ) ;
  assign n8771 = n454 & ~n8455 ;
  assign n8772 = ( n8460 & n8770 ) | ( n8460 & n8771 ) | ( n8770 & n8771 ) ;
  assign n8773 = ( ~n8460 & n8770 ) | ( ~n8460 & n8771 ) | ( n8770 & n8771 ) ;
  assign n8774 = ( n8460 & ~n8772 ) | ( n8460 & n8773 ) | ( ~n8772 & n8773 ) ;
  assign n8775 = ( ~n396 & n8769 ) | ( ~n396 & n8774 ) | ( n8769 & n8774 ) ;
  assign n8776 = ( n396 & ~n8461 ) | ( n396 & n8517 ) | ( ~n8461 & n8517 ) ;
  assign n8777 = n396 & ~n8461 ;
  assign n8778 = ( n8466 & n8776 ) | ( n8466 & n8777 ) | ( n8776 & n8777 ) ;
  assign n8779 = ( ~n8466 & n8776 ) | ( ~n8466 & n8777 ) | ( n8776 & n8777 ) ;
  assign n8780 = ( n8466 & ~n8778 ) | ( n8466 & n8779 ) | ( ~n8778 & n8779 ) ;
  assign n8781 = ( ~n344 & n8775 ) | ( ~n344 & n8780 ) | ( n8775 & n8780 ) ;
  assign n8782 = ( n344 & ~n8467 ) | ( n344 & n8517 ) | ( ~n8467 & n8517 ) ;
  assign n8783 = n344 & ~n8467 ;
  assign n8784 = ( n8472 & n8782 ) | ( n8472 & n8783 ) | ( n8782 & n8783 ) ;
  assign n8785 = ( ~n8472 & n8782 ) | ( ~n8472 & n8783 ) | ( n8782 & n8783 ) ;
  assign n8786 = ( n8472 & ~n8784 ) | ( n8472 & n8785 ) | ( ~n8784 & n8785 ) ;
  assign n8787 = ( ~n298 & n8781 ) | ( ~n298 & n8786 ) | ( n8781 & n8786 ) ;
  assign n8788 = ~n298 & n8473 ;
  assign n8789 = ( ~n298 & n8473 ) | ( ~n298 & n8517 ) | ( n8473 & n8517 ) ;
  assign n8790 = ( n8478 & n8788 ) | ( n8478 & n8789 ) | ( n8788 & n8789 ) ;
  assign n8791 = ( ~n8478 & n8788 ) | ( ~n8478 & n8789 ) | ( n8788 & n8789 ) ;
  assign n8792 = ( n8478 & ~n8790 ) | ( n8478 & n8791 ) | ( ~n8790 & n8791 ) ;
  assign n8793 = ( ~n258 & n8787 ) | ( ~n258 & n8792 ) | ( n8787 & n8792 ) ;
  assign n8794 = n258 & ~n8479 ;
  assign n8795 = ( n258 & ~n8479 ) | ( n258 & n8517 ) | ( ~n8479 & n8517 ) ;
  assign n8796 = ( n8484 & n8794 ) | ( n8484 & n8795 ) | ( n8794 & n8795 ) ;
  assign n8797 = ( ~n8484 & n8794 ) | ( ~n8484 & n8795 ) | ( n8794 & n8795 ) ;
  assign n8798 = ( n8484 & ~n8796 ) | ( n8484 & n8797 ) | ( ~n8796 & n8797 ) ;
  assign n8799 = ( ~n225 & n8793 ) | ( ~n225 & n8798 ) | ( n8793 & n8798 ) ;
  assign n8800 = ~n225 & n8485 ;
  assign n8801 = ( ~n225 & n8485 ) | ( ~n225 & n8517 ) | ( n8485 & n8517 ) ;
  assign n8802 = ( ~n8490 & n8800 ) | ( ~n8490 & n8801 ) | ( n8800 & n8801 ) ;
  assign n8803 = ( n8490 & n8800 ) | ( n8490 & n8801 ) | ( n8800 & n8801 ) ;
  assign n8804 = ( n8490 & n8802 ) | ( n8490 & ~n8803 ) | ( n8802 & ~n8803 ) ;
  assign n8805 = ( ~n197 & n8799 ) | ( ~n197 & n8804 ) | ( n8799 & n8804 ) ;
  assign n8806 = ( n197 & ~n8491 ) | ( n197 & n8517 ) | ( ~n8491 & n8517 ) ;
  assign n8807 = n197 & ~n8491 ;
  assign n8808 = ( n8496 & n8806 ) | ( n8496 & n8807 ) | ( n8806 & n8807 ) ;
  assign n8809 = ( ~n8496 & n8806 ) | ( ~n8496 & n8807 ) | ( n8806 & n8807 ) ;
  assign n8810 = ( n8496 & ~n8808 ) | ( n8496 & n8809 ) | ( ~n8808 & n8809 ) ;
  assign n8811 = ( ~n170 & n8805 ) | ( ~n170 & n8810 ) | ( n8805 & n8810 ) ;
  assign n8812 = ( n170 & ~n8497 ) | ( n170 & n8517 ) | ( ~n8497 & n8517 ) ;
  assign n8813 = n170 & ~n8497 ;
  assign n8814 = ( n8502 & n8812 ) | ( n8502 & n8813 ) | ( n8812 & n8813 ) ;
  assign n8815 = ( ~n8502 & n8812 ) | ( ~n8502 & n8813 ) | ( n8812 & n8813 ) ;
  assign n8816 = ( n8502 & ~n8814 ) | ( n8502 & n8815 ) | ( ~n8814 & n8815 ) ;
  assign n8817 = ( ~n142 & n8811 ) | ( ~n142 & n8816 ) | ( n8811 & n8816 ) ;
  assign n8818 = ( n142 & ~n8503 ) | ( n142 & n8517 ) | ( ~n8503 & n8517 ) ;
  assign n8819 = n142 & ~n8503 ;
  assign n8820 = ( n8508 & n8818 ) | ( n8508 & n8819 ) | ( n8818 & n8819 ) ;
  assign n8821 = ( ~n8508 & n8818 ) | ( ~n8508 & n8819 ) | ( n8818 & n8819 ) ;
  assign n8822 = ( n8508 & ~n8820 ) | ( n8508 & n8821 ) | ( ~n8820 & n8821 ) ;
  assign n8823 = ( ~n132 & n8817 ) | ( ~n132 & n8822 ) | ( n8817 & n8822 ) ;
  assign n8824 = ( n132 & ~n8509 ) | ( n132 & n8517 ) | ( ~n8509 & n8517 ) ;
  assign n8825 = n132 & ~n8509 ;
  assign n8826 = ( n8514 & n8824 ) | ( n8514 & n8825 ) | ( n8824 & n8825 ) ;
  assign n8827 = ( ~n8514 & n8824 ) | ( ~n8514 & n8825 ) | ( n8824 & n8825 ) ;
  assign n8828 = ( n8514 & ~n8826 ) | ( n8514 & n8827 ) | ( ~n8826 & n8827 ) ;
  assign n8829 = ( ~n131 & n8823 ) | ( ~n131 & n8828 ) | ( n8823 & n8828 ) ;
  assign n8830 = n8215 & n8515 ;
  assign n8831 = ~n131 & n8830 ;
  assign n8832 = ( ~n8206 & n8209 ) | ( ~n8206 & n8215 ) | ( n8209 & n8215 ) ;
  assign n8833 = n131 & ~n8832 ;
  assign n8834 = ( n8215 & n8515 ) | ( n8215 & ~n8833 ) | ( n8515 & ~n8833 ) ;
  assign n8835 = n8210 | n8832 ;
  assign n8836 = ( ~n131 & n8834 ) | ( ~n131 & n8835 ) | ( n8834 & n8835 ) ;
  assign n8837 = ( ~n8516 & n8831 ) | ( ~n8516 & n8836 ) | ( n8831 & n8836 ) ;
  assign n8838 = n8829 | n8837 ;
  assign n8839 = ( n132 & ~n8817 ) | ( n132 & n8838 ) | ( ~n8817 & n8838 ) ;
  assign n8840 = n132 & ~n8817 ;
  assign n8841 = ( n8822 & ~n8839 ) | ( n8822 & n8840 ) | ( ~n8839 & n8840 ) ;
  assign n8842 = ( n8822 & n8839 ) | ( n8822 & n8840 ) | ( n8839 & n8840 ) ;
  assign n8843 = ( n8839 & n8841 ) | ( n8839 & ~n8842 ) | ( n8841 & ~n8842 ) ;
  assign n8844 = ~n8519 & n8838 ;
  assign n8845 = x18 | x19 ;
  assign n8846 = x20 | n8845 ;
  assign n8847 = n8517 & ~n8846 ;
  assign n8848 = ~n8517 & n8846 ;
  assign n8849 = ( x21 & ~n8838 ) | ( x21 & n8848 ) | ( ~n8838 & n8848 ) ;
  assign n8850 = ( n8844 & ~n8847 ) | ( n8844 & n8849 ) | ( ~n8847 & n8849 ) ;
  assign n8851 = n8517 & ~n8838 ;
  assign n8852 = ( x22 & n8844 ) | ( x22 & n8851 ) | ( n8844 & n8851 ) ;
  assign n8853 = ( ~x22 & n8844 ) | ( ~x22 & n8851 ) | ( n8844 & n8851 ) ;
  assign n8854 = ( x22 & ~n8852 ) | ( x22 & n8853 ) | ( ~n8852 & n8853 ) ;
  assign n8855 = ( ~n8201 & n8850 ) | ( ~n8201 & n8854 ) | ( n8850 & n8854 ) ;
  assign n8856 = ~n8201 & n8517 ;
  assign n8857 = ( n8525 & n8838 ) | ( n8525 & n8856 ) | ( n8838 & n8856 ) ;
  assign n8858 = ( ~x23 & n8853 ) | ( ~x23 & n8857 ) | ( n8853 & n8857 ) ;
  assign n8859 = ( x23 & n8853 ) | ( x23 & n8857 ) | ( n8853 & n8857 ) ;
  assign n8860 = ( x23 & n8858 ) | ( x23 & ~n8859 ) | ( n8858 & ~n8859 ) ;
  assign n8861 = ( ~n7897 & n8855 ) | ( ~n7897 & n8860 ) | ( n8855 & n8860 ) ;
  assign n8862 = n7897 & ~n8524 ;
  assign n8863 = ( n7897 & ~n8524 ) | ( n7897 & n8838 ) | ( ~n8524 & n8838 ) ;
  assign n8864 = ( ~n8528 & n8862 ) | ( ~n8528 & n8863 ) | ( n8862 & n8863 ) ;
  assign n8865 = ( n8528 & n8862 ) | ( n8528 & n8863 ) | ( n8862 & n8863 ) ;
  assign n8866 = ( n8528 & n8864 ) | ( n8528 & ~n8865 ) | ( n8864 & ~n8865 ) ;
  assign n8867 = ( ~n7594 & n8861 ) | ( ~n7594 & n8866 ) | ( n8861 & n8866 ) ;
  assign n8868 = ~n7594 & n8529 ;
  assign n8869 = ( ~n7594 & n8529 ) | ( ~n7594 & n8838 ) | ( n8529 & n8838 ) ;
  assign n8870 = ( ~n8534 & n8868 ) | ( ~n8534 & n8869 ) | ( n8868 & n8869 ) ;
  assign n8871 = ( n8534 & n8868 ) | ( n8534 & n8869 ) | ( n8868 & n8869 ) ;
  assign n8872 = ( n8534 & n8870 ) | ( n8534 & ~n8871 ) | ( n8870 & ~n8871 ) ;
  assign n8873 = ( ~n7296 & n8867 ) | ( ~n7296 & n8872 ) | ( n8867 & n8872 ) ;
  assign n8874 = ( n7296 & ~n8535 ) | ( n7296 & n8838 ) | ( ~n8535 & n8838 ) ;
  assign n8875 = n7296 & ~n8535 ;
  assign n8876 = ( n8540 & n8874 ) | ( n8540 & n8875 ) | ( n8874 & n8875 ) ;
  assign n8877 = ( ~n8540 & n8874 ) | ( ~n8540 & n8875 ) | ( n8874 & n8875 ) ;
  assign n8878 = ( n8540 & ~n8876 ) | ( n8540 & n8877 ) | ( ~n8876 & n8877 ) ;
  assign n8879 = ( ~n7006 & n8873 ) | ( ~n7006 & n8878 ) | ( n8873 & n8878 ) ;
  assign n8880 = n7006 & ~n8541 ;
  assign n8881 = ( n7006 & ~n8541 ) | ( n7006 & n8838 ) | ( ~n8541 & n8838 ) ;
  assign n8882 = ( n8546 & n8880 ) | ( n8546 & n8881 ) | ( n8880 & n8881 ) ;
  assign n8883 = ( ~n8546 & n8880 ) | ( ~n8546 & n8881 ) | ( n8880 & n8881 ) ;
  assign n8884 = ( n8546 & ~n8882 ) | ( n8546 & n8883 ) | ( ~n8882 & n8883 ) ;
  assign n8885 = ( ~n6723 & n8879 ) | ( ~n6723 & n8884 ) | ( n8879 & n8884 ) ;
  assign n8886 = ( n6723 & ~n8547 ) | ( n6723 & n8838 ) | ( ~n8547 & n8838 ) ;
  assign n8887 = n6723 & ~n8547 ;
  assign n8888 = ( n8552 & n8886 ) | ( n8552 & n8887 ) | ( n8886 & n8887 ) ;
  assign n8889 = ( ~n8552 & n8886 ) | ( ~n8552 & n8887 ) | ( n8886 & n8887 ) ;
  assign n8890 = ( n8552 & ~n8888 ) | ( n8552 & n8889 ) | ( ~n8888 & n8889 ) ;
  assign n8891 = ( ~n6442 & n8885 ) | ( ~n6442 & n8890 ) | ( n8885 & n8890 ) ;
  assign n8892 = ( n6442 & ~n8553 ) | ( n6442 & n8838 ) | ( ~n8553 & n8838 ) ;
  assign n8893 = n6442 & ~n8553 ;
  assign n8894 = ( n8558 & n8892 ) | ( n8558 & n8893 ) | ( n8892 & n8893 ) ;
  assign n8895 = ( ~n8558 & n8892 ) | ( ~n8558 & n8893 ) | ( n8892 & n8893 ) ;
  assign n8896 = ( n8558 & ~n8894 ) | ( n8558 & n8895 ) | ( ~n8894 & n8895 ) ;
  assign n8897 = ( ~n6172 & n8891 ) | ( ~n6172 & n8896 ) | ( n8891 & n8896 ) ;
  assign n8898 = ( n6172 & ~n8559 ) | ( n6172 & n8838 ) | ( ~n8559 & n8838 ) ;
  assign n8899 = n6172 & ~n8559 ;
  assign n8900 = ( n8564 & n8898 ) | ( n8564 & n8899 ) | ( n8898 & n8899 ) ;
  assign n8901 = ( ~n8564 & n8898 ) | ( ~n8564 & n8899 ) | ( n8898 & n8899 ) ;
  assign n8902 = ( n8564 & ~n8900 ) | ( n8564 & n8901 ) | ( ~n8900 & n8901 ) ;
  assign n8903 = ( ~n5905 & n8897 ) | ( ~n5905 & n8902 ) | ( n8897 & n8902 ) ;
  assign n8904 = ~n5905 & n8565 ;
  assign n8905 = ( ~n5905 & n8565 ) | ( ~n5905 & n8838 ) | ( n8565 & n8838 ) ;
  assign n8906 = ( ~n8570 & n8904 ) | ( ~n8570 & n8905 ) | ( n8904 & n8905 ) ;
  assign n8907 = ( n8570 & n8904 ) | ( n8570 & n8905 ) | ( n8904 & n8905 ) ;
  assign n8908 = ( n8570 & n8906 ) | ( n8570 & ~n8907 ) | ( n8906 & ~n8907 ) ;
  assign n8909 = ( ~n5642 & n8903 ) | ( ~n5642 & n8908 ) | ( n8903 & n8908 ) ;
  assign n8910 = ( n5642 & ~n8571 ) | ( n5642 & n8838 ) | ( ~n8571 & n8838 ) ;
  assign n8911 = n5642 & ~n8571 ;
  assign n8912 = ( n8576 & n8910 ) | ( n8576 & n8911 ) | ( n8910 & n8911 ) ;
  assign n8913 = ( ~n8576 & n8910 ) | ( ~n8576 & n8911 ) | ( n8910 & n8911 ) ;
  assign n8914 = ( n8576 & ~n8912 ) | ( n8576 & n8913 ) | ( ~n8912 & n8913 ) ;
  assign n8915 = ( ~n5386 & n8909 ) | ( ~n5386 & n8914 ) | ( n8909 & n8914 ) ;
  assign n8916 = ( n5386 & ~n8577 ) | ( n5386 & n8838 ) | ( ~n8577 & n8838 ) ;
  assign n8917 = n5386 & ~n8577 ;
  assign n8918 = ( n8582 & n8916 ) | ( n8582 & n8917 ) | ( n8916 & n8917 ) ;
  assign n8919 = ( ~n8582 & n8916 ) | ( ~n8582 & n8917 ) | ( n8916 & n8917 ) ;
  assign n8920 = ( n8582 & ~n8918 ) | ( n8582 & n8919 ) | ( ~n8918 & n8919 ) ;
  assign n8921 = ( ~n5139 & n8915 ) | ( ~n5139 & n8920 ) | ( n8915 & n8920 ) ;
  assign n8922 = ( n5139 & ~n8583 ) | ( n5139 & n8838 ) | ( ~n8583 & n8838 ) ;
  assign n8923 = n5139 & ~n8583 ;
  assign n8924 = ( n8588 & n8922 ) | ( n8588 & n8923 ) | ( n8922 & n8923 ) ;
  assign n8925 = ( ~n8588 & n8922 ) | ( ~n8588 & n8923 ) | ( n8922 & n8923 ) ;
  assign n8926 = ( n8588 & ~n8924 ) | ( n8588 & n8925 ) | ( ~n8924 & n8925 ) ;
  assign n8927 = ( ~n4898 & n8921 ) | ( ~n4898 & n8926 ) | ( n8921 & n8926 ) ;
  assign n8928 = ( n4898 & ~n8589 ) | ( n4898 & n8838 ) | ( ~n8589 & n8838 ) ;
  assign n8929 = n4898 & ~n8589 ;
  assign n8930 = ( n8594 & n8928 ) | ( n8594 & n8929 ) | ( n8928 & n8929 ) ;
  assign n8931 = ( ~n8594 & n8928 ) | ( ~n8594 & n8929 ) | ( n8928 & n8929 ) ;
  assign n8932 = ( n8594 & ~n8930 ) | ( n8594 & n8931 ) | ( ~n8930 & n8931 ) ;
  assign n8933 = ( ~n4661 & n8927 ) | ( ~n4661 & n8932 ) | ( n8927 & n8932 ) ;
  assign n8934 = ( n4661 & ~n8595 ) | ( n4661 & n8838 ) | ( ~n8595 & n8838 ) ;
  assign n8935 = n4661 & ~n8595 ;
  assign n8936 = ( n8600 & n8934 ) | ( n8600 & n8935 ) | ( n8934 & n8935 ) ;
  assign n8937 = ( ~n8600 & n8934 ) | ( ~n8600 & n8935 ) | ( n8934 & n8935 ) ;
  assign n8938 = ( n8600 & ~n8936 ) | ( n8600 & n8937 ) | ( ~n8936 & n8937 ) ;
  assign n8939 = ( ~n4432 & n8933 ) | ( ~n4432 & n8938 ) | ( n8933 & n8938 ) ;
  assign n8940 = ( n4432 & ~n8601 ) | ( n4432 & n8838 ) | ( ~n8601 & n8838 ) ;
  assign n8941 = n4432 & ~n8601 ;
  assign n8942 = ( n8606 & n8940 ) | ( n8606 & n8941 ) | ( n8940 & n8941 ) ;
  assign n8943 = ( ~n8606 & n8940 ) | ( ~n8606 & n8941 ) | ( n8940 & n8941 ) ;
  assign n8944 = ( n8606 & ~n8942 ) | ( n8606 & n8943 ) | ( ~n8942 & n8943 ) ;
  assign n8945 = ( ~n4203 & n8939 ) | ( ~n4203 & n8944 ) | ( n8939 & n8944 ) ;
  assign n8946 = ~n4203 & n8607 ;
  assign n8947 = ( ~n4203 & n8607 ) | ( ~n4203 & n8838 ) | ( n8607 & n8838 ) ;
  assign n8948 = ( n8612 & n8946 ) | ( n8612 & n8947 ) | ( n8946 & n8947 ) ;
  assign n8949 = ( ~n8612 & n8946 ) | ( ~n8612 & n8947 ) | ( n8946 & n8947 ) ;
  assign n8950 = ( n8612 & ~n8948 ) | ( n8612 & n8949 ) | ( ~n8948 & n8949 ) ;
  assign n8951 = ( ~n3985 & n8945 ) | ( ~n3985 & n8950 ) | ( n8945 & n8950 ) ;
  assign n8952 = ~n3985 & n8613 ;
  assign n8953 = ( ~n3985 & n8613 ) | ( ~n3985 & n8838 ) | ( n8613 & n8838 ) ;
  assign n8954 = ( ~n8618 & n8952 ) | ( ~n8618 & n8953 ) | ( n8952 & n8953 ) ;
  assign n8955 = ( n8618 & n8952 ) | ( n8618 & n8953 ) | ( n8952 & n8953 ) ;
  assign n8956 = ( n8618 & n8954 ) | ( n8618 & ~n8955 ) | ( n8954 & ~n8955 ) ;
  assign n8957 = ( ~n3772 & n8951 ) | ( ~n3772 & n8956 ) | ( n8951 & n8956 ) ;
  assign n8958 = n3772 & ~n8619 ;
  assign n8959 = ( n3772 & ~n8619 ) | ( n3772 & n8838 ) | ( ~n8619 & n8838 ) ;
  assign n8960 = ( n8624 & n8958 ) | ( n8624 & n8959 ) | ( n8958 & n8959 ) ;
  assign n8961 = ( ~n8624 & n8958 ) | ( ~n8624 & n8959 ) | ( n8958 & n8959 ) ;
  assign n8962 = ( n8624 & ~n8960 ) | ( n8624 & n8961 ) | ( ~n8960 & n8961 ) ;
  assign n8963 = ( ~n3567 & n8957 ) | ( ~n3567 & n8962 ) | ( n8957 & n8962 ) ;
  assign n8964 = ~n3567 & n8625 ;
  assign n8965 = ( ~n3567 & n8625 ) | ( ~n3567 & n8838 ) | ( n8625 & n8838 ) ;
  assign n8966 = ( ~n8630 & n8964 ) | ( ~n8630 & n8965 ) | ( n8964 & n8965 ) ;
  assign n8967 = ( n8630 & n8964 ) | ( n8630 & n8965 ) | ( n8964 & n8965 ) ;
  assign n8968 = ( n8630 & n8966 ) | ( n8630 & ~n8967 ) | ( n8966 & ~n8967 ) ;
  assign n8969 = ( ~n3362 & n8963 ) | ( ~n3362 & n8968 ) | ( n8963 & n8968 ) ;
  assign n8970 = n3362 & ~n8631 ;
  assign n8971 = ( n3362 & ~n8631 ) | ( n3362 & n8838 ) | ( ~n8631 & n8838 ) ;
  assign n8972 = ( n8636 & n8970 ) | ( n8636 & n8971 ) | ( n8970 & n8971 ) ;
  assign n8973 = ( ~n8636 & n8970 ) | ( ~n8636 & n8971 ) | ( n8970 & n8971 ) ;
  assign n8974 = ( n8636 & ~n8972 ) | ( n8636 & n8973 ) | ( ~n8972 & n8973 ) ;
  assign n8975 = ( ~n3169 & n8969 ) | ( ~n3169 & n8974 ) | ( n8969 & n8974 ) ;
  assign n8976 = ( n3169 & ~n8637 ) | ( n3169 & n8838 ) | ( ~n8637 & n8838 ) ;
  assign n8977 = n3169 & ~n8637 ;
  assign n8978 = ( n8642 & n8976 ) | ( n8642 & n8977 ) | ( n8976 & n8977 ) ;
  assign n8979 = ( ~n8642 & n8976 ) | ( ~n8642 & n8977 ) | ( n8976 & n8977 ) ;
  assign n8980 = ( n8642 & ~n8978 ) | ( n8642 & n8979 ) | ( ~n8978 & n8979 ) ;
  assign n8981 = ( ~n2979 & n8975 ) | ( ~n2979 & n8980 ) | ( n8975 & n8980 ) ;
  assign n8982 = ~n2979 & n8643 ;
  assign n8983 = ( ~n2979 & n8643 ) | ( ~n2979 & n8838 ) | ( n8643 & n8838 ) ;
  assign n8984 = ( ~n8648 & n8982 ) | ( ~n8648 & n8983 ) | ( n8982 & n8983 ) ;
  assign n8985 = ( n8648 & n8982 ) | ( n8648 & n8983 ) | ( n8982 & n8983 ) ;
  assign n8986 = ( n8648 & n8984 ) | ( n8648 & ~n8985 ) | ( n8984 & ~n8985 ) ;
  assign n8987 = ( ~n2791 & n8981 ) | ( ~n2791 & n8986 ) | ( n8981 & n8986 ) ;
  assign n8988 = ( n2791 & ~n8649 ) | ( n2791 & n8838 ) | ( ~n8649 & n8838 ) ;
  assign n8989 = n2791 & ~n8649 ;
  assign n8990 = ( n8654 & n8988 ) | ( n8654 & n8989 ) | ( n8988 & n8989 ) ;
  assign n8991 = ( ~n8654 & n8988 ) | ( ~n8654 & n8989 ) | ( n8988 & n8989 ) ;
  assign n8992 = ( n8654 & ~n8990 ) | ( n8654 & n8991 ) | ( ~n8990 & n8991 ) ;
  assign n8993 = ( ~n2615 & n8987 ) | ( ~n2615 & n8992 ) | ( n8987 & n8992 ) ;
  assign n8994 = ~n2615 & n8655 ;
  assign n8995 = ( ~n2615 & n8655 ) | ( ~n2615 & n8838 ) | ( n8655 & n8838 ) ;
  assign n8996 = ( ~n8660 & n8994 ) | ( ~n8660 & n8995 ) | ( n8994 & n8995 ) ;
  assign n8997 = ( n8660 & n8994 ) | ( n8660 & n8995 ) | ( n8994 & n8995 ) ;
  assign n8998 = ( n8660 & n8996 ) | ( n8660 & ~n8997 ) | ( n8996 & ~n8997 ) ;
  assign n8999 = ( ~n2443 & n8993 ) | ( ~n2443 & n8998 ) | ( n8993 & n8998 ) ;
  assign n9000 = ( n2443 & ~n8661 ) | ( n2443 & n8838 ) | ( ~n8661 & n8838 ) ;
  assign n9001 = n2443 & ~n8661 ;
  assign n9002 = ( n8666 & n9000 ) | ( n8666 & n9001 ) | ( n9000 & n9001 ) ;
  assign n9003 = ( ~n8666 & n9000 ) | ( ~n8666 & n9001 ) | ( n9000 & n9001 ) ;
  assign n9004 = ( n8666 & ~n9002 ) | ( n8666 & n9003 ) | ( ~n9002 & n9003 ) ;
  assign n9005 = ( ~n2277 & n8999 ) | ( ~n2277 & n9004 ) | ( n8999 & n9004 ) ;
  assign n9006 = ( n2277 & ~n8667 ) | ( n2277 & n8838 ) | ( ~n8667 & n8838 ) ;
  assign n9007 = n2277 & ~n8667 ;
  assign n9008 = ( n8672 & n9006 ) | ( n8672 & n9007 ) | ( n9006 & n9007 ) ;
  assign n9009 = ( ~n8672 & n9006 ) | ( ~n8672 & n9007 ) | ( n9006 & n9007 ) ;
  assign n9010 = ( n8672 & ~n9008 ) | ( n8672 & n9009 ) | ( ~n9008 & n9009 ) ;
  assign n9011 = ( ~n2111 & n9005 ) | ( ~n2111 & n9010 ) | ( n9005 & n9010 ) ;
  assign n9012 = ( n2111 & ~n8673 ) | ( n2111 & n8838 ) | ( ~n8673 & n8838 ) ;
  assign n9013 = n2111 & ~n8673 ;
  assign n9014 = ( n8678 & n9012 ) | ( n8678 & n9013 ) | ( n9012 & n9013 ) ;
  assign n9015 = ( ~n8678 & n9012 ) | ( ~n8678 & n9013 ) | ( n9012 & n9013 ) ;
  assign n9016 = ( n8678 & ~n9014 ) | ( n8678 & n9015 ) | ( ~n9014 & n9015 ) ;
  assign n9017 = ( ~n1949 & n9011 ) | ( ~n1949 & n9016 ) | ( n9011 & n9016 ) ;
  assign n9018 = ( n1949 & ~n8679 ) | ( n1949 & n8838 ) | ( ~n8679 & n8838 ) ;
  assign n9019 = n1949 & ~n8679 ;
  assign n9020 = ( n8684 & n9018 ) | ( n8684 & n9019 ) | ( n9018 & n9019 ) ;
  assign n9021 = ( ~n8684 & n9018 ) | ( ~n8684 & n9019 ) | ( n9018 & n9019 ) ;
  assign n9022 = ( n8684 & ~n9020 ) | ( n8684 & n9021 ) | ( ~n9020 & n9021 ) ;
  assign n9023 = ( ~n1802 & n9017 ) | ( ~n1802 & n9022 ) | ( n9017 & n9022 ) ;
  assign n9024 = n1802 & ~n8685 ;
  assign n9025 = ( n1802 & ~n8685 ) | ( n1802 & n8838 ) | ( ~n8685 & n8838 ) ;
  assign n9026 = ( n8690 & n9024 ) | ( n8690 & n9025 ) | ( n9024 & n9025 ) ;
  assign n9027 = ( ~n8690 & n9024 ) | ( ~n8690 & n9025 ) | ( n9024 & n9025 ) ;
  assign n9028 = ( n8690 & ~n9026 ) | ( n8690 & n9027 ) | ( ~n9026 & n9027 ) ;
  assign n9029 = ( ~n1661 & n9023 ) | ( ~n1661 & n9028 ) | ( n9023 & n9028 ) ;
  assign n9030 = ~n1661 & n8691 ;
  assign n9031 = ( ~n1661 & n8691 ) | ( ~n1661 & n8838 ) | ( n8691 & n8838 ) ;
  assign n9032 = ( ~n8696 & n9030 ) | ( ~n8696 & n9031 ) | ( n9030 & n9031 ) ;
  assign n9033 = ( n8696 & n9030 ) | ( n8696 & n9031 ) | ( n9030 & n9031 ) ;
  assign n9034 = ( n8696 & n9032 ) | ( n8696 & ~n9033 ) | ( n9032 & ~n9033 ) ;
  assign n9035 = ( ~n1523 & n9029 ) | ( ~n1523 & n9034 ) | ( n9029 & n9034 ) ;
  assign n9036 = ~n1523 & n8697 ;
  assign n9037 = ( ~n1523 & n8697 ) | ( ~n1523 & n8838 ) | ( n8697 & n8838 ) ;
  assign n9038 = ( ~n8702 & n9036 ) | ( ~n8702 & n9037 ) | ( n9036 & n9037 ) ;
  assign n9039 = ( n8702 & n9036 ) | ( n8702 & n9037 ) | ( n9036 & n9037 ) ;
  assign n9040 = ( n8702 & n9038 ) | ( n8702 & ~n9039 ) | ( n9038 & ~n9039 ) ;
  assign n9041 = ( ~n1393 & n9035 ) | ( ~n1393 & n9040 ) | ( n9035 & n9040 ) ;
  assign n9042 = ~n1393 & n8703 ;
  assign n9043 = ( ~n1393 & n8703 ) | ( ~n1393 & n8838 ) | ( n8703 & n8838 ) ;
  assign n9044 = ( n8708 & n9042 ) | ( n8708 & n9043 ) | ( n9042 & n9043 ) ;
  assign n9045 = ( ~n8708 & n9042 ) | ( ~n8708 & n9043 ) | ( n9042 & n9043 ) ;
  assign n9046 = ( n8708 & ~n9044 ) | ( n8708 & n9045 ) | ( ~n9044 & n9045 ) ;
  assign n9047 = ( ~n1266 & n9041 ) | ( ~n1266 & n9046 ) | ( n9041 & n9046 ) ;
  assign n9048 = ( n1266 & ~n8709 ) | ( n1266 & n8838 ) | ( ~n8709 & n8838 ) ;
  assign n9049 = n1266 & ~n8709 ;
  assign n9050 = ( n8714 & n9048 ) | ( n8714 & n9049 ) | ( n9048 & n9049 ) ;
  assign n9051 = ( ~n8714 & n9048 ) | ( ~n8714 & n9049 ) | ( n9048 & n9049 ) ;
  assign n9052 = ( n8714 & ~n9050 ) | ( n8714 & n9051 ) | ( ~n9050 & n9051 ) ;
  assign n9053 = ( ~n1150 & n9047 ) | ( ~n1150 & n9052 ) | ( n9047 & n9052 ) ;
  assign n9054 = ~n1150 & n8715 ;
  assign n9055 = ( ~n1150 & n8715 ) | ( ~n1150 & n8838 ) | ( n8715 & n8838 ) ;
  assign n9056 = ( n8720 & n9054 ) | ( n8720 & n9055 ) | ( n9054 & n9055 ) ;
  assign n9057 = ( ~n8720 & n9054 ) | ( ~n8720 & n9055 ) | ( n9054 & n9055 ) ;
  assign n9058 = ( n8720 & ~n9056 ) | ( n8720 & n9057 ) | ( ~n9056 & n9057 ) ;
  assign n9059 = ( ~n1038 & n9053 ) | ( ~n1038 & n9058 ) | ( n9053 & n9058 ) ;
  assign n9060 = ~n1038 & n8721 ;
  assign n9061 = ( ~n1038 & n8721 ) | ( ~n1038 & n8838 ) | ( n8721 & n8838 ) ;
  assign n9062 = ( ~n8726 & n9060 ) | ( ~n8726 & n9061 ) | ( n9060 & n9061 ) ;
  assign n9063 = ( n8726 & n9060 ) | ( n8726 & n9061 ) | ( n9060 & n9061 ) ;
  assign n9064 = ( n8726 & n9062 ) | ( n8726 & ~n9063 ) | ( n9062 & ~n9063 ) ;
  assign n9065 = ( ~n933 & n9059 ) | ( ~n933 & n9064 ) | ( n9059 & n9064 ) ;
  assign n9066 = ( n933 & ~n8727 ) | ( n933 & n8838 ) | ( ~n8727 & n8838 ) ;
  assign n9067 = n933 & ~n8727 ;
  assign n9068 = ( n8732 & n9066 ) | ( n8732 & n9067 ) | ( n9066 & n9067 ) ;
  assign n9069 = ( ~n8732 & n9066 ) | ( ~n8732 & n9067 ) | ( n9066 & n9067 ) ;
  assign n9070 = ( n8732 & ~n9068 ) | ( n8732 & n9069 ) | ( ~n9068 & n9069 ) ;
  assign n9071 = ( ~n839 & n9065 ) | ( ~n839 & n9070 ) | ( n9065 & n9070 ) ;
  assign n9072 = ( n839 & ~n8733 ) | ( n839 & n8838 ) | ( ~n8733 & n8838 ) ;
  assign n9073 = n839 & ~n8733 ;
  assign n9074 = ( n8738 & n9072 ) | ( n8738 & n9073 ) | ( n9072 & n9073 ) ;
  assign n9075 = ( ~n8738 & n9072 ) | ( ~n8738 & n9073 ) | ( n9072 & n9073 ) ;
  assign n9076 = ( n8738 & ~n9074 ) | ( n8738 & n9075 ) | ( ~n9074 & n9075 ) ;
  assign n9077 = ( ~n746 & n9071 ) | ( ~n746 & n9076 ) | ( n9071 & n9076 ) ;
  assign n9078 = ~n746 & n8739 ;
  assign n9079 = ( ~n746 & n8739 ) | ( ~n746 & n8838 ) | ( n8739 & n8838 ) ;
  assign n9080 = ( n8744 & n9078 ) | ( n8744 & n9079 ) | ( n9078 & n9079 ) ;
  assign n9081 = ( ~n8744 & n9078 ) | ( ~n8744 & n9079 ) | ( n9078 & n9079 ) ;
  assign n9082 = ( n8744 & ~n9080 ) | ( n8744 & n9081 ) | ( ~n9080 & n9081 ) ;
  assign n9083 = ( ~n664 & n9077 ) | ( ~n664 & n9082 ) | ( n9077 & n9082 ) ;
  assign n9084 = ~n664 & n8745 ;
  assign n9085 = ( ~n664 & n8745 ) | ( ~n664 & n8838 ) | ( n8745 & n8838 ) ;
  assign n9086 = ( n8750 & n9084 ) | ( n8750 & n9085 ) | ( n9084 & n9085 ) ;
  assign n9087 = ( ~n8750 & n9084 ) | ( ~n8750 & n9085 ) | ( n9084 & n9085 ) ;
  assign n9088 = ( n8750 & ~n9086 ) | ( n8750 & n9087 ) | ( ~n9086 & n9087 ) ;
  assign n9089 = ( ~n588 & n9083 ) | ( ~n588 & n9088 ) | ( n9083 & n9088 ) ;
  assign n9090 = ~n588 & n8751 ;
  assign n9091 = ( ~n588 & n8751 ) | ( ~n588 & n8838 ) | ( n8751 & n8838 ) ;
  assign n9092 = ( n8756 & n9090 ) | ( n8756 & n9091 ) | ( n9090 & n9091 ) ;
  assign n9093 = ( ~n8756 & n9090 ) | ( ~n8756 & n9091 ) | ( n9090 & n9091 ) ;
  assign n9094 = ( n8756 & ~n9092 ) | ( n8756 & n9093 ) | ( ~n9092 & n9093 ) ;
  assign n9095 = ( ~n518 & n9089 ) | ( ~n518 & n9094 ) | ( n9089 & n9094 ) ;
  assign n9096 = ( n518 & ~n8757 ) | ( n518 & n8838 ) | ( ~n8757 & n8838 ) ;
  assign n9097 = n518 & ~n8757 ;
  assign n9098 = ( n8762 & n9096 ) | ( n8762 & n9097 ) | ( n9096 & n9097 ) ;
  assign n9099 = ( ~n8762 & n9096 ) | ( ~n8762 & n9097 ) | ( n9096 & n9097 ) ;
  assign n9100 = ( n8762 & ~n9098 ) | ( n8762 & n9099 ) | ( ~n9098 & n9099 ) ;
  assign n9101 = ( ~n454 & n9095 ) | ( ~n454 & n9100 ) | ( n9095 & n9100 ) ;
  assign n9102 = ~n454 & n8763 ;
  assign n9103 = ( ~n454 & n8763 ) | ( ~n454 & n8838 ) | ( n8763 & n8838 ) ;
  assign n9104 = ( ~n8768 & n9102 ) | ( ~n8768 & n9103 ) | ( n9102 & n9103 ) ;
  assign n9105 = ( n8768 & n9102 ) | ( n8768 & n9103 ) | ( n9102 & n9103 ) ;
  assign n9106 = ( n8768 & n9104 ) | ( n8768 & ~n9105 ) | ( n9104 & ~n9105 ) ;
  assign n9107 = ( ~n396 & n9101 ) | ( ~n396 & n9106 ) | ( n9101 & n9106 ) ;
  assign n9108 = ~n396 & n8769 ;
  assign n9109 = ( ~n396 & n8769 ) | ( ~n396 & n8838 ) | ( n8769 & n8838 ) ;
  assign n9110 = ( ~n8774 & n9108 ) | ( ~n8774 & n9109 ) | ( n9108 & n9109 ) ;
  assign n9111 = ( n8774 & n9108 ) | ( n8774 & n9109 ) | ( n9108 & n9109 ) ;
  assign n9112 = ( n8774 & n9110 ) | ( n8774 & ~n9111 ) | ( n9110 & ~n9111 ) ;
  assign n9113 = ( ~n344 & n9107 ) | ( ~n344 & n9112 ) | ( n9107 & n9112 ) ;
  assign n9114 = ( n344 & ~n8775 ) | ( n344 & n8838 ) | ( ~n8775 & n8838 ) ;
  assign n9115 = n344 & ~n8775 ;
  assign n9116 = ( n8780 & n9114 ) | ( n8780 & n9115 ) | ( n9114 & n9115 ) ;
  assign n9117 = ( ~n8780 & n9114 ) | ( ~n8780 & n9115 ) | ( n9114 & n9115 ) ;
  assign n9118 = ( n8780 & ~n9116 ) | ( n8780 & n9117 ) | ( ~n9116 & n9117 ) ;
  assign n9119 = ( ~n298 & n9113 ) | ( ~n298 & n9118 ) | ( n9113 & n9118 ) ;
  assign n9120 = ( n298 & ~n8781 ) | ( n298 & n8838 ) | ( ~n8781 & n8838 ) ;
  assign n9121 = n298 & ~n8781 ;
  assign n9122 = ( n8786 & n9120 ) | ( n8786 & n9121 ) | ( n9120 & n9121 ) ;
  assign n9123 = ( ~n8786 & n9120 ) | ( ~n8786 & n9121 ) | ( n9120 & n9121 ) ;
  assign n9124 = ( n8786 & ~n9122 ) | ( n8786 & n9123 ) | ( ~n9122 & n9123 ) ;
  assign n9125 = ( ~n258 & n9119 ) | ( ~n258 & n9124 ) | ( n9119 & n9124 ) ;
  assign n9126 = n258 & ~n8787 ;
  assign n9127 = ( n258 & ~n8787 ) | ( n258 & n8838 ) | ( ~n8787 & n8838 ) ;
  assign n9128 = ( ~n8792 & n9126 ) | ( ~n8792 & n9127 ) | ( n9126 & n9127 ) ;
  assign n9129 = ( n8792 & n9126 ) | ( n8792 & n9127 ) | ( n9126 & n9127 ) ;
  assign n9130 = ( n8792 & n9128 ) | ( n8792 & ~n9129 ) | ( n9128 & ~n9129 ) ;
  assign n9131 = ( ~n225 & n9125 ) | ( ~n225 & n9130 ) | ( n9125 & n9130 ) ;
  assign n9132 = ( n225 & ~n8793 ) | ( n225 & n8838 ) | ( ~n8793 & n8838 ) ;
  assign n9133 = n225 & ~n8793 ;
  assign n9134 = ( n8798 & n9132 ) | ( n8798 & n9133 ) | ( n9132 & n9133 ) ;
  assign n9135 = ( ~n8798 & n9132 ) | ( ~n8798 & n9133 ) | ( n9132 & n9133 ) ;
  assign n9136 = ( n8798 & ~n9134 ) | ( n8798 & n9135 ) | ( ~n9134 & n9135 ) ;
  assign n9137 = ( ~n197 & n9131 ) | ( ~n197 & n9136 ) | ( n9131 & n9136 ) ;
  assign n9138 = ~n197 & n8799 ;
  assign n9139 = ( ~n197 & n8799 ) | ( ~n197 & n8838 ) | ( n8799 & n8838 ) ;
  assign n9140 = ( n8804 & n9138 ) | ( n8804 & n9139 ) | ( n9138 & n9139 ) ;
  assign n9141 = ( ~n8804 & n9138 ) | ( ~n8804 & n9139 ) | ( n9138 & n9139 ) ;
  assign n9142 = ( n8804 & ~n9140 ) | ( n8804 & n9141 ) | ( ~n9140 & n9141 ) ;
  assign n9143 = ( ~n170 & n9137 ) | ( ~n170 & n9142 ) | ( n9137 & n9142 ) ;
  assign n9144 = ~n170 & n8805 ;
  assign n9145 = ( ~n170 & n8805 ) | ( ~n170 & n8838 ) | ( n8805 & n8838 ) ;
  assign n9146 = ( ~n8810 & n9144 ) | ( ~n8810 & n9145 ) | ( n9144 & n9145 ) ;
  assign n9147 = ( n8810 & n9144 ) | ( n8810 & n9145 ) | ( n9144 & n9145 ) ;
  assign n9148 = ( n8810 & n9146 ) | ( n8810 & ~n9147 ) | ( n9146 & ~n9147 ) ;
  assign n9149 = ( ~n142 & n9143 ) | ( ~n142 & n9148 ) | ( n9143 & n9148 ) ;
  assign n9150 = ( n142 & ~n8811 ) | ( n142 & n8838 ) | ( ~n8811 & n8838 ) ;
  assign n9151 = n142 & ~n8811 ;
  assign n9152 = ( n8816 & n9150 ) | ( n8816 & n9151 ) | ( n9150 & n9151 ) ;
  assign n9153 = ( ~n8816 & n9150 ) | ( ~n8816 & n9151 ) | ( n9150 & n9151 ) ;
  assign n9154 = ( n8816 & ~n9152 ) | ( n8816 & n9153 ) | ( ~n9152 & n9153 ) ;
  assign n9155 = ( ~n132 & n9149 ) | ( ~n132 & n9154 ) | ( n9149 & n9154 ) ;
  assign n9156 = n8843 & n9155 ;
  assign n9157 = ( n8828 & ~n8830 ) | ( n8828 & n8834 ) | ( ~n8830 & n8834 ) ;
  assign n9158 = ( n8823 & n8828 ) | ( n8823 & n9157 ) | ( n8828 & n9157 ) ;
  assign n9159 = ~n8829 & n9158 ;
  assign n9160 = n9156 | n9159 ;
  assign n9161 = n8843 | n9155 ;
  assign n9162 = n8823 & n8828 ;
  assign n9163 = ~n8828 & n8837 ;
  assign n9164 = ~n8823 & n9163 ;
  assign n9165 = ( ~n9161 & n9162 ) | ( ~n9161 & n9164 ) | ( n9162 & n9164 ) ;
  assign n9166 = ( ~n131 & n9161 ) | ( ~n131 & n9165 ) | ( n9161 & n9165 ) ;
  assign n9167 = n9160 | n9166 ;
  assign n9168 = ( n132 & ~n9149 ) | ( n132 & n9167 ) | ( ~n9149 & n9167 ) ;
  assign n9169 = n132 & ~n9149 ;
  assign n9170 = ( n9154 & n9168 ) | ( n9154 & n9169 ) | ( n9168 & n9169 ) ;
  assign n9171 = ( n9154 & ~n9168 ) | ( n9154 & n9169 ) | ( ~n9168 & n9169 ) ;
  assign n9172 = ( n9168 & ~n9170 ) | ( n9168 & n9171 ) | ( ~n9170 & n9171 ) ;
  assign n9173 = ~n518 & n9089 ;
  assign n9174 = ( ~n518 & n9089 ) | ( ~n518 & n9167 ) | ( n9089 & n9167 ) ;
  assign n9175 = ( n9094 & n9173 ) | ( n9094 & n9174 ) | ( n9173 & n9174 ) ;
  assign n9176 = ( ~n9094 & n9173 ) | ( ~n9094 & n9174 ) | ( n9173 & n9174 ) ;
  assign n9177 = ( n9094 & ~n9175 ) | ( n9094 & n9176 ) | ( ~n9175 & n9176 ) ;
  assign n9178 = ~n8845 & n9167 ;
  assign n9179 = x16 | x17 ;
  assign n9180 = x18 | n9179 ;
  assign n9181 = n8838 & ~n9180 ;
  assign n9182 = ~n8838 & n9180 ;
  assign n9183 = ( x19 & ~n9167 ) | ( x19 & n9182 ) | ( ~n9167 & n9182 ) ;
  assign n9184 = ( n9178 & ~n9181 ) | ( n9178 & n9183 ) | ( ~n9181 & n9183 ) ;
  assign n9185 = n8838 & ~n9167 ;
  assign n9186 = ( x20 & n9178 ) | ( x20 & n9185 ) | ( n9178 & n9185 ) ;
  assign n9187 = ( ~x20 & n9178 ) | ( ~x20 & n9185 ) | ( n9178 & n9185 ) ;
  assign n9188 = ( x20 & ~n9186 ) | ( x20 & n9187 ) | ( ~n9186 & n9187 ) ;
  assign n9189 = ( ~n8517 & n9184 ) | ( ~n8517 & n9188 ) | ( n9184 & n9188 ) ;
  assign n9190 = ~n8517 & n8838 ;
  assign n9191 = ( n8851 & n9167 ) | ( n8851 & n9190 ) | ( n9167 & n9190 ) ;
  assign n9192 = ( x21 & n9187 ) | ( x21 & n9191 ) | ( n9187 & n9191 ) ;
  assign n9193 = ( ~x21 & n9187 ) | ( ~x21 & n9191 ) | ( n9187 & n9191 ) ;
  assign n9194 = ( x21 & ~n9192 ) | ( x21 & n9193 ) | ( ~n9192 & n9193 ) ;
  assign n9195 = ( ~n8201 & n9189 ) | ( ~n8201 & n9194 ) | ( n9189 & n9194 ) ;
  assign n9196 = ( n8201 & ~n8850 ) | ( n8201 & n9167 ) | ( ~n8850 & n9167 ) ;
  assign n9197 = n8201 & ~n8850 ;
  assign n9198 = ( n8854 & n9196 ) | ( n8854 & n9197 ) | ( n9196 & n9197 ) ;
  assign n9199 = ( ~n8854 & n9196 ) | ( ~n8854 & n9197 ) | ( n9196 & n9197 ) ;
  assign n9200 = ( n8854 & ~n9198 ) | ( n8854 & n9199 ) | ( ~n9198 & n9199 ) ;
  assign n9201 = ( ~n7897 & n9195 ) | ( ~n7897 & n9200 ) | ( n9195 & n9200 ) ;
  assign n9202 = ( n7897 & ~n8855 ) | ( n7897 & n9167 ) | ( ~n8855 & n9167 ) ;
  assign n9203 = n7897 & ~n8855 ;
  assign n9204 = ( n8860 & n9202 ) | ( n8860 & n9203 ) | ( n9202 & n9203 ) ;
  assign n9205 = ( ~n8860 & n9202 ) | ( ~n8860 & n9203 ) | ( n9202 & n9203 ) ;
  assign n9206 = ( n8860 & ~n9204 ) | ( n8860 & n9205 ) | ( ~n9204 & n9205 ) ;
  assign n9207 = ( ~n7594 & n9201 ) | ( ~n7594 & n9206 ) | ( n9201 & n9206 ) ;
  assign n9208 = ( n7594 & ~n8861 ) | ( n7594 & n9167 ) | ( ~n8861 & n9167 ) ;
  assign n9209 = n7594 & ~n8861 ;
  assign n9210 = ( n8866 & n9208 ) | ( n8866 & n9209 ) | ( n9208 & n9209 ) ;
  assign n9211 = ( ~n8866 & n9208 ) | ( ~n8866 & n9209 ) | ( n9208 & n9209 ) ;
  assign n9212 = ( n8866 & ~n9210 ) | ( n8866 & n9211 ) | ( ~n9210 & n9211 ) ;
  assign n9213 = ( ~n7296 & n9207 ) | ( ~n7296 & n9212 ) | ( n9207 & n9212 ) ;
  assign n9214 = ~n7296 & n8867 ;
  assign n9215 = ( ~n7296 & n8867 ) | ( ~n7296 & n9167 ) | ( n8867 & n9167 ) ;
  assign n9216 = ( ~n8872 & n9214 ) | ( ~n8872 & n9215 ) | ( n9214 & n9215 ) ;
  assign n9217 = ( n8872 & n9214 ) | ( n8872 & n9215 ) | ( n9214 & n9215 ) ;
  assign n9218 = ( n8872 & n9216 ) | ( n8872 & ~n9217 ) | ( n9216 & ~n9217 ) ;
  assign n9219 = ( ~n7006 & n9213 ) | ( ~n7006 & n9218 ) | ( n9213 & n9218 ) ;
  assign n9220 = ~n7006 & n8873 ;
  assign n9221 = ( ~n7006 & n8873 ) | ( ~n7006 & n9167 ) | ( n8873 & n9167 ) ;
  assign n9222 = ( n8878 & n9220 ) | ( n8878 & n9221 ) | ( n9220 & n9221 ) ;
  assign n9223 = ( ~n8878 & n9220 ) | ( ~n8878 & n9221 ) | ( n9220 & n9221 ) ;
  assign n9224 = ( n8878 & ~n9222 ) | ( n8878 & n9223 ) | ( ~n9222 & n9223 ) ;
  assign n9225 = ( ~n6723 & n9219 ) | ( ~n6723 & n9224 ) | ( n9219 & n9224 ) ;
  assign n9226 = ~n6723 & n8879 ;
  assign n9227 = ( ~n6723 & n8879 ) | ( ~n6723 & n9167 ) | ( n8879 & n9167 ) ;
  assign n9228 = ( ~n8884 & n9226 ) | ( ~n8884 & n9227 ) | ( n9226 & n9227 ) ;
  assign n9229 = ( n8884 & n9226 ) | ( n8884 & n9227 ) | ( n9226 & n9227 ) ;
  assign n9230 = ( n8884 & n9228 ) | ( n8884 & ~n9229 ) | ( n9228 & ~n9229 ) ;
  assign n9231 = ( ~n6442 & n9225 ) | ( ~n6442 & n9230 ) | ( n9225 & n9230 ) ;
  assign n9232 = ( n6442 & ~n8885 ) | ( n6442 & n9167 ) | ( ~n8885 & n9167 ) ;
  assign n9233 = n6442 & ~n8885 ;
  assign n9234 = ( n8890 & n9232 ) | ( n8890 & n9233 ) | ( n9232 & n9233 ) ;
  assign n9235 = ( ~n8890 & n9232 ) | ( ~n8890 & n9233 ) | ( n9232 & n9233 ) ;
  assign n9236 = ( n8890 & ~n9234 ) | ( n8890 & n9235 ) | ( ~n9234 & n9235 ) ;
  assign n9237 = ( ~n6172 & n9231 ) | ( ~n6172 & n9236 ) | ( n9231 & n9236 ) ;
  assign n9238 = ~n6172 & n8891 ;
  assign n9239 = ( ~n6172 & n8891 ) | ( ~n6172 & n9167 ) | ( n8891 & n9167 ) ;
  assign n9240 = ( ~n8896 & n9238 ) | ( ~n8896 & n9239 ) | ( n9238 & n9239 ) ;
  assign n9241 = ( n8896 & n9238 ) | ( n8896 & n9239 ) | ( n9238 & n9239 ) ;
  assign n9242 = ( n8896 & n9240 ) | ( n8896 & ~n9241 ) | ( n9240 & ~n9241 ) ;
  assign n9243 = ( ~n5905 & n9237 ) | ( ~n5905 & n9242 ) | ( n9237 & n9242 ) ;
  assign n9244 = ( n5905 & ~n8897 ) | ( n5905 & n9167 ) | ( ~n8897 & n9167 ) ;
  assign n9245 = n5905 & ~n8897 ;
  assign n9246 = ( n8902 & n9244 ) | ( n8902 & n9245 ) | ( n9244 & n9245 ) ;
  assign n9247 = ( ~n8902 & n9244 ) | ( ~n8902 & n9245 ) | ( n9244 & n9245 ) ;
  assign n9248 = ( n8902 & ~n9246 ) | ( n8902 & n9247 ) | ( ~n9246 & n9247 ) ;
  assign n9249 = ( ~n5642 & n9243 ) | ( ~n5642 & n9248 ) | ( n9243 & n9248 ) ;
  assign n9250 = n5642 & ~n8903 ;
  assign n9251 = ( n5642 & ~n8903 ) | ( n5642 & n9167 ) | ( ~n8903 & n9167 ) ;
  assign n9252 = ( ~n8908 & n9250 ) | ( ~n8908 & n9251 ) | ( n9250 & n9251 ) ;
  assign n9253 = ( n8908 & n9250 ) | ( n8908 & n9251 ) | ( n9250 & n9251 ) ;
  assign n9254 = ( n8908 & n9252 ) | ( n8908 & ~n9253 ) | ( n9252 & ~n9253 ) ;
  assign n9255 = ( ~n5386 & n9249 ) | ( ~n5386 & n9254 ) | ( n9249 & n9254 ) ;
  assign n9256 = ( n5386 & ~n8909 ) | ( n5386 & n9167 ) | ( ~n8909 & n9167 ) ;
  assign n9257 = n5386 & ~n8909 ;
  assign n9258 = ( n8914 & n9256 ) | ( n8914 & n9257 ) | ( n9256 & n9257 ) ;
  assign n9259 = ( ~n8914 & n9256 ) | ( ~n8914 & n9257 ) | ( n9256 & n9257 ) ;
  assign n9260 = ( n8914 & ~n9258 ) | ( n8914 & n9259 ) | ( ~n9258 & n9259 ) ;
  assign n9261 = ( ~n5139 & n9255 ) | ( ~n5139 & n9260 ) | ( n9255 & n9260 ) ;
  assign n9262 = n5139 & ~n8915 ;
  assign n9263 = ( n5139 & ~n8915 ) | ( n5139 & n9167 ) | ( ~n8915 & n9167 ) ;
  assign n9264 = ( ~n8920 & n9262 ) | ( ~n8920 & n9263 ) | ( n9262 & n9263 ) ;
  assign n9265 = ( n8920 & n9262 ) | ( n8920 & n9263 ) | ( n9262 & n9263 ) ;
  assign n9266 = ( n8920 & n9264 ) | ( n8920 & ~n9265 ) | ( n9264 & ~n9265 ) ;
  assign n9267 = ( ~n4898 & n9261 ) | ( ~n4898 & n9266 ) | ( n9261 & n9266 ) ;
  assign n9268 = ( n4898 & ~n8921 ) | ( n4898 & n9167 ) | ( ~n8921 & n9167 ) ;
  assign n9269 = n4898 & ~n8921 ;
  assign n9270 = ( n8926 & n9268 ) | ( n8926 & n9269 ) | ( n9268 & n9269 ) ;
  assign n9271 = ( ~n8926 & n9268 ) | ( ~n8926 & n9269 ) | ( n9268 & n9269 ) ;
  assign n9272 = ( n8926 & ~n9270 ) | ( n8926 & n9271 ) | ( ~n9270 & n9271 ) ;
  assign n9273 = ( ~n4661 & n9267 ) | ( ~n4661 & n9272 ) | ( n9267 & n9272 ) ;
  assign n9274 = ( n4661 & ~n8927 ) | ( n4661 & n9167 ) | ( ~n8927 & n9167 ) ;
  assign n9275 = n4661 & ~n8927 ;
  assign n9276 = ( n8932 & n9274 ) | ( n8932 & n9275 ) | ( n9274 & n9275 ) ;
  assign n9277 = ( ~n8932 & n9274 ) | ( ~n8932 & n9275 ) | ( n9274 & n9275 ) ;
  assign n9278 = ( n8932 & ~n9276 ) | ( n8932 & n9277 ) | ( ~n9276 & n9277 ) ;
  assign n9279 = ( ~n4432 & n9273 ) | ( ~n4432 & n9278 ) | ( n9273 & n9278 ) ;
  assign n9280 = ( n4432 & ~n8933 ) | ( n4432 & n9167 ) | ( ~n8933 & n9167 ) ;
  assign n9281 = n4432 & ~n8933 ;
  assign n9282 = ( n8938 & n9280 ) | ( n8938 & n9281 ) | ( n9280 & n9281 ) ;
  assign n9283 = ( ~n8938 & n9280 ) | ( ~n8938 & n9281 ) | ( n9280 & n9281 ) ;
  assign n9284 = ( n8938 & ~n9282 ) | ( n8938 & n9283 ) | ( ~n9282 & n9283 ) ;
  assign n9285 = ( ~n4203 & n9279 ) | ( ~n4203 & n9284 ) | ( n9279 & n9284 ) ;
  assign n9286 = ~n4203 & n8939 ;
  assign n9287 = ( ~n4203 & n8939 ) | ( ~n4203 & n9167 ) | ( n8939 & n9167 ) ;
  assign n9288 = ( ~n8944 & n9286 ) | ( ~n8944 & n9287 ) | ( n9286 & n9287 ) ;
  assign n9289 = ( n8944 & n9286 ) | ( n8944 & n9287 ) | ( n9286 & n9287 ) ;
  assign n9290 = ( n8944 & n9288 ) | ( n8944 & ~n9289 ) | ( n9288 & ~n9289 ) ;
  assign n9291 = ( ~n3985 & n9285 ) | ( ~n3985 & n9290 ) | ( n9285 & n9290 ) ;
  assign n9292 = ( n3985 & ~n8945 ) | ( n3985 & n9167 ) | ( ~n8945 & n9167 ) ;
  assign n9293 = n3985 & ~n8945 ;
  assign n9294 = ( n8950 & n9292 ) | ( n8950 & n9293 ) | ( n9292 & n9293 ) ;
  assign n9295 = ( ~n8950 & n9292 ) | ( ~n8950 & n9293 ) | ( n9292 & n9293 ) ;
  assign n9296 = ( n8950 & ~n9294 ) | ( n8950 & n9295 ) | ( ~n9294 & n9295 ) ;
  assign n9297 = ( ~n3772 & n9291 ) | ( ~n3772 & n9296 ) | ( n9291 & n9296 ) ;
  assign n9298 = ~n3772 & n8951 ;
  assign n9299 = ( ~n3772 & n8951 ) | ( ~n3772 & n9167 ) | ( n8951 & n9167 ) ;
  assign n9300 = ( ~n8956 & n9298 ) | ( ~n8956 & n9299 ) | ( n9298 & n9299 ) ;
  assign n9301 = ( n8956 & n9298 ) | ( n8956 & n9299 ) | ( n9298 & n9299 ) ;
  assign n9302 = ( n8956 & n9300 ) | ( n8956 & ~n9301 ) | ( n9300 & ~n9301 ) ;
  assign n9303 = ( ~n3567 & n9297 ) | ( ~n3567 & n9302 ) | ( n9297 & n9302 ) ;
  assign n9304 = ( n3567 & ~n8957 ) | ( n3567 & n9167 ) | ( ~n8957 & n9167 ) ;
  assign n9305 = n3567 & ~n8957 ;
  assign n9306 = ( n8962 & n9304 ) | ( n8962 & n9305 ) | ( n9304 & n9305 ) ;
  assign n9307 = ( ~n8962 & n9304 ) | ( ~n8962 & n9305 ) | ( n9304 & n9305 ) ;
  assign n9308 = ( n8962 & ~n9306 ) | ( n8962 & n9307 ) | ( ~n9306 & n9307 ) ;
  assign n9309 = ( ~n3362 & n9303 ) | ( ~n3362 & n9308 ) | ( n9303 & n9308 ) ;
  assign n9310 = ( n3362 & ~n8963 ) | ( n3362 & n9167 ) | ( ~n8963 & n9167 ) ;
  assign n9311 = n3362 & ~n8963 ;
  assign n9312 = ( n8968 & n9310 ) | ( n8968 & n9311 ) | ( n9310 & n9311 ) ;
  assign n9313 = ( ~n8968 & n9310 ) | ( ~n8968 & n9311 ) | ( n9310 & n9311 ) ;
  assign n9314 = ( n8968 & ~n9312 ) | ( n8968 & n9313 ) | ( ~n9312 & n9313 ) ;
  assign n9315 = ( ~n3169 & n9309 ) | ( ~n3169 & n9314 ) | ( n9309 & n9314 ) ;
  assign n9316 = ( n3169 & ~n8969 ) | ( n3169 & n9167 ) | ( ~n8969 & n9167 ) ;
  assign n9317 = n3169 & ~n8969 ;
  assign n9318 = ( n8974 & n9316 ) | ( n8974 & n9317 ) | ( n9316 & n9317 ) ;
  assign n9319 = ( ~n8974 & n9316 ) | ( ~n8974 & n9317 ) | ( n9316 & n9317 ) ;
  assign n9320 = ( n8974 & ~n9318 ) | ( n8974 & n9319 ) | ( ~n9318 & n9319 ) ;
  assign n9321 = ( ~n2979 & n9315 ) | ( ~n2979 & n9320 ) | ( n9315 & n9320 ) ;
  assign n9322 = ~n2979 & n8975 ;
  assign n9323 = ( ~n2979 & n8975 ) | ( ~n2979 & n9167 ) | ( n8975 & n9167 ) ;
  assign n9324 = ( n8980 & n9322 ) | ( n8980 & n9323 ) | ( n9322 & n9323 ) ;
  assign n9325 = ( ~n8980 & n9322 ) | ( ~n8980 & n9323 ) | ( n9322 & n9323 ) ;
  assign n9326 = ( n8980 & ~n9324 ) | ( n8980 & n9325 ) | ( ~n9324 & n9325 ) ;
  assign n9327 = ( ~n2791 & n9321 ) | ( ~n2791 & n9326 ) | ( n9321 & n9326 ) ;
  assign n9328 = n2791 & ~n8981 ;
  assign n9329 = ( n2791 & ~n8981 ) | ( n2791 & n9167 ) | ( ~n8981 & n9167 ) ;
  assign n9330 = ( ~n8986 & n9328 ) | ( ~n8986 & n9329 ) | ( n9328 & n9329 ) ;
  assign n9331 = ( n8986 & n9328 ) | ( n8986 & n9329 ) | ( n9328 & n9329 ) ;
  assign n9332 = ( n8986 & n9330 ) | ( n8986 & ~n9331 ) | ( n9330 & ~n9331 ) ;
  assign n9333 = ( ~n2615 & n9327 ) | ( ~n2615 & n9332 ) | ( n9327 & n9332 ) ;
  assign n9334 = ~n2615 & n8987 ;
  assign n9335 = ( ~n2615 & n8987 ) | ( ~n2615 & n9167 ) | ( n8987 & n9167 ) ;
  assign n9336 = ( ~n8992 & n9334 ) | ( ~n8992 & n9335 ) | ( n9334 & n9335 ) ;
  assign n9337 = ( n8992 & n9334 ) | ( n8992 & n9335 ) | ( n9334 & n9335 ) ;
  assign n9338 = ( n8992 & n9336 ) | ( n8992 & ~n9337 ) | ( n9336 & ~n9337 ) ;
  assign n9339 = ( ~n2443 & n9333 ) | ( ~n2443 & n9338 ) | ( n9333 & n9338 ) ;
  assign n9340 = ( n2443 & ~n8993 ) | ( n2443 & n9167 ) | ( ~n8993 & n9167 ) ;
  assign n9341 = n2443 & ~n8993 ;
  assign n9342 = ( n8998 & n9340 ) | ( n8998 & n9341 ) | ( n9340 & n9341 ) ;
  assign n9343 = ( ~n8998 & n9340 ) | ( ~n8998 & n9341 ) | ( n9340 & n9341 ) ;
  assign n9344 = ( n8998 & ~n9342 ) | ( n8998 & n9343 ) | ( ~n9342 & n9343 ) ;
  assign n9345 = ( ~n2277 & n9339 ) | ( ~n2277 & n9344 ) | ( n9339 & n9344 ) ;
  assign n9346 = ( n2277 & ~n8999 ) | ( n2277 & n9167 ) | ( ~n8999 & n9167 ) ;
  assign n9347 = n2277 & ~n8999 ;
  assign n9348 = ( n9004 & n9346 ) | ( n9004 & n9347 ) | ( n9346 & n9347 ) ;
  assign n9349 = ( ~n9004 & n9346 ) | ( ~n9004 & n9347 ) | ( n9346 & n9347 ) ;
  assign n9350 = ( n9004 & ~n9348 ) | ( n9004 & n9349 ) | ( ~n9348 & n9349 ) ;
  assign n9351 = ( ~n2111 & n9345 ) | ( ~n2111 & n9350 ) | ( n9345 & n9350 ) ;
  assign n9352 = ~n2111 & n9005 ;
  assign n9353 = ( ~n2111 & n9005 ) | ( ~n2111 & n9167 ) | ( n9005 & n9167 ) ;
  assign n9354 = ( n9010 & n9352 ) | ( n9010 & n9353 ) | ( n9352 & n9353 ) ;
  assign n9355 = ( ~n9010 & n9352 ) | ( ~n9010 & n9353 ) | ( n9352 & n9353 ) ;
  assign n9356 = ( n9010 & ~n9354 ) | ( n9010 & n9355 ) | ( ~n9354 & n9355 ) ;
  assign n9357 = ( ~n1949 & n9351 ) | ( ~n1949 & n9356 ) | ( n9351 & n9356 ) ;
  assign n9358 = ~n1949 & n9011 ;
  assign n9359 = ( ~n1949 & n9011 ) | ( ~n1949 & n9167 ) | ( n9011 & n9167 ) ;
  assign n9360 = ( ~n9016 & n9358 ) | ( ~n9016 & n9359 ) | ( n9358 & n9359 ) ;
  assign n9361 = ( n9016 & n9358 ) | ( n9016 & n9359 ) | ( n9358 & n9359 ) ;
  assign n9362 = ( n9016 & n9360 ) | ( n9016 & ~n9361 ) | ( n9360 & ~n9361 ) ;
  assign n9363 = ( ~n1802 & n9357 ) | ( ~n1802 & n9362 ) | ( n9357 & n9362 ) ;
  assign n9364 = ( n1802 & ~n9017 ) | ( n1802 & n9167 ) | ( ~n9017 & n9167 ) ;
  assign n9365 = n1802 & ~n9017 ;
  assign n9366 = ( n9022 & n9364 ) | ( n9022 & n9365 ) | ( n9364 & n9365 ) ;
  assign n9367 = ( ~n9022 & n9364 ) | ( ~n9022 & n9365 ) | ( n9364 & n9365 ) ;
  assign n9368 = ( n9022 & ~n9366 ) | ( n9022 & n9367 ) | ( ~n9366 & n9367 ) ;
  assign n9369 = ( ~n1661 & n9363 ) | ( ~n1661 & n9368 ) | ( n9363 & n9368 ) ;
  assign n9370 = ( n1661 & ~n9023 ) | ( n1661 & n9167 ) | ( ~n9023 & n9167 ) ;
  assign n9371 = n1661 & ~n9023 ;
  assign n9372 = ( n9028 & n9370 ) | ( n9028 & n9371 ) | ( n9370 & n9371 ) ;
  assign n9373 = ( ~n9028 & n9370 ) | ( ~n9028 & n9371 ) | ( n9370 & n9371 ) ;
  assign n9374 = ( n9028 & ~n9372 ) | ( n9028 & n9373 ) | ( ~n9372 & n9373 ) ;
  assign n9375 = ( ~n1523 & n9369 ) | ( ~n1523 & n9374 ) | ( n9369 & n9374 ) ;
  assign n9376 = ~n1523 & n9029 ;
  assign n9377 = ( ~n1523 & n9029 ) | ( ~n1523 & n9167 ) | ( n9029 & n9167 ) ;
  assign n9378 = ( ~n9034 & n9376 ) | ( ~n9034 & n9377 ) | ( n9376 & n9377 ) ;
  assign n9379 = ( n9034 & n9376 ) | ( n9034 & n9377 ) | ( n9376 & n9377 ) ;
  assign n9380 = ( n9034 & n9378 ) | ( n9034 & ~n9379 ) | ( n9378 & ~n9379 ) ;
  assign n9381 = ( ~n1393 & n9375 ) | ( ~n1393 & n9380 ) | ( n9375 & n9380 ) ;
  assign n9382 = n1393 & ~n9035 ;
  assign n9383 = ( n1393 & ~n9035 ) | ( n1393 & n9167 ) | ( ~n9035 & n9167 ) ;
  assign n9384 = ( n9040 & n9382 ) | ( n9040 & n9383 ) | ( n9382 & n9383 ) ;
  assign n9385 = ( ~n9040 & n9382 ) | ( ~n9040 & n9383 ) | ( n9382 & n9383 ) ;
  assign n9386 = ( n9040 & ~n9384 ) | ( n9040 & n9385 ) | ( ~n9384 & n9385 ) ;
  assign n9387 = ( ~n1266 & n9381 ) | ( ~n1266 & n9386 ) | ( n9381 & n9386 ) ;
  assign n9388 = ~n1266 & n9041 ;
  assign n9389 = ( ~n1266 & n9041 ) | ( ~n1266 & n9167 ) | ( n9041 & n9167 ) ;
  assign n9390 = ( n9046 & n9388 ) | ( n9046 & n9389 ) | ( n9388 & n9389 ) ;
  assign n9391 = ( ~n9046 & n9388 ) | ( ~n9046 & n9389 ) | ( n9388 & n9389 ) ;
  assign n9392 = ( n9046 & ~n9390 ) | ( n9046 & n9391 ) | ( ~n9390 & n9391 ) ;
  assign n9393 = ( ~n1150 & n9387 ) | ( ~n1150 & n9392 ) | ( n9387 & n9392 ) ;
  assign n9394 = n1150 & ~n9047 ;
  assign n9395 = ( n1150 & ~n9047 ) | ( n1150 & n9167 ) | ( ~n9047 & n9167 ) ;
  assign n9396 = ( n9052 & n9394 ) | ( n9052 & n9395 ) | ( n9394 & n9395 ) ;
  assign n9397 = ( ~n9052 & n9394 ) | ( ~n9052 & n9395 ) | ( n9394 & n9395 ) ;
  assign n9398 = ( n9052 & ~n9396 ) | ( n9052 & n9397 ) | ( ~n9396 & n9397 ) ;
  assign n9399 = ( ~n1038 & n9393 ) | ( ~n1038 & n9398 ) | ( n9393 & n9398 ) ;
  assign n9400 = ( n1038 & ~n9053 ) | ( n1038 & n9167 ) | ( ~n9053 & n9167 ) ;
  assign n9401 = n1038 & ~n9053 ;
  assign n9402 = ( n9058 & n9400 ) | ( n9058 & n9401 ) | ( n9400 & n9401 ) ;
  assign n9403 = ( ~n9058 & n9400 ) | ( ~n9058 & n9401 ) | ( n9400 & n9401 ) ;
  assign n9404 = ( n9058 & ~n9402 ) | ( n9058 & n9403 ) | ( ~n9402 & n9403 ) ;
  assign n9405 = ( ~n933 & n9399 ) | ( ~n933 & n9404 ) | ( n9399 & n9404 ) ;
  assign n9406 = ~n933 & n9059 ;
  assign n9407 = ( ~n933 & n9059 ) | ( ~n933 & n9167 ) | ( n9059 & n9167 ) ;
  assign n9408 = ( ~n9064 & n9406 ) | ( ~n9064 & n9407 ) | ( n9406 & n9407 ) ;
  assign n9409 = ( n9064 & n9406 ) | ( n9064 & n9407 ) | ( n9406 & n9407 ) ;
  assign n9410 = ( n9064 & n9408 ) | ( n9064 & ~n9409 ) | ( n9408 & ~n9409 ) ;
  assign n9411 = ( ~n839 & n9405 ) | ( ~n839 & n9410 ) | ( n9405 & n9410 ) ;
  assign n9412 = ( ~n839 & n9065 ) | ( ~n839 & n9167 ) | ( n9065 & n9167 ) ;
  assign n9413 = ~n839 & n9065 ;
  assign n9414 = ( ~n9070 & n9412 ) | ( ~n9070 & n9413 ) | ( n9412 & n9413 ) ;
  assign n9415 = ( n9070 & n9412 ) | ( n9070 & n9413 ) | ( n9412 & n9413 ) ;
  assign n9416 = ( n9070 & n9414 ) | ( n9070 & ~n9415 ) | ( n9414 & ~n9415 ) ;
  assign n9417 = ( ~n746 & n9411 ) | ( ~n746 & n9416 ) | ( n9411 & n9416 ) ;
  assign n9418 = n746 & ~n9071 ;
  assign n9419 = ( n746 & ~n9071 ) | ( n746 & n9167 ) | ( ~n9071 & n9167 ) ;
  assign n9420 = ( n9076 & n9418 ) | ( n9076 & n9419 ) | ( n9418 & n9419 ) ;
  assign n9421 = ( ~n9076 & n9418 ) | ( ~n9076 & n9419 ) | ( n9418 & n9419 ) ;
  assign n9422 = ( n9076 & ~n9420 ) | ( n9076 & n9421 ) | ( ~n9420 & n9421 ) ;
  assign n9423 = ( ~n664 & n9417 ) | ( ~n664 & n9422 ) | ( n9417 & n9422 ) ;
  assign n9424 = ( n664 & ~n9077 ) | ( n664 & n9167 ) | ( ~n9077 & n9167 ) ;
  assign n9425 = n664 & ~n9077 ;
  assign n9426 = ( n9082 & n9424 ) | ( n9082 & n9425 ) | ( n9424 & n9425 ) ;
  assign n9427 = ( ~n9082 & n9424 ) | ( ~n9082 & n9425 ) | ( n9424 & n9425 ) ;
  assign n9428 = ( n9082 & ~n9426 ) | ( n9082 & n9427 ) | ( ~n9426 & n9427 ) ;
  assign n9429 = ( ~n588 & n9423 ) | ( ~n588 & n9428 ) | ( n9423 & n9428 ) ;
  assign n9430 = ~n588 & n9083 ;
  assign n9431 = ( ~n588 & n9083 ) | ( ~n588 & n9167 ) | ( n9083 & n9167 ) ;
  assign n9432 = ( ~n9088 & n9430 ) | ( ~n9088 & n9431 ) | ( n9430 & n9431 ) ;
  assign n9433 = ( n9088 & n9430 ) | ( n9088 & n9431 ) | ( n9430 & n9431 ) ;
  assign n9434 = ( n9088 & n9432 ) | ( n9088 & ~n9433 ) | ( n9432 & ~n9433 ) ;
  assign n9435 = ( ~n518 & n9429 ) | ( ~n518 & n9434 ) | ( n9429 & n9434 ) ;
  assign n9436 = ( ~n454 & n9177 ) | ( ~n454 & n9435 ) | ( n9177 & n9435 ) ;
  assign n9437 = ( n454 & ~n9095 ) | ( n454 & n9167 ) | ( ~n9095 & n9167 ) ;
  assign n9438 = n454 & ~n9095 ;
  assign n9439 = ( n9100 & n9437 ) | ( n9100 & n9438 ) | ( n9437 & n9438 ) ;
  assign n9440 = ( ~n9100 & n9437 ) | ( ~n9100 & n9438 ) | ( n9437 & n9438 ) ;
  assign n9441 = ( n9100 & ~n9439 ) | ( n9100 & n9440 ) | ( ~n9439 & n9440 ) ;
  assign n9442 = ( ~n396 & n9436 ) | ( ~n396 & n9441 ) | ( n9436 & n9441 ) ;
  assign n9443 = ( n396 & ~n9101 ) | ( n396 & n9167 ) | ( ~n9101 & n9167 ) ;
  assign n9444 = n396 & ~n9101 ;
  assign n9445 = ( n9106 & n9443 ) | ( n9106 & n9444 ) | ( n9443 & n9444 ) ;
  assign n9446 = ( ~n9106 & n9443 ) | ( ~n9106 & n9444 ) | ( n9443 & n9444 ) ;
  assign n9447 = ( n9106 & ~n9445 ) | ( n9106 & n9446 ) | ( ~n9445 & n9446 ) ;
  assign n9448 = ( ~n344 & n9442 ) | ( ~n344 & n9447 ) | ( n9442 & n9447 ) ;
  assign n9449 = ( n344 & ~n9107 ) | ( n344 & n9167 ) | ( ~n9107 & n9167 ) ;
  assign n9450 = n344 & ~n9107 ;
  assign n9451 = ( n9112 & n9449 ) | ( n9112 & n9450 ) | ( n9449 & n9450 ) ;
  assign n9452 = ( ~n9112 & n9449 ) | ( ~n9112 & n9450 ) | ( n9449 & n9450 ) ;
  assign n9453 = ( n9112 & ~n9451 ) | ( n9112 & n9452 ) | ( ~n9451 & n9452 ) ;
  assign n9454 = ( ~n298 & n9448 ) | ( ~n298 & n9453 ) | ( n9448 & n9453 ) ;
  assign n9455 = ( n298 & ~n9113 ) | ( n298 & n9167 ) | ( ~n9113 & n9167 ) ;
  assign n9456 = n298 & ~n9113 ;
  assign n9457 = ( n9118 & n9455 ) | ( n9118 & n9456 ) | ( n9455 & n9456 ) ;
  assign n9458 = ( ~n9118 & n9455 ) | ( ~n9118 & n9456 ) | ( n9455 & n9456 ) ;
  assign n9459 = ( n9118 & ~n9457 ) | ( n9118 & n9458 ) | ( ~n9457 & n9458 ) ;
  assign n9460 = ( ~n258 & n9454 ) | ( ~n258 & n9459 ) | ( n9454 & n9459 ) ;
  assign n9461 = ( n258 & ~n9119 ) | ( n258 & n9167 ) | ( ~n9119 & n9167 ) ;
  assign n9462 = n258 & ~n9119 ;
  assign n9463 = ( n9124 & n9461 ) | ( n9124 & n9462 ) | ( n9461 & n9462 ) ;
  assign n9464 = ( ~n9124 & n9461 ) | ( ~n9124 & n9462 ) | ( n9461 & n9462 ) ;
  assign n9465 = ( n9124 & ~n9463 ) | ( n9124 & n9464 ) | ( ~n9463 & n9464 ) ;
  assign n9466 = ( ~n225 & n9460 ) | ( ~n225 & n9465 ) | ( n9460 & n9465 ) ;
  assign n9467 = ~n225 & n9125 ;
  assign n9468 = ( ~n225 & n9125 ) | ( ~n225 & n9167 ) | ( n9125 & n9167 ) ;
  assign n9469 = ( ~n9130 & n9467 ) | ( ~n9130 & n9468 ) | ( n9467 & n9468 ) ;
  assign n9470 = ( n9130 & n9467 ) | ( n9130 & n9468 ) | ( n9467 & n9468 ) ;
  assign n9471 = ( n9130 & n9469 ) | ( n9130 & ~n9470 ) | ( n9469 & ~n9470 ) ;
  assign n9472 = ( ~n197 & n9466 ) | ( ~n197 & n9471 ) | ( n9466 & n9471 ) ;
  assign n9473 = ~n197 & n9131 ;
  assign n9474 = ( ~n197 & n9131 ) | ( ~n197 & n9167 ) | ( n9131 & n9167 ) ;
  assign n9475 = ( ~n9136 & n9473 ) | ( ~n9136 & n9474 ) | ( n9473 & n9474 ) ;
  assign n9476 = ( n9136 & n9473 ) | ( n9136 & n9474 ) | ( n9473 & n9474 ) ;
  assign n9477 = ( n9136 & n9475 ) | ( n9136 & ~n9476 ) | ( n9475 & ~n9476 ) ;
  assign n9478 = ( ~n170 & n9472 ) | ( ~n170 & n9477 ) | ( n9472 & n9477 ) ;
  assign n9479 = ( n170 & ~n9137 ) | ( n170 & n9167 ) | ( ~n9137 & n9167 ) ;
  assign n9480 = n170 & ~n9137 ;
  assign n9481 = ( n9142 & n9479 ) | ( n9142 & n9480 ) | ( n9479 & n9480 ) ;
  assign n9482 = ( ~n9142 & n9479 ) | ( ~n9142 & n9480 ) | ( n9479 & n9480 ) ;
  assign n9483 = ( n9142 & ~n9481 ) | ( n9142 & n9482 ) | ( ~n9481 & n9482 ) ;
  assign n9484 = ( ~n142 & n9478 ) | ( ~n142 & n9483 ) | ( n9478 & n9483 ) ;
  assign n9485 = ( n142 & ~n9143 ) | ( n142 & n9167 ) | ( ~n9143 & n9167 ) ;
  assign n9486 = n142 & ~n9143 ;
  assign n9487 = ( n9148 & n9485 ) | ( n9148 & n9486 ) | ( n9485 & n9486 ) ;
  assign n9488 = ( ~n9148 & n9485 ) | ( ~n9148 & n9486 ) | ( n9485 & n9486 ) ;
  assign n9489 = ( n9148 & ~n9487 ) | ( n9148 & n9488 ) | ( ~n9487 & n9488 ) ;
  assign n9490 = ( ~n132 & n9484 ) | ( ~n132 & n9489 ) | ( n9484 & n9489 ) ;
  assign n9491 = ( ~n131 & n9172 ) | ( ~n131 & n9490 ) | ( n9172 & n9490 ) ;
  assign n9492 = ~n8843 & n9159 ;
  assign n9493 = ( n131 & ~n9155 ) | ( n131 & n9492 ) | ( ~n9155 & n9492 ) ;
  assign n9494 = n9161 & n9493 ;
  assign n9495 = ( ~n131 & n9156 ) | ( ~n131 & n9165 ) | ( n9156 & n9165 ) ;
  assign n9496 = n9494 | n9495 ;
  assign n9497 = n9491 | n9496 ;
  assign n9498 = ( n131 & ~n9172 ) | ( n131 & n9490 ) | ( ~n9172 & n9490 ) ;
  assign n9499 = ( n9160 & n9165 ) | ( n9160 & ~n9172 ) | ( n9165 & ~n9172 ) ;
  assign n9500 = ( ~n9172 & n9490 ) | ( ~n9172 & n9499 ) | ( n9490 & n9499 ) ;
  assign n9501 = ( n131 & n9172 ) | ( n131 & n9494 ) | ( n9172 & n9494 ) ;
  assign n9502 = ( n9172 & n9490 ) | ( n9172 & n9501 ) | ( n9490 & n9501 ) ;
  assign n9503 = ( ~n9498 & n9500 ) | ( ~n9498 & n9502 ) | ( n9500 & n9502 ) ;
  assign n9504 = x14 | x15 ;
  assign n9505 = x16 | n9504 ;
  assign n9506 = n9167 & ~n9505 ;
  assign n9507 = ~n9179 & n9497 ;
  assign n9508 = ~n9167 & n9505 ;
  assign n9509 = ( x17 & ~n9497 ) | ( x17 & n9508 ) | ( ~n9497 & n9508 ) ;
  assign n9510 = ( ~n9506 & n9507 ) | ( ~n9506 & n9509 ) | ( n9507 & n9509 ) ;
  assign n9511 = n9167 & ~n9497 ;
  assign n9512 = ( ~x18 & n9507 ) | ( ~x18 & n9511 ) | ( n9507 & n9511 ) ;
  assign n9513 = ( x18 & n9507 ) | ( x18 & n9511 ) | ( n9507 & n9511 ) ;
  assign n9514 = ( x18 & n9512 ) | ( x18 & ~n9513 ) | ( n9512 & ~n9513 ) ;
  assign n9515 = ( ~n8838 & n9510 ) | ( ~n8838 & n9514 ) | ( n9510 & n9514 ) ;
  assign n9516 = ~n8838 & n9167 ;
  assign n9517 = ( n9185 & n9497 ) | ( n9185 & n9516 ) | ( n9497 & n9516 ) ;
  assign n9518 = ( x19 & n9512 ) | ( x19 & n9517 ) | ( n9512 & n9517 ) ;
  assign n9519 = ( ~x19 & n9512 ) | ( ~x19 & n9517 ) | ( n9512 & n9517 ) ;
  assign n9520 = ( x19 & ~n9518 ) | ( x19 & n9519 ) | ( ~n9518 & n9519 ) ;
  assign n9521 = ( ~n8517 & n9515 ) | ( ~n8517 & n9520 ) | ( n9515 & n9520 ) ;
  assign n9522 = ( n8517 & ~n9184 ) | ( n8517 & n9497 ) | ( ~n9184 & n9497 ) ;
  assign n9523 = n8517 & ~n9184 ;
  assign n9524 = ( n9188 & n9522 ) | ( n9188 & n9523 ) | ( n9522 & n9523 ) ;
  assign n9525 = ( ~n9188 & n9522 ) | ( ~n9188 & n9523 ) | ( n9522 & n9523 ) ;
  assign n9526 = ( n9188 & ~n9524 ) | ( n9188 & n9525 ) | ( ~n9524 & n9525 ) ;
  assign n9527 = ( ~n8201 & n9521 ) | ( ~n8201 & n9526 ) | ( n9521 & n9526 ) ;
  assign n9528 = ( n8201 & ~n9189 ) | ( n8201 & n9497 ) | ( ~n9189 & n9497 ) ;
  assign n9529 = n8201 & ~n9189 ;
  assign n9530 = ( n9194 & n9528 ) | ( n9194 & n9529 ) | ( n9528 & n9529 ) ;
  assign n9531 = ( ~n9194 & n9528 ) | ( ~n9194 & n9529 ) | ( n9528 & n9529 ) ;
  assign n9532 = ( n9194 & ~n9530 ) | ( n9194 & n9531 ) | ( ~n9530 & n9531 ) ;
  assign n9533 = ( ~n7897 & n9527 ) | ( ~n7897 & n9532 ) | ( n9527 & n9532 ) ;
  assign n9534 = ( n7897 & ~n9195 ) | ( n7897 & n9497 ) | ( ~n9195 & n9497 ) ;
  assign n9535 = n7897 & ~n9195 ;
  assign n9536 = ( n9200 & n9534 ) | ( n9200 & n9535 ) | ( n9534 & n9535 ) ;
  assign n9537 = ( ~n9200 & n9534 ) | ( ~n9200 & n9535 ) | ( n9534 & n9535 ) ;
  assign n9538 = ( n9200 & ~n9536 ) | ( n9200 & n9537 ) | ( ~n9536 & n9537 ) ;
  assign n9539 = ( ~n7594 & n9533 ) | ( ~n7594 & n9538 ) | ( n9533 & n9538 ) ;
  assign n9540 = ~n7594 & n9201 ;
  assign n9541 = ( ~n7594 & n9201 ) | ( ~n7594 & n9497 ) | ( n9201 & n9497 ) ;
  assign n9542 = ( n9206 & n9540 ) | ( n9206 & n9541 ) | ( n9540 & n9541 ) ;
  assign n9543 = ( ~n9206 & n9540 ) | ( ~n9206 & n9541 ) | ( n9540 & n9541 ) ;
  assign n9544 = ( n9206 & ~n9542 ) | ( n9206 & n9543 ) | ( ~n9542 & n9543 ) ;
  assign n9545 = ( ~n7296 & n9539 ) | ( ~n7296 & n9544 ) | ( n9539 & n9544 ) ;
  assign n9546 = ( n7296 & ~n9207 ) | ( n7296 & n9497 ) | ( ~n9207 & n9497 ) ;
  assign n9547 = n7296 & ~n9207 ;
  assign n9548 = ( n9212 & n9546 ) | ( n9212 & n9547 ) | ( n9546 & n9547 ) ;
  assign n9549 = ( ~n9212 & n9546 ) | ( ~n9212 & n9547 ) | ( n9546 & n9547 ) ;
  assign n9550 = ( n9212 & ~n9548 ) | ( n9212 & n9549 ) | ( ~n9548 & n9549 ) ;
  assign n9551 = ( ~n7006 & n9545 ) | ( ~n7006 & n9550 ) | ( n9545 & n9550 ) ;
  assign n9552 = ( n7006 & ~n9213 ) | ( n7006 & n9497 ) | ( ~n9213 & n9497 ) ;
  assign n9553 = n7006 & ~n9213 ;
  assign n9554 = ( n9218 & n9552 ) | ( n9218 & n9553 ) | ( n9552 & n9553 ) ;
  assign n9555 = ( ~n9218 & n9552 ) | ( ~n9218 & n9553 ) | ( n9552 & n9553 ) ;
  assign n9556 = ( n9218 & ~n9554 ) | ( n9218 & n9555 ) | ( ~n9554 & n9555 ) ;
  assign n9557 = ( ~n6723 & n9551 ) | ( ~n6723 & n9556 ) | ( n9551 & n9556 ) ;
  assign n9558 = ( n6723 & ~n9219 ) | ( n6723 & n9497 ) | ( ~n9219 & n9497 ) ;
  assign n9559 = n6723 & ~n9219 ;
  assign n9560 = ( n9224 & n9558 ) | ( n9224 & n9559 ) | ( n9558 & n9559 ) ;
  assign n9561 = ( ~n9224 & n9558 ) | ( ~n9224 & n9559 ) | ( n9558 & n9559 ) ;
  assign n9562 = ( n9224 & ~n9560 ) | ( n9224 & n9561 ) | ( ~n9560 & n9561 ) ;
  assign n9563 = ( ~n6442 & n9557 ) | ( ~n6442 & n9562 ) | ( n9557 & n9562 ) ;
  assign n9564 = ~n6442 & n9225 ;
  assign n9565 = ( ~n6442 & n9225 ) | ( ~n6442 & n9497 ) | ( n9225 & n9497 ) ;
  assign n9566 = ( ~n9230 & n9564 ) | ( ~n9230 & n9565 ) | ( n9564 & n9565 ) ;
  assign n9567 = ( n9230 & n9564 ) | ( n9230 & n9565 ) | ( n9564 & n9565 ) ;
  assign n9568 = ( n9230 & n9566 ) | ( n9230 & ~n9567 ) | ( n9566 & ~n9567 ) ;
  assign n9569 = ( ~n6172 & n9563 ) | ( ~n6172 & n9568 ) | ( n9563 & n9568 ) ;
  assign n9570 = ~n6172 & n9231 ;
  assign n9571 = ( ~n6172 & n9231 ) | ( ~n6172 & n9497 ) | ( n9231 & n9497 ) ;
  assign n9572 = ( ~n9236 & n9570 ) | ( ~n9236 & n9571 ) | ( n9570 & n9571 ) ;
  assign n9573 = ( n9236 & n9570 ) | ( n9236 & n9571 ) | ( n9570 & n9571 ) ;
  assign n9574 = ( n9236 & n9572 ) | ( n9236 & ~n9573 ) | ( n9572 & ~n9573 ) ;
  assign n9575 = ( ~n5905 & n9569 ) | ( ~n5905 & n9574 ) | ( n9569 & n9574 ) ;
  assign n9576 = ~n5905 & n9237 ;
  assign n9577 = ( ~n5905 & n9237 ) | ( ~n5905 & n9497 ) | ( n9237 & n9497 ) ;
  assign n9578 = ( ~n9242 & n9576 ) | ( ~n9242 & n9577 ) | ( n9576 & n9577 ) ;
  assign n9579 = ( n9242 & n9576 ) | ( n9242 & n9577 ) | ( n9576 & n9577 ) ;
  assign n9580 = ( n9242 & n9578 ) | ( n9242 & ~n9579 ) | ( n9578 & ~n9579 ) ;
  assign n9581 = ( ~n5642 & n9575 ) | ( ~n5642 & n9580 ) | ( n9575 & n9580 ) ;
  assign n9582 = ~n5642 & n9243 ;
  assign n9583 = ( ~n5642 & n9243 ) | ( ~n5642 & n9497 ) | ( n9243 & n9497 ) ;
  assign n9584 = ( ~n9248 & n9582 ) | ( ~n9248 & n9583 ) | ( n9582 & n9583 ) ;
  assign n9585 = ( n9248 & n9582 ) | ( n9248 & n9583 ) | ( n9582 & n9583 ) ;
  assign n9586 = ( n9248 & n9584 ) | ( n9248 & ~n9585 ) | ( n9584 & ~n9585 ) ;
  assign n9587 = ( ~n5386 & n9581 ) | ( ~n5386 & n9586 ) | ( n9581 & n9586 ) ;
  assign n9588 = ( n5386 & ~n9249 ) | ( n5386 & n9497 ) | ( ~n9249 & n9497 ) ;
  assign n9589 = n5386 & ~n9249 ;
  assign n9590 = ( n9254 & n9588 ) | ( n9254 & n9589 ) | ( n9588 & n9589 ) ;
  assign n9591 = ( ~n9254 & n9588 ) | ( ~n9254 & n9589 ) | ( n9588 & n9589 ) ;
  assign n9592 = ( n9254 & ~n9590 ) | ( n9254 & n9591 ) | ( ~n9590 & n9591 ) ;
  assign n9593 = ( ~n5139 & n9587 ) | ( ~n5139 & n9592 ) | ( n9587 & n9592 ) ;
  assign n9594 = ( n5139 & ~n9255 ) | ( n5139 & n9497 ) | ( ~n9255 & n9497 ) ;
  assign n9595 = n5139 & ~n9255 ;
  assign n9596 = ( n9260 & n9594 ) | ( n9260 & n9595 ) | ( n9594 & n9595 ) ;
  assign n9597 = ( ~n9260 & n9594 ) | ( ~n9260 & n9595 ) | ( n9594 & n9595 ) ;
  assign n9598 = ( n9260 & ~n9596 ) | ( n9260 & n9597 ) | ( ~n9596 & n9597 ) ;
  assign n9599 = ( ~n4898 & n9593 ) | ( ~n4898 & n9598 ) | ( n9593 & n9598 ) ;
  assign n9600 = n4898 & ~n9261 ;
  assign n9601 = ( n4898 & ~n9261 ) | ( n4898 & n9497 ) | ( ~n9261 & n9497 ) ;
  assign n9602 = ( n9266 & n9600 ) | ( n9266 & n9601 ) | ( n9600 & n9601 ) ;
  assign n9603 = ( ~n9266 & n9600 ) | ( ~n9266 & n9601 ) | ( n9600 & n9601 ) ;
  assign n9604 = ( n9266 & ~n9602 ) | ( n9266 & n9603 ) | ( ~n9602 & n9603 ) ;
  assign n9605 = ( ~n4661 & n9599 ) | ( ~n4661 & n9604 ) | ( n9599 & n9604 ) ;
  assign n9606 = ( n4661 & ~n9267 ) | ( n4661 & n9497 ) | ( ~n9267 & n9497 ) ;
  assign n9607 = n4661 & ~n9267 ;
  assign n9608 = ( n9272 & n9606 ) | ( n9272 & n9607 ) | ( n9606 & n9607 ) ;
  assign n9609 = ( ~n9272 & n9606 ) | ( ~n9272 & n9607 ) | ( n9606 & n9607 ) ;
  assign n9610 = ( n9272 & ~n9608 ) | ( n9272 & n9609 ) | ( ~n9608 & n9609 ) ;
  assign n9611 = ( ~n4432 & n9605 ) | ( ~n4432 & n9610 ) | ( n9605 & n9610 ) ;
  assign n9612 = ~n4432 & n9273 ;
  assign n9613 = ( ~n4432 & n9273 ) | ( ~n4432 & n9497 ) | ( n9273 & n9497 ) ;
  assign n9614 = ( ~n9278 & n9612 ) | ( ~n9278 & n9613 ) | ( n9612 & n9613 ) ;
  assign n9615 = ( n9278 & n9612 ) | ( n9278 & n9613 ) | ( n9612 & n9613 ) ;
  assign n9616 = ( n9278 & n9614 ) | ( n9278 & ~n9615 ) | ( n9614 & ~n9615 ) ;
  assign n9617 = ( ~n4203 & n9611 ) | ( ~n4203 & n9616 ) | ( n9611 & n9616 ) ;
  assign n9618 = ( n4203 & ~n9279 ) | ( n4203 & n9497 ) | ( ~n9279 & n9497 ) ;
  assign n9619 = n4203 & ~n9279 ;
  assign n9620 = ( n9284 & n9618 ) | ( n9284 & n9619 ) | ( n9618 & n9619 ) ;
  assign n9621 = ( ~n9284 & n9618 ) | ( ~n9284 & n9619 ) | ( n9618 & n9619 ) ;
  assign n9622 = ( n9284 & ~n9620 ) | ( n9284 & n9621 ) | ( ~n9620 & n9621 ) ;
  assign n9623 = ( ~n3985 & n9617 ) | ( ~n3985 & n9622 ) | ( n9617 & n9622 ) ;
  assign n9624 = ~n3985 & n9285 ;
  assign n9625 = ( ~n3985 & n9285 ) | ( ~n3985 & n9497 ) | ( n9285 & n9497 ) ;
  assign n9626 = ( ~n9290 & n9624 ) | ( ~n9290 & n9625 ) | ( n9624 & n9625 ) ;
  assign n9627 = ( n9290 & n9624 ) | ( n9290 & n9625 ) | ( n9624 & n9625 ) ;
  assign n9628 = ( n9290 & n9626 ) | ( n9290 & ~n9627 ) | ( n9626 & ~n9627 ) ;
  assign n9629 = ( ~n3772 & n9623 ) | ( ~n3772 & n9628 ) | ( n9623 & n9628 ) ;
  assign n9630 = ( n3772 & ~n9291 ) | ( n3772 & n9497 ) | ( ~n9291 & n9497 ) ;
  assign n9631 = n3772 & ~n9291 ;
  assign n9632 = ( n9296 & n9630 ) | ( n9296 & n9631 ) | ( n9630 & n9631 ) ;
  assign n9633 = ( ~n9296 & n9630 ) | ( ~n9296 & n9631 ) | ( n9630 & n9631 ) ;
  assign n9634 = ( n9296 & ~n9632 ) | ( n9296 & n9633 ) | ( ~n9632 & n9633 ) ;
  assign n9635 = ( ~n3567 & n9629 ) | ( ~n3567 & n9634 ) | ( n9629 & n9634 ) ;
  assign n9636 = n3567 & ~n9297 ;
  assign n9637 = ( n3567 & ~n9297 ) | ( n3567 & n9497 ) | ( ~n9297 & n9497 ) ;
  assign n9638 = ( n9302 & n9636 ) | ( n9302 & n9637 ) | ( n9636 & n9637 ) ;
  assign n9639 = ( ~n9302 & n9636 ) | ( ~n9302 & n9637 ) | ( n9636 & n9637 ) ;
  assign n9640 = ( n9302 & ~n9638 ) | ( n9302 & n9639 ) | ( ~n9638 & n9639 ) ;
  assign n9641 = ( ~n3362 & n9635 ) | ( ~n3362 & n9640 ) | ( n9635 & n9640 ) ;
  assign n9642 = ( n3362 & ~n9303 ) | ( n3362 & n9497 ) | ( ~n9303 & n9497 ) ;
  assign n9643 = n3362 & ~n9303 ;
  assign n9644 = ( n9308 & n9642 ) | ( n9308 & n9643 ) | ( n9642 & n9643 ) ;
  assign n9645 = ( ~n9308 & n9642 ) | ( ~n9308 & n9643 ) | ( n9642 & n9643 ) ;
  assign n9646 = ( n9308 & ~n9644 ) | ( n9308 & n9645 ) | ( ~n9644 & n9645 ) ;
  assign n9647 = ( ~n3169 & n9641 ) | ( ~n3169 & n9646 ) | ( n9641 & n9646 ) ;
  assign n9648 = ( n3169 & ~n9309 ) | ( n3169 & n9497 ) | ( ~n9309 & n9497 ) ;
  assign n9649 = n3169 & ~n9309 ;
  assign n9650 = ( n9314 & n9648 ) | ( n9314 & n9649 ) | ( n9648 & n9649 ) ;
  assign n9651 = ( ~n9314 & n9648 ) | ( ~n9314 & n9649 ) | ( n9648 & n9649 ) ;
  assign n9652 = ( n9314 & ~n9650 ) | ( n9314 & n9651 ) | ( ~n9650 & n9651 ) ;
  assign n9653 = ( ~n2979 & n9647 ) | ( ~n2979 & n9652 ) | ( n9647 & n9652 ) ;
  assign n9654 = ( n2979 & ~n9315 ) | ( n2979 & n9497 ) | ( ~n9315 & n9497 ) ;
  assign n9655 = n2979 & ~n9315 ;
  assign n9656 = ( n9320 & n9654 ) | ( n9320 & n9655 ) | ( n9654 & n9655 ) ;
  assign n9657 = ( ~n9320 & n9654 ) | ( ~n9320 & n9655 ) | ( n9654 & n9655 ) ;
  assign n9658 = ( n9320 & ~n9656 ) | ( n9320 & n9657 ) | ( ~n9656 & n9657 ) ;
  assign n9659 = ( ~n2791 & n9653 ) | ( ~n2791 & n9658 ) | ( n9653 & n9658 ) ;
  assign n9660 = ~n2791 & n9321 ;
  assign n9661 = ( ~n2791 & n9321 ) | ( ~n2791 & n9497 ) | ( n9321 & n9497 ) ;
  assign n9662 = ( ~n9326 & n9660 ) | ( ~n9326 & n9661 ) | ( n9660 & n9661 ) ;
  assign n9663 = ( n9326 & n9660 ) | ( n9326 & n9661 ) | ( n9660 & n9661 ) ;
  assign n9664 = ( n9326 & n9662 ) | ( n9326 & ~n9663 ) | ( n9662 & ~n9663 ) ;
  assign n9665 = ( ~n2615 & n9659 ) | ( ~n2615 & n9664 ) | ( n9659 & n9664 ) ;
  assign n9666 = ~n2615 & n9327 ;
  assign n9667 = ( ~n2615 & n9327 ) | ( ~n2615 & n9497 ) | ( n9327 & n9497 ) ;
  assign n9668 = ( ~n9332 & n9666 ) | ( ~n9332 & n9667 ) | ( n9666 & n9667 ) ;
  assign n9669 = ( n9332 & n9666 ) | ( n9332 & n9667 ) | ( n9666 & n9667 ) ;
  assign n9670 = ( n9332 & n9668 ) | ( n9332 & ~n9669 ) | ( n9668 & ~n9669 ) ;
  assign n9671 = ( ~n2443 & n9665 ) | ( ~n2443 & n9670 ) | ( n9665 & n9670 ) ;
  assign n9672 = ( n2443 & ~n9333 ) | ( n2443 & n9497 ) | ( ~n9333 & n9497 ) ;
  assign n9673 = n2443 & ~n9333 ;
  assign n9674 = ( n9338 & n9672 ) | ( n9338 & n9673 ) | ( n9672 & n9673 ) ;
  assign n9675 = ( ~n9338 & n9672 ) | ( ~n9338 & n9673 ) | ( n9672 & n9673 ) ;
  assign n9676 = ( n9338 & ~n9674 ) | ( n9338 & n9675 ) | ( ~n9674 & n9675 ) ;
  assign n9677 = ( ~n2277 & n9671 ) | ( ~n2277 & n9676 ) | ( n9671 & n9676 ) ;
  assign n9678 = ~n2277 & n9339 ;
  assign n9679 = ( ~n2277 & n9339 ) | ( ~n2277 & n9497 ) | ( n9339 & n9497 ) ;
  assign n9680 = ( ~n9344 & n9678 ) | ( ~n9344 & n9679 ) | ( n9678 & n9679 ) ;
  assign n9681 = ( n9344 & n9678 ) | ( n9344 & n9679 ) | ( n9678 & n9679 ) ;
  assign n9682 = ( n9344 & n9680 ) | ( n9344 & ~n9681 ) | ( n9680 & ~n9681 ) ;
  assign n9683 = ( ~n2111 & n9677 ) | ( ~n2111 & n9682 ) | ( n9677 & n9682 ) ;
  assign n9684 = ( n2111 & ~n9345 ) | ( n2111 & n9497 ) | ( ~n9345 & n9497 ) ;
  assign n9685 = n2111 & ~n9345 ;
  assign n9686 = ( n9350 & n9684 ) | ( n9350 & n9685 ) | ( n9684 & n9685 ) ;
  assign n9687 = ( ~n9350 & n9684 ) | ( ~n9350 & n9685 ) | ( n9684 & n9685 ) ;
  assign n9688 = ( n9350 & ~n9686 ) | ( n9350 & n9687 ) | ( ~n9686 & n9687 ) ;
  assign n9689 = ( ~n1949 & n9683 ) | ( ~n1949 & n9688 ) | ( n9683 & n9688 ) ;
  assign n9690 = ( n1949 & ~n9351 ) | ( n1949 & n9497 ) | ( ~n9351 & n9497 ) ;
  assign n9691 = n1949 & ~n9351 ;
  assign n9692 = ( n9356 & n9690 ) | ( n9356 & n9691 ) | ( n9690 & n9691 ) ;
  assign n9693 = ( ~n9356 & n9690 ) | ( ~n9356 & n9691 ) | ( n9690 & n9691 ) ;
  assign n9694 = ( n9356 & ~n9692 ) | ( n9356 & n9693 ) | ( ~n9692 & n9693 ) ;
  assign n9695 = ( ~n1802 & n9689 ) | ( ~n1802 & n9694 ) | ( n9689 & n9694 ) ;
  assign n9696 = ( n1802 & ~n9357 ) | ( n1802 & n9497 ) | ( ~n9357 & n9497 ) ;
  assign n9697 = n1802 & ~n9357 ;
  assign n9698 = ( n9362 & n9696 ) | ( n9362 & n9697 ) | ( n9696 & n9697 ) ;
  assign n9699 = ( ~n9362 & n9696 ) | ( ~n9362 & n9697 ) | ( n9696 & n9697 ) ;
  assign n9700 = ( n9362 & ~n9698 ) | ( n9362 & n9699 ) | ( ~n9698 & n9699 ) ;
  assign n9701 = ( ~n1661 & n9695 ) | ( ~n1661 & n9700 ) | ( n9695 & n9700 ) ;
  assign n9702 = ~n1661 & n9363 ;
  assign n9703 = ( ~n1661 & n9363 ) | ( ~n1661 & n9497 ) | ( n9363 & n9497 ) ;
  assign n9704 = ( ~n9368 & n9702 ) | ( ~n9368 & n9703 ) | ( n9702 & n9703 ) ;
  assign n9705 = ( n9368 & n9702 ) | ( n9368 & n9703 ) | ( n9702 & n9703 ) ;
  assign n9706 = ( n9368 & n9704 ) | ( n9368 & ~n9705 ) | ( n9704 & ~n9705 ) ;
  assign n9707 = ( ~n1523 & n9701 ) | ( ~n1523 & n9706 ) | ( n9701 & n9706 ) ;
  assign n9708 = ( n1523 & ~n9369 ) | ( n1523 & n9497 ) | ( ~n9369 & n9497 ) ;
  assign n9709 = n1523 & ~n9369 ;
  assign n9710 = ( n9374 & n9708 ) | ( n9374 & n9709 ) | ( n9708 & n9709 ) ;
  assign n9711 = ( ~n9374 & n9708 ) | ( ~n9374 & n9709 ) | ( n9708 & n9709 ) ;
  assign n9712 = ( n9374 & ~n9710 ) | ( n9374 & n9711 ) | ( ~n9710 & n9711 ) ;
  assign n9713 = ( ~n1393 & n9707 ) | ( ~n1393 & n9712 ) | ( n9707 & n9712 ) ;
  assign n9714 = ( n1393 & ~n9375 ) | ( n1393 & n9497 ) | ( ~n9375 & n9497 ) ;
  assign n9715 = n1393 & ~n9375 ;
  assign n9716 = ( n9380 & n9714 ) | ( n9380 & n9715 ) | ( n9714 & n9715 ) ;
  assign n9717 = ( ~n9380 & n9714 ) | ( ~n9380 & n9715 ) | ( n9714 & n9715 ) ;
  assign n9718 = ( n9380 & ~n9716 ) | ( n9380 & n9717 ) | ( ~n9716 & n9717 ) ;
  assign n9719 = ( ~n1266 & n9713 ) | ( ~n1266 & n9718 ) | ( n9713 & n9718 ) ;
  assign n9720 = ~n1266 & n9381 ;
  assign n9721 = ( ~n1266 & n9381 ) | ( ~n1266 & n9497 ) | ( n9381 & n9497 ) ;
  assign n9722 = ( ~n9386 & n9720 ) | ( ~n9386 & n9721 ) | ( n9720 & n9721 ) ;
  assign n9723 = ( n9386 & n9720 ) | ( n9386 & n9721 ) | ( n9720 & n9721 ) ;
  assign n9724 = ( n9386 & n9722 ) | ( n9386 & ~n9723 ) | ( n9722 & ~n9723 ) ;
  assign n9725 = ( ~n1150 & n9719 ) | ( ~n1150 & n9724 ) | ( n9719 & n9724 ) ;
  assign n9726 = ~n1150 & n9387 ;
  assign n9727 = ( ~n1150 & n9387 ) | ( ~n1150 & n9497 ) | ( n9387 & n9497 ) ;
  assign n9728 = ( ~n9392 & n9726 ) | ( ~n9392 & n9727 ) | ( n9726 & n9727 ) ;
  assign n9729 = ( n9392 & n9726 ) | ( n9392 & n9727 ) | ( n9726 & n9727 ) ;
  assign n9730 = ( n9392 & n9728 ) | ( n9392 & ~n9729 ) | ( n9728 & ~n9729 ) ;
  assign n9731 = ( ~n1038 & n9725 ) | ( ~n1038 & n9730 ) | ( n9725 & n9730 ) ;
  assign n9732 = ( n1038 & ~n9393 ) | ( n1038 & n9497 ) | ( ~n9393 & n9497 ) ;
  assign n9733 = n1038 & ~n9393 ;
  assign n9734 = ( n9398 & n9732 ) | ( n9398 & n9733 ) | ( n9732 & n9733 ) ;
  assign n9735 = ( ~n9398 & n9732 ) | ( ~n9398 & n9733 ) | ( n9732 & n9733 ) ;
  assign n9736 = ( n9398 & ~n9734 ) | ( n9398 & n9735 ) | ( ~n9734 & n9735 ) ;
  assign n9737 = ( ~n933 & n9731 ) | ( ~n933 & n9736 ) | ( n9731 & n9736 ) ;
  assign n9738 = ( n933 & ~n9399 ) | ( n933 & n9497 ) | ( ~n9399 & n9497 ) ;
  assign n9739 = n933 & ~n9399 ;
  assign n9740 = ( n9404 & n9738 ) | ( n9404 & n9739 ) | ( n9738 & n9739 ) ;
  assign n9741 = ( ~n9404 & n9738 ) | ( ~n9404 & n9739 ) | ( n9738 & n9739 ) ;
  assign n9742 = ( n9404 & ~n9740 ) | ( n9404 & n9741 ) | ( ~n9740 & n9741 ) ;
  assign n9743 = ( ~n839 & n9737 ) | ( ~n839 & n9742 ) | ( n9737 & n9742 ) ;
  assign n9744 = ( n839 & ~n9405 ) | ( n839 & n9497 ) | ( ~n9405 & n9497 ) ;
  assign n9745 = n839 & ~n9405 ;
  assign n9746 = ( n9410 & n9744 ) | ( n9410 & n9745 ) | ( n9744 & n9745 ) ;
  assign n9747 = ( ~n9410 & n9744 ) | ( ~n9410 & n9745 ) | ( n9744 & n9745 ) ;
  assign n9748 = ( n9410 & ~n9746 ) | ( n9410 & n9747 ) | ( ~n9746 & n9747 ) ;
  assign n9749 = ( ~n746 & n9743 ) | ( ~n746 & n9748 ) | ( n9743 & n9748 ) ;
  assign n9750 = ( n746 & ~n9411 ) | ( n746 & n9497 ) | ( ~n9411 & n9497 ) ;
  assign n9751 = n746 & ~n9411 ;
  assign n9752 = ( n9416 & n9750 ) | ( n9416 & n9751 ) | ( n9750 & n9751 ) ;
  assign n9753 = ( ~n9416 & n9750 ) | ( ~n9416 & n9751 ) | ( n9750 & n9751 ) ;
  assign n9754 = ( n9416 & ~n9752 ) | ( n9416 & n9753 ) | ( ~n9752 & n9753 ) ;
  assign n9755 = ( ~n664 & n9749 ) | ( ~n664 & n9754 ) | ( n9749 & n9754 ) ;
  assign n9756 = ( n664 & ~n9417 ) | ( n664 & n9497 ) | ( ~n9417 & n9497 ) ;
  assign n9757 = n664 & ~n9417 ;
  assign n9758 = ( n9422 & n9756 ) | ( n9422 & n9757 ) | ( n9756 & n9757 ) ;
  assign n9759 = ( ~n9422 & n9756 ) | ( ~n9422 & n9757 ) | ( n9756 & n9757 ) ;
  assign n9760 = ( n9422 & ~n9758 ) | ( n9422 & n9759 ) | ( ~n9758 & n9759 ) ;
  assign n9761 = ( ~n588 & n9755 ) | ( ~n588 & n9760 ) | ( n9755 & n9760 ) ;
  assign n9762 = ( n588 & ~n9423 ) | ( n588 & n9497 ) | ( ~n9423 & n9497 ) ;
  assign n9763 = n588 & ~n9423 ;
  assign n9764 = ( n9428 & n9762 ) | ( n9428 & n9763 ) | ( n9762 & n9763 ) ;
  assign n9765 = ( ~n9428 & n9762 ) | ( ~n9428 & n9763 ) | ( n9762 & n9763 ) ;
  assign n9766 = ( n9428 & ~n9764 ) | ( n9428 & n9765 ) | ( ~n9764 & n9765 ) ;
  assign n9767 = ( ~n518 & n9761 ) | ( ~n518 & n9766 ) | ( n9761 & n9766 ) ;
  assign n9768 = ( n518 & ~n9429 ) | ( n518 & n9497 ) | ( ~n9429 & n9497 ) ;
  assign n9769 = n518 & ~n9429 ;
  assign n9770 = ( n9434 & n9768 ) | ( n9434 & n9769 ) | ( n9768 & n9769 ) ;
  assign n9771 = ( ~n9434 & n9768 ) | ( ~n9434 & n9769 ) | ( n9768 & n9769 ) ;
  assign n9772 = ( n9434 & ~n9770 ) | ( n9434 & n9771 ) | ( ~n9770 & n9771 ) ;
  assign n9773 = ( ~n454 & n9767 ) | ( ~n454 & n9772 ) | ( n9767 & n9772 ) ;
  assign n9774 = ~n454 & n9435 ;
  assign n9775 = ( ~n454 & n9435 ) | ( ~n454 & n9497 ) | ( n9435 & n9497 ) ;
  assign n9776 = ( ~n9177 & n9774 ) | ( ~n9177 & n9775 ) | ( n9774 & n9775 ) ;
  assign n9777 = ( n9177 & n9774 ) | ( n9177 & n9775 ) | ( n9774 & n9775 ) ;
  assign n9778 = ( n9177 & n9776 ) | ( n9177 & ~n9777 ) | ( n9776 & ~n9777 ) ;
  assign n9779 = ( ~n396 & n9773 ) | ( ~n396 & n9778 ) | ( n9773 & n9778 ) ;
  assign n9780 = ~n396 & n9436 ;
  assign n9781 = ( ~n396 & n9436 ) | ( ~n396 & n9497 ) | ( n9436 & n9497 ) ;
  assign n9782 = ( ~n9441 & n9780 ) | ( ~n9441 & n9781 ) | ( n9780 & n9781 ) ;
  assign n9783 = ( n9441 & n9780 ) | ( n9441 & n9781 ) | ( n9780 & n9781 ) ;
  assign n9784 = ( n9441 & n9782 ) | ( n9441 & ~n9783 ) | ( n9782 & ~n9783 ) ;
  assign n9785 = ( ~n344 & n9779 ) | ( ~n344 & n9784 ) | ( n9779 & n9784 ) ;
  assign n9786 = n344 & ~n9442 ;
  assign n9787 = ( n344 & ~n9442 ) | ( n344 & n9497 ) | ( ~n9442 & n9497 ) ;
  assign n9788 = ( ~n9447 & n9786 ) | ( ~n9447 & n9787 ) | ( n9786 & n9787 ) ;
  assign n9789 = ( n9447 & n9786 ) | ( n9447 & n9787 ) | ( n9786 & n9787 ) ;
  assign n9790 = ( n9447 & n9788 ) | ( n9447 & ~n9789 ) | ( n9788 & ~n9789 ) ;
  assign n9791 = ( ~n298 & n9785 ) | ( ~n298 & n9790 ) | ( n9785 & n9790 ) ;
  assign n9792 = ~n298 & n9448 ;
  assign n9793 = ( ~n298 & n9448 ) | ( ~n298 & n9497 ) | ( n9448 & n9497 ) ;
  assign n9794 = ( n9453 & n9792 ) | ( n9453 & n9793 ) | ( n9792 & n9793 ) ;
  assign n9795 = ( ~n9453 & n9792 ) | ( ~n9453 & n9793 ) | ( n9792 & n9793 ) ;
  assign n9796 = ( n9453 & ~n9794 ) | ( n9453 & n9795 ) | ( ~n9794 & n9795 ) ;
  assign n9797 = ( ~n258 & n9791 ) | ( ~n258 & n9796 ) | ( n9791 & n9796 ) ;
  assign n9798 = ( n258 & ~n9454 ) | ( n258 & n9497 ) | ( ~n9454 & n9497 ) ;
  assign n9799 = n258 & ~n9454 ;
  assign n9800 = ( n9459 & n9798 ) | ( n9459 & n9799 ) | ( n9798 & n9799 ) ;
  assign n9801 = ( ~n9459 & n9798 ) | ( ~n9459 & n9799 ) | ( n9798 & n9799 ) ;
  assign n9802 = ( n9459 & ~n9800 ) | ( n9459 & n9801 ) | ( ~n9800 & n9801 ) ;
  assign n9803 = ( ~n225 & n9797 ) | ( ~n225 & n9802 ) | ( n9797 & n9802 ) ;
  assign n9804 = ( n225 & ~n9460 ) | ( n225 & n9497 ) | ( ~n9460 & n9497 ) ;
  assign n9805 = n225 & ~n9460 ;
  assign n9806 = ( n9465 & n9804 ) | ( n9465 & n9805 ) | ( n9804 & n9805 ) ;
  assign n9807 = ( ~n9465 & n9804 ) | ( ~n9465 & n9805 ) | ( n9804 & n9805 ) ;
  assign n9808 = ( n9465 & ~n9806 ) | ( n9465 & n9807 ) | ( ~n9806 & n9807 ) ;
  assign n9809 = ( ~n197 & n9803 ) | ( ~n197 & n9808 ) | ( n9803 & n9808 ) ;
  assign n9810 = ~n197 & n9466 ;
  assign n9811 = ( ~n197 & n9466 ) | ( ~n197 & n9497 ) | ( n9466 & n9497 ) ;
  assign n9812 = ( ~n9471 & n9810 ) | ( ~n9471 & n9811 ) | ( n9810 & n9811 ) ;
  assign n9813 = ( n9471 & n9810 ) | ( n9471 & n9811 ) | ( n9810 & n9811 ) ;
  assign n9814 = ( n9471 & n9812 ) | ( n9471 & ~n9813 ) | ( n9812 & ~n9813 ) ;
  assign n9815 = ( ~n170 & n9809 ) | ( ~n170 & n9814 ) | ( n9809 & n9814 ) ;
  assign n9816 = ( n170 & ~n9472 ) | ( n170 & n9497 ) | ( ~n9472 & n9497 ) ;
  assign n9817 = n170 & ~n9472 ;
  assign n9818 = ( n9477 & n9816 ) | ( n9477 & n9817 ) | ( n9816 & n9817 ) ;
  assign n9819 = ( ~n9477 & n9816 ) | ( ~n9477 & n9817 ) | ( n9816 & n9817 ) ;
  assign n9820 = ( n9477 & ~n9818 ) | ( n9477 & n9819 ) | ( ~n9818 & n9819 ) ;
  assign n9821 = ( ~n142 & n9815 ) | ( ~n142 & n9820 ) | ( n9815 & n9820 ) ;
  assign n9822 = ~n142 & n9478 ;
  assign n9823 = ( ~n142 & n9478 ) | ( ~n142 & n9497 ) | ( n9478 & n9497 ) ;
  assign n9824 = ( ~n9483 & n9822 ) | ( ~n9483 & n9823 ) | ( n9822 & n9823 ) ;
  assign n9825 = ( n9483 & n9822 ) | ( n9483 & n9823 ) | ( n9822 & n9823 ) ;
  assign n9826 = ( n9483 & n9824 ) | ( n9483 & ~n9825 ) | ( n9824 & ~n9825 ) ;
  assign n9827 = ( ~n132 & n9821 ) | ( ~n132 & n9826 ) | ( n9821 & n9826 ) ;
  assign n9828 = ( n132 & ~n9484 ) | ( n132 & n9497 ) | ( ~n9484 & n9497 ) ;
  assign n9829 = n132 & ~n9484 ;
  assign n9830 = ( n9489 & n9828 ) | ( n9489 & n9829 ) | ( n9828 & n9829 ) ;
  assign n9831 = ( ~n9489 & n9828 ) | ( ~n9489 & n9829 ) | ( n9828 & n9829 ) ;
  assign n9832 = ( n9489 & ~n9830 ) | ( n9489 & n9831 ) | ( ~n9830 & n9831 ) ;
  assign n9833 = ( ~n131 & n9827 ) | ( ~n131 & n9832 ) | ( n9827 & n9832 ) ;
  assign n9834 = n9503 | n9833 ;
  assign n9835 = n9172 & n9490 ;
  assign n9836 = ( ~n9498 & n9500 ) | ( ~n9498 & n9835 ) | ( n9500 & n9835 ) ;
  assign n9837 = ~n9832 & n9836 ;
  assign n9838 = ~n9827 & n9837 ;
  assign n9839 = n9502 & ~n9835 ;
  assign n9840 = ~n9832 & n9839 ;
  assign n9841 = ( ~n131 & n9827 ) | ( ~n131 & n9840 ) | ( n9827 & n9840 ) ;
  assign n9842 = ( n9832 & ~n9833 ) | ( n9832 & n9841 ) | ( ~n9833 & n9841 ) ;
  assign n9843 = n9838 | n9842 ;
  assign n9844 = ( n132 & ~n9821 ) | ( n132 & n9834 ) | ( ~n9821 & n9834 ) ;
  assign n9845 = n132 & ~n9821 ;
  assign n9846 = ( n9826 & ~n9844 ) | ( n9826 & n9845 ) | ( ~n9844 & n9845 ) ;
  assign n9847 = ( n9826 & n9844 ) | ( n9826 & n9845 ) | ( n9844 & n9845 ) ;
  assign n9848 = ( n9844 & n9846 ) | ( n9844 & ~n9847 ) | ( n9846 & ~n9847 ) ;
  assign n9849 = x12 | x13 ;
  assign n9850 = x14 | n9849 ;
  assign n9851 = ~n9497 & n9850 ;
  assign n9852 = ( x15 & ~n9834 ) | ( x15 & n9851 ) | ( ~n9834 & n9851 ) ;
  assign n9853 = n9497 & ~n9850 ;
  assign n9854 = ~n9504 & n9834 ;
  assign n9855 = ( n9852 & ~n9853 ) | ( n9852 & n9854 ) | ( ~n9853 & n9854 ) ;
  assign n9856 = n9497 & ~n9834 ;
  assign n9857 = ( x16 & n9854 ) | ( x16 & n9856 ) | ( n9854 & n9856 ) ;
  assign n9858 = ( ~x16 & n9854 ) | ( ~x16 & n9856 ) | ( n9854 & n9856 ) ;
  assign n9859 = ( x16 & ~n9857 ) | ( x16 & n9858 ) | ( ~n9857 & n9858 ) ;
  assign n9860 = ( ~n9167 & n9855 ) | ( ~n9167 & n9859 ) | ( n9855 & n9859 ) ;
  assign n9861 = ~n9167 & n9497 ;
  assign n9862 = ( n9511 & n9834 ) | ( n9511 & n9861 ) | ( n9834 & n9861 ) ;
  assign n9863 = ( ~x17 & n9858 ) | ( ~x17 & n9862 ) | ( n9858 & n9862 ) ;
  assign n9864 = ( x17 & n9858 ) | ( x17 & n9862 ) | ( n9858 & n9862 ) ;
  assign n9865 = ( x17 & n9863 ) | ( x17 & ~n9864 ) | ( n9863 & ~n9864 ) ;
  assign n9866 = ( ~n8838 & n9860 ) | ( ~n8838 & n9865 ) | ( n9860 & n9865 ) ;
  assign n9867 = ( n8838 & ~n9510 ) | ( n8838 & n9834 ) | ( ~n9510 & n9834 ) ;
  assign n9868 = n8838 & ~n9510 ;
  assign n9869 = ( n9514 & n9867 ) | ( n9514 & n9868 ) | ( n9867 & n9868 ) ;
  assign n9870 = ( ~n9514 & n9867 ) | ( ~n9514 & n9868 ) | ( n9867 & n9868 ) ;
  assign n9871 = ( n9514 & ~n9869 ) | ( n9514 & n9870 ) | ( ~n9869 & n9870 ) ;
  assign n9872 = ( ~n8517 & n9866 ) | ( ~n8517 & n9871 ) | ( n9866 & n9871 ) ;
  assign n9873 = ( n8517 & ~n9515 ) | ( n8517 & n9834 ) | ( ~n9515 & n9834 ) ;
  assign n9874 = n8517 & ~n9515 ;
  assign n9875 = ( n9520 & n9873 ) | ( n9520 & n9874 ) | ( n9873 & n9874 ) ;
  assign n9876 = ( ~n9520 & n9873 ) | ( ~n9520 & n9874 ) | ( n9873 & n9874 ) ;
  assign n9877 = ( n9520 & ~n9875 ) | ( n9520 & n9876 ) | ( ~n9875 & n9876 ) ;
  assign n9878 = ( ~n8201 & n9872 ) | ( ~n8201 & n9877 ) | ( n9872 & n9877 ) ;
  assign n9879 = ( n8201 & ~n9521 ) | ( n8201 & n9834 ) | ( ~n9521 & n9834 ) ;
  assign n9880 = n8201 & ~n9521 ;
  assign n9881 = ( n9526 & n9879 ) | ( n9526 & n9880 ) | ( n9879 & n9880 ) ;
  assign n9882 = ( ~n9526 & n9879 ) | ( ~n9526 & n9880 ) | ( n9879 & n9880 ) ;
  assign n9883 = ( n9526 & ~n9881 ) | ( n9526 & n9882 ) | ( ~n9881 & n9882 ) ;
  assign n9884 = ( ~n7897 & n9878 ) | ( ~n7897 & n9883 ) | ( n9878 & n9883 ) ;
  assign n9885 = ( n7897 & ~n9527 ) | ( n7897 & n9834 ) | ( ~n9527 & n9834 ) ;
  assign n9886 = n7897 & ~n9527 ;
  assign n9887 = ( n9532 & n9885 ) | ( n9532 & n9886 ) | ( n9885 & n9886 ) ;
  assign n9888 = ( ~n9532 & n9885 ) | ( ~n9532 & n9886 ) | ( n9885 & n9886 ) ;
  assign n9889 = ( n9532 & ~n9887 ) | ( n9532 & n9888 ) | ( ~n9887 & n9888 ) ;
  assign n9890 = ( ~n7594 & n9884 ) | ( ~n7594 & n9889 ) | ( n9884 & n9889 ) ;
  assign n9891 = ~n7594 & n9533 ;
  assign n9892 = ( ~n7594 & n9533 ) | ( ~n7594 & n9834 ) | ( n9533 & n9834 ) ;
  assign n9893 = ( ~n9538 & n9891 ) | ( ~n9538 & n9892 ) | ( n9891 & n9892 ) ;
  assign n9894 = ( n9538 & n9891 ) | ( n9538 & n9892 ) | ( n9891 & n9892 ) ;
  assign n9895 = ( n9538 & n9893 ) | ( n9538 & ~n9894 ) | ( n9893 & ~n9894 ) ;
  assign n9896 = ( ~n7296 & n9890 ) | ( ~n7296 & n9895 ) | ( n9890 & n9895 ) ;
  assign n9897 = n7296 & ~n9539 ;
  assign n9898 = ( n7296 & ~n9539 ) | ( n7296 & n9834 ) | ( ~n9539 & n9834 ) ;
  assign n9899 = ( ~n9544 & n9897 ) | ( ~n9544 & n9898 ) | ( n9897 & n9898 ) ;
  assign n9900 = ( n9544 & n9897 ) | ( n9544 & n9898 ) | ( n9897 & n9898 ) ;
  assign n9901 = ( n9544 & n9899 ) | ( n9544 & ~n9900 ) | ( n9899 & ~n9900 ) ;
  assign n9902 = ( ~n7006 & n9896 ) | ( ~n7006 & n9901 ) | ( n9896 & n9901 ) ;
  assign n9903 = ~n7006 & n9545 ;
  assign n9904 = ( ~n7006 & n9545 ) | ( ~n7006 & n9834 ) | ( n9545 & n9834 ) ;
  assign n9905 = ( ~n9550 & n9903 ) | ( ~n9550 & n9904 ) | ( n9903 & n9904 ) ;
  assign n9906 = ( n9550 & n9903 ) | ( n9550 & n9904 ) | ( n9903 & n9904 ) ;
  assign n9907 = ( n9550 & n9905 ) | ( n9550 & ~n9906 ) | ( n9905 & ~n9906 ) ;
  assign n9908 = ( ~n6723 & n9902 ) | ( ~n6723 & n9907 ) | ( n9902 & n9907 ) ;
  assign n9909 = ( n6723 & ~n9551 ) | ( n6723 & n9834 ) | ( ~n9551 & n9834 ) ;
  assign n9910 = n6723 & ~n9551 ;
  assign n9911 = ( n9556 & n9909 ) | ( n9556 & n9910 ) | ( n9909 & n9910 ) ;
  assign n9912 = ( ~n9556 & n9909 ) | ( ~n9556 & n9910 ) | ( n9909 & n9910 ) ;
  assign n9913 = ( n9556 & ~n9911 ) | ( n9556 & n9912 ) | ( ~n9911 & n9912 ) ;
  assign n9914 = ( ~n6442 & n9908 ) | ( ~n6442 & n9913 ) | ( n9908 & n9913 ) ;
  assign n9915 = ~n6442 & n9557 ;
  assign n9916 = ( ~n6442 & n9557 ) | ( ~n6442 & n9834 ) | ( n9557 & n9834 ) ;
  assign n9917 = ( ~n9562 & n9915 ) | ( ~n9562 & n9916 ) | ( n9915 & n9916 ) ;
  assign n9918 = ( n9562 & n9915 ) | ( n9562 & n9916 ) | ( n9915 & n9916 ) ;
  assign n9919 = ( n9562 & n9917 ) | ( n9562 & ~n9918 ) | ( n9917 & ~n9918 ) ;
  assign n9920 = ( ~n6172 & n9914 ) | ( ~n6172 & n9919 ) | ( n9914 & n9919 ) ;
  assign n9921 = ( n6172 & ~n9563 ) | ( n6172 & n9834 ) | ( ~n9563 & n9834 ) ;
  assign n9922 = n6172 & ~n9563 ;
  assign n9923 = ( n9568 & n9921 ) | ( n9568 & n9922 ) | ( n9921 & n9922 ) ;
  assign n9924 = ( ~n9568 & n9921 ) | ( ~n9568 & n9922 ) | ( n9921 & n9922 ) ;
  assign n9925 = ( n9568 & ~n9923 ) | ( n9568 & n9924 ) | ( ~n9923 & n9924 ) ;
  assign n9926 = ( ~n5905 & n9920 ) | ( ~n5905 & n9925 ) | ( n9920 & n9925 ) ;
  assign n9927 = ~n5905 & n9569 ;
  assign n9928 = ( ~n5905 & n9569 ) | ( ~n5905 & n9834 ) | ( n9569 & n9834 ) ;
  assign n9929 = ( ~n9574 & n9927 ) | ( ~n9574 & n9928 ) | ( n9927 & n9928 ) ;
  assign n9930 = ( n9574 & n9927 ) | ( n9574 & n9928 ) | ( n9927 & n9928 ) ;
  assign n9931 = ( n9574 & n9929 ) | ( n9574 & ~n9930 ) | ( n9929 & ~n9930 ) ;
  assign n9932 = ( ~n5642 & n9926 ) | ( ~n5642 & n9931 ) | ( n9926 & n9931 ) ;
  assign n9933 = ~n5642 & n9575 ;
  assign n9934 = ( ~n5642 & n9575 ) | ( ~n5642 & n9834 ) | ( n9575 & n9834 ) ;
  assign n9935 = ( ~n9580 & n9933 ) | ( ~n9580 & n9934 ) | ( n9933 & n9934 ) ;
  assign n9936 = ( n9580 & n9933 ) | ( n9580 & n9934 ) | ( n9933 & n9934 ) ;
  assign n9937 = ( n9580 & n9935 ) | ( n9580 & ~n9936 ) | ( n9935 & ~n9936 ) ;
  assign n9938 = ( ~n5386 & n9932 ) | ( ~n5386 & n9937 ) | ( n9932 & n9937 ) ;
  assign n9939 = ~n5386 & n9581 ;
  assign n9940 = ( ~n5386 & n9581 ) | ( ~n5386 & n9834 ) | ( n9581 & n9834 ) ;
  assign n9941 = ( ~n9586 & n9939 ) | ( ~n9586 & n9940 ) | ( n9939 & n9940 ) ;
  assign n9942 = ( n9586 & n9939 ) | ( n9586 & n9940 ) | ( n9939 & n9940 ) ;
  assign n9943 = ( n9586 & n9941 ) | ( n9586 & ~n9942 ) | ( n9941 & ~n9942 ) ;
  assign n9944 = ( ~n5139 & n9938 ) | ( ~n5139 & n9943 ) | ( n9938 & n9943 ) ;
  assign n9945 = ~n5139 & n9587 ;
  assign n9946 = ( ~n5139 & n9587 ) | ( ~n5139 & n9834 ) | ( n9587 & n9834 ) ;
  assign n9947 = ( ~n9592 & n9945 ) | ( ~n9592 & n9946 ) | ( n9945 & n9946 ) ;
  assign n9948 = ( n9592 & n9945 ) | ( n9592 & n9946 ) | ( n9945 & n9946 ) ;
  assign n9949 = ( n9592 & n9947 ) | ( n9592 & ~n9948 ) | ( n9947 & ~n9948 ) ;
  assign n9950 = ( ~n4898 & n9944 ) | ( ~n4898 & n9949 ) | ( n9944 & n9949 ) ;
  assign n9951 = ( n4898 & ~n9593 ) | ( n4898 & n9834 ) | ( ~n9593 & n9834 ) ;
  assign n9952 = n4898 & ~n9593 ;
  assign n9953 = ( n9598 & n9951 ) | ( n9598 & n9952 ) | ( n9951 & n9952 ) ;
  assign n9954 = ( ~n9598 & n9951 ) | ( ~n9598 & n9952 ) | ( n9951 & n9952 ) ;
  assign n9955 = ( n9598 & ~n9953 ) | ( n9598 & n9954 ) | ( ~n9953 & n9954 ) ;
  assign n9956 = ( ~n4661 & n9950 ) | ( ~n4661 & n9955 ) | ( n9950 & n9955 ) ;
  assign n9957 = ~n4661 & n9599 ;
  assign n9958 = ( ~n4661 & n9599 ) | ( ~n4661 & n9834 ) | ( n9599 & n9834 ) ;
  assign n9959 = ( ~n9604 & n9957 ) | ( ~n9604 & n9958 ) | ( n9957 & n9958 ) ;
  assign n9960 = ( n9604 & n9957 ) | ( n9604 & n9958 ) | ( n9957 & n9958 ) ;
  assign n9961 = ( n9604 & n9959 ) | ( n9604 & ~n9960 ) | ( n9959 & ~n9960 ) ;
  assign n9962 = ( ~n4432 & n9956 ) | ( ~n4432 & n9961 ) | ( n9956 & n9961 ) ;
  assign n9963 = ~n4432 & n9605 ;
  assign n9964 = ( ~n4432 & n9605 ) | ( ~n4432 & n9834 ) | ( n9605 & n9834 ) ;
  assign n9965 = ( n9610 & n9963 ) | ( n9610 & n9964 ) | ( n9963 & n9964 ) ;
  assign n9966 = ( ~n9610 & n9963 ) | ( ~n9610 & n9964 ) | ( n9963 & n9964 ) ;
  assign n9967 = ( n9610 & ~n9965 ) | ( n9610 & n9966 ) | ( ~n9965 & n9966 ) ;
  assign n9968 = ( ~n4203 & n9962 ) | ( ~n4203 & n9967 ) | ( n9962 & n9967 ) ;
  assign n9969 = ~n4203 & n9611 ;
  assign n9970 = ( ~n4203 & n9611 ) | ( ~n4203 & n9834 ) | ( n9611 & n9834 ) ;
  assign n9971 = ( ~n9616 & n9969 ) | ( ~n9616 & n9970 ) | ( n9969 & n9970 ) ;
  assign n9972 = ( n9616 & n9969 ) | ( n9616 & n9970 ) | ( n9969 & n9970 ) ;
  assign n9973 = ( n9616 & n9971 ) | ( n9616 & ~n9972 ) | ( n9971 & ~n9972 ) ;
  assign n9974 = ( ~n3985 & n9968 ) | ( ~n3985 & n9973 ) | ( n9968 & n9973 ) ;
  assign n9975 = ( n3985 & ~n9617 ) | ( n3985 & n9834 ) | ( ~n9617 & n9834 ) ;
  assign n9976 = n3985 & ~n9617 ;
  assign n9977 = ( n9622 & n9975 ) | ( n9622 & n9976 ) | ( n9975 & n9976 ) ;
  assign n9978 = ( ~n9622 & n9975 ) | ( ~n9622 & n9976 ) | ( n9975 & n9976 ) ;
  assign n9979 = ( n9622 & ~n9977 ) | ( n9622 & n9978 ) | ( ~n9977 & n9978 ) ;
  assign n9980 = ( ~n3772 & n9974 ) | ( ~n3772 & n9979 ) | ( n9974 & n9979 ) ;
  assign n9981 = ( n3772 & ~n9623 ) | ( n3772 & n9834 ) | ( ~n9623 & n9834 ) ;
  assign n9982 = n3772 & ~n9623 ;
  assign n9983 = ( n9628 & n9981 ) | ( n9628 & n9982 ) | ( n9981 & n9982 ) ;
  assign n9984 = ( ~n9628 & n9981 ) | ( ~n9628 & n9982 ) | ( n9981 & n9982 ) ;
  assign n9985 = ( n9628 & ~n9983 ) | ( n9628 & n9984 ) | ( ~n9983 & n9984 ) ;
  assign n9986 = ( ~n3567 & n9980 ) | ( ~n3567 & n9985 ) | ( n9980 & n9985 ) ;
  assign n9987 = ( n3567 & ~n9629 ) | ( n3567 & n9834 ) | ( ~n9629 & n9834 ) ;
  assign n9988 = n3567 & ~n9629 ;
  assign n9989 = ( n9634 & n9987 ) | ( n9634 & n9988 ) | ( n9987 & n9988 ) ;
  assign n9990 = ( ~n9634 & n9987 ) | ( ~n9634 & n9988 ) | ( n9987 & n9988 ) ;
  assign n9991 = ( n9634 & ~n9989 ) | ( n9634 & n9990 ) | ( ~n9989 & n9990 ) ;
  assign n9992 = ( ~n3362 & n9986 ) | ( ~n3362 & n9991 ) | ( n9986 & n9991 ) ;
  assign n9993 = ~n3362 & n9635 ;
  assign n9994 = ( ~n3362 & n9635 ) | ( ~n3362 & n9834 ) | ( n9635 & n9834 ) ;
  assign n9995 = ( ~n9640 & n9993 ) | ( ~n9640 & n9994 ) | ( n9993 & n9994 ) ;
  assign n9996 = ( n9640 & n9993 ) | ( n9640 & n9994 ) | ( n9993 & n9994 ) ;
  assign n9997 = ( n9640 & n9995 ) | ( n9640 & ~n9996 ) | ( n9995 & ~n9996 ) ;
  assign n9998 = ( ~n3169 & n9992 ) | ( ~n3169 & n9997 ) | ( n9992 & n9997 ) ;
  assign n9999 = ~n3169 & n9641 ;
  assign n10000 = ( ~n3169 & n9641 ) | ( ~n3169 & n9834 ) | ( n9641 & n9834 ) ;
  assign n10001 = ( ~n9646 & n9999 ) | ( ~n9646 & n10000 ) | ( n9999 & n10000 ) ;
  assign n10002 = ( n9646 & n9999 ) | ( n9646 & n10000 ) | ( n9999 & n10000 ) ;
  assign n10003 = ( n9646 & n10001 ) | ( n9646 & ~n10002 ) | ( n10001 & ~n10002 ) ;
  assign n10004 = ( ~n2979 & n9998 ) | ( ~n2979 & n10003 ) | ( n9998 & n10003 ) ;
  assign n10005 = n2979 & ~n9647 ;
  assign n10006 = ( n2979 & ~n9647 ) | ( n2979 & n9834 ) | ( ~n9647 & n9834 ) ;
  assign n10007 = ( ~n9652 & n10005 ) | ( ~n9652 & n10006 ) | ( n10005 & n10006 ) ;
  assign n10008 = ( n9652 & n10005 ) | ( n9652 & n10006 ) | ( n10005 & n10006 ) ;
  assign n10009 = ( n9652 & n10007 ) | ( n9652 & ~n10008 ) | ( n10007 & ~n10008 ) ;
  assign n10010 = ( ~n2791 & n10004 ) | ( ~n2791 & n10009 ) | ( n10004 & n10009 ) ;
  assign n10011 = ( n2791 & ~n9653 ) | ( n2791 & n9834 ) | ( ~n9653 & n9834 ) ;
  assign n10012 = n2791 & ~n9653 ;
  assign n10013 = ( n9658 & n10011 ) | ( n9658 & n10012 ) | ( n10011 & n10012 ) ;
  assign n10014 = ( ~n9658 & n10011 ) | ( ~n9658 & n10012 ) | ( n10011 & n10012 ) ;
  assign n10015 = ( n9658 & ~n10013 ) | ( n9658 & n10014 ) | ( ~n10013 & n10014 ) ;
  assign n10016 = ( ~n2615 & n10010 ) | ( ~n2615 & n10015 ) | ( n10010 & n10015 ) ;
  assign n10017 = ~n2615 & n9659 ;
  assign n10018 = ( ~n2615 & n9659 ) | ( ~n2615 & n9834 ) | ( n9659 & n9834 ) ;
  assign n10019 = ( n9664 & n10017 ) | ( n9664 & n10018 ) | ( n10017 & n10018 ) ;
  assign n10020 = ( ~n9664 & n10017 ) | ( ~n9664 & n10018 ) | ( n10017 & n10018 ) ;
  assign n10021 = ( n9664 & ~n10019 ) | ( n9664 & n10020 ) | ( ~n10019 & n10020 ) ;
  assign n10022 = ( ~n2443 & n10016 ) | ( ~n2443 & n10021 ) | ( n10016 & n10021 ) ;
  assign n10023 = n2443 & ~n9665 ;
  assign n10024 = ( n2443 & ~n9665 ) | ( n2443 & n9834 ) | ( ~n9665 & n9834 ) ;
  assign n10025 = ( n9670 & n10023 ) | ( n9670 & n10024 ) | ( n10023 & n10024 ) ;
  assign n10026 = ( ~n9670 & n10023 ) | ( ~n9670 & n10024 ) | ( n10023 & n10024 ) ;
  assign n10027 = ( n9670 & ~n10025 ) | ( n9670 & n10026 ) | ( ~n10025 & n10026 ) ;
  assign n10028 = ( ~n2277 & n10022 ) | ( ~n2277 & n10027 ) | ( n10022 & n10027 ) ;
  assign n10029 = ( n2277 & ~n9671 ) | ( n2277 & n9834 ) | ( ~n9671 & n9834 ) ;
  assign n10030 = n2277 & ~n9671 ;
  assign n10031 = ( n9676 & n10029 ) | ( n9676 & n10030 ) | ( n10029 & n10030 ) ;
  assign n10032 = ( ~n9676 & n10029 ) | ( ~n9676 & n10030 ) | ( n10029 & n10030 ) ;
  assign n10033 = ( n9676 & ~n10031 ) | ( n9676 & n10032 ) | ( ~n10031 & n10032 ) ;
  assign n10034 = ( ~n2111 & n10028 ) | ( ~n2111 & n10033 ) | ( n10028 & n10033 ) ;
  assign n10035 = ( n2111 & ~n9677 ) | ( n2111 & n9834 ) | ( ~n9677 & n9834 ) ;
  assign n10036 = n2111 & ~n9677 ;
  assign n10037 = ( n9682 & n10035 ) | ( n9682 & n10036 ) | ( n10035 & n10036 ) ;
  assign n10038 = ( ~n9682 & n10035 ) | ( ~n9682 & n10036 ) | ( n10035 & n10036 ) ;
  assign n10039 = ( n9682 & ~n10037 ) | ( n9682 & n10038 ) | ( ~n10037 & n10038 ) ;
  assign n10040 = ( ~n1949 & n10034 ) | ( ~n1949 & n10039 ) | ( n10034 & n10039 ) ;
  assign n10041 = ~n1949 & n9683 ;
  assign n10042 = ( ~n1949 & n9683 ) | ( ~n1949 & n9834 ) | ( n9683 & n9834 ) ;
  assign n10043 = ( ~n9688 & n10041 ) | ( ~n9688 & n10042 ) | ( n10041 & n10042 ) ;
  assign n10044 = ( n9688 & n10041 ) | ( n9688 & n10042 ) | ( n10041 & n10042 ) ;
  assign n10045 = ( n9688 & n10043 ) | ( n9688 & ~n10044 ) | ( n10043 & ~n10044 ) ;
  assign n10046 = ( ~n1802 & n10040 ) | ( ~n1802 & n10045 ) | ( n10040 & n10045 ) ;
  assign n10047 = ( n1802 & ~n9689 ) | ( n1802 & n9834 ) | ( ~n9689 & n9834 ) ;
  assign n10048 = n1802 & ~n9689 ;
  assign n10049 = ( n9694 & n10047 ) | ( n9694 & n10048 ) | ( n10047 & n10048 ) ;
  assign n10050 = ( ~n9694 & n10047 ) | ( ~n9694 & n10048 ) | ( n10047 & n10048 ) ;
  assign n10051 = ( n9694 & ~n10049 ) | ( n9694 & n10050 ) | ( ~n10049 & n10050 ) ;
  assign n10052 = ( ~n1661 & n10046 ) | ( ~n1661 & n10051 ) | ( n10046 & n10051 ) ;
  assign n10053 = n1661 & ~n9695 ;
  assign n10054 = ( n1661 & ~n9695 ) | ( n1661 & n9834 ) | ( ~n9695 & n9834 ) ;
  assign n10055 = ( ~n9700 & n10053 ) | ( ~n9700 & n10054 ) | ( n10053 & n10054 ) ;
  assign n10056 = ( n9700 & n10053 ) | ( n9700 & n10054 ) | ( n10053 & n10054 ) ;
  assign n10057 = ( n9700 & n10055 ) | ( n9700 & ~n10056 ) | ( n10055 & ~n10056 ) ;
  assign n10058 = ( ~n1523 & n10052 ) | ( ~n1523 & n10057 ) | ( n10052 & n10057 ) ;
  assign n10059 = ( n1523 & ~n9701 ) | ( n1523 & n9834 ) | ( ~n9701 & n9834 ) ;
  assign n10060 = n1523 & ~n9701 ;
  assign n10061 = ( n9706 & n10059 ) | ( n9706 & n10060 ) | ( n10059 & n10060 ) ;
  assign n10062 = ( ~n9706 & n10059 ) | ( ~n9706 & n10060 ) | ( n10059 & n10060 ) ;
  assign n10063 = ( n9706 & ~n10061 ) | ( n9706 & n10062 ) | ( ~n10061 & n10062 ) ;
  assign n10064 = ( ~n1393 & n10058 ) | ( ~n1393 & n10063 ) | ( n10058 & n10063 ) ;
  assign n10065 = ( n1393 & ~n9707 ) | ( n1393 & n9834 ) | ( ~n9707 & n9834 ) ;
  assign n10066 = n1393 & ~n9707 ;
  assign n10067 = ( n9712 & n10065 ) | ( n9712 & n10066 ) | ( n10065 & n10066 ) ;
  assign n10068 = ( ~n9712 & n10065 ) | ( ~n9712 & n10066 ) | ( n10065 & n10066 ) ;
  assign n10069 = ( n9712 & ~n10067 ) | ( n9712 & n10068 ) | ( ~n10067 & n10068 ) ;
  assign n10070 = ( ~n1266 & n10064 ) | ( ~n1266 & n10069 ) | ( n10064 & n10069 ) ;
  assign n10071 = ( n1266 & ~n9713 ) | ( n1266 & n9834 ) | ( ~n9713 & n9834 ) ;
  assign n10072 = n1266 & ~n9713 ;
  assign n10073 = ( n9718 & n10071 ) | ( n9718 & n10072 ) | ( n10071 & n10072 ) ;
  assign n10074 = ( ~n9718 & n10071 ) | ( ~n9718 & n10072 ) | ( n10071 & n10072 ) ;
  assign n10075 = ( n9718 & ~n10073 ) | ( n9718 & n10074 ) | ( ~n10073 & n10074 ) ;
  assign n10076 = ( ~n1150 & n10070 ) | ( ~n1150 & n10075 ) | ( n10070 & n10075 ) ;
  assign n10077 = ~n1150 & n9719 ;
  assign n10078 = ( ~n1150 & n9719 ) | ( ~n1150 & n9834 ) | ( n9719 & n9834 ) ;
  assign n10079 = ( ~n9724 & n10077 ) | ( ~n9724 & n10078 ) | ( n10077 & n10078 ) ;
  assign n10080 = ( n9724 & n10077 ) | ( n9724 & n10078 ) | ( n10077 & n10078 ) ;
  assign n10081 = ( n9724 & n10079 ) | ( n9724 & ~n10080 ) | ( n10079 & ~n10080 ) ;
  assign n10082 = ( ~n1038 & n10076 ) | ( ~n1038 & n10081 ) | ( n10076 & n10081 ) ;
  assign n10083 = ~n1038 & n9725 ;
  assign n10084 = ( ~n1038 & n9725 ) | ( ~n1038 & n9834 ) | ( n9725 & n9834 ) ;
  assign n10085 = ( ~n9730 & n10083 ) | ( ~n9730 & n10084 ) | ( n10083 & n10084 ) ;
  assign n10086 = ( n9730 & n10083 ) | ( n9730 & n10084 ) | ( n10083 & n10084 ) ;
  assign n10087 = ( n9730 & n10085 ) | ( n9730 & ~n10086 ) | ( n10085 & ~n10086 ) ;
  assign n10088 = ( ~n933 & n10082 ) | ( ~n933 & n10087 ) | ( n10082 & n10087 ) ;
  assign n10089 = ~n933 & n9731 ;
  assign n10090 = ( ~n933 & n9731 ) | ( ~n933 & n9834 ) | ( n9731 & n9834 ) ;
  assign n10091 = ( ~n9736 & n10089 ) | ( ~n9736 & n10090 ) | ( n10089 & n10090 ) ;
  assign n10092 = ( n9736 & n10089 ) | ( n9736 & n10090 ) | ( n10089 & n10090 ) ;
  assign n10093 = ( n9736 & n10091 ) | ( n9736 & ~n10092 ) | ( n10091 & ~n10092 ) ;
  assign n10094 = ( ~n839 & n10088 ) | ( ~n839 & n10093 ) | ( n10088 & n10093 ) ;
  assign n10095 = n839 & ~n9737 ;
  assign n10096 = ( n839 & ~n9737 ) | ( n839 & n9834 ) | ( ~n9737 & n9834 ) ;
  assign n10097 = ( ~n9742 & n10095 ) | ( ~n9742 & n10096 ) | ( n10095 & n10096 ) ;
  assign n10098 = ( n9742 & n10095 ) | ( n9742 & n10096 ) | ( n10095 & n10096 ) ;
  assign n10099 = ( n9742 & n10097 ) | ( n9742 & ~n10098 ) | ( n10097 & ~n10098 ) ;
  assign n10100 = ( ~n746 & n10094 ) | ( ~n746 & n10099 ) | ( n10094 & n10099 ) ;
  assign n10101 = ( n746 & ~n9743 ) | ( n746 & n9834 ) | ( ~n9743 & n9834 ) ;
  assign n10102 = n746 & ~n9743 ;
  assign n10103 = ( n9748 & n10101 ) | ( n9748 & n10102 ) | ( n10101 & n10102 ) ;
  assign n10104 = ( ~n9748 & n10101 ) | ( ~n9748 & n10102 ) | ( n10101 & n10102 ) ;
  assign n10105 = ( n9748 & ~n10103 ) | ( n9748 & n10104 ) | ( ~n10103 & n10104 ) ;
  assign n10106 = ( ~n664 & n10100 ) | ( ~n664 & n10105 ) | ( n10100 & n10105 ) ;
  assign n10107 = ( n664 & ~n9749 ) | ( n664 & n9834 ) | ( ~n9749 & n9834 ) ;
  assign n10108 = n664 & ~n9749 ;
  assign n10109 = ( n9754 & n10107 ) | ( n9754 & n10108 ) | ( n10107 & n10108 ) ;
  assign n10110 = ( ~n9754 & n10107 ) | ( ~n9754 & n10108 ) | ( n10107 & n10108 ) ;
  assign n10111 = ( n9754 & ~n10109 ) | ( n9754 & n10110 ) | ( ~n10109 & n10110 ) ;
  assign n10112 = ( ~n588 & n10106 ) | ( ~n588 & n10111 ) | ( n10106 & n10111 ) ;
  assign n10113 = ( n588 & ~n9755 ) | ( n588 & n9834 ) | ( ~n9755 & n9834 ) ;
  assign n10114 = n588 & ~n9755 ;
  assign n10115 = ( n9760 & n10113 ) | ( n9760 & n10114 ) | ( n10113 & n10114 ) ;
  assign n10116 = ( ~n9760 & n10113 ) | ( ~n9760 & n10114 ) | ( n10113 & n10114 ) ;
  assign n10117 = ( n9760 & ~n10115 ) | ( n9760 & n10116 ) | ( ~n10115 & n10116 ) ;
  assign n10118 = ( ~n518 & n10112 ) | ( ~n518 & n10117 ) | ( n10112 & n10117 ) ;
  assign n10119 = n518 & ~n9761 ;
  assign n10120 = ( n518 & ~n9761 ) | ( n518 & n9834 ) | ( ~n9761 & n9834 ) ;
  assign n10121 = ( ~n9766 & n10119 ) | ( ~n9766 & n10120 ) | ( n10119 & n10120 ) ;
  assign n10122 = ( n9766 & n10119 ) | ( n9766 & n10120 ) | ( n10119 & n10120 ) ;
  assign n10123 = ( n9766 & n10121 ) | ( n9766 & ~n10122 ) | ( n10121 & ~n10122 ) ;
  assign n10124 = ( ~n454 & n10118 ) | ( ~n454 & n10123 ) | ( n10118 & n10123 ) ;
  assign n10125 = ~n454 & n9767 ;
  assign n10126 = ( ~n454 & n9767 ) | ( ~n454 & n9834 ) | ( n9767 & n9834 ) ;
  assign n10127 = ( ~n9772 & n10125 ) | ( ~n9772 & n10126 ) | ( n10125 & n10126 ) ;
  assign n10128 = ( n9772 & n10125 ) | ( n9772 & n10126 ) | ( n10125 & n10126 ) ;
  assign n10129 = ( n9772 & n10127 ) | ( n9772 & ~n10128 ) | ( n10127 & ~n10128 ) ;
  assign n10130 = ( ~n396 & n10124 ) | ( ~n396 & n10129 ) | ( n10124 & n10129 ) ;
  assign n10131 = n396 & ~n9773 ;
  assign n10132 = ( n396 & ~n9773 ) | ( n396 & n9834 ) | ( ~n9773 & n9834 ) ;
  assign n10133 = ( n9778 & n10131 ) | ( n9778 & n10132 ) | ( n10131 & n10132 ) ;
  assign n10134 = ( ~n9778 & n10131 ) | ( ~n9778 & n10132 ) | ( n10131 & n10132 ) ;
  assign n10135 = ( n9778 & ~n10133 ) | ( n9778 & n10134 ) | ( ~n10133 & n10134 ) ;
  assign n10136 = ( ~n344 & n10130 ) | ( ~n344 & n10135 ) | ( n10130 & n10135 ) ;
  assign n10137 = ( n344 & ~n9779 ) | ( n344 & n9834 ) | ( ~n9779 & n9834 ) ;
  assign n10138 = n344 & ~n9779 ;
  assign n10139 = ( n9784 & n10137 ) | ( n9784 & n10138 ) | ( n10137 & n10138 ) ;
  assign n10140 = ( ~n9784 & n10137 ) | ( ~n9784 & n10138 ) | ( n10137 & n10138 ) ;
  assign n10141 = ( n9784 & ~n10139 ) | ( n9784 & n10140 ) | ( ~n10139 & n10140 ) ;
  assign n10142 = ( ~n298 & n10136 ) | ( ~n298 & n10141 ) | ( n10136 & n10141 ) ;
  assign n10143 = ~n298 & n9785 ;
  assign n10144 = ( ~n298 & n9785 ) | ( ~n298 & n9834 ) | ( n9785 & n9834 ) ;
  assign n10145 = ( n9790 & n10143 ) | ( n9790 & n10144 ) | ( n10143 & n10144 ) ;
  assign n10146 = ( ~n9790 & n10143 ) | ( ~n9790 & n10144 ) | ( n10143 & n10144 ) ;
  assign n10147 = ( n9790 & ~n10145 ) | ( n9790 & n10146 ) | ( ~n10145 & n10146 ) ;
  assign n10148 = ( ~n258 & n10142 ) | ( ~n258 & n10147 ) | ( n10142 & n10147 ) ;
  assign n10149 = ( n258 & ~n9791 ) | ( n258 & n9834 ) | ( ~n9791 & n9834 ) ;
  assign n10150 = n258 & ~n9791 ;
  assign n10151 = ( n9796 & n10149 ) | ( n9796 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10152 = ( ~n9796 & n10149 ) | ( ~n9796 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10153 = ( n9796 & ~n10151 ) | ( n9796 & n10152 ) | ( ~n10151 & n10152 ) ;
  assign n10154 = ( ~n225 & n10148 ) | ( ~n225 & n10153 ) | ( n10148 & n10153 ) ;
  assign n10155 = ( n225 & ~n9797 ) | ( n225 & n9834 ) | ( ~n9797 & n9834 ) ;
  assign n10156 = n225 & ~n9797 ;
  assign n10157 = ( n9802 & n10155 ) | ( n9802 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10158 = ( ~n9802 & n10155 ) | ( ~n9802 & n10156 ) | ( n10155 & n10156 ) ;
  assign n10159 = ( n9802 & ~n10157 ) | ( n9802 & n10158 ) | ( ~n10157 & n10158 ) ;
  assign n10160 = ( ~n197 & n10154 ) | ( ~n197 & n10159 ) | ( n10154 & n10159 ) ;
  assign n10161 = ( n197 & ~n9803 ) | ( n197 & n9834 ) | ( ~n9803 & n9834 ) ;
  assign n10162 = n197 & ~n9803 ;
  assign n10163 = ( n9808 & n10161 ) | ( n9808 & n10162 ) | ( n10161 & n10162 ) ;
  assign n10164 = ( ~n9808 & n10161 ) | ( ~n9808 & n10162 ) | ( n10161 & n10162 ) ;
  assign n10165 = ( n9808 & ~n10163 ) | ( n9808 & n10164 ) | ( ~n10163 & n10164 ) ;
  assign n10166 = ( ~n170 & n10160 ) | ( ~n170 & n10165 ) | ( n10160 & n10165 ) ;
  assign n10167 = ~n170 & n9809 ;
  assign n10168 = ( ~n170 & n9809 ) | ( ~n170 & n9834 ) | ( n9809 & n9834 ) ;
  assign n10169 = ( ~n9814 & n10167 ) | ( ~n9814 & n10168 ) | ( n10167 & n10168 ) ;
  assign n10170 = ( n9814 & n10167 ) | ( n9814 & n10168 ) | ( n10167 & n10168 ) ;
  assign n10171 = ( n9814 & n10169 ) | ( n9814 & ~n10170 ) | ( n10169 & ~n10170 ) ;
  assign n10172 = ( ~n142 & n10166 ) | ( ~n142 & n10171 ) | ( n10166 & n10171 ) ;
  assign n10173 = ( n142 & ~n9815 ) | ( n142 & n9834 ) | ( ~n9815 & n9834 ) ;
  assign n10174 = n142 & ~n9815 ;
  assign n10175 = ( n9820 & n10173 ) | ( n9820 & n10174 ) | ( n10173 & n10174 ) ;
  assign n10176 = ( ~n9820 & n10173 ) | ( ~n9820 & n10174 ) | ( n10173 & n10174 ) ;
  assign n10177 = ( n9820 & ~n10175 ) | ( n9820 & n10176 ) | ( ~n10175 & n10176 ) ;
  assign n10178 = ( ~n132 & n10172 ) | ( ~n132 & n10177 ) | ( n10172 & n10177 ) ;
  assign n10179 = ( ~n131 & n9848 ) | ( ~n131 & n10178 ) | ( n9848 & n10178 ) ;
  assign n10180 = n9843 | n10179 ;
  assign n10181 = n9834 & ~n10180 ;
  assign n10182 = ~n9849 & n10180 ;
  assign n10183 = ( x14 & n10181 ) | ( x14 & n10182 ) | ( n10181 & n10182 ) ;
  assign n10184 = ( ~x14 & n10181 ) | ( ~x14 & n10182 ) | ( n10181 & n10182 ) ;
  assign n10185 = ( x14 & ~n10183 ) | ( x14 & n10184 ) | ( ~n10183 & n10184 ) ;
  assign n10186 = x10 | x11 ;
  assign n10187 = x12 | n10186 ;
  assign n10188 = n9834 & ~n10187 ;
  assign n10189 = ~n9834 & n10187 ;
  assign n10190 = ( x13 & ~n10180 ) | ( x13 & n10189 ) | ( ~n10180 & n10189 ) ;
  assign n10191 = ( n10182 & ~n10188 ) | ( n10182 & n10190 ) | ( ~n10188 & n10190 ) ;
  assign n10192 = ( ~n9497 & n10185 ) | ( ~n9497 & n10191 ) | ( n10185 & n10191 ) ;
  assign n10193 = ~n9497 & n9834 ;
  assign n10194 = ( n9856 & n10180 ) | ( n9856 & n10193 ) | ( n10180 & n10193 ) ;
  assign n10195 = ( ~x15 & n10184 ) | ( ~x15 & n10194 ) | ( n10184 & n10194 ) ;
  assign n10196 = ( x15 & n10184 ) | ( x15 & n10194 ) | ( n10184 & n10194 ) ;
  assign n10197 = ( x15 & n10195 ) | ( x15 & ~n10196 ) | ( n10195 & ~n10196 ) ;
  assign n10198 = ( ~n9167 & n10192 ) | ( ~n9167 & n10197 ) | ( n10192 & n10197 ) ;
  assign n10199 = ( n9167 & ~n9855 ) | ( n9167 & n10180 ) | ( ~n9855 & n10180 ) ;
  assign n10200 = n9167 & ~n9855 ;
  assign n10201 = ( n9859 & n10199 ) | ( n9859 & n10200 ) | ( n10199 & n10200 ) ;
  assign n10202 = ( ~n9859 & n10199 ) | ( ~n9859 & n10200 ) | ( n10199 & n10200 ) ;
  assign n10203 = ( n9859 & ~n10201 ) | ( n9859 & n10202 ) | ( ~n10201 & n10202 ) ;
  assign n10204 = ( ~n8838 & n10198 ) | ( ~n8838 & n10203 ) | ( n10198 & n10203 ) ;
  assign n10205 = ( n8838 & ~n9860 ) | ( n8838 & n10180 ) | ( ~n9860 & n10180 ) ;
  assign n10206 = n8838 & ~n9860 ;
  assign n10207 = ( n9865 & n10205 ) | ( n9865 & n10206 ) | ( n10205 & n10206 ) ;
  assign n10208 = ( ~n9865 & n10205 ) | ( ~n9865 & n10206 ) | ( n10205 & n10206 ) ;
  assign n10209 = ( n9865 & ~n10207 ) | ( n9865 & n10208 ) | ( ~n10207 & n10208 ) ;
  assign n10210 = ( ~n8517 & n10204 ) | ( ~n8517 & n10209 ) | ( n10204 & n10209 ) ;
  assign n10211 = ( n8517 & ~n9866 ) | ( n8517 & n10180 ) | ( ~n9866 & n10180 ) ;
  assign n10212 = n8517 & ~n9866 ;
  assign n10213 = ( n9871 & n10211 ) | ( n9871 & n10212 ) | ( n10211 & n10212 ) ;
  assign n10214 = ( ~n9871 & n10211 ) | ( ~n9871 & n10212 ) | ( n10211 & n10212 ) ;
  assign n10215 = ( n9871 & ~n10213 ) | ( n9871 & n10214 ) | ( ~n10213 & n10214 ) ;
  assign n10216 = ( ~n8201 & n10210 ) | ( ~n8201 & n10215 ) | ( n10210 & n10215 ) ;
  assign n10217 = n8201 & ~n9872 ;
  assign n10218 = ( n8201 & ~n9872 ) | ( n8201 & n10180 ) | ( ~n9872 & n10180 ) ;
  assign n10219 = ( n9877 & n10217 ) | ( n9877 & n10218 ) | ( n10217 & n10218 ) ;
  assign n10220 = ( ~n9877 & n10217 ) | ( ~n9877 & n10218 ) | ( n10217 & n10218 ) ;
  assign n10221 = ( n9877 & ~n10219 ) | ( n9877 & n10220 ) | ( ~n10219 & n10220 ) ;
  assign n10222 = ( ~n7897 & n10216 ) | ( ~n7897 & n10221 ) | ( n10216 & n10221 ) ;
  assign n10223 = ( n7897 & ~n9878 ) | ( n7897 & n10180 ) | ( ~n9878 & n10180 ) ;
  assign n10224 = n7897 & ~n9878 ;
  assign n10225 = ( n9883 & n10223 ) | ( n9883 & n10224 ) | ( n10223 & n10224 ) ;
  assign n10226 = ( ~n9883 & n10223 ) | ( ~n9883 & n10224 ) | ( n10223 & n10224 ) ;
  assign n10227 = ( n9883 & ~n10225 ) | ( n9883 & n10226 ) | ( ~n10225 & n10226 ) ;
  assign n10228 = ( ~n7594 & n10222 ) | ( ~n7594 & n10227 ) | ( n10222 & n10227 ) ;
  assign n10229 = ( n7594 & ~n9884 ) | ( n7594 & n10180 ) | ( ~n9884 & n10180 ) ;
  assign n10230 = n7594 & ~n9884 ;
  assign n10231 = ( n9889 & n10229 ) | ( n9889 & n10230 ) | ( n10229 & n10230 ) ;
  assign n10232 = ( ~n9889 & n10229 ) | ( ~n9889 & n10230 ) | ( n10229 & n10230 ) ;
  assign n10233 = ( n9889 & ~n10231 ) | ( n9889 & n10232 ) | ( ~n10231 & n10232 ) ;
  assign n10234 = ( ~n7296 & n10228 ) | ( ~n7296 & n10233 ) | ( n10228 & n10233 ) ;
  assign n10235 = ( n7296 & ~n9890 ) | ( n7296 & n10180 ) | ( ~n9890 & n10180 ) ;
  assign n10236 = n7296 & ~n9890 ;
  assign n10237 = ( n9895 & n10235 ) | ( n9895 & n10236 ) | ( n10235 & n10236 ) ;
  assign n10238 = ( ~n9895 & n10235 ) | ( ~n9895 & n10236 ) | ( n10235 & n10236 ) ;
  assign n10239 = ( n9895 & ~n10237 ) | ( n9895 & n10238 ) | ( ~n10237 & n10238 ) ;
  assign n10240 = ( ~n7006 & n10234 ) | ( ~n7006 & n10239 ) | ( n10234 & n10239 ) ;
  assign n10241 = ~n7006 & n9896 ;
  assign n10242 = ( ~n7006 & n9896 ) | ( ~n7006 & n10180 ) | ( n9896 & n10180 ) ;
  assign n10243 = ( ~n9901 & n10241 ) | ( ~n9901 & n10242 ) | ( n10241 & n10242 ) ;
  assign n10244 = ( n9901 & n10241 ) | ( n9901 & n10242 ) | ( n10241 & n10242 ) ;
  assign n10245 = ( n9901 & n10243 ) | ( n9901 & ~n10244 ) | ( n10243 & ~n10244 ) ;
  assign n10246 = ( ~n6723 & n10240 ) | ( ~n6723 & n10245 ) | ( n10240 & n10245 ) ;
  assign n10247 = ~n6723 & n9902 ;
  assign n10248 = ( ~n6723 & n9902 ) | ( ~n6723 & n10180 ) | ( n9902 & n10180 ) ;
  assign n10249 = ( ~n9907 & n10247 ) | ( ~n9907 & n10248 ) | ( n10247 & n10248 ) ;
  assign n10250 = ( n9907 & n10247 ) | ( n9907 & n10248 ) | ( n10247 & n10248 ) ;
  assign n10251 = ( n9907 & n10249 ) | ( n9907 & ~n10250 ) | ( n10249 & ~n10250 ) ;
  assign n10252 = ( ~n6442 & n10246 ) | ( ~n6442 & n10251 ) | ( n10246 & n10251 ) ;
  assign n10253 = ~n6442 & n9908 ;
  assign n10254 = ( ~n6442 & n9908 ) | ( ~n6442 & n10180 ) | ( n9908 & n10180 ) ;
  assign n10255 = ( ~n9913 & n10253 ) | ( ~n9913 & n10254 ) | ( n10253 & n10254 ) ;
  assign n10256 = ( n9913 & n10253 ) | ( n9913 & n10254 ) | ( n10253 & n10254 ) ;
  assign n10257 = ( n9913 & n10255 ) | ( n9913 & ~n10256 ) | ( n10255 & ~n10256 ) ;
  assign n10258 = ( ~n6172 & n10252 ) | ( ~n6172 & n10257 ) | ( n10252 & n10257 ) ;
  assign n10259 = ( n6172 & ~n9914 ) | ( n6172 & n10180 ) | ( ~n9914 & n10180 ) ;
  assign n10260 = n6172 & ~n9914 ;
  assign n10261 = ( n9919 & n10259 ) | ( n9919 & n10260 ) | ( n10259 & n10260 ) ;
  assign n10262 = ( ~n9919 & n10259 ) | ( ~n9919 & n10260 ) | ( n10259 & n10260 ) ;
  assign n10263 = ( n9919 & ~n10261 ) | ( n9919 & n10262 ) | ( ~n10261 & n10262 ) ;
  assign n10264 = ( ~n5905 & n10258 ) | ( ~n5905 & n10263 ) | ( n10258 & n10263 ) ;
  assign n10265 = n5905 & ~n9920 ;
  assign n10266 = ( n5905 & ~n9920 ) | ( n5905 & n10180 ) | ( ~n9920 & n10180 ) ;
  assign n10267 = ( n9925 & n10265 ) | ( n9925 & n10266 ) | ( n10265 & n10266 ) ;
  assign n10268 = ( ~n9925 & n10265 ) | ( ~n9925 & n10266 ) | ( n10265 & n10266 ) ;
  assign n10269 = ( n9925 & ~n10267 ) | ( n9925 & n10268 ) | ( ~n10267 & n10268 ) ;
  assign n10270 = ( ~n5642 & n10264 ) | ( ~n5642 & n10269 ) | ( n10264 & n10269 ) ;
  assign n10271 = ~n5642 & n9926 ;
  assign n10272 = ( ~n5642 & n9926 ) | ( ~n5642 & n10180 ) | ( n9926 & n10180 ) ;
  assign n10273 = ( n9931 & n10271 ) | ( n9931 & n10272 ) | ( n10271 & n10272 ) ;
  assign n10274 = ( ~n9931 & n10271 ) | ( ~n9931 & n10272 ) | ( n10271 & n10272 ) ;
  assign n10275 = ( n9931 & ~n10273 ) | ( n9931 & n10274 ) | ( ~n10273 & n10274 ) ;
  assign n10276 = ( ~n5386 & n10270 ) | ( ~n5386 & n10275 ) | ( n10270 & n10275 ) ;
  assign n10277 = ( n5386 & ~n9932 ) | ( n5386 & n10180 ) | ( ~n9932 & n10180 ) ;
  assign n10278 = n5386 & ~n9932 ;
  assign n10279 = ( n9937 & n10277 ) | ( n9937 & n10278 ) | ( n10277 & n10278 ) ;
  assign n10280 = ( ~n9937 & n10277 ) | ( ~n9937 & n10278 ) | ( n10277 & n10278 ) ;
  assign n10281 = ( n9937 & ~n10279 ) | ( n9937 & n10280 ) | ( ~n10279 & n10280 ) ;
  assign n10282 = ( ~n5139 & n10276 ) | ( ~n5139 & n10281 ) | ( n10276 & n10281 ) ;
  assign n10283 = ~n5139 & n9938 ;
  assign n10284 = ( ~n5139 & n9938 ) | ( ~n5139 & n10180 ) | ( n9938 & n10180 ) ;
  assign n10285 = ( n9943 & n10283 ) | ( n9943 & n10284 ) | ( n10283 & n10284 ) ;
  assign n10286 = ( ~n9943 & n10283 ) | ( ~n9943 & n10284 ) | ( n10283 & n10284 ) ;
  assign n10287 = ( n9943 & ~n10285 ) | ( n9943 & n10286 ) | ( ~n10285 & n10286 ) ;
  assign n10288 = ( ~n4898 & n10282 ) | ( ~n4898 & n10287 ) | ( n10282 & n10287 ) ;
  assign n10289 = n4898 & ~n9944 ;
  assign n10290 = ( n4898 & ~n9944 ) | ( n4898 & n10180 ) | ( ~n9944 & n10180 ) ;
  assign n10291 = ( n9949 & n10289 ) | ( n9949 & n10290 ) | ( n10289 & n10290 ) ;
  assign n10292 = ( ~n9949 & n10289 ) | ( ~n9949 & n10290 ) | ( n10289 & n10290 ) ;
  assign n10293 = ( n9949 & ~n10291 ) | ( n9949 & n10292 ) | ( ~n10291 & n10292 ) ;
  assign n10294 = ( ~n4661 & n10288 ) | ( ~n4661 & n10293 ) | ( n10288 & n10293 ) ;
  assign n10295 = ~n4661 & n9950 ;
  assign n10296 = ( ~n4661 & n9950 ) | ( ~n4661 & n10180 ) | ( n9950 & n10180 ) ;
  assign n10297 = ( ~n9955 & n10295 ) | ( ~n9955 & n10296 ) | ( n10295 & n10296 ) ;
  assign n10298 = ( n9955 & n10295 ) | ( n9955 & n10296 ) | ( n10295 & n10296 ) ;
  assign n10299 = ( n9955 & n10297 ) | ( n9955 & ~n10298 ) | ( n10297 & ~n10298 ) ;
  assign n10300 = ( ~n4432 & n10294 ) | ( ~n4432 & n10299 ) | ( n10294 & n10299 ) ;
  assign n10301 = ~n4432 & n9956 ;
  assign n10302 = ( ~n4432 & n9956 ) | ( ~n4432 & n10180 ) | ( n9956 & n10180 ) ;
  assign n10303 = ( n9961 & n10301 ) | ( n9961 & n10302 ) | ( n10301 & n10302 ) ;
  assign n10304 = ( ~n9961 & n10301 ) | ( ~n9961 & n10302 ) | ( n10301 & n10302 ) ;
  assign n10305 = ( n9961 & ~n10303 ) | ( n9961 & n10304 ) | ( ~n10303 & n10304 ) ;
  assign n10306 = ( ~n4203 & n10300 ) | ( ~n4203 & n10305 ) | ( n10300 & n10305 ) ;
  assign n10307 = ( n4203 & ~n9962 ) | ( n4203 & n10180 ) | ( ~n9962 & n10180 ) ;
  assign n10308 = n4203 & ~n9962 ;
  assign n10309 = ( n9967 & n10307 ) | ( n9967 & n10308 ) | ( n10307 & n10308 ) ;
  assign n10310 = ( ~n9967 & n10307 ) | ( ~n9967 & n10308 ) | ( n10307 & n10308 ) ;
  assign n10311 = ( n9967 & ~n10309 ) | ( n9967 & n10310 ) | ( ~n10309 & n10310 ) ;
  assign n10312 = ( ~n3985 & n10306 ) | ( ~n3985 & n10311 ) | ( n10306 & n10311 ) ;
  assign n10313 = ( n3985 & ~n9968 ) | ( n3985 & n10180 ) | ( ~n9968 & n10180 ) ;
  assign n10314 = n3985 & ~n9968 ;
  assign n10315 = ( n9973 & n10313 ) | ( n9973 & n10314 ) | ( n10313 & n10314 ) ;
  assign n10316 = ( ~n9973 & n10313 ) | ( ~n9973 & n10314 ) | ( n10313 & n10314 ) ;
  assign n10317 = ( n9973 & ~n10315 ) | ( n9973 & n10316 ) | ( ~n10315 & n10316 ) ;
  assign n10318 = ( ~n3772 & n10312 ) | ( ~n3772 & n10317 ) | ( n10312 & n10317 ) ;
  assign n10319 = ( n3772 & ~n9974 ) | ( n3772 & n10180 ) | ( ~n9974 & n10180 ) ;
  assign n10320 = n3772 & ~n9974 ;
  assign n10321 = ( n9979 & n10319 ) | ( n9979 & n10320 ) | ( n10319 & n10320 ) ;
  assign n10322 = ( ~n9979 & n10319 ) | ( ~n9979 & n10320 ) | ( n10319 & n10320 ) ;
  assign n10323 = ( n9979 & ~n10321 ) | ( n9979 & n10322 ) | ( ~n10321 & n10322 ) ;
  assign n10324 = ( ~n3567 & n10318 ) | ( ~n3567 & n10323 ) | ( n10318 & n10323 ) ;
  assign n10325 = ~n3567 & n9980 ;
  assign n10326 = ( ~n3567 & n9980 ) | ( ~n3567 & n10180 ) | ( n9980 & n10180 ) ;
  assign n10327 = ( n9985 & n10325 ) | ( n9985 & n10326 ) | ( n10325 & n10326 ) ;
  assign n10328 = ( ~n9985 & n10325 ) | ( ~n9985 & n10326 ) | ( n10325 & n10326 ) ;
  assign n10329 = ( n9985 & ~n10327 ) | ( n9985 & n10328 ) | ( ~n10327 & n10328 ) ;
  assign n10330 = ( ~n3362 & n10324 ) | ( ~n3362 & n10329 ) | ( n10324 & n10329 ) ;
  assign n10331 = ( n3362 & ~n9986 ) | ( n3362 & n10180 ) | ( ~n9986 & n10180 ) ;
  assign n10332 = n3362 & ~n9986 ;
  assign n10333 = ( n9991 & n10331 ) | ( n9991 & n10332 ) | ( n10331 & n10332 ) ;
  assign n10334 = ( ~n9991 & n10331 ) | ( ~n9991 & n10332 ) | ( n10331 & n10332 ) ;
  assign n10335 = ( n9991 & ~n10333 ) | ( n9991 & n10334 ) | ( ~n10333 & n10334 ) ;
  assign n10336 = ( ~n3169 & n10330 ) | ( ~n3169 & n10335 ) | ( n10330 & n10335 ) ;
  assign n10337 = ( n3169 & ~n9992 ) | ( n3169 & n10180 ) | ( ~n9992 & n10180 ) ;
  assign n10338 = n3169 & ~n9992 ;
  assign n10339 = ( n9997 & n10337 ) | ( n9997 & n10338 ) | ( n10337 & n10338 ) ;
  assign n10340 = ( ~n9997 & n10337 ) | ( ~n9997 & n10338 ) | ( n10337 & n10338 ) ;
  assign n10341 = ( n9997 & ~n10339 ) | ( n9997 & n10340 ) | ( ~n10339 & n10340 ) ;
  assign n10342 = ( ~n2979 & n10336 ) | ( ~n2979 & n10341 ) | ( n10336 & n10341 ) ;
  assign n10343 = ~n2979 & n9998 ;
  assign n10344 = ( ~n2979 & n9998 ) | ( ~n2979 & n10180 ) | ( n9998 & n10180 ) ;
  assign n10345 = ( n10003 & n10343 ) | ( n10003 & n10344 ) | ( n10343 & n10344 ) ;
  assign n10346 = ( ~n10003 & n10343 ) | ( ~n10003 & n10344 ) | ( n10343 & n10344 ) ;
  assign n10347 = ( n10003 & ~n10345 ) | ( n10003 & n10346 ) | ( ~n10345 & n10346 ) ;
  assign n10348 = ( ~n2791 & n10342 ) | ( ~n2791 & n10347 ) | ( n10342 & n10347 ) ;
  assign n10349 = ( n2791 & ~n10004 ) | ( n2791 & n10180 ) | ( ~n10004 & n10180 ) ;
  assign n10350 = n2791 & ~n10004 ;
  assign n10351 = ( n10009 & n10349 ) | ( n10009 & n10350 ) | ( n10349 & n10350 ) ;
  assign n10352 = ( ~n10009 & n10349 ) | ( ~n10009 & n10350 ) | ( n10349 & n10350 ) ;
  assign n10353 = ( n10009 & ~n10351 ) | ( n10009 & n10352 ) | ( ~n10351 & n10352 ) ;
  assign n10354 = ( ~n2615 & n10348 ) | ( ~n2615 & n10353 ) | ( n10348 & n10353 ) ;
  assign n10355 = ( n2615 & ~n10010 ) | ( n2615 & n10180 ) | ( ~n10010 & n10180 ) ;
  assign n10356 = n2615 & ~n10010 ;
  assign n10357 = ( n10015 & n10355 ) | ( n10015 & n10356 ) | ( n10355 & n10356 ) ;
  assign n10358 = ( ~n10015 & n10355 ) | ( ~n10015 & n10356 ) | ( n10355 & n10356 ) ;
  assign n10359 = ( n10015 & ~n10357 ) | ( n10015 & n10358 ) | ( ~n10357 & n10358 ) ;
  assign n10360 = ( ~n2443 & n10354 ) | ( ~n2443 & n10359 ) | ( n10354 & n10359 ) ;
  assign n10361 = ( n2443 & ~n10016 ) | ( n2443 & n10180 ) | ( ~n10016 & n10180 ) ;
  assign n10362 = n2443 & ~n10016 ;
  assign n10363 = ( n10021 & n10361 ) | ( n10021 & n10362 ) | ( n10361 & n10362 ) ;
  assign n10364 = ( ~n10021 & n10361 ) | ( ~n10021 & n10362 ) | ( n10361 & n10362 ) ;
  assign n10365 = ( n10021 & ~n10363 ) | ( n10021 & n10364 ) | ( ~n10363 & n10364 ) ;
  assign n10366 = ( ~n2277 & n10360 ) | ( ~n2277 & n10365 ) | ( n10360 & n10365 ) ;
  assign n10367 = ~n2277 & n10022 ;
  assign n10368 = ( ~n2277 & n10022 ) | ( ~n2277 & n10180 ) | ( n10022 & n10180 ) ;
  assign n10369 = ( n10027 & n10367 ) | ( n10027 & n10368 ) | ( n10367 & n10368 ) ;
  assign n10370 = ( ~n10027 & n10367 ) | ( ~n10027 & n10368 ) | ( n10367 & n10368 ) ;
  assign n10371 = ( n10027 & ~n10369 ) | ( n10027 & n10370 ) | ( ~n10369 & n10370 ) ;
  assign n10372 = ( ~n2111 & n10366 ) | ( ~n2111 & n10371 ) | ( n10366 & n10371 ) ;
  assign n10373 = ( n2111 & ~n10028 ) | ( n2111 & n10180 ) | ( ~n10028 & n10180 ) ;
  assign n10374 = n2111 & ~n10028 ;
  assign n10375 = ( n10033 & n10373 ) | ( n10033 & n10374 ) | ( n10373 & n10374 ) ;
  assign n10376 = ( ~n10033 & n10373 ) | ( ~n10033 & n10374 ) | ( n10373 & n10374 ) ;
  assign n10377 = ( n10033 & ~n10375 ) | ( n10033 & n10376 ) | ( ~n10375 & n10376 ) ;
  assign n10378 = ( ~n1949 & n10372 ) | ( ~n1949 & n10377 ) | ( n10372 & n10377 ) ;
  assign n10379 = ( n1949 & ~n10034 ) | ( n1949 & n10180 ) | ( ~n10034 & n10180 ) ;
  assign n10380 = n1949 & ~n10034 ;
  assign n10381 = ( n10039 & n10379 ) | ( n10039 & n10380 ) | ( n10379 & n10380 ) ;
  assign n10382 = ( ~n10039 & n10379 ) | ( ~n10039 & n10380 ) | ( n10379 & n10380 ) ;
  assign n10383 = ( n10039 & ~n10381 ) | ( n10039 & n10382 ) | ( ~n10381 & n10382 ) ;
  assign n10384 = ( ~n1802 & n10378 ) | ( ~n1802 & n10383 ) | ( n10378 & n10383 ) ;
  assign n10385 = ( n1802 & ~n10040 ) | ( n1802 & n10180 ) | ( ~n10040 & n10180 ) ;
  assign n10386 = n1802 & ~n10040 ;
  assign n10387 = ( n10045 & n10385 ) | ( n10045 & n10386 ) | ( n10385 & n10386 ) ;
  assign n10388 = ( ~n10045 & n10385 ) | ( ~n10045 & n10386 ) | ( n10385 & n10386 ) ;
  assign n10389 = ( n10045 & ~n10387 ) | ( n10045 & n10388 ) | ( ~n10387 & n10388 ) ;
  assign n10390 = ( ~n1661 & n10384 ) | ( ~n1661 & n10389 ) | ( n10384 & n10389 ) ;
  assign n10391 = ~n1661 & n10046 ;
  assign n10392 = ( ~n1661 & n10046 ) | ( ~n1661 & n10180 ) | ( n10046 & n10180 ) ;
  assign n10393 = ( n10051 & n10391 ) | ( n10051 & n10392 ) | ( n10391 & n10392 ) ;
  assign n10394 = ( ~n10051 & n10391 ) | ( ~n10051 & n10392 ) | ( n10391 & n10392 ) ;
  assign n10395 = ( n10051 & ~n10393 ) | ( n10051 & n10394 ) | ( ~n10393 & n10394 ) ;
  assign n10396 = ( ~n1523 & n10390 ) | ( ~n1523 & n10395 ) | ( n10390 & n10395 ) ;
  assign n10397 = ~n1523 & n10052 ;
  assign n10398 = ( ~n1523 & n10052 ) | ( ~n1523 & n10180 ) | ( n10052 & n10180 ) ;
  assign n10399 = ( n10057 & n10397 ) | ( n10057 & n10398 ) | ( n10397 & n10398 ) ;
  assign n10400 = ( ~n10057 & n10397 ) | ( ~n10057 & n10398 ) | ( n10397 & n10398 ) ;
  assign n10401 = ( n10057 & ~n10399 ) | ( n10057 & n10400 ) | ( ~n10399 & n10400 ) ;
  assign n10402 = ( ~n1393 & n10396 ) | ( ~n1393 & n10401 ) | ( n10396 & n10401 ) ;
  assign n10403 = ~n1393 & n10058 ;
  assign n10404 = ( ~n1393 & n10058 ) | ( ~n1393 & n10180 ) | ( n10058 & n10180 ) ;
  assign n10405 = ( n10063 & n10403 ) | ( n10063 & n10404 ) | ( n10403 & n10404 ) ;
  assign n10406 = ( ~n10063 & n10403 ) | ( ~n10063 & n10404 ) | ( n10403 & n10404 ) ;
  assign n10407 = ( n10063 & ~n10405 ) | ( n10063 & n10406 ) | ( ~n10405 & n10406 ) ;
  assign n10408 = ( ~n1266 & n10402 ) | ( ~n1266 & n10407 ) | ( n10402 & n10407 ) ;
  assign n10409 = ( n1266 & ~n10064 ) | ( n1266 & n10180 ) | ( ~n10064 & n10180 ) ;
  assign n10410 = n1266 & ~n10064 ;
  assign n10411 = ( n10069 & n10409 ) | ( n10069 & n10410 ) | ( n10409 & n10410 ) ;
  assign n10412 = ( ~n10069 & n10409 ) | ( ~n10069 & n10410 ) | ( n10409 & n10410 ) ;
  assign n10413 = ( n10069 & ~n10411 ) | ( n10069 & n10412 ) | ( ~n10411 & n10412 ) ;
  assign n10414 = ( ~n1150 & n10408 ) | ( ~n1150 & n10413 ) | ( n10408 & n10413 ) ;
  assign n10415 = ( n1150 & ~n10070 ) | ( n1150 & n10180 ) | ( ~n10070 & n10180 ) ;
  assign n10416 = n1150 & ~n10070 ;
  assign n10417 = ( n10075 & n10415 ) | ( n10075 & n10416 ) | ( n10415 & n10416 ) ;
  assign n10418 = ( ~n10075 & n10415 ) | ( ~n10075 & n10416 ) | ( n10415 & n10416 ) ;
  assign n10419 = ( n10075 & ~n10417 ) | ( n10075 & n10418 ) | ( ~n10417 & n10418 ) ;
  assign n10420 = ( ~n1038 & n10414 ) | ( ~n1038 & n10419 ) | ( n10414 & n10419 ) ;
  assign n10421 = ~n1038 & n10076 ;
  assign n10422 = ( ~n1038 & n10076 ) | ( ~n1038 & n10180 ) | ( n10076 & n10180 ) ;
  assign n10423 = ( ~n10081 & n10421 ) | ( ~n10081 & n10422 ) | ( n10421 & n10422 ) ;
  assign n10424 = ( n10081 & n10421 ) | ( n10081 & n10422 ) | ( n10421 & n10422 ) ;
  assign n10425 = ( n10081 & n10423 ) | ( n10081 & ~n10424 ) | ( n10423 & ~n10424 ) ;
  assign n10426 = ( ~n933 & n10420 ) | ( ~n933 & n10425 ) | ( n10420 & n10425 ) ;
  assign n10427 = ( n933 & ~n10082 ) | ( n933 & n10180 ) | ( ~n10082 & n10180 ) ;
  assign n10428 = n933 & ~n10082 ;
  assign n10429 = ( n10087 & n10427 ) | ( n10087 & n10428 ) | ( n10427 & n10428 ) ;
  assign n10430 = ( ~n10087 & n10427 ) | ( ~n10087 & n10428 ) | ( n10427 & n10428 ) ;
  assign n10431 = ( n10087 & ~n10429 ) | ( n10087 & n10430 ) | ( ~n10429 & n10430 ) ;
  assign n10432 = ( ~n839 & n10426 ) | ( ~n839 & n10431 ) | ( n10426 & n10431 ) ;
  assign n10433 = ( n839 & ~n10088 ) | ( n839 & n10180 ) | ( ~n10088 & n10180 ) ;
  assign n10434 = n839 & ~n10088 ;
  assign n10435 = ( n10093 & n10433 ) | ( n10093 & n10434 ) | ( n10433 & n10434 ) ;
  assign n10436 = ( ~n10093 & n10433 ) | ( ~n10093 & n10434 ) | ( n10433 & n10434 ) ;
  assign n10437 = ( n10093 & ~n10435 ) | ( n10093 & n10436 ) | ( ~n10435 & n10436 ) ;
  assign n10438 = ( ~n746 & n10432 ) | ( ~n746 & n10437 ) | ( n10432 & n10437 ) ;
  assign n10439 = ( n746 & ~n10094 ) | ( n746 & n10180 ) | ( ~n10094 & n10180 ) ;
  assign n10440 = n746 & ~n10094 ;
  assign n10441 = ( n10099 & n10439 ) | ( n10099 & n10440 ) | ( n10439 & n10440 ) ;
  assign n10442 = ( ~n10099 & n10439 ) | ( ~n10099 & n10440 ) | ( n10439 & n10440 ) ;
  assign n10443 = ( n10099 & ~n10441 ) | ( n10099 & n10442 ) | ( ~n10441 & n10442 ) ;
  assign n10444 = ( ~n664 & n10438 ) | ( ~n664 & n10443 ) | ( n10438 & n10443 ) ;
  assign n10445 = ( n664 & ~n10100 ) | ( n664 & n10180 ) | ( ~n10100 & n10180 ) ;
  assign n10446 = n664 & ~n10100 ;
  assign n10447 = ( n10105 & n10445 ) | ( n10105 & n10446 ) | ( n10445 & n10446 ) ;
  assign n10448 = ( ~n10105 & n10445 ) | ( ~n10105 & n10446 ) | ( n10445 & n10446 ) ;
  assign n10449 = ( n10105 & ~n10447 ) | ( n10105 & n10448 ) | ( ~n10447 & n10448 ) ;
  assign n10450 = ( ~n588 & n10444 ) | ( ~n588 & n10449 ) | ( n10444 & n10449 ) ;
  assign n10451 = ( n588 & ~n10106 ) | ( n588 & n10180 ) | ( ~n10106 & n10180 ) ;
  assign n10452 = n588 & ~n10106 ;
  assign n10453 = ( n10111 & n10451 ) | ( n10111 & n10452 ) | ( n10451 & n10452 ) ;
  assign n10454 = ( ~n10111 & n10451 ) | ( ~n10111 & n10452 ) | ( n10451 & n10452 ) ;
  assign n10455 = ( n10111 & ~n10453 ) | ( n10111 & n10454 ) | ( ~n10453 & n10454 ) ;
  assign n10456 = ( ~n518 & n10450 ) | ( ~n518 & n10455 ) | ( n10450 & n10455 ) ;
  assign n10457 = ( n518 & ~n10112 ) | ( n518 & n10180 ) | ( ~n10112 & n10180 ) ;
  assign n10458 = n518 & ~n10112 ;
  assign n10459 = ( n10117 & n10457 ) | ( n10117 & n10458 ) | ( n10457 & n10458 ) ;
  assign n10460 = ( ~n10117 & n10457 ) | ( ~n10117 & n10458 ) | ( n10457 & n10458 ) ;
  assign n10461 = ( n10117 & ~n10459 ) | ( n10117 & n10460 ) | ( ~n10459 & n10460 ) ;
  assign n10462 = ( ~n454 & n10456 ) | ( ~n454 & n10461 ) | ( n10456 & n10461 ) ;
  assign n10463 = ( n454 & ~n10118 ) | ( n454 & n10180 ) | ( ~n10118 & n10180 ) ;
  assign n10464 = n454 & ~n10118 ;
  assign n10465 = ( n10123 & n10463 ) | ( n10123 & n10464 ) | ( n10463 & n10464 ) ;
  assign n10466 = ( ~n10123 & n10463 ) | ( ~n10123 & n10464 ) | ( n10463 & n10464 ) ;
  assign n10467 = ( n10123 & ~n10465 ) | ( n10123 & n10466 ) | ( ~n10465 & n10466 ) ;
  assign n10468 = ( ~n396 & n10462 ) | ( ~n396 & n10467 ) | ( n10462 & n10467 ) ;
  assign n10469 = ( n396 & ~n10124 ) | ( n396 & n10180 ) | ( ~n10124 & n10180 ) ;
  assign n10470 = n396 & ~n10124 ;
  assign n10471 = ( n10129 & n10469 ) | ( n10129 & n10470 ) | ( n10469 & n10470 ) ;
  assign n10472 = ( ~n10129 & n10469 ) | ( ~n10129 & n10470 ) | ( n10469 & n10470 ) ;
  assign n10473 = ( n10129 & ~n10471 ) | ( n10129 & n10472 ) | ( ~n10471 & n10472 ) ;
  assign n10474 = ( ~n344 & n10468 ) | ( ~n344 & n10473 ) | ( n10468 & n10473 ) ;
  assign n10475 = n344 & ~n10130 ;
  assign n10476 = ( n344 & ~n10130 ) | ( n344 & n10180 ) | ( ~n10130 & n10180 ) ;
  assign n10477 = ( n10135 & n10475 ) | ( n10135 & n10476 ) | ( n10475 & n10476 ) ;
  assign n10478 = ( ~n10135 & n10475 ) | ( ~n10135 & n10476 ) | ( n10475 & n10476 ) ;
  assign n10479 = ( n10135 & ~n10477 ) | ( n10135 & n10478 ) | ( ~n10477 & n10478 ) ;
  assign n10480 = ( ~n298 & n10474 ) | ( ~n298 & n10479 ) | ( n10474 & n10479 ) ;
  assign n10481 = ~n298 & n10136 ;
  assign n10482 = ( ~n298 & n10136 ) | ( ~n298 & n10180 ) | ( n10136 & n10180 ) ;
  assign n10483 = ( ~n10141 & n10481 ) | ( ~n10141 & n10482 ) | ( n10481 & n10482 ) ;
  assign n10484 = ( n10141 & n10481 ) | ( n10141 & n10482 ) | ( n10481 & n10482 ) ;
  assign n10485 = ( n10141 & n10483 ) | ( n10141 & ~n10484 ) | ( n10483 & ~n10484 ) ;
  assign n10486 = ( ~n258 & n10480 ) | ( ~n258 & n10485 ) | ( n10480 & n10485 ) ;
  assign n10487 = ( n258 & ~n10142 ) | ( n258 & n10180 ) | ( ~n10142 & n10180 ) ;
  assign n10488 = n258 & ~n10142 ;
  assign n10489 = ( n10147 & n10487 ) | ( n10147 & n10488 ) | ( n10487 & n10488 ) ;
  assign n10490 = ( ~n10147 & n10487 ) | ( ~n10147 & n10488 ) | ( n10487 & n10488 ) ;
  assign n10491 = ( n10147 & ~n10489 ) | ( n10147 & n10490 ) | ( ~n10489 & n10490 ) ;
  assign n10492 = ( ~n225 & n10486 ) | ( ~n225 & n10491 ) | ( n10486 & n10491 ) ;
  assign n10493 = n225 & ~n10148 ;
  assign n10494 = ( n225 & ~n10148 ) | ( n225 & n10180 ) | ( ~n10148 & n10180 ) ;
  assign n10495 = ( n10153 & n10493 ) | ( n10153 & n10494 ) | ( n10493 & n10494 ) ;
  assign n10496 = ( ~n10153 & n10493 ) | ( ~n10153 & n10494 ) | ( n10493 & n10494 ) ;
  assign n10497 = ( n10153 & ~n10495 ) | ( n10153 & n10496 ) | ( ~n10495 & n10496 ) ;
  assign n10498 = ( ~n197 & n10492 ) | ( ~n197 & n10497 ) | ( n10492 & n10497 ) ;
  assign n10499 = ( n197 & ~n10154 ) | ( n197 & n10180 ) | ( ~n10154 & n10180 ) ;
  assign n10500 = n197 & ~n10154 ;
  assign n10501 = ( n10159 & n10499 ) | ( n10159 & n10500 ) | ( n10499 & n10500 ) ;
  assign n10502 = ( ~n10159 & n10499 ) | ( ~n10159 & n10500 ) | ( n10499 & n10500 ) ;
  assign n10503 = ( n10159 & ~n10501 ) | ( n10159 & n10502 ) | ( ~n10501 & n10502 ) ;
  assign n10504 = ( ~n170 & n10498 ) | ( ~n170 & n10503 ) | ( n10498 & n10503 ) ;
  assign n10505 = ( n170 & ~n10160 ) | ( n170 & n10180 ) | ( ~n10160 & n10180 ) ;
  assign n10506 = n170 & ~n10160 ;
  assign n10507 = ( n10165 & n10505 ) | ( n10165 & n10506 ) | ( n10505 & n10506 ) ;
  assign n10508 = ( ~n10165 & n10505 ) | ( ~n10165 & n10506 ) | ( n10505 & n10506 ) ;
  assign n10509 = ( n10165 & ~n10507 ) | ( n10165 & n10508 ) | ( ~n10507 & n10508 ) ;
  assign n10510 = ( ~n142 & n10504 ) | ( ~n142 & n10509 ) | ( n10504 & n10509 ) ;
  assign n10511 = ( n142 & ~n10166 ) | ( n142 & n10180 ) | ( ~n10166 & n10180 ) ;
  assign n10512 = n142 & ~n10166 ;
  assign n10513 = ( n10171 & n10511 ) | ( n10171 & n10512 ) | ( n10511 & n10512 ) ;
  assign n10514 = ( ~n10171 & n10511 ) | ( ~n10171 & n10512 ) | ( n10511 & n10512 ) ;
  assign n10515 = ( n10171 & ~n10513 ) | ( n10171 & n10514 ) | ( ~n10513 & n10514 ) ;
  assign n10516 = ( ~n132 & n10510 ) | ( ~n132 & n10515 ) | ( n10510 & n10515 ) ;
  assign n10517 = n9842 | n9848 ;
  assign n10518 = ( n9848 & n10178 ) | ( n9848 & n10517 ) | ( n10178 & n10517 ) ;
  assign n10519 = ~n10179 & n10518 ;
  assign n10520 = ( n132 & ~n10172 ) | ( n132 & n10180 ) | ( ~n10172 & n10180 ) ;
  assign n10521 = n132 & ~n10172 ;
  assign n10522 = ( n10177 & n10520 ) | ( n10177 & n10521 ) | ( n10520 & n10521 ) ;
  assign n10523 = ( ~n10177 & n10520 ) | ( ~n10177 & n10521 ) | ( n10520 & n10521 ) ;
  assign n10524 = ( n10177 & ~n10522 ) | ( n10177 & n10523 ) | ( ~n10522 & n10523 ) ;
  assign n10525 = n10519 | n10524 ;
  assign n10526 = ( n10516 & n10519 ) | ( n10516 & n10525 ) | ( n10519 & n10525 ) ;
  assign n10527 = n10516 | n10524 ;
  assign n10528 = n9848 & n10178 ;
  assign n10529 = n9843 & ~n9848 ;
  assign n10530 = ~n10178 & n10529 ;
  assign n10531 = ( ~n10527 & n10528 ) | ( ~n10527 & n10530 ) | ( n10528 & n10530 ) ;
  assign n10532 = ( ~n131 & n10527 ) | ( ~n131 & n10531 ) | ( n10527 & n10531 ) ;
  assign n10533 = n10526 | n10532 ;
  assign n10534 = ( n132 & ~n10510 ) | ( n132 & n10533 ) | ( ~n10510 & n10533 ) ;
  assign n10535 = n132 & ~n10510 ;
  assign n10536 = ( n10515 & n10534 ) | ( n10515 & n10535 ) | ( n10534 & n10535 ) ;
  assign n10537 = ( ~n10515 & n10534 ) | ( ~n10515 & n10535 ) | ( n10534 & n10535 ) ;
  assign n10538 = ( n10515 & ~n10536 ) | ( n10515 & n10537 ) | ( ~n10536 & n10537 ) ;
  assign n10539 = n131 | n10538 ;
  assign n10540 = ( n10516 & n10524 ) | ( n10516 & ~n10525 ) | ( n10524 & ~n10525 ) ;
  assign n10541 = ( n131 & ~n10527 ) | ( n131 & n10540 ) | ( ~n10527 & n10540 ) ;
  assign n10542 = x8 | x9 ;
  assign n10543 = x10 | n10542 ;
  assign n10544 = ~n10180 & n10543 ;
  assign n10545 = ( x11 & ~n10533 ) | ( x11 & n10544 ) | ( ~n10533 & n10544 ) ;
  assign n10546 = n10180 & ~n10543 ;
  assign n10547 = ~n10186 & n10533 ;
  assign n10548 = ( n10545 & ~n10546 ) | ( n10545 & n10547 ) | ( ~n10546 & n10547 ) ;
  assign n10549 = n10180 & ~n10533 ;
  assign n10550 = ( ~x12 & n10547 ) | ( ~x12 & n10549 ) | ( n10547 & n10549 ) ;
  assign n10551 = ( x12 & n10547 ) | ( x12 & n10549 ) | ( n10547 & n10549 ) ;
  assign n10552 = ( x12 & n10550 ) | ( x12 & ~n10551 ) | ( n10550 & ~n10551 ) ;
  assign n10553 = ( ~n9834 & n10548 ) | ( ~n9834 & n10552 ) | ( n10548 & n10552 ) ;
  assign n10554 = ~n9834 & n10180 ;
  assign n10555 = ( n10181 & n10533 ) | ( n10181 & n10554 ) | ( n10533 & n10554 ) ;
  assign n10556 = ( ~x13 & n10550 ) | ( ~x13 & n10555 ) | ( n10550 & n10555 ) ;
  assign n10557 = ( x13 & n10550 ) | ( x13 & n10555 ) | ( n10550 & n10555 ) ;
  assign n10558 = ( x13 & n10556 ) | ( x13 & ~n10557 ) | ( n10556 & ~n10557 ) ;
  assign n10559 = ( ~n9497 & n10553 ) | ( ~n9497 & n10558 ) | ( n10553 & n10558 ) ;
  assign n10560 = n9497 & ~n10191 ;
  assign n10561 = ( n9497 & ~n10191 ) | ( n9497 & n10533 ) | ( ~n10191 & n10533 ) ;
  assign n10562 = ( n10185 & n10560 ) | ( n10185 & n10561 ) | ( n10560 & n10561 ) ;
  assign n10563 = ( ~n10185 & n10560 ) | ( ~n10185 & n10561 ) | ( n10560 & n10561 ) ;
  assign n10564 = ( n10185 & ~n10562 ) | ( n10185 & n10563 ) | ( ~n10562 & n10563 ) ;
  assign n10565 = ( ~n9167 & n10559 ) | ( ~n9167 & n10564 ) | ( n10559 & n10564 ) ;
  assign n10566 = n9167 & ~n10192 ;
  assign n10567 = ( n9167 & ~n10192 ) | ( n9167 & n10533 ) | ( ~n10192 & n10533 ) ;
  assign n10568 = ( n10197 & n10566 ) | ( n10197 & n10567 ) | ( n10566 & n10567 ) ;
  assign n10569 = ( ~n10197 & n10566 ) | ( ~n10197 & n10567 ) | ( n10566 & n10567 ) ;
  assign n10570 = ( n10197 & ~n10568 ) | ( n10197 & n10569 ) | ( ~n10568 & n10569 ) ;
  assign n10571 = ( ~n8838 & n10565 ) | ( ~n8838 & n10570 ) | ( n10565 & n10570 ) ;
  assign n10572 = n8838 & ~n10198 ;
  assign n10573 = ( n8838 & ~n10198 ) | ( n8838 & n10533 ) | ( ~n10198 & n10533 ) ;
  assign n10574 = ( n10203 & n10572 ) | ( n10203 & n10573 ) | ( n10572 & n10573 ) ;
  assign n10575 = ( ~n10203 & n10572 ) | ( ~n10203 & n10573 ) | ( n10572 & n10573 ) ;
  assign n10576 = ( n10203 & ~n10574 ) | ( n10203 & n10575 ) | ( ~n10574 & n10575 ) ;
  assign n10577 = ( ~n8517 & n10571 ) | ( ~n8517 & n10576 ) | ( n10571 & n10576 ) ;
  assign n10578 = ( n8517 & ~n10204 ) | ( n8517 & n10533 ) | ( ~n10204 & n10533 ) ;
  assign n10579 = n8517 & ~n10204 ;
  assign n10580 = ( n10209 & n10578 ) | ( n10209 & n10579 ) | ( n10578 & n10579 ) ;
  assign n10581 = ( ~n10209 & n10578 ) | ( ~n10209 & n10579 ) | ( n10578 & n10579 ) ;
  assign n10582 = ( n10209 & ~n10580 ) | ( n10209 & n10581 ) | ( ~n10580 & n10581 ) ;
  assign n10583 = ( ~n8201 & n10577 ) | ( ~n8201 & n10582 ) | ( n10577 & n10582 ) ;
  assign n10584 = ~n8201 & n10210 ;
  assign n10585 = ( ~n8201 & n10210 ) | ( ~n8201 & n10533 ) | ( n10210 & n10533 ) ;
  assign n10586 = ( ~n10215 & n10584 ) | ( ~n10215 & n10585 ) | ( n10584 & n10585 ) ;
  assign n10587 = ( n10215 & n10584 ) | ( n10215 & n10585 ) | ( n10584 & n10585 ) ;
  assign n10588 = ( n10215 & n10586 ) | ( n10215 & ~n10587 ) | ( n10586 & ~n10587 ) ;
  assign n10589 = ( ~n7897 & n10583 ) | ( ~n7897 & n10588 ) | ( n10583 & n10588 ) ;
  assign n10590 = ( n7897 & ~n10216 ) | ( n7897 & n10533 ) | ( ~n10216 & n10533 ) ;
  assign n10591 = n7897 & ~n10216 ;
  assign n10592 = ( n10221 & n10590 ) | ( n10221 & n10591 ) | ( n10590 & n10591 ) ;
  assign n10593 = ( ~n10221 & n10590 ) | ( ~n10221 & n10591 ) | ( n10590 & n10591 ) ;
  assign n10594 = ( n10221 & ~n10592 ) | ( n10221 & n10593 ) | ( ~n10592 & n10593 ) ;
  assign n10595 = ( ~n7594 & n10589 ) | ( ~n7594 & n10594 ) | ( n10589 & n10594 ) ;
  assign n10596 = ~n7594 & n10222 ;
  assign n10597 = ( ~n7594 & n10222 ) | ( ~n7594 & n10533 ) | ( n10222 & n10533 ) ;
  assign n10598 = ( ~n10227 & n10596 ) | ( ~n10227 & n10597 ) | ( n10596 & n10597 ) ;
  assign n10599 = ( n10227 & n10596 ) | ( n10227 & n10597 ) | ( n10596 & n10597 ) ;
  assign n10600 = ( n10227 & n10598 ) | ( n10227 & ~n10599 ) | ( n10598 & ~n10599 ) ;
  assign n10601 = ( ~n7296 & n10595 ) | ( ~n7296 & n10600 ) | ( n10595 & n10600 ) ;
  assign n10602 = ~n7296 & n10228 ;
  assign n10603 = ( ~n7296 & n10228 ) | ( ~n7296 & n10533 ) | ( n10228 & n10533 ) ;
  assign n10604 = ( n10233 & n10602 ) | ( n10233 & n10603 ) | ( n10602 & n10603 ) ;
  assign n10605 = ( ~n10233 & n10602 ) | ( ~n10233 & n10603 ) | ( n10602 & n10603 ) ;
  assign n10606 = ( n10233 & ~n10604 ) | ( n10233 & n10605 ) | ( ~n10604 & n10605 ) ;
  assign n10607 = ( ~n7006 & n10601 ) | ( ~n7006 & n10606 ) | ( n10601 & n10606 ) ;
  assign n10608 = ( n7006 & ~n10234 ) | ( n7006 & n10533 ) | ( ~n10234 & n10533 ) ;
  assign n10609 = n7006 & ~n10234 ;
  assign n10610 = ( n10239 & n10608 ) | ( n10239 & n10609 ) | ( n10608 & n10609 ) ;
  assign n10611 = ( ~n10239 & n10608 ) | ( ~n10239 & n10609 ) | ( n10608 & n10609 ) ;
  assign n10612 = ( n10239 & ~n10610 ) | ( n10239 & n10611 ) | ( ~n10610 & n10611 ) ;
  assign n10613 = ( ~n6723 & n10607 ) | ( ~n6723 & n10612 ) | ( n10607 & n10612 ) ;
  assign n10614 = n6723 & ~n10240 ;
  assign n10615 = ( n6723 & ~n10240 ) | ( n6723 & n10533 ) | ( ~n10240 & n10533 ) ;
  assign n10616 = ( ~n10245 & n10614 ) | ( ~n10245 & n10615 ) | ( n10614 & n10615 ) ;
  assign n10617 = ( n10245 & n10614 ) | ( n10245 & n10615 ) | ( n10614 & n10615 ) ;
  assign n10618 = ( n10245 & n10616 ) | ( n10245 & ~n10617 ) | ( n10616 & ~n10617 ) ;
  assign n10619 = ( ~n6442 & n10613 ) | ( ~n6442 & n10618 ) | ( n10613 & n10618 ) ;
  assign n10620 = ~n6442 & n10246 ;
  assign n10621 = ( ~n6442 & n10246 ) | ( ~n6442 & n10533 ) | ( n10246 & n10533 ) ;
  assign n10622 = ( ~n10251 & n10620 ) | ( ~n10251 & n10621 ) | ( n10620 & n10621 ) ;
  assign n10623 = ( n10251 & n10620 ) | ( n10251 & n10621 ) | ( n10620 & n10621 ) ;
  assign n10624 = ( n10251 & n10622 ) | ( n10251 & ~n10623 ) | ( n10622 & ~n10623 ) ;
  assign n10625 = ( ~n6172 & n10619 ) | ( ~n6172 & n10624 ) | ( n10619 & n10624 ) ;
  assign n10626 = ( n6172 & ~n10252 ) | ( n6172 & n10533 ) | ( ~n10252 & n10533 ) ;
  assign n10627 = n6172 & ~n10252 ;
  assign n10628 = ( n10257 & n10626 ) | ( n10257 & n10627 ) | ( n10626 & n10627 ) ;
  assign n10629 = ( ~n10257 & n10626 ) | ( ~n10257 & n10627 ) | ( n10626 & n10627 ) ;
  assign n10630 = ( n10257 & ~n10628 ) | ( n10257 & n10629 ) | ( ~n10628 & n10629 ) ;
  assign n10631 = ( ~n5905 & n10625 ) | ( ~n5905 & n10630 ) | ( n10625 & n10630 ) ;
  assign n10632 = ( n5905 & ~n10258 ) | ( n5905 & n10533 ) | ( ~n10258 & n10533 ) ;
  assign n10633 = n5905 & ~n10258 ;
  assign n10634 = ( n10263 & n10632 ) | ( n10263 & n10633 ) | ( n10632 & n10633 ) ;
  assign n10635 = ( ~n10263 & n10632 ) | ( ~n10263 & n10633 ) | ( n10632 & n10633 ) ;
  assign n10636 = ( n10263 & ~n10634 ) | ( n10263 & n10635 ) | ( ~n10634 & n10635 ) ;
  assign n10637 = ( ~n5642 & n10631 ) | ( ~n5642 & n10636 ) | ( n10631 & n10636 ) ;
  assign n10638 = ( n5642 & ~n10264 ) | ( n5642 & n10533 ) | ( ~n10264 & n10533 ) ;
  assign n10639 = n5642 & ~n10264 ;
  assign n10640 = ( n10269 & n10638 ) | ( n10269 & n10639 ) | ( n10638 & n10639 ) ;
  assign n10641 = ( ~n10269 & n10638 ) | ( ~n10269 & n10639 ) | ( n10638 & n10639 ) ;
  assign n10642 = ( n10269 & ~n10640 ) | ( n10269 & n10641 ) | ( ~n10640 & n10641 ) ;
  assign n10643 = ( ~n5386 & n10637 ) | ( ~n5386 & n10642 ) | ( n10637 & n10642 ) ;
  assign n10644 = ~n5386 & n10270 ;
  assign n10645 = ( ~n5386 & n10270 ) | ( ~n5386 & n10533 ) | ( n10270 & n10533 ) ;
  assign n10646 = ( ~n10275 & n10644 ) | ( ~n10275 & n10645 ) | ( n10644 & n10645 ) ;
  assign n10647 = ( n10275 & n10644 ) | ( n10275 & n10645 ) | ( n10644 & n10645 ) ;
  assign n10648 = ( n10275 & n10646 ) | ( n10275 & ~n10647 ) | ( n10646 & ~n10647 ) ;
  assign n10649 = ( ~n5139 & n10643 ) | ( ~n5139 & n10648 ) | ( n10643 & n10648 ) ;
  assign n10650 = ( n5139 & ~n10276 ) | ( n5139 & n10533 ) | ( ~n10276 & n10533 ) ;
  assign n10651 = n5139 & ~n10276 ;
  assign n10652 = ( n10281 & n10650 ) | ( n10281 & n10651 ) | ( n10650 & n10651 ) ;
  assign n10653 = ( ~n10281 & n10650 ) | ( ~n10281 & n10651 ) | ( n10650 & n10651 ) ;
  assign n10654 = ( n10281 & ~n10652 ) | ( n10281 & n10653 ) | ( ~n10652 & n10653 ) ;
  assign n10655 = ( ~n4898 & n10649 ) | ( ~n4898 & n10654 ) | ( n10649 & n10654 ) ;
  assign n10656 = ( n4898 & ~n10282 ) | ( n4898 & n10533 ) | ( ~n10282 & n10533 ) ;
  assign n10657 = n4898 & ~n10282 ;
  assign n10658 = ( n10287 & n10656 ) | ( n10287 & n10657 ) | ( n10656 & n10657 ) ;
  assign n10659 = ( ~n10287 & n10656 ) | ( ~n10287 & n10657 ) | ( n10656 & n10657 ) ;
  assign n10660 = ( n10287 & ~n10658 ) | ( n10287 & n10659 ) | ( ~n10658 & n10659 ) ;
  assign n10661 = ( ~n4661 & n10655 ) | ( ~n4661 & n10660 ) | ( n10655 & n10660 ) ;
  assign n10662 = ( n4661 & ~n10288 ) | ( n4661 & n10533 ) | ( ~n10288 & n10533 ) ;
  assign n10663 = n4661 & ~n10288 ;
  assign n10664 = ( n10293 & n10662 ) | ( n10293 & n10663 ) | ( n10662 & n10663 ) ;
  assign n10665 = ( ~n10293 & n10662 ) | ( ~n10293 & n10663 ) | ( n10662 & n10663 ) ;
  assign n10666 = ( n10293 & ~n10664 ) | ( n10293 & n10665 ) | ( ~n10664 & n10665 ) ;
  assign n10667 = ( ~n4432 & n10661 ) | ( ~n4432 & n10666 ) | ( n10661 & n10666 ) ;
  assign n10668 = ( n4432 & ~n10294 ) | ( n4432 & n10533 ) | ( ~n10294 & n10533 ) ;
  assign n10669 = n4432 & ~n10294 ;
  assign n10670 = ( n10299 & n10668 ) | ( n10299 & n10669 ) | ( n10668 & n10669 ) ;
  assign n10671 = ( ~n10299 & n10668 ) | ( ~n10299 & n10669 ) | ( n10668 & n10669 ) ;
  assign n10672 = ( n10299 & ~n10670 ) | ( n10299 & n10671 ) | ( ~n10670 & n10671 ) ;
  assign n10673 = ( ~n4203 & n10667 ) | ( ~n4203 & n10672 ) | ( n10667 & n10672 ) ;
  assign n10674 = ~n4203 & n10300 ;
  assign n10675 = ( ~n4203 & n10300 ) | ( ~n4203 & n10533 ) | ( n10300 & n10533 ) ;
  assign n10676 = ( n10305 & n10674 ) | ( n10305 & n10675 ) | ( n10674 & n10675 ) ;
  assign n10677 = ( ~n10305 & n10674 ) | ( ~n10305 & n10675 ) | ( n10674 & n10675 ) ;
  assign n10678 = ( n10305 & ~n10676 ) | ( n10305 & n10677 ) | ( ~n10676 & n10677 ) ;
  assign n10679 = ( ~n3985 & n10673 ) | ( ~n3985 & n10678 ) | ( n10673 & n10678 ) ;
  assign n10680 = ( n3985 & ~n10306 ) | ( n3985 & n10533 ) | ( ~n10306 & n10533 ) ;
  assign n10681 = n3985 & ~n10306 ;
  assign n10682 = ( n10311 & n10680 ) | ( n10311 & n10681 ) | ( n10680 & n10681 ) ;
  assign n10683 = ( ~n10311 & n10680 ) | ( ~n10311 & n10681 ) | ( n10680 & n10681 ) ;
  assign n10684 = ( n10311 & ~n10682 ) | ( n10311 & n10683 ) | ( ~n10682 & n10683 ) ;
  assign n10685 = ( ~n3772 & n10679 ) | ( ~n3772 & n10684 ) | ( n10679 & n10684 ) ;
  assign n10686 = ( n3772 & ~n10312 ) | ( n3772 & n10533 ) | ( ~n10312 & n10533 ) ;
  assign n10687 = n3772 & ~n10312 ;
  assign n10688 = ( n10317 & n10686 ) | ( n10317 & n10687 ) | ( n10686 & n10687 ) ;
  assign n10689 = ( ~n10317 & n10686 ) | ( ~n10317 & n10687 ) | ( n10686 & n10687 ) ;
  assign n10690 = ( n10317 & ~n10688 ) | ( n10317 & n10689 ) | ( ~n10688 & n10689 ) ;
  assign n10691 = ( ~n3567 & n10685 ) | ( ~n3567 & n10690 ) | ( n10685 & n10690 ) ;
  assign n10692 = ( n3567 & ~n10318 ) | ( n3567 & n10533 ) | ( ~n10318 & n10533 ) ;
  assign n10693 = n3567 & ~n10318 ;
  assign n10694 = ( n10323 & n10692 ) | ( n10323 & n10693 ) | ( n10692 & n10693 ) ;
  assign n10695 = ( ~n10323 & n10692 ) | ( ~n10323 & n10693 ) | ( n10692 & n10693 ) ;
  assign n10696 = ( n10323 & ~n10694 ) | ( n10323 & n10695 ) | ( ~n10694 & n10695 ) ;
  assign n10697 = ( ~n3362 & n10691 ) | ( ~n3362 & n10696 ) | ( n10691 & n10696 ) ;
  assign n10698 = ( n3362 & ~n10324 ) | ( n3362 & n10533 ) | ( ~n10324 & n10533 ) ;
  assign n10699 = n3362 & ~n10324 ;
  assign n10700 = ( n10329 & n10698 ) | ( n10329 & n10699 ) | ( n10698 & n10699 ) ;
  assign n10701 = ( ~n10329 & n10698 ) | ( ~n10329 & n10699 ) | ( n10698 & n10699 ) ;
  assign n10702 = ( n10329 & ~n10700 ) | ( n10329 & n10701 ) | ( ~n10700 & n10701 ) ;
  assign n10703 = ( ~n3169 & n10697 ) | ( ~n3169 & n10702 ) | ( n10697 & n10702 ) ;
  assign n10704 = ~n3169 & n10330 ;
  assign n10705 = ( ~n3169 & n10330 ) | ( ~n3169 & n10533 ) | ( n10330 & n10533 ) ;
  assign n10706 = ( ~n10335 & n10704 ) | ( ~n10335 & n10705 ) | ( n10704 & n10705 ) ;
  assign n10707 = ( n10335 & n10704 ) | ( n10335 & n10705 ) | ( n10704 & n10705 ) ;
  assign n10708 = ( n10335 & n10706 ) | ( n10335 & ~n10707 ) | ( n10706 & ~n10707 ) ;
  assign n10709 = ( ~n2979 & n10703 ) | ( ~n2979 & n10708 ) | ( n10703 & n10708 ) ;
  assign n10710 = ~n2979 & n10336 ;
  assign n10711 = ( ~n2979 & n10336 ) | ( ~n2979 & n10533 ) | ( n10336 & n10533 ) ;
  assign n10712 = ( ~n10341 & n10710 ) | ( ~n10341 & n10711 ) | ( n10710 & n10711 ) ;
  assign n10713 = ( n10341 & n10710 ) | ( n10341 & n10711 ) | ( n10710 & n10711 ) ;
  assign n10714 = ( n10341 & n10712 ) | ( n10341 & ~n10713 ) | ( n10712 & ~n10713 ) ;
  assign n10715 = ( ~n2791 & n10709 ) | ( ~n2791 & n10714 ) | ( n10709 & n10714 ) ;
  assign n10716 = ~n2791 & n10342 ;
  assign n10717 = ( ~n2791 & n10342 ) | ( ~n2791 & n10533 ) | ( n10342 & n10533 ) ;
  assign n10718 = ( n10347 & n10716 ) | ( n10347 & n10717 ) | ( n10716 & n10717 ) ;
  assign n10719 = ( ~n10347 & n10716 ) | ( ~n10347 & n10717 ) | ( n10716 & n10717 ) ;
  assign n10720 = ( n10347 & ~n10718 ) | ( n10347 & n10719 ) | ( ~n10718 & n10719 ) ;
  assign n10721 = ( ~n2615 & n10715 ) | ( ~n2615 & n10720 ) | ( n10715 & n10720 ) ;
  assign n10722 = ( n2615 & ~n10348 ) | ( n2615 & n10533 ) | ( ~n10348 & n10533 ) ;
  assign n10723 = n2615 & ~n10348 ;
  assign n10724 = ( n10353 & n10722 ) | ( n10353 & n10723 ) | ( n10722 & n10723 ) ;
  assign n10725 = ( ~n10353 & n10722 ) | ( ~n10353 & n10723 ) | ( n10722 & n10723 ) ;
  assign n10726 = ( n10353 & ~n10724 ) | ( n10353 & n10725 ) | ( ~n10724 & n10725 ) ;
  assign n10727 = ( ~n2443 & n10721 ) | ( ~n2443 & n10726 ) | ( n10721 & n10726 ) ;
  assign n10728 = ~n2443 & n10354 ;
  assign n10729 = ( ~n2443 & n10354 ) | ( ~n2443 & n10533 ) | ( n10354 & n10533 ) ;
  assign n10730 = ( n10359 & n10728 ) | ( n10359 & n10729 ) | ( n10728 & n10729 ) ;
  assign n10731 = ( ~n10359 & n10728 ) | ( ~n10359 & n10729 ) | ( n10728 & n10729 ) ;
  assign n10732 = ( n10359 & ~n10730 ) | ( n10359 & n10731 ) | ( ~n10730 & n10731 ) ;
  assign n10733 = ( ~n2277 & n10727 ) | ( ~n2277 & n10732 ) | ( n10727 & n10732 ) ;
  assign n10734 = ( n2277 & ~n10360 ) | ( n2277 & n10533 ) | ( ~n10360 & n10533 ) ;
  assign n10735 = n2277 & ~n10360 ;
  assign n10736 = ( n10365 & n10734 ) | ( n10365 & n10735 ) | ( n10734 & n10735 ) ;
  assign n10737 = ( ~n10365 & n10734 ) | ( ~n10365 & n10735 ) | ( n10734 & n10735 ) ;
  assign n10738 = ( n10365 & ~n10736 ) | ( n10365 & n10737 ) | ( ~n10736 & n10737 ) ;
  assign n10739 = ( ~n2111 & n10733 ) | ( ~n2111 & n10738 ) | ( n10733 & n10738 ) ;
  assign n10740 = ~n2111 & n10366 ;
  assign n10741 = ( ~n2111 & n10366 ) | ( ~n2111 & n10533 ) | ( n10366 & n10533 ) ;
  assign n10742 = ( n10371 & n10740 ) | ( n10371 & n10741 ) | ( n10740 & n10741 ) ;
  assign n10743 = ( ~n10371 & n10740 ) | ( ~n10371 & n10741 ) | ( n10740 & n10741 ) ;
  assign n10744 = ( n10371 & ~n10742 ) | ( n10371 & n10743 ) | ( ~n10742 & n10743 ) ;
  assign n10745 = ( ~n1949 & n10739 ) | ( ~n1949 & n10744 ) | ( n10739 & n10744 ) ;
  assign n10746 = ~n1949 & n10372 ;
  assign n10747 = ( ~n1949 & n10372 ) | ( ~n1949 & n10533 ) | ( n10372 & n10533 ) ;
  assign n10748 = ( ~n10377 & n10746 ) | ( ~n10377 & n10747 ) | ( n10746 & n10747 ) ;
  assign n10749 = ( n10377 & n10746 ) | ( n10377 & n10747 ) | ( n10746 & n10747 ) ;
  assign n10750 = ( n10377 & n10748 ) | ( n10377 & ~n10749 ) | ( n10748 & ~n10749 ) ;
  assign n10751 = ( ~n1802 & n10745 ) | ( ~n1802 & n10750 ) | ( n10745 & n10750 ) ;
  assign n10752 = ~n1802 & n10378 ;
  assign n10753 = ( ~n1802 & n10378 ) | ( ~n1802 & n10533 ) | ( n10378 & n10533 ) ;
  assign n10754 = ( ~n10383 & n10752 ) | ( ~n10383 & n10753 ) | ( n10752 & n10753 ) ;
  assign n10755 = ( n10383 & n10752 ) | ( n10383 & n10753 ) | ( n10752 & n10753 ) ;
  assign n10756 = ( n10383 & n10754 ) | ( n10383 & ~n10755 ) | ( n10754 & ~n10755 ) ;
  assign n10757 = ( ~n1661 & n10751 ) | ( ~n1661 & n10756 ) | ( n10751 & n10756 ) ;
  assign n10758 = ( n1661 & ~n10384 ) | ( n1661 & n10533 ) | ( ~n10384 & n10533 ) ;
  assign n10759 = n1661 & ~n10384 ;
  assign n10760 = ( n10389 & n10758 ) | ( n10389 & n10759 ) | ( n10758 & n10759 ) ;
  assign n10761 = ( ~n10389 & n10758 ) | ( ~n10389 & n10759 ) | ( n10758 & n10759 ) ;
  assign n10762 = ( n10389 & ~n10760 ) | ( n10389 & n10761 ) | ( ~n10760 & n10761 ) ;
  assign n10763 = ( ~n1523 & n10757 ) | ( ~n1523 & n10762 ) | ( n10757 & n10762 ) ;
  assign n10764 = ( n1523 & ~n10390 ) | ( n1523 & n10533 ) | ( ~n10390 & n10533 ) ;
  assign n10765 = n1523 & ~n10390 ;
  assign n10766 = ( n10395 & n10764 ) | ( n10395 & n10765 ) | ( n10764 & n10765 ) ;
  assign n10767 = ( ~n10395 & n10764 ) | ( ~n10395 & n10765 ) | ( n10764 & n10765 ) ;
  assign n10768 = ( n10395 & ~n10766 ) | ( n10395 & n10767 ) | ( ~n10766 & n10767 ) ;
  assign n10769 = ( ~n1393 & n10763 ) | ( ~n1393 & n10768 ) | ( n10763 & n10768 ) ;
  assign n10770 = ~n1393 & n10396 ;
  assign n10771 = ( ~n1393 & n10396 ) | ( ~n1393 & n10533 ) | ( n10396 & n10533 ) ;
  assign n10772 = ( n10401 & n10770 ) | ( n10401 & n10771 ) | ( n10770 & n10771 ) ;
  assign n10773 = ( ~n10401 & n10770 ) | ( ~n10401 & n10771 ) | ( n10770 & n10771 ) ;
  assign n10774 = ( n10401 & ~n10772 ) | ( n10401 & n10773 ) | ( ~n10772 & n10773 ) ;
  assign n10775 = ( ~n1266 & n10769 ) | ( ~n1266 & n10774 ) | ( n10769 & n10774 ) ;
  assign n10776 = n1266 & ~n10402 ;
  assign n10777 = ( n1266 & ~n10402 ) | ( n1266 & n10533 ) | ( ~n10402 & n10533 ) ;
  assign n10778 = ( ~n10407 & n10776 ) | ( ~n10407 & n10777 ) | ( n10776 & n10777 ) ;
  assign n10779 = ( n10407 & n10776 ) | ( n10407 & n10777 ) | ( n10776 & n10777 ) ;
  assign n10780 = ( n10407 & n10778 ) | ( n10407 & ~n10779 ) | ( n10778 & ~n10779 ) ;
  assign n10781 = ( ~n1150 & n10775 ) | ( ~n1150 & n10780 ) | ( n10775 & n10780 ) ;
  assign n10782 = ( n1150 & ~n10408 ) | ( n1150 & n10533 ) | ( ~n10408 & n10533 ) ;
  assign n10783 = n1150 & ~n10408 ;
  assign n10784 = ( n10413 & n10782 ) | ( n10413 & n10783 ) | ( n10782 & n10783 ) ;
  assign n10785 = ( ~n10413 & n10782 ) | ( ~n10413 & n10783 ) | ( n10782 & n10783 ) ;
  assign n10786 = ( n10413 & ~n10784 ) | ( n10413 & n10785 ) | ( ~n10784 & n10785 ) ;
  assign n10787 = ( ~n1038 & n10781 ) | ( ~n1038 & n10786 ) | ( n10781 & n10786 ) ;
  assign n10788 = ( n1038 & ~n10414 ) | ( n1038 & n10533 ) | ( ~n10414 & n10533 ) ;
  assign n10789 = n1038 & ~n10414 ;
  assign n10790 = ( n10419 & n10788 ) | ( n10419 & n10789 ) | ( n10788 & n10789 ) ;
  assign n10791 = ( ~n10419 & n10788 ) | ( ~n10419 & n10789 ) | ( n10788 & n10789 ) ;
  assign n10792 = ( n10419 & ~n10790 ) | ( n10419 & n10791 ) | ( ~n10790 & n10791 ) ;
  assign n10793 = ( ~n933 & n10787 ) | ( ~n933 & n10792 ) | ( n10787 & n10792 ) ;
  assign n10794 = ~n933 & n10420 ;
  assign n10795 = ( ~n933 & n10420 ) | ( ~n933 & n10533 ) | ( n10420 & n10533 ) ;
  assign n10796 = ( n10425 & n10794 ) | ( n10425 & n10795 ) | ( n10794 & n10795 ) ;
  assign n10797 = ( ~n10425 & n10794 ) | ( ~n10425 & n10795 ) | ( n10794 & n10795 ) ;
  assign n10798 = ( n10425 & ~n10796 ) | ( n10425 & n10797 ) | ( ~n10796 & n10797 ) ;
  assign n10799 = ( ~n839 & n10793 ) | ( ~n839 & n10798 ) | ( n10793 & n10798 ) ;
  assign n10800 = ( n839 & ~n10426 ) | ( n839 & n10533 ) | ( ~n10426 & n10533 ) ;
  assign n10801 = n839 & ~n10426 ;
  assign n10802 = ( n10431 & n10800 ) | ( n10431 & n10801 ) | ( n10800 & n10801 ) ;
  assign n10803 = ( ~n10431 & n10800 ) | ( ~n10431 & n10801 ) | ( n10800 & n10801 ) ;
  assign n10804 = ( n10431 & ~n10802 ) | ( n10431 & n10803 ) | ( ~n10802 & n10803 ) ;
  assign n10805 = ( ~n746 & n10799 ) | ( ~n746 & n10804 ) | ( n10799 & n10804 ) ;
  assign n10806 = ( n746 & ~n10432 ) | ( n746 & n10533 ) | ( ~n10432 & n10533 ) ;
  assign n10807 = n746 & ~n10432 ;
  assign n10808 = ( n10437 & n10806 ) | ( n10437 & n10807 ) | ( n10806 & n10807 ) ;
  assign n10809 = ( ~n10437 & n10806 ) | ( ~n10437 & n10807 ) | ( n10806 & n10807 ) ;
  assign n10810 = ( n10437 & ~n10808 ) | ( n10437 & n10809 ) | ( ~n10808 & n10809 ) ;
  assign n10811 = ( ~n664 & n10805 ) | ( ~n664 & n10810 ) | ( n10805 & n10810 ) ;
  assign n10812 = ( n664 & ~n10438 ) | ( n664 & n10533 ) | ( ~n10438 & n10533 ) ;
  assign n10813 = n664 & ~n10438 ;
  assign n10814 = ( n10443 & n10812 ) | ( n10443 & n10813 ) | ( n10812 & n10813 ) ;
  assign n10815 = ( ~n10443 & n10812 ) | ( ~n10443 & n10813 ) | ( n10812 & n10813 ) ;
  assign n10816 = ( n10443 & ~n10814 ) | ( n10443 & n10815 ) | ( ~n10814 & n10815 ) ;
  assign n10817 = ( ~n588 & n10811 ) | ( ~n588 & n10816 ) | ( n10811 & n10816 ) ;
  assign n10818 = ~n588 & n10444 ;
  assign n10819 = ( ~n588 & n10444 ) | ( ~n588 & n10533 ) | ( n10444 & n10533 ) ;
  assign n10820 = ( ~n10449 & n10818 ) | ( ~n10449 & n10819 ) | ( n10818 & n10819 ) ;
  assign n10821 = ( n10449 & n10818 ) | ( n10449 & n10819 ) | ( n10818 & n10819 ) ;
  assign n10822 = ( n10449 & n10820 ) | ( n10449 & ~n10821 ) | ( n10820 & ~n10821 ) ;
  assign n10823 = ( ~n518 & n10817 ) | ( ~n518 & n10822 ) | ( n10817 & n10822 ) ;
  assign n10824 = ( n518 & ~n10450 ) | ( n518 & n10533 ) | ( ~n10450 & n10533 ) ;
  assign n10825 = n518 & ~n10450 ;
  assign n10826 = ( n10455 & n10824 ) | ( n10455 & n10825 ) | ( n10824 & n10825 ) ;
  assign n10827 = ( ~n10455 & n10824 ) | ( ~n10455 & n10825 ) | ( n10824 & n10825 ) ;
  assign n10828 = ( n10455 & ~n10826 ) | ( n10455 & n10827 ) | ( ~n10826 & n10827 ) ;
  assign n10829 = ( ~n454 & n10823 ) | ( ~n454 & n10828 ) | ( n10823 & n10828 ) ;
  assign n10830 = ( n454 & ~n10456 ) | ( n454 & n10533 ) | ( ~n10456 & n10533 ) ;
  assign n10831 = n454 & ~n10456 ;
  assign n10832 = ( n10461 & n10830 ) | ( n10461 & n10831 ) | ( n10830 & n10831 ) ;
  assign n10833 = ( ~n10461 & n10830 ) | ( ~n10461 & n10831 ) | ( n10830 & n10831 ) ;
  assign n10834 = ( n10461 & ~n10832 ) | ( n10461 & n10833 ) | ( ~n10832 & n10833 ) ;
  assign n10835 = ( ~n396 & n10829 ) | ( ~n396 & n10834 ) | ( n10829 & n10834 ) ;
  assign n10836 = ~n396 & n10462 ;
  assign n10837 = ( ~n396 & n10462 ) | ( ~n396 & n10533 ) | ( n10462 & n10533 ) ;
  assign n10838 = ( n10467 & n10836 ) | ( n10467 & n10837 ) | ( n10836 & n10837 ) ;
  assign n10839 = ( ~n10467 & n10836 ) | ( ~n10467 & n10837 ) | ( n10836 & n10837 ) ;
  assign n10840 = ( n10467 & ~n10838 ) | ( n10467 & n10839 ) | ( ~n10838 & n10839 ) ;
  assign n10841 = ( ~n344 & n10835 ) | ( ~n344 & n10840 ) | ( n10835 & n10840 ) ;
  assign n10842 = ( n344 & ~n10468 ) | ( n344 & n10533 ) | ( ~n10468 & n10533 ) ;
  assign n10843 = n344 & ~n10468 ;
  assign n10844 = ( n10473 & n10842 ) | ( n10473 & n10843 ) | ( n10842 & n10843 ) ;
  assign n10845 = ( ~n10473 & n10842 ) | ( ~n10473 & n10843 ) | ( n10842 & n10843 ) ;
  assign n10846 = ( n10473 & ~n10844 ) | ( n10473 & n10845 ) | ( ~n10844 & n10845 ) ;
  assign n10847 = ( ~n298 & n10841 ) | ( ~n298 & n10846 ) | ( n10841 & n10846 ) ;
  assign n10848 = ( n298 & ~n10474 ) | ( n298 & n10533 ) | ( ~n10474 & n10533 ) ;
  assign n10849 = n298 & ~n10474 ;
  assign n10850 = ( n10479 & n10848 ) | ( n10479 & n10849 ) | ( n10848 & n10849 ) ;
  assign n10851 = ( ~n10479 & n10848 ) | ( ~n10479 & n10849 ) | ( n10848 & n10849 ) ;
  assign n10852 = ( n10479 & ~n10850 ) | ( n10479 & n10851 ) | ( ~n10850 & n10851 ) ;
  assign n10853 = ( ~n258 & n10847 ) | ( ~n258 & n10852 ) | ( n10847 & n10852 ) ;
  assign n10854 = ~n258 & n10480 ;
  assign n10855 = ( ~n258 & n10480 ) | ( ~n258 & n10533 ) | ( n10480 & n10533 ) ;
  assign n10856 = ( ~n10485 & n10854 ) | ( ~n10485 & n10855 ) | ( n10854 & n10855 ) ;
  assign n10857 = ( n10485 & n10854 ) | ( n10485 & n10855 ) | ( n10854 & n10855 ) ;
  assign n10858 = ( n10485 & n10856 ) | ( n10485 & ~n10857 ) | ( n10856 & ~n10857 ) ;
  assign n10859 = ( ~n225 & n10853 ) | ( ~n225 & n10858 ) | ( n10853 & n10858 ) ;
  assign n10860 = n225 & ~n10486 ;
  assign n10861 = ( n225 & ~n10486 ) | ( n225 & n10533 ) | ( ~n10486 & n10533 ) ;
  assign n10862 = ( n10491 & n10860 ) | ( n10491 & n10861 ) | ( n10860 & n10861 ) ;
  assign n10863 = ( ~n10491 & n10860 ) | ( ~n10491 & n10861 ) | ( n10860 & n10861 ) ;
  assign n10864 = ( n10491 & ~n10862 ) | ( n10491 & n10863 ) | ( ~n10862 & n10863 ) ;
  assign n10865 = ( ~n197 & n10859 ) | ( ~n197 & n10864 ) | ( n10859 & n10864 ) ;
  assign n10866 = ~n197 & n10492 ;
  assign n10867 = ( ~n197 & n10492 ) | ( ~n197 & n10533 ) | ( n10492 & n10533 ) ;
  assign n10868 = ( ~n10497 & n10866 ) | ( ~n10497 & n10867 ) | ( n10866 & n10867 ) ;
  assign n10869 = ( n10497 & n10866 ) | ( n10497 & n10867 ) | ( n10866 & n10867 ) ;
  assign n10870 = ( n10497 & n10868 ) | ( n10497 & ~n10869 ) | ( n10868 & ~n10869 ) ;
  assign n10871 = ( ~n170 & n10865 ) | ( ~n170 & n10870 ) | ( n10865 & n10870 ) ;
  assign n10872 = ( n170 & ~n10498 ) | ( n170 & n10533 ) | ( ~n10498 & n10533 ) ;
  assign n10873 = n170 & ~n10498 ;
  assign n10874 = ( n10503 & n10872 ) | ( n10503 & n10873 ) | ( n10872 & n10873 ) ;
  assign n10875 = ( ~n10503 & n10872 ) | ( ~n10503 & n10873 ) | ( n10872 & n10873 ) ;
  assign n10876 = ( n10503 & ~n10874 ) | ( n10503 & n10875 ) | ( ~n10874 & n10875 ) ;
  assign n10877 = ( ~n142 & n10871 ) | ( ~n142 & n10876 ) | ( n10871 & n10876 ) ;
  assign n10878 = ~n142 & n10504 ;
  assign n10879 = ( ~n142 & n10504 ) | ( ~n142 & n10533 ) | ( n10504 & n10533 ) ;
  assign n10880 = ( n10509 & n10878 ) | ( n10509 & n10879 ) | ( n10878 & n10879 ) ;
  assign n10881 = ( ~n10509 & n10878 ) | ( ~n10509 & n10879 ) | ( n10878 & n10879 ) ;
  assign n10882 = ( n10509 & ~n10880 ) | ( n10509 & n10881 ) | ( ~n10880 & n10881 ) ;
  assign n10883 = ( ~n132 & n10877 ) | ( ~n132 & n10882 ) | ( n10877 & n10882 ) ;
  assign n10884 = n10538 & n10883 ;
  assign n10885 = n10526 | n10531 ;
  assign n10886 = n10883 | n10885 ;
  assign n10887 = ( ~n131 & n10884 ) | ( ~n131 & n10886 ) | ( n10884 & n10886 ) ;
  assign n10888 = ( n10539 & ~n10541 ) | ( n10539 & n10887 ) | ( ~n10541 & n10887 ) ;
  assign n10889 = ( n131 & n10538 ) | ( n131 & n10883 ) | ( n10538 & n10883 ) ;
  assign n10890 = n10527 & ~n10540 ;
  assign n10891 = ( n10883 & n10884 ) | ( n10883 & ~n10890 ) | ( n10884 & ~n10890 ) ;
  assign n10892 = n10889 & ~n10891 ;
  assign n10893 = ( n10527 & n10538 ) | ( n10527 & ~n10540 ) | ( n10538 & ~n10540 ) ;
  assign n10894 = n10883 | n10893 ;
  assign n10895 = ~n131 & n10889 ;
  assign n10896 = ( n10887 & ~n10894 ) | ( n10887 & n10895 ) | ( ~n10894 & n10895 ) ;
  assign n10897 = n10892 | n10896 ;
  assign n10898 = x6 | x7 ;
  assign n10899 = x8 | n10898 ;
  assign n10900 = n10533 & ~n10899 ;
  assign n10901 = ~n10542 & n10888 ;
  assign n10902 = ~n10533 & n10899 ;
  assign n10903 = ( x9 & ~n10888 ) | ( x9 & n10902 ) | ( ~n10888 & n10902 ) ;
  assign n10904 = ( ~n10900 & n10901 ) | ( ~n10900 & n10903 ) | ( n10901 & n10903 ) ;
  assign n10905 = n10533 & ~n10888 ;
  assign n10906 = ( x10 & n10901 ) | ( x10 & n10905 ) | ( n10901 & n10905 ) ;
  assign n10907 = ( ~x10 & n10901 ) | ( ~x10 & n10905 ) | ( n10901 & n10905 ) ;
  assign n10908 = ( x10 & ~n10906 ) | ( x10 & n10907 ) | ( ~n10906 & n10907 ) ;
  assign n10909 = ( ~n10180 & n10904 ) | ( ~n10180 & n10908 ) | ( n10904 & n10908 ) ;
  assign n10910 = ~n10180 & n10533 ;
  assign n10911 = ( n10549 & n10888 ) | ( n10549 & n10910 ) | ( n10888 & n10910 ) ;
  assign n10912 = ( ~x11 & n10907 ) | ( ~x11 & n10911 ) | ( n10907 & n10911 ) ;
  assign n10913 = ( x11 & n10907 ) | ( x11 & n10911 ) | ( n10907 & n10911 ) ;
  assign n10914 = ( x11 & n10912 ) | ( x11 & ~n10913 ) | ( n10912 & ~n10913 ) ;
  assign n10915 = ( ~n9834 & n10909 ) | ( ~n9834 & n10914 ) | ( n10909 & n10914 ) ;
  assign n10916 = n9834 & ~n10548 ;
  assign n10917 = ( n9834 & ~n10548 ) | ( n9834 & n10888 ) | ( ~n10548 & n10888 ) ;
  assign n10918 = ( n10552 & n10916 ) | ( n10552 & n10917 ) | ( n10916 & n10917 ) ;
  assign n10919 = ( ~n10552 & n10916 ) | ( ~n10552 & n10917 ) | ( n10916 & n10917 ) ;
  assign n10920 = ( n10552 & ~n10918 ) | ( n10552 & n10919 ) | ( ~n10918 & n10919 ) ;
  assign n10921 = ( ~n9497 & n10915 ) | ( ~n9497 & n10920 ) | ( n10915 & n10920 ) ;
  assign n10922 = n9497 & ~n10553 ;
  assign n10923 = ( n9497 & ~n10553 ) | ( n9497 & n10888 ) | ( ~n10553 & n10888 ) ;
  assign n10924 = ( ~n10558 & n10922 ) | ( ~n10558 & n10923 ) | ( n10922 & n10923 ) ;
  assign n10925 = ( n10558 & n10922 ) | ( n10558 & n10923 ) | ( n10922 & n10923 ) ;
  assign n10926 = ( n10558 & n10924 ) | ( n10558 & ~n10925 ) | ( n10924 & ~n10925 ) ;
  assign n10927 = ( ~n9167 & n10921 ) | ( ~n9167 & n10926 ) | ( n10921 & n10926 ) ;
  assign n10928 = ( n9167 & ~n10559 ) | ( n9167 & n10888 ) | ( ~n10559 & n10888 ) ;
  assign n10929 = n9167 & ~n10559 ;
  assign n10930 = ( n10564 & n10928 ) | ( n10564 & n10929 ) | ( n10928 & n10929 ) ;
  assign n10931 = ( ~n10564 & n10928 ) | ( ~n10564 & n10929 ) | ( n10928 & n10929 ) ;
  assign n10932 = ( n10564 & ~n10930 ) | ( n10564 & n10931 ) | ( ~n10930 & n10931 ) ;
  assign n10933 = ( ~n8838 & n10927 ) | ( ~n8838 & n10932 ) | ( n10927 & n10932 ) ;
  assign n10934 = ~n8838 & n10565 ;
  assign n10935 = ( ~n8838 & n10565 ) | ( ~n8838 & n10888 ) | ( n10565 & n10888 ) ;
  assign n10936 = ( n10570 & n10934 ) | ( n10570 & n10935 ) | ( n10934 & n10935 ) ;
  assign n10937 = ( ~n10570 & n10934 ) | ( ~n10570 & n10935 ) | ( n10934 & n10935 ) ;
  assign n10938 = ( n10570 & ~n10936 ) | ( n10570 & n10937 ) | ( ~n10936 & n10937 ) ;
  assign n10939 = ( ~n8517 & n10933 ) | ( ~n8517 & n10938 ) | ( n10933 & n10938 ) ;
  assign n10940 = ~n8517 & n10571 ;
  assign n10941 = ( ~n8517 & n10571 ) | ( ~n8517 & n10888 ) | ( n10571 & n10888 ) ;
  assign n10942 = ( ~n10576 & n10940 ) | ( ~n10576 & n10941 ) | ( n10940 & n10941 ) ;
  assign n10943 = ( n10576 & n10940 ) | ( n10576 & n10941 ) | ( n10940 & n10941 ) ;
  assign n10944 = ( n10576 & n10942 ) | ( n10576 & ~n10943 ) | ( n10942 & ~n10943 ) ;
  assign n10945 = ( ~n8201 & n10939 ) | ( ~n8201 & n10944 ) | ( n10939 & n10944 ) ;
  assign n10946 = ( n8201 & ~n10577 ) | ( n8201 & n10888 ) | ( ~n10577 & n10888 ) ;
  assign n10947 = n8201 & ~n10577 ;
  assign n10948 = ( n10582 & n10946 ) | ( n10582 & n10947 ) | ( n10946 & n10947 ) ;
  assign n10949 = ( ~n10582 & n10946 ) | ( ~n10582 & n10947 ) | ( n10946 & n10947 ) ;
  assign n10950 = ( n10582 & ~n10948 ) | ( n10582 & n10949 ) | ( ~n10948 & n10949 ) ;
  assign n10951 = ( ~n7897 & n10945 ) | ( ~n7897 & n10950 ) | ( n10945 & n10950 ) ;
  assign n10952 = n7897 & ~n10583 ;
  assign n10953 = ( n7897 & ~n10583 ) | ( n7897 & n10888 ) | ( ~n10583 & n10888 ) ;
  assign n10954 = ( n10588 & n10952 ) | ( n10588 & n10953 ) | ( n10952 & n10953 ) ;
  assign n10955 = ( ~n10588 & n10952 ) | ( ~n10588 & n10953 ) | ( n10952 & n10953 ) ;
  assign n10956 = ( n10588 & ~n10954 ) | ( n10588 & n10955 ) | ( ~n10954 & n10955 ) ;
  assign n10957 = ( ~n7594 & n10951 ) | ( ~n7594 & n10956 ) | ( n10951 & n10956 ) ;
  assign n10958 = ( n7594 & ~n10589 ) | ( n7594 & n10888 ) | ( ~n10589 & n10888 ) ;
  assign n10959 = n7594 & ~n10589 ;
  assign n10960 = ( n10594 & n10958 ) | ( n10594 & n10959 ) | ( n10958 & n10959 ) ;
  assign n10961 = ( ~n10594 & n10958 ) | ( ~n10594 & n10959 ) | ( n10958 & n10959 ) ;
  assign n10962 = ( n10594 & ~n10960 ) | ( n10594 & n10961 ) | ( ~n10960 & n10961 ) ;
  assign n10963 = ( ~n7296 & n10957 ) | ( ~n7296 & n10962 ) | ( n10957 & n10962 ) ;
  assign n10964 = ( n7296 & ~n10595 ) | ( n7296 & n10888 ) | ( ~n10595 & n10888 ) ;
  assign n10965 = n7296 & ~n10595 ;
  assign n10966 = ( n10600 & n10964 ) | ( n10600 & n10965 ) | ( n10964 & n10965 ) ;
  assign n10967 = ( ~n10600 & n10964 ) | ( ~n10600 & n10965 ) | ( n10964 & n10965 ) ;
  assign n10968 = ( n10600 & ~n10966 ) | ( n10600 & n10967 ) | ( ~n10966 & n10967 ) ;
  assign n10969 = ( ~n7006 & n10963 ) | ( ~n7006 & n10968 ) | ( n10963 & n10968 ) ;
  assign n10970 = ( n7006 & ~n10601 ) | ( n7006 & n10888 ) | ( ~n10601 & n10888 ) ;
  assign n10971 = n7006 & ~n10601 ;
  assign n10972 = ( n10606 & n10970 ) | ( n10606 & n10971 ) | ( n10970 & n10971 ) ;
  assign n10973 = ( ~n10606 & n10970 ) | ( ~n10606 & n10971 ) | ( n10970 & n10971 ) ;
  assign n10974 = ( n10606 & ~n10972 ) | ( n10606 & n10973 ) | ( ~n10972 & n10973 ) ;
  assign n10975 = ( ~n6723 & n10969 ) | ( ~n6723 & n10974 ) | ( n10969 & n10974 ) ;
  assign n10976 = ( n6723 & ~n10607 ) | ( n6723 & n10888 ) | ( ~n10607 & n10888 ) ;
  assign n10977 = n6723 & ~n10607 ;
  assign n10978 = ( n10612 & n10976 ) | ( n10612 & n10977 ) | ( n10976 & n10977 ) ;
  assign n10979 = ( ~n10612 & n10976 ) | ( ~n10612 & n10977 ) | ( n10976 & n10977 ) ;
  assign n10980 = ( n10612 & ~n10978 ) | ( n10612 & n10979 ) | ( ~n10978 & n10979 ) ;
  assign n10981 = ( ~n6442 & n10975 ) | ( ~n6442 & n10980 ) | ( n10975 & n10980 ) ;
  assign n10982 = ( n6442 & ~n10613 ) | ( n6442 & n10888 ) | ( ~n10613 & n10888 ) ;
  assign n10983 = n6442 & ~n10613 ;
  assign n10984 = ( n10618 & n10982 ) | ( n10618 & n10983 ) | ( n10982 & n10983 ) ;
  assign n10985 = ( ~n10618 & n10982 ) | ( ~n10618 & n10983 ) | ( n10982 & n10983 ) ;
  assign n10986 = ( n10618 & ~n10984 ) | ( n10618 & n10985 ) | ( ~n10984 & n10985 ) ;
  assign n10987 = ( ~n6172 & n10981 ) | ( ~n6172 & n10986 ) | ( n10981 & n10986 ) ;
  assign n10988 = ~n6172 & n10619 ;
  assign n10989 = ( ~n6172 & n10619 ) | ( ~n6172 & n10888 ) | ( n10619 & n10888 ) ;
  assign n10990 = ( ~n10624 & n10988 ) | ( ~n10624 & n10989 ) | ( n10988 & n10989 ) ;
  assign n10991 = ( n10624 & n10988 ) | ( n10624 & n10989 ) | ( n10988 & n10989 ) ;
  assign n10992 = ( n10624 & n10990 ) | ( n10624 & ~n10991 ) | ( n10990 & ~n10991 ) ;
  assign n10993 = ( ~n5905 & n10987 ) | ( ~n5905 & n10992 ) | ( n10987 & n10992 ) ;
  assign n10994 = ( n5905 & ~n10625 ) | ( n5905 & n10888 ) | ( ~n10625 & n10888 ) ;
  assign n10995 = n5905 & ~n10625 ;
  assign n10996 = ( n10630 & n10994 ) | ( n10630 & n10995 ) | ( n10994 & n10995 ) ;
  assign n10997 = ( ~n10630 & n10994 ) | ( ~n10630 & n10995 ) | ( n10994 & n10995 ) ;
  assign n10998 = ( n10630 & ~n10996 ) | ( n10630 & n10997 ) | ( ~n10996 & n10997 ) ;
  assign n10999 = ( ~n5642 & n10993 ) | ( ~n5642 & n10998 ) | ( n10993 & n10998 ) ;
  assign n11000 = ( n5642 & ~n10631 ) | ( n5642 & n10888 ) | ( ~n10631 & n10888 ) ;
  assign n11001 = n5642 & ~n10631 ;
  assign n11002 = ( n10636 & n11000 ) | ( n10636 & n11001 ) | ( n11000 & n11001 ) ;
  assign n11003 = ( ~n10636 & n11000 ) | ( ~n10636 & n11001 ) | ( n11000 & n11001 ) ;
  assign n11004 = ( n10636 & ~n11002 ) | ( n10636 & n11003 ) | ( ~n11002 & n11003 ) ;
  assign n11005 = ( ~n5386 & n10999 ) | ( ~n5386 & n11004 ) | ( n10999 & n11004 ) ;
  assign n11006 = ~n5386 & n10637 ;
  assign n11007 = ( ~n5386 & n10637 ) | ( ~n5386 & n10888 ) | ( n10637 & n10888 ) ;
  assign n11008 = ( ~n10642 & n11006 ) | ( ~n10642 & n11007 ) | ( n11006 & n11007 ) ;
  assign n11009 = ( n10642 & n11006 ) | ( n10642 & n11007 ) | ( n11006 & n11007 ) ;
  assign n11010 = ( n10642 & n11008 ) | ( n10642 & ~n11009 ) | ( n11008 & ~n11009 ) ;
  assign n11011 = ( ~n5139 & n11005 ) | ( ~n5139 & n11010 ) | ( n11005 & n11010 ) ;
  assign n11012 = ~n5139 & n10643 ;
  assign n11013 = ( ~n5139 & n10643 ) | ( ~n5139 & n10888 ) | ( n10643 & n10888 ) ;
  assign n11014 = ( ~n10648 & n11012 ) | ( ~n10648 & n11013 ) | ( n11012 & n11013 ) ;
  assign n11015 = ( n10648 & n11012 ) | ( n10648 & n11013 ) | ( n11012 & n11013 ) ;
  assign n11016 = ( n10648 & n11014 ) | ( n10648 & ~n11015 ) | ( n11014 & ~n11015 ) ;
  assign n11017 = ( ~n4898 & n11011 ) | ( ~n4898 & n11016 ) | ( n11011 & n11016 ) ;
  assign n11018 = ( n4898 & ~n10649 ) | ( n4898 & n10888 ) | ( ~n10649 & n10888 ) ;
  assign n11019 = n4898 & ~n10649 ;
  assign n11020 = ( n10654 & n11018 ) | ( n10654 & n11019 ) | ( n11018 & n11019 ) ;
  assign n11021 = ( ~n10654 & n11018 ) | ( ~n10654 & n11019 ) | ( n11018 & n11019 ) ;
  assign n11022 = ( n10654 & ~n11020 ) | ( n10654 & n11021 ) | ( ~n11020 & n11021 ) ;
  assign n11023 = ( ~n4661 & n11017 ) | ( ~n4661 & n11022 ) | ( n11017 & n11022 ) ;
  assign n11024 = ( n4661 & ~n10655 ) | ( n4661 & n10888 ) | ( ~n10655 & n10888 ) ;
  assign n11025 = n4661 & ~n10655 ;
  assign n11026 = ( n10660 & n11024 ) | ( n10660 & n11025 ) | ( n11024 & n11025 ) ;
  assign n11027 = ( ~n10660 & n11024 ) | ( ~n10660 & n11025 ) | ( n11024 & n11025 ) ;
  assign n11028 = ( n10660 & ~n11026 ) | ( n10660 & n11027 ) | ( ~n11026 & n11027 ) ;
  assign n11029 = ( ~n4432 & n11023 ) | ( ~n4432 & n11028 ) | ( n11023 & n11028 ) ;
  assign n11030 = ( n4432 & ~n10661 ) | ( n4432 & n10888 ) | ( ~n10661 & n10888 ) ;
  assign n11031 = n4432 & ~n10661 ;
  assign n11032 = ( n10666 & n11030 ) | ( n10666 & n11031 ) | ( n11030 & n11031 ) ;
  assign n11033 = ( ~n10666 & n11030 ) | ( ~n10666 & n11031 ) | ( n11030 & n11031 ) ;
  assign n11034 = ( n10666 & ~n11032 ) | ( n10666 & n11033 ) | ( ~n11032 & n11033 ) ;
  assign n11035 = ( ~n4203 & n11029 ) | ( ~n4203 & n11034 ) | ( n11029 & n11034 ) ;
  assign n11036 = ( n4203 & ~n10667 ) | ( n4203 & n10888 ) | ( ~n10667 & n10888 ) ;
  assign n11037 = n4203 & ~n10667 ;
  assign n11038 = ( n10672 & n11036 ) | ( n10672 & n11037 ) | ( n11036 & n11037 ) ;
  assign n11039 = ( ~n10672 & n11036 ) | ( ~n10672 & n11037 ) | ( n11036 & n11037 ) ;
  assign n11040 = ( n10672 & ~n11038 ) | ( n10672 & n11039 ) | ( ~n11038 & n11039 ) ;
  assign n11041 = ( ~n3985 & n11035 ) | ( ~n3985 & n11040 ) | ( n11035 & n11040 ) ;
  assign n11042 = ~n3985 & n10673 ;
  assign n11043 = ( ~n3985 & n10673 ) | ( ~n3985 & n10888 ) | ( n10673 & n10888 ) ;
  assign n11044 = ( n10678 & n11042 ) | ( n10678 & n11043 ) | ( n11042 & n11043 ) ;
  assign n11045 = ( ~n10678 & n11042 ) | ( ~n10678 & n11043 ) | ( n11042 & n11043 ) ;
  assign n11046 = ( n10678 & ~n11044 ) | ( n10678 & n11045 ) | ( ~n11044 & n11045 ) ;
  assign n11047 = ( ~n3772 & n11041 ) | ( ~n3772 & n11046 ) | ( n11041 & n11046 ) ;
  assign n11048 = ( n3772 & ~n10679 ) | ( n3772 & n10888 ) | ( ~n10679 & n10888 ) ;
  assign n11049 = n3772 & ~n10679 ;
  assign n11050 = ( n10684 & n11048 ) | ( n10684 & n11049 ) | ( n11048 & n11049 ) ;
  assign n11051 = ( ~n10684 & n11048 ) | ( ~n10684 & n11049 ) | ( n11048 & n11049 ) ;
  assign n11052 = ( n10684 & ~n11050 ) | ( n10684 & n11051 ) | ( ~n11050 & n11051 ) ;
  assign n11053 = ( ~n3567 & n11047 ) | ( ~n3567 & n11052 ) | ( n11047 & n11052 ) ;
  assign n11054 = ( n3567 & ~n10685 ) | ( n3567 & n10888 ) | ( ~n10685 & n10888 ) ;
  assign n11055 = n3567 & ~n10685 ;
  assign n11056 = ( n10690 & n11054 ) | ( n10690 & n11055 ) | ( n11054 & n11055 ) ;
  assign n11057 = ( ~n10690 & n11054 ) | ( ~n10690 & n11055 ) | ( n11054 & n11055 ) ;
  assign n11058 = ( n10690 & ~n11056 ) | ( n10690 & n11057 ) | ( ~n11056 & n11057 ) ;
  assign n11059 = ( ~n3362 & n11053 ) | ( ~n3362 & n11058 ) | ( n11053 & n11058 ) ;
  assign n11060 = ( n3362 & ~n10691 ) | ( n3362 & n10888 ) | ( ~n10691 & n10888 ) ;
  assign n11061 = n3362 & ~n10691 ;
  assign n11062 = ( n10696 & n11060 ) | ( n10696 & n11061 ) | ( n11060 & n11061 ) ;
  assign n11063 = ( ~n10696 & n11060 ) | ( ~n10696 & n11061 ) | ( n11060 & n11061 ) ;
  assign n11064 = ( n10696 & ~n11062 ) | ( n10696 & n11063 ) | ( ~n11062 & n11063 ) ;
  assign n11065 = ( ~n3169 & n11059 ) | ( ~n3169 & n11064 ) | ( n11059 & n11064 ) ;
  assign n11066 = ~n3169 & n10697 ;
  assign n11067 = ( ~n3169 & n10697 ) | ( ~n3169 & n10888 ) | ( n10697 & n10888 ) ;
  assign n11068 = ( ~n10702 & n11066 ) | ( ~n10702 & n11067 ) | ( n11066 & n11067 ) ;
  assign n11069 = ( n10702 & n11066 ) | ( n10702 & n11067 ) | ( n11066 & n11067 ) ;
  assign n11070 = ( n10702 & n11068 ) | ( n10702 & ~n11069 ) | ( n11068 & ~n11069 ) ;
  assign n11071 = ( ~n2979 & n11065 ) | ( ~n2979 & n11070 ) | ( n11065 & n11070 ) ;
  assign n11072 = ( n2979 & ~n10703 ) | ( n2979 & n10888 ) | ( ~n10703 & n10888 ) ;
  assign n11073 = n2979 & ~n10703 ;
  assign n11074 = ( n10708 & n11072 ) | ( n10708 & n11073 ) | ( n11072 & n11073 ) ;
  assign n11075 = ( ~n10708 & n11072 ) | ( ~n10708 & n11073 ) | ( n11072 & n11073 ) ;
  assign n11076 = ( n10708 & ~n11074 ) | ( n10708 & n11075 ) | ( ~n11074 & n11075 ) ;
  assign n11077 = ( ~n2791 & n11071 ) | ( ~n2791 & n11076 ) | ( n11071 & n11076 ) ;
  assign n11078 = ~n2791 & n10709 ;
  assign n11079 = ( ~n2791 & n10709 ) | ( ~n2791 & n10888 ) | ( n10709 & n10888 ) ;
  assign n11080 = ( ~n10714 & n11078 ) | ( ~n10714 & n11079 ) | ( n11078 & n11079 ) ;
  assign n11081 = ( n10714 & n11078 ) | ( n10714 & n11079 ) | ( n11078 & n11079 ) ;
  assign n11082 = ( n10714 & n11080 ) | ( n10714 & ~n11081 ) | ( n11080 & ~n11081 ) ;
  assign n11083 = ( ~n2615 & n11077 ) | ( ~n2615 & n11082 ) | ( n11077 & n11082 ) ;
  assign n11084 = ( n2615 & ~n10715 ) | ( n2615 & n10888 ) | ( ~n10715 & n10888 ) ;
  assign n11085 = n2615 & ~n10715 ;
  assign n11086 = ( n10720 & n11084 ) | ( n10720 & n11085 ) | ( n11084 & n11085 ) ;
  assign n11087 = ( ~n10720 & n11084 ) | ( ~n10720 & n11085 ) | ( n11084 & n11085 ) ;
  assign n11088 = ( n10720 & ~n11086 ) | ( n10720 & n11087 ) | ( ~n11086 & n11087 ) ;
  assign n11089 = ( ~n2443 & n11083 ) | ( ~n2443 & n11088 ) | ( n11083 & n11088 ) ;
  assign n11090 = ( n2443 & ~n10721 ) | ( n2443 & n10888 ) | ( ~n10721 & n10888 ) ;
  assign n11091 = n2443 & ~n10721 ;
  assign n11092 = ( n10726 & n11090 ) | ( n10726 & n11091 ) | ( n11090 & n11091 ) ;
  assign n11093 = ( ~n10726 & n11090 ) | ( ~n10726 & n11091 ) | ( n11090 & n11091 ) ;
  assign n11094 = ( n10726 & ~n11092 ) | ( n10726 & n11093 ) | ( ~n11092 & n11093 ) ;
  assign n11095 = ( ~n2277 & n11089 ) | ( ~n2277 & n11094 ) | ( n11089 & n11094 ) ;
  assign n11096 = ( n2277 & ~n10727 ) | ( n2277 & n10888 ) | ( ~n10727 & n10888 ) ;
  assign n11097 = n2277 & ~n10727 ;
  assign n11098 = ( n10732 & n11096 ) | ( n10732 & n11097 ) | ( n11096 & n11097 ) ;
  assign n11099 = ( ~n10732 & n11096 ) | ( ~n10732 & n11097 ) | ( n11096 & n11097 ) ;
  assign n11100 = ( n10732 & ~n11098 ) | ( n10732 & n11099 ) | ( ~n11098 & n11099 ) ;
  assign n11101 = ( ~n2111 & n11095 ) | ( ~n2111 & n11100 ) | ( n11095 & n11100 ) ;
  assign n11102 = ~n2111 & n10733 ;
  assign n11103 = ( ~n2111 & n10733 ) | ( ~n2111 & n10888 ) | ( n10733 & n10888 ) ;
  assign n11104 = ( ~n10738 & n11102 ) | ( ~n10738 & n11103 ) | ( n11102 & n11103 ) ;
  assign n11105 = ( n10738 & n11102 ) | ( n10738 & n11103 ) | ( n11102 & n11103 ) ;
  assign n11106 = ( n10738 & n11104 ) | ( n10738 & ~n11105 ) | ( n11104 & ~n11105 ) ;
  assign n11107 = ( ~n1949 & n11101 ) | ( ~n1949 & n11106 ) | ( n11101 & n11106 ) ;
  assign n11108 = ( n1949 & ~n10739 ) | ( n1949 & n10888 ) | ( ~n10739 & n10888 ) ;
  assign n11109 = n1949 & ~n10739 ;
  assign n11110 = ( n10744 & n11108 ) | ( n10744 & n11109 ) | ( n11108 & n11109 ) ;
  assign n11111 = ( ~n10744 & n11108 ) | ( ~n10744 & n11109 ) | ( n11108 & n11109 ) ;
  assign n11112 = ( n10744 & ~n11110 ) | ( n10744 & n11111 ) | ( ~n11110 & n11111 ) ;
  assign n11113 = ( ~n1802 & n11107 ) | ( ~n1802 & n11112 ) | ( n11107 & n11112 ) ;
  assign n11114 = ( n1802 & ~n10745 ) | ( n1802 & n10888 ) | ( ~n10745 & n10888 ) ;
  assign n11115 = n1802 & ~n10745 ;
  assign n11116 = ( n10750 & n11114 ) | ( n10750 & n11115 ) | ( n11114 & n11115 ) ;
  assign n11117 = ( ~n10750 & n11114 ) | ( ~n10750 & n11115 ) | ( n11114 & n11115 ) ;
  assign n11118 = ( n10750 & ~n11116 ) | ( n10750 & n11117 ) | ( ~n11116 & n11117 ) ;
  assign n11119 = ( ~n1661 & n11113 ) | ( ~n1661 & n11118 ) | ( n11113 & n11118 ) ;
  assign n11120 = ( n1661 & ~n10751 ) | ( n1661 & n10888 ) | ( ~n10751 & n10888 ) ;
  assign n11121 = n1661 & ~n10751 ;
  assign n11122 = ( n10756 & n11120 ) | ( n10756 & n11121 ) | ( n11120 & n11121 ) ;
  assign n11123 = ( ~n10756 & n11120 ) | ( ~n10756 & n11121 ) | ( n11120 & n11121 ) ;
  assign n11124 = ( n10756 & ~n11122 ) | ( n10756 & n11123 ) | ( ~n11122 & n11123 ) ;
  assign n11125 = ( ~n1523 & n11119 ) | ( ~n1523 & n11124 ) | ( n11119 & n11124 ) ;
  assign n11126 = ( n1523 & ~n10757 ) | ( n1523 & n10888 ) | ( ~n10757 & n10888 ) ;
  assign n11127 = n1523 & ~n10757 ;
  assign n11128 = ( n10762 & n11126 ) | ( n10762 & n11127 ) | ( n11126 & n11127 ) ;
  assign n11129 = ( ~n10762 & n11126 ) | ( ~n10762 & n11127 ) | ( n11126 & n11127 ) ;
  assign n11130 = ( n10762 & ~n11128 ) | ( n10762 & n11129 ) | ( ~n11128 & n11129 ) ;
  assign n11131 = ( ~n1393 & n11125 ) | ( ~n1393 & n11130 ) | ( n11125 & n11130 ) ;
  assign n11132 = ~n1393 & n10763 ;
  assign n11133 = ( ~n1393 & n10763 ) | ( ~n1393 & n10888 ) | ( n10763 & n10888 ) ;
  assign n11134 = ( ~n10768 & n11132 ) | ( ~n10768 & n11133 ) | ( n11132 & n11133 ) ;
  assign n11135 = ( n10768 & n11132 ) | ( n10768 & n11133 ) | ( n11132 & n11133 ) ;
  assign n11136 = ( n10768 & n11134 ) | ( n10768 & ~n11135 ) | ( n11134 & ~n11135 ) ;
  assign n11137 = ( ~n1266 & n11131 ) | ( ~n1266 & n11136 ) | ( n11131 & n11136 ) ;
  assign n11138 = ( n1266 & ~n10769 ) | ( n1266 & n10888 ) | ( ~n10769 & n10888 ) ;
  assign n11139 = n1266 & ~n10769 ;
  assign n11140 = ( n10774 & n11138 ) | ( n10774 & n11139 ) | ( n11138 & n11139 ) ;
  assign n11141 = ( ~n10774 & n11138 ) | ( ~n10774 & n11139 ) | ( n11138 & n11139 ) ;
  assign n11142 = ( n10774 & ~n11140 ) | ( n10774 & n11141 ) | ( ~n11140 & n11141 ) ;
  assign n11143 = ( ~n1150 & n11137 ) | ( ~n1150 & n11142 ) | ( n11137 & n11142 ) ;
  assign n11144 = ( n1150 & ~n10775 ) | ( n1150 & n10888 ) | ( ~n10775 & n10888 ) ;
  assign n11145 = n1150 & ~n10775 ;
  assign n11146 = ( n10780 & n11144 ) | ( n10780 & n11145 ) | ( n11144 & n11145 ) ;
  assign n11147 = ( ~n10780 & n11144 ) | ( ~n10780 & n11145 ) | ( n11144 & n11145 ) ;
  assign n11148 = ( n10780 & ~n11146 ) | ( n10780 & n11147 ) | ( ~n11146 & n11147 ) ;
  assign n11149 = ( ~n1038 & n11143 ) | ( ~n1038 & n11148 ) | ( n11143 & n11148 ) ;
  assign n11150 = ~n1038 & n10781 ;
  assign n11151 = ( ~n1038 & n10781 ) | ( ~n1038 & n10888 ) | ( n10781 & n10888 ) ;
  assign n11152 = ( ~n10786 & n11150 ) | ( ~n10786 & n11151 ) | ( n11150 & n11151 ) ;
  assign n11153 = ( n10786 & n11150 ) | ( n10786 & n11151 ) | ( n11150 & n11151 ) ;
  assign n11154 = ( n10786 & n11152 ) | ( n10786 & ~n11153 ) | ( n11152 & ~n11153 ) ;
  assign n11155 = ( ~n933 & n11149 ) | ( ~n933 & n11154 ) | ( n11149 & n11154 ) ;
  assign n11156 = ~n933 & n10787 ;
  assign n11157 = ( ~n933 & n10787 ) | ( ~n933 & n10888 ) | ( n10787 & n10888 ) ;
  assign n11158 = ( ~n10792 & n11156 ) | ( ~n10792 & n11157 ) | ( n11156 & n11157 ) ;
  assign n11159 = ( n10792 & n11156 ) | ( n10792 & n11157 ) | ( n11156 & n11157 ) ;
  assign n11160 = ( n10792 & n11158 ) | ( n10792 & ~n11159 ) | ( n11158 & ~n11159 ) ;
  assign n11161 = ( ~n839 & n11155 ) | ( ~n839 & n11160 ) | ( n11155 & n11160 ) ;
  assign n11162 = ~n839 & n10793 ;
  assign n11163 = ( ~n839 & n10793 ) | ( ~n839 & n10888 ) | ( n10793 & n10888 ) ;
  assign n11164 = ( ~n10798 & n11162 ) | ( ~n10798 & n11163 ) | ( n11162 & n11163 ) ;
  assign n11165 = ( n10798 & n11162 ) | ( n10798 & n11163 ) | ( n11162 & n11163 ) ;
  assign n11166 = ( n10798 & n11164 ) | ( n10798 & ~n11165 ) | ( n11164 & ~n11165 ) ;
  assign n11167 = ( ~n746 & n11161 ) | ( ~n746 & n11166 ) | ( n11161 & n11166 ) ;
  assign n11168 = ( n746 & ~n10799 ) | ( n746 & n10888 ) | ( ~n10799 & n10888 ) ;
  assign n11169 = n746 & ~n10799 ;
  assign n11170 = ( n10804 & n11168 ) | ( n10804 & n11169 ) | ( n11168 & n11169 ) ;
  assign n11171 = ( ~n10804 & n11168 ) | ( ~n10804 & n11169 ) | ( n11168 & n11169 ) ;
  assign n11172 = ( n10804 & ~n11170 ) | ( n10804 & n11171 ) | ( ~n11170 & n11171 ) ;
  assign n11173 = ( ~n664 & n11167 ) | ( ~n664 & n11172 ) | ( n11167 & n11172 ) ;
  assign n11174 = ( n664 & ~n10805 ) | ( n664 & n10888 ) | ( ~n10805 & n10888 ) ;
  assign n11175 = n664 & ~n10805 ;
  assign n11176 = ( n10810 & n11174 ) | ( n10810 & n11175 ) | ( n11174 & n11175 ) ;
  assign n11177 = ( ~n10810 & n11174 ) | ( ~n10810 & n11175 ) | ( n11174 & n11175 ) ;
  assign n11178 = ( n10810 & ~n11176 ) | ( n10810 & n11177 ) | ( ~n11176 & n11177 ) ;
  assign n11179 = ( ~n588 & n11173 ) | ( ~n588 & n11178 ) | ( n11173 & n11178 ) ;
  assign n11180 = ~n588 & n10811 ;
  assign n11181 = ( ~n588 & n10811 ) | ( ~n588 & n10888 ) | ( n10811 & n10888 ) ;
  assign n11182 = ( ~n10816 & n11180 ) | ( ~n10816 & n11181 ) | ( n11180 & n11181 ) ;
  assign n11183 = ( n10816 & n11180 ) | ( n10816 & n11181 ) | ( n11180 & n11181 ) ;
  assign n11184 = ( n10816 & n11182 ) | ( n10816 & ~n11183 ) | ( n11182 & ~n11183 ) ;
  assign n11185 = ( ~n518 & n11179 ) | ( ~n518 & n11184 ) | ( n11179 & n11184 ) ;
  assign n11186 = ( n518 & ~n10817 ) | ( n518 & n10888 ) | ( ~n10817 & n10888 ) ;
  assign n11187 = n518 & ~n10817 ;
  assign n11188 = ( n10822 & n11186 ) | ( n10822 & n11187 ) | ( n11186 & n11187 ) ;
  assign n11189 = ( ~n10822 & n11186 ) | ( ~n10822 & n11187 ) | ( n11186 & n11187 ) ;
  assign n11190 = ( n10822 & ~n11188 ) | ( n10822 & n11189 ) | ( ~n11188 & n11189 ) ;
  assign n11191 = ( ~n454 & n11185 ) | ( ~n454 & n11190 ) | ( n11185 & n11190 ) ;
  assign n11192 = ( n454 & ~n10823 ) | ( n454 & n10888 ) | ( ~n10823 & n10888 ) ;
  assign n11193 = n454 & ~n10823 ;
  assign n11194 = ( n10828 & n11192 ) | ( n10828 & n11193 ) | ( n11192 & n11193 ) ;
  assign n11195 = ( ~n10828 & n11192 ) | ( ~n10828 & n11193 ) | ( n11192 & n11193 ) ;
  assign n11196 = ( n10828 & ~n11194 ) | ( n10828 & n11195 ) | ( ~n11194 & n11195 ) ;
  assign n11197 = ( ~n396 & n11191 ) | ( ~n396 & n11196 ) | ( n11191 & n11196 ) ;
  assign n11198 = ~n396 & n10829 ;
  assign n11199 = ( ~n396 & n10829 ) | ( ~n396 & n10888 ) | ( n10829 & n10888 ) ;
  assign n11200 = ( n10834 & n11198 ) | ( n10834 & n11199 ) | ( n11198 & n11199 ) ;
  assign n11201 = ( ~n10834 & n11198 ) | ( ~n10834 & n11199 ) | ( n11198 & n11199 ) ;
  assign n11202 = ( n10834 & ~n11200 ) | ( n10834 & n11201 ) | ( ~n11200 & n11201 ) ;
  assign n11203 = ( ~n344 & n11197 ) | ( ~n344 & n11202 ) | ( n11197 & n11202 ) ;
  assign n11204 = ( n344 & ~n10835 ) | ( n344 & n10888 ) | ( ~n10835 & n10888 ) ;
  assign n11205 = n344 & ~n10835 ;
  assign n11206 = ( n10840 & n11204 ) | ( n10840 & n11205 ) | ( n11204 & n11205 ) ;
  assign n11207 = ( ~n10840 & n11204 ) | ( ~n10840 & n11205 ) | ( n11204 & n11205 ) ;
  assign n11208 = ( n10840 & ~n11206 ) | ( n10840 & n11207 ) | ( ~n11206 & n11207 ) ;
  assign n11209 = ( ~n298 & n11203 ) | ( ~n298 & n11208 ) | ( n11203 & n11208 ) ;
  assign n11210 = ( n298 & ~n10841 ) | ( n298 & n10888 ) | ( ~n10841 & n10888 ) ;
  assign n11211 = n298 & ~n10841 ;
  assign n11212 = ( n10846 & n11210 ) | ( n10846 & n11211 ) | ( n11210 & n11211 ) ;
  assign n11213 = ( ~n10846 & n11210 ) | ( ~n10846 & n11211 ) | ( n11210 & n11211 ) ;
  assign n11214 = ( n10846 & ~n11212 ) | ( n10846 & n11213 ) | ( ~n11212 & n11213 ) ;
  assign n11215 = ( ~n258 & n11209 ) | ( ~n258 & n11214 ) | ( n11209 & n11214 ) ;
  assign n11216 = n258 & ~n10847 ;
  assign n11217 = ( n258 & ~n10847 ) | ( n258 & n10888 ) | ( ~n10847 & n10888 ) ;
  assign n11218 = ( n10852 & n11216 ) | ( n10852 & n11217 ) | ( n11216 & n11217 ) ;
  assign n11219 = ( ~n10852 & n11216 ) | ( ~n10852 & n11217 ) | ( n11216 & n11217 ) ;
  assign n11220 = ( n10852 & ~n11218 ) | ( n10852 & n11219 ) | ( ~n11218 & n11219 ) ;
  assign n11221 = ( ~n225 & n11215 ) | ( ~n225 & n11220 ) | ( n11215 & n11220 ) ;
  assign n11222 = ( n225 & ~n10853 ) | ( n225 & n10888 ) | ( ~n10853 & n10888 ) ;
  assign n11223 = n225 & ~n10853 ;
  assign n11224 = ( n10858 & n11222 ) | ( n10858 & n11223 ) | ( n11222 & n11223 ) ;
  assign n11225 = ( ~n10858 & n11222 ) | ( ~n10858 & n11223 ) | ( n11222 & n11223 ) ;
  assign n11226 = ( n10858 & ~n11224 ) | ( n10858 & n11225 ) | ( ~n11224 & n11225 ) ;
  assign n11227 = ( ~n197 & n11221 ) | ( ~n197 & n11226 ) | ( n11221 & n11226 ) ;
  assign n11228 = ~n197 & n10859 ;
  assign n11229 = ( ~n197 & n10859 ) | ( ~n197 & n10888 ) | ( n10859 & n10888 ) ;
  assign n11230 = ( ~n10864 & n11228 ) | ( ~n10864 & n11229 ) | ( n11228 & n11229 ) ;
  assign n11231 = ( n10864 & n11228 ) | ( n10864 & n11229 ) | ( n11228 & n11229 ) ;
  assign n11232 = ( n10864 & n11230 ) | ( n10864 & ~n11231 ) | ( n11230 & ~n11231 ) ;
  assign n11233 = ( ~n170 & n11227 ) | ( ~n170 & n11232 ) | ( n11227 & n11232 ) ;
  assign n11234 = ~n170 & n10865 ;
  assign n11235 = ( ~n170 & n10865 ) | ( ~n170 & n10888 ) | ( n10865 & n10888 ) ;
  assign n11236 = ( n10870 & n11234 ) | ( n10870 & n11235 ) | ( n11234 & n11235 ) ;
  assign n11237 = ( ~n10870 & n11234 ) | ( ~n10870 & n11235 ) | ( n11234 & n11235 ) ;
  assign n11238 = ( n10870 & ~n11236 ) | ( n10870 & n11237 ) | ( ~n11236 & n11237 ) ;
  assign n11239 = ( ~n142 & n11233 ) | ( ~n142 & n11238 ) | ( n11233 & n11238 ) ;
  assign n11240 = ( n142 & ~n10871 ) | ( n142 & n10888 ) | ( ~n10871 & n10888 ) ;
  assign n11241 = n142 & ~n10871 ;
  assign n11242 = ( n10876 & n11240 ) | ( n10876 & n11241 ) | ( n11240 & n11241 ) ;
  assign n11243 = ( ~n10876 & n11240 ) | ( ~n10876 & n11241 ) | ( n11240 & n11241 ) ;
  assign n11244 = ( n10876 & ~n11242 ) | ( n10876 & n11243 ) | ( ~n11242 & n11243 ) ;
  assign n11245 = ( ~n132 & n11239 ) | ( ~n132 & n11244 ) | ( n11239 & n11244 ) ;
  assign n11246 = ~n132 & n10877 ;
  assign n11247 = ( ~n132 & n10877 ) | ( ~n132 & n10888 ) | ( n10877 & n10888 ) ;
  assign n11248 = ( ~n10882 & n11246 ) | ( ~n10882 & n11247 ) | ( n11246 & n11247 ) ;
  assign n11249 = ( n10882 & n11246 ) | ( n10882 & n11247 ) | ( n11246 & n11247 ) ;
  assign n11250 = ( n10882 & n11248 ) | ( n10882 & ~n11249 ) | ( n11248 & ~n11249 ) ;
  assign n11251 = ( ~n131 & n11245 ) | ( ~n131 & n11250 ) | ( n11245 & n11250 ) ;
  assign n11252 = n10897 | n11251 ;
  assign n11253 = n10888 & ~n11252 ;
  assign n11254 = ~n10898 & n11252 ;
  assign n11255 = ( x8 & n11253 ) | ( x8 & n11254 ) | ( n11253 & n11254 ) ;
  assign n11256 = ( ~x8 & n11253 ) | ( ~x8 & n11254 ) | ( n11253 & n11254 ) ;
  assign n11257 = ( x8 & ~n11255 ) | ( x8 & n11256 ) | ( ~n11255 & n11256 ) ;
  assign n11258 = x4 | x5 ;
  assign n11259 = x6 | n11258 ;
  assign n11260 = ~n10888 & n11259 ;
  assign n11261 = ( x7 & ~n11252 ) | ( x7 & n11260 ) | ( ~n11252 & n11260 ) ;
  assign n11262 = n10888 & ~n11259 ;
  assign n11263 = ( n11254 & n11261 ) | ( n11254 & ~n11262 ) | ( n11261 & ~n11262 ) ;
  assign n11264 = ( ~n10533 & n11257 ) | ( ~n10533 & n11263 ) | ( n11257 & n11263 ) ;
  assign n11265 = ~n10533 & n10888 ;
  assign n11266 = ( n10905 & n11252 ) | ( n10905 & n11265 ) | ( n11252 & n11265 ) ;
  assign n11267 = ( x9 & n11256 ) | ( x9 & n11266 ) | ( n11256 & n11266 ) ;
  assign n11268 = ( ~x9 & n11256 ) | ( ~x9 & n11266 ) | ( n11256 & n11266 ) ;
  assign n11269 = ( x9 & ~n11267 ) | ( x9 & n11268 ) | ( ~n11267 & n11268 ) ;
  assign n11270 = ( ~n10180 & n11264 ) | ( ~n10180 & n11269 ) | ( n11264 & n11269 ) ;
  assign n11271 = n10180 & ~n10904 ;
  assign n11272 = ( n10180 & ~n10904 ) | ( n10180 & n11252 ) | ( ~n10904 & n11252 ) ;
  assign n11273 = ( n10908 & n11271 ) | ( n10908 & n11272 ) | ( n11271 & n11272 ) ;
  assign n11274 = ( ~n10908 & n11271 ) | ( ~n10908 & n11272 ) | ( n11271 & n11272 ) ;
  assign n11275 = ( n10908 & ~n11273 ) | ( n10908 & n11274 ) | ( ~n11273 & n11274 ) ;
  assign n11276 = ( ~n9834 & n11270 ) | ( ~n9834 & n11275 ) | ( n11270 & n11275 ) ;
  assign n11277 = ( n9834 & ~n10909 ) | ( n9834 & n11252 ) | ( ~n10909 & n11252 ) ;
  assign n11278 = n9834 & ~n10909 ;
  assign n11279 = ( n10914 & n11277 ) | ( n10914 & n11278 ) | ( n11277 & n11278 ) ;
  assign n11280 = ( ~n10914 & n11277 ) | ( ~n10914 & n11278 ) | ( n11277 & n11278 ) ;
  assign n11281 = ( n10914 & ~n11279 ) | ( n10914 & n11280 ) | ( ~n11279 & n11280 ) ;
  assign n11282 = ( ~n9497 & n11276 ) | ( ~n9497 & n11281 ) | ( n11276 & n11281 ) ;
  assign n11283 = n9497 & ~n10915 ;
  assign n11284 = ( n9497 & ~n10915 ) | ( n9497 & n11252 ) | ( ~n10915 & n11252 ) ;
  assign n11285 = ( n10920 & n11283 ) | ( n10920 & n11284 ) | ( n11283 & n11284 ) ;
  assign n11286 = ( ~n10920 & n11283 ) | ( ~n10920 & n11284 ) | ( n11283 & n11284 ) ;
  assign n11287 = ( n10920 & ~n11285 ) | ( n10920 & n11286 ) | ( ~n11285 & n11286 ) ;
  assign n11288 = ( ~n9167 & n11282 ) | ( ~n9167 & n11287 ) | ( n11282 & n11287 ) ;
  assign n11289 = n9167 & ~n10921 ;
  assign n11290 = ( n9167 & ~n10921 ) | ( n9167 & n11252 ) | ( ~n10921 & n11252 ) ;
  assign n11291 = ( n10926 & n11289 ) | ( n10926 & n11290 ) | ( n11289 & n11290 ) ;
  assign n11292 = ( ~n10926 & n11289 ) | ( ~n10926 & n11290 ) | ( n11289 & n11290 ) ;
  assign n11293 = ( n10926 & ~n11291 ) | ( n10926 & n11292 ) | ( ~n11291 & n11292 ) ;
  assign n11294 = ( ~n8838 & n11288 ) | ( ~n8838 & n11293 ) | ( n11288 & n11293 ) ;
  assign n11295 = ( n8838 & ~n10927 ) | ( n8838 & n11252 ) | ( ~n10927 & n11252 ) ;
  assign n11296 = n8838 & ~n10927 ;
  assign n11297 = ( n10932 & n11295 ) | ( n10932 & n11296 ) | ( n11295 & n11296 ) ;
  assign n11298 = ( ~n10932 & n11295 ) | ( ~n10932 & n11296 ) | ( n11295 & n11296 ) ;
  assign n11299 = ( n10932 & ~n11297 ) | ( n10932 & n11298 ) | ( ~n11297 & n11298 ) ;
  assign n11300 = ( ~n8517 & n11294 ) | ( ~n8517 & n11299 ) | ( n11294 & n11299 ) ;
  assign n11301 = ~n8517 & n10933 ;
  assign n11302 = ( ~n8517 & n10933 ) | ( ~n8517 & n11252 ) | ( n10933 & n11252 ) ;
  assign n11303 = ( ~n10938 & n11301 ) | ( ~n10938 & n11302 ) | ( n11301 & n11302 ) ;
  assign n11304 = ( n10938 & n11301 ) | ( n10938 & n11302 ) | ( n11301 & n11302 ) ;
  assign n11305 = ( n10938 & n11303 ) | ( n10938 & ~n11304 ) | ( n11303 & ~n11304 ) ;
  assign n11306 = ( ~n8201 & n11300 ) | ( ~n8201 & n11305 ) | ( n11300 & n11305 ) ;
  assign n11307 = ( n8201 & ~n10939 ) | ( n8201 & n11252 ) | ( ~n10939 & n11252 ) ;
  assign n11308 = n8201 & ~n10939 ;
  assign n11309 = ( n10944 & n11307 ) | ( n10944 & n11308 ) | ( n11307 & n11308 ) ;
  assign n11310 = ( ~n10944 & n11307 ) | ( ~n10944 & n11308 ) | ( n11307 & n11308 ) ;
  assign n11311 = ( n10944 & ~n11309 ) | ( n10944 & n11310 ) | ( ~n11309 & n11310 ) ;
  assign n11312 = ( ~n7897 & n11306 ) | ( ~n7897 & n11311 ) | ( n11306 & n11311 ) ;
  assign n11313 = ( n7897 & ~n10945 ) | ( n7897 & n11252 ) | ( ~n10945 & n11252 ) ;
  assign n11314 = n7897 & ~n10945 ;
  assign n11315 = ( n10950 & n11313 ) | ( n10950 & n11314 ) | ( n11313 & n11314 ) ;
  assign n11316 = ( ~n10950 & n11313 ) | ( ~n10950 & n11314 ) | ( n11313 & n11314 ) ;
  assign n11317 = ( n10950 & ~n11315 ) | ( n10950 & n11316 ) | ( ~n11315 & n11316 ) ;
  assign n11318 = ( ~n7594 & n11312 ) | ( ~n7594 & n11317 ) | ( n11312 & n11317 ) ;
  assign n11319 = ~n7594 & n10951 ;
  assign n11320 = ( ~n7594 & n10951 ) | ( ~n7594 & n11252 ) | ( n10951 & n11252 ) ;
  assign n11321 = ( n10956 & n11319 ) | ( n10956 & n11320 ) | ( n11319 & n11320 ) ;
  assign n11322 = ( ~n10956 & n11319 ) | ( ~n10956 & n11320 ) | ( n11319 & n11320 ) ;
  assign n11323 = ( n10956 & ~n11321 ) | ( n10956 & n11322 ) | ( ~n11321 & n11322 ) ;
  assign n11324 = ( ~n7296 & n11318 ) | ( ~n7296 & n11323 ) | ( n11318 & n11323 ) ;
  assign n11325 = ~n7296 & n10957 ;
  assign n11326 = ( ~n7296 & n10957 ) | ( ~n7296 & n11252 ) | ( n10957 & n11252 ) ;
  assign n11327 = ( n10962 & n11325 ) | ( n10962 & n11326 ) | ( n11325 & n11326 ) ;
  assign n11328 = ( ~n10962 & n11325 ) | ( ~n10962 & n11326 ) | ( n11325 & n11326 ) ;
  assign n11329 = ( n10962 & ~n11327 ) | ( n10962 & n11328 ) | ( ~n11327 & n11328 ) ;
  assign n11330 = ( ~n7006 & n11324 ) | ( ~n7006 & n11329 ) | ( n11324 & n11329 ) ;
  assign n11331 = ( n7006 & ~n10963 ) | ( n7006 & n11252 ) | ( ~n10963 & n11252 ) ;
  assign n11332 = n7006 & ~n10963 ;
  assign n11333 = ( n10968 & n11331 ) | ( n10968 & n11332 ) | ( n11331 & n11332 ) ;
  assign n11334 = ( ~n10968 & n11331 ) | ( ~n10968 & n11332 ) | ( n11331 & n11332 ) ;
  assign n11335 = ( n10968 & ~n11333 ) | ( n10968 & n11334 ) | ( ~n11333 & n11334 ) ;
  assign n11336 = ( ~n6723 & n11330 ) | ( ~n6723 & n11335 ) | ( n11330 & n11335 ) ;
  assign n11337 = n6723 & ~n10969 ;
  assign n11338 = ( n6723 & ~n10969 ) | ( n6723 & n11252 ) | ( ~n10969 & n11252 ) ;
  assign n11339 = ( ~n10974 & n11337 ) | ( ~n10974 & n11338 ) | ( n11337 & n11338 ) ;
  assign n11340 = ( n10974 & n11337 ) | ( n10974 & n11338 ) | ( n11337 & n11338 ) ;
  assign n11341 = ( n10974 & n11339 ) | ( n10974 & ~n11340 ) | ( n11339 & ~n11340 ) ;
  assign n11342 = ( ~n6442 & n11336 ) | ( ~n6442 & n11341 ) | ( n11336 & n11341 ) ;
  assign n11343 = ( n6442 & ~n10975 ) | ( n6442 & n11252 ) | ( ~n10975 & n11252 ) ;
  assign n11344 = n6442 & ~n10975 ;
  assign n11345 = ( n10980 & n11343 ) | ( n10980 & n11344 ) | ( n11343 & n11344 ) ;
  assign n11346 = ( ~n10980 & n11343 ) | ( ~n10980 & n11344 ) | ( n11343 & n11344 ) ;
  assign n11347 = ( n10980 & ~n11345 ) | ( n10980 & n11346 ) | ( ~n11345 & n11346 ) ;
  assign n11348 = ( ~n6172 & n11342 ) | ( ~n6172 & n11347 ) | ( n11342 & n11347 ) ;
  assign n11349 = ~n6172 & n10981 ;
  assign n11350 = ( ~n6172 & n10981 ) | ( ~n6172 & n11252 ) | ( n10981 & n11252 ) ;
  assign n11351 = ( n10986 & n11349 ) | ( n10986 & n11350 ) | ( n11349 & n11350 ) ;
  assign n11352 = ( ~n10986 & n11349 ) | ( ~n10986 & n11350 ) | ( n11349 & n11350 ) ;
  assign n11353 = ( n10986 & ~n11351 ) | ( n10986 & n11352 ) | ( ~n11351 & n11352 ) ;
  assign n11354 = ( ~n5905 & n11348 ) | ( ~n5905 & n11353 ) | ( n11348 & n11353 ) ;
  assign n11355 = ( n5905 & ~n10987 ) | ( n5905 & n11252 ) | ( ~n10987 & n11252 ) ;
  assign n11356 = n5905 & ~n10987 ;
  assign n11357 = ( n10992 & n11355 ) | ( n10992 & n11356 ) | ( n11355 & n11356 ) ;
  assign n11358 = ( ~n10992 & n11355 ) | ( ~n10992 & n11356 ) | ( n11355 & n11356 ) ;
  assign n11359 = ( n10992 & ~n11357 ) | ( n10992 & n11358 ) | ( ~n11357 & n11358 ) ;
  assign n11360 = ( ~n5642 & n11354 ) | ( ~n5642 & n11359 ) | ( n11354 & n11359 ) ;
  assign n11361 = ( n5642 & ~n10993 ) | ( n5642 & n11252 ) | ( ~n10993 & n11252 ) ;
  assign n11362 = n5642 & ~n10993 ;
  assign n11363 = ( n10998 & n11361 ) | ( n10998 & n11362 ) | ( n11361 & n11362 ) ;
  assign n11364 = ( ~n10998 & n11361 ) | ( ~n10998 & n11362 ) | ( n11361 & n11362 ) ;
  assign n11365 = ( n10998 & ~n11363 ) | ( n10998 & n11364 ) | ( ~n11363 & n11364 ) ;
  assign n11366 = ( ~n5386 & n11360 ) | ( ~n5386 & n11365 ) | ( n11360 & n11365 ) ;
  assign n11367 = ( n5386 & ~n10999 ) | ( n5386 & n11252 ) | ( ~n10999 & n11252 ) ;
  assign n11368 = n5386 & ~n10999 ;
  assign n11369 = ( n11004 & n11367 ) | ( n11004 & n11368 ) | ( n11367 & n11368 ) ;
  assign n11370 = ( ~n11004 & n11367 ) | ( ~n11004 & n11368 ) | ( n11367 & n11368 ) ;
  assign n11371 = ( n11004 & ~n11369 ) | ( n11004 & n11370 ) | ( ~n11369 & n11370 ) ;
  assign n11372 = ( ~n5139 & n11366 ) | ( ~n5139 & n11371 ) | ( n11366 & n11371 ) ;
  assign n11373 = ( n5139 & ~n11005 ) | ( n5139 & n11252 ) | ( ~n11005 & n11252 ) ;
  assign n11374 = n5139 & ~n11005 ;
  assign n11375 = ( n11010 & n11373 ) | ( n11010 & n11374 ) | ( n11373 & n11374 ) ;
  assign n11376 = ( ~n11010 & n11373 ) | ( ~n11010 & n11374 ) | ( n11373 & n11374 ) ;
  assign n11377 = ( n11010 & ~n11375 ) | ( n11010 & n11376 ) | ( ~n11375 & n11376 ) ;
  assign n11378 = ( ~n4898 & n11372 ) | ( ~n4898 & n11377 ) | ( n11372 & n11377 ) ;
  assign n11379 = ( n4898 & ~n11011 ) | ( n4898 & n11252 ) | ( ~n11011 & n11252 ) ;
  assign n11380 = n4898 & ~n11011 ;
  assign n11381 = ( n11016 & n11379 ) | ( n11016 & n11380 ) | ( n11379 & n11380 ) ;
  assign n11382 = ( ~n11016 & n11379 ) | ( ~n11016 & n11380 ) | ( n11379 & n11380 ) ;
  assign n11383 = ( n11016 & ~n11381 ) | ( n11016 & n11382 ) | ( ~n11381 & n11382 ) ;
  assign n11384 = ( ~n4661 & n11378 ) | ( ~n4661 & n11383 ) | ( n11378 & n11383 ) ;
  assign n11385 = ~n4661 & n11017 ;
  assign n11386 = ( ~n4661 & n11017 ) | ( ~n4661 & n11252 ) | ( n11017 & n11252 ) ;
  assign n11387 = ( n11022 & n11385 ) | ( n11022 & n11386 ) | ( n11385 & n11386 ) ;
  assign n11388 = ( ~n11022 & n11385 ) | ( ~n11022 & n11386 ) | ( n11385 & n11386 ) ;
  assign n11389 = ( n11022 & ~n11387 ) | ( n11022 & n11388 ) | ( ~n11387 & n11388 ) ;
  assign n11390 = ( ~n4432 & n11384 ) | ( ~n4432 & n11389 ) | ( n11384 & n11389 ) ;
  assign n11391 = ( n4432 & ~n11023 ) | ( n4432 & n11252 ) | ( ~n11023 & n11252 ) ;
  assign n11392 = n4432 & ~n11023 ;
  assign n11393 = ( n11028 & n11391 ) | ( n11028 & n11392 ) | ( n11391 & n11392 ) ;
  assign n11394 = ( ~n11028 & n11391 ) | ( ~n11028 & n11392 ) | ( n11391 & n11392 ) ;
  assign n11395 = ( n11028 & ~n11393 ) | ( n11028 & n11394 ) | ( ~n11393 & n11394 ) ;
  assign n11396 = ( ~n4203 & n11390 ) | ( ~n4203 & n11395 ) | ( n11390 & n11395 ) ;
  assign n11397 = ~n4203 & n11029 ;
  assign n11398 = ( ~n4203 & n11029 ) | ( ~n4203 & n11252 ) | ( n11029 & n11252 ) ;
  assign n11399 = ( ~n11034 & n11397 ) | ( ~n11034 & n11398 ) | ( n11397 & n11398 ) ;
  assign n11400 = ( n11034 & n11397 ) | ( n11034 & n11398 ) | ( n11397 & n11398 ) ;
  assign n11401 = ( n11034 & n11399 ) | ( n11034 & ~n11400 ) | ( n11399 & ~n11400 ) ;
  assign n11402 = ( ~n3985 & n11396 ) | ( ~n3985 & n11401 ) | ( n11396 & n11401 ) ;
  assign n11403 = ~n3985 & n11035 ;
  assign n11404 = ( ~n3985 & n11035 ) | ( ~n3985 & n11252 ) | ( n11035 & n11252 ) ;
  assign n11405 = ( n11040 & n11403 ) | ( n11040 & n11404 ) | ( n11403 & n11404 ) ;
  assign n11406 = ( ~n11040 & n11403 ) | ( ~n11040 & n11404 ) | ( n11403 & n11404 ) ;
  assign n11407 = ( n11040 & ~n11405 ) | ( n11040 & n11406 ) | ( ~n11405 & n11406 ) ;
  assign n11408 = ( ~n3772 & n11402 ) | ( ~n3772 & n11407 ) | ( n11402 & n11407 ) ;
  assign n11409 = ~n3772 & n11041 ;
  assign n11410 = ( ~n3772 & n11041 ) | ( ~n3772 & n11252 ) | ( n11041 & n11252 ) ;
  assign n11411 = ( n11046 & n11409 ) | ( n11046 & n11410 ) | ( n11409 & n11410 ) ;
  assign n11412 = ( ~n11046 & n11409 ) | ( ~n11046 & n11410 ) | ( n11409 & n11410 ) ;
  assign n11413 = ( n11046 & ~n11411 ) | ( n11046 & n11412 ) | ( ~n11411 & n11412 ) ;
  assign n11414 = ( ~n3567 & n11408 ) | ( ~n3567 & n11413 ) | ( n11408 & n11413 ) ;
  assign n11415 = ~n3567 & n11047 ;
  assign n11416 = ( ~n3567 & n11047 ) | ( ~n3567 & n11252 ) | ( n11047 & n11252 ) ;
  assign n11417 = ( n11052 & n11415 ) | ( n11052 & n11416 ) | ( n11415 & n11416 ) ;
  assign n11418 = ( ~n11052 & n11415 ) | ( ~n11052 & n11416 ) | ( n11415 & n11416 ) ;
  assign n11419 = ( n11052 & ~n11417 ) | ( n11052 & n11418 ) | ( ~n11417 & n11418 ) ;
  assign n11420 = ( ~n3362 & n11414 ) | ( ~n3362 & n11419 ) | ( n11414 & n11419 ) ;
  assign n11421 = ~n3362 & n11053 ;
  assign n11422 = ( ~n3362 & n11053 ) | ( ~n3362 & n11252 ) | ( n11053 & n11252 ) ;
  assign n11423 = ( n11058 & n11421 ) | ( n11058 & n11422 ) | ( n11421 & n11422 ) ;
  assign n11424 = ( ~n11058 & n11421 ) | ( ~n11058 & n11422 ) | ( n11421 & n11422 ) ;
  assign n11425 = ( n11058 & ~n11423 ) | ( n11058 & n11424 ) | ( ~n11423 & n11424 ) ;
  assign n11426 = ( ~n3169 & n11420 ) | ( ~n3169 & n11425 ) | ( n11420 & n11425 ) ;
  assign n11427 = ( n3169 & ~n11059 ) | ( n3169 & n11252 ) | ( ~n11059 & n11252 ) ;
  assign n11428 = n3169 & ~n11059 ;
  assign n11429 = ( n11064 & n11427 ) | ( n11064 & n11428 ) | ( n11427 & n11428 ) ;
  assign n11430 = ( ~n11064 & n11427 ) | ( ~n11064 & n11428 ) | ( n11427 & n11428 ) ;
  assign n11431 = ( n11064 & ~n11429 ) | ( n11064 & n11430 ) | ( ~n11429 & n11430 ) ;
  assign n11432 = ( ~n2979 & n11426 ) | ( ~n2979 & n11431 ) | ( n11426 & n11431 ) ;
  assign n11433 = ~n2979 & n11065 ;
  assign n11434 = ( ~n2979 & n11065 ) | ( ~n2979 & n11252 ) | ( n11065 & n11252 ) ;
  assign n11435 = ( n11070 & n11433 ) | ( n11070 & n11434 ) | ( n11433 & n11434 ) ;
  assign n11436 = ( ~n11070 & n11433 ) | ( ~n11070 & n11434 ) | ( n11433 & n11434 ) ;
  assign n11437 = ( n11070 & ~n11435 ) | ( n11070 & n11436 ) | ( ~n11435 & n11436 ) ;
  assign n11438 = ( ~n2791 & n11432 ) | ( ~n2791 & n11437 ) | ( n11432 & n11437 ) ;
  assign n11439 = ( n2791 & ~n11071 ) | ( n2791 & n11252 ) | ( ~n11071 & n11252 ) ;
  assign n11440 = n2791 & ~n11071 ;
  assign n11441 = ( n11076 & n11439 ) | ( n11076 & n11440 ) | ( n11439 & n11440 ) ;
  assign n11442 = ( ~n11076 & n11439 ) | ( ~n11076 & n11440 ) | ( n11439 & n11440 ) ;
  assign n11443 = ( n11076 & ~n11441 ) | ( n11076 & n11442 ) | ( ~n11441 & n11442 ) ;
  assign n11444 = ( ~n2615 & n11438 ) | ( ~n2615 & n11443 ) | ( n11438 & n11443 ) ;
  assign n11445 = ( n2615 & ~n11077 ) | ( n2615 & n11252 ) | ( ~n11077 & n11252 ) ;
  assign n11446 = n2615 & ~n11077 ;
  assign n11447 = ( n11082 & n11445 ) | ( n11082 & n11446 ) | ( n11445 & n11446 ) ;
  assign n11448 = ( ~n11082 & n11445 ) | ( ~n11082 & n11446 ) | ( n11445 & n11446 ) ;
  assign n11449 = ( n11082 & ~n11447 ) | ( n11082 & n11448 ) | ( ~n11447 & n11448 ) ;
  assign n11450 = ( ~n2443 & n11444 ) | ( ~n2443 & n11449 ) | ( n11444 & n11449 ) ;
  assign n11451 = ~n2443 & n11083 ;
  assign n11452 = ( ~n2443 & n11083 ) | ( ~n2443 & n11252 ) | ( n11083 & n11252 ) ;
  assign n11453 = ( n11088 & n11451 ) | ( n11088 & n11452 ) | ( n11451 & n11452 ) ;
  assign n11454 = ( ~n11088 & n11451 ) | ( ~n11088 & n11452 ) | ( n11451 & n11452 ) ;
  assign n11455 = ( n11088 & ~n11453 ) | ( n11088 & n11454 ) | ( ~n11453 & n11454 ) ;
  assign n11456 = ( ~n2277 & n11450 ) | ( ~n2277 & n11455 ) | ( n11450 & n11455 ) ;
  assign n11457 = ( n2277 & ~n11089 ) | ( n2277 & n11252 ) | ( ~n11089 & n11252 ) ;
  assign n11458 = n2277 & ~n11089 ;
  assign n11459 = ( n11094 & n11457 ) | ( n11094 & n11458 ) | ( n11457 & n11458 ) ;
  assign n11460 = ( ~n11094 & n11457 ) | ( ~n11094 & n11458 ) | ( n11457 & n11458 ) ;
  assign n11461 = ( n11094 & ~n11459 ) | ( n11094 & n11460 ) | ( ~n11459 & n11460 ) ;
  assign n11462 = ( ~n2111 & n11456 ) | ( ~n2111 & n11461 ) | ( n11456 & n11461 ) ;
  assign n11463 = ( n2111 & ~n11095 ) | ( n2111 & n11252 ) | ( ~n11095 & n11252 ) ;
  assign n11464 = n2111 & ~n11095 ;
  assign n11465 = ( n11100 & n11463 ) | ( n11100 & n11464 ) | ( n11463 & n11464 ) ;
  assign n11466 = ( ~n11100 & n11463 ) | ( ~n11100 & n11464 ) | ( n11463 & n11464 ) ;
  assign n11467 = ( n11100 & ~n11465 ) | ( n11100 & n11466 ) | ( ~n11465 & n11466 ) ;
  assign n11468 = ( ~n1949 & n11462 ) | ( ~n1949 & n11467 ) | ( n11462 & n11467 ) ;
  assign n11469 = ~n1949 & n11101 ;
  assign n11470 = ( ~n1949 & n11101 ) | ( ~n1949 & n11252 ) | ( n11101 & n11252 ) ;
  assign n11471 = ( ~n11106 & n11469 ) | ( ~n11106 & n11470 ) | ( n11469 & n11470 ) ;
  assign n11472 = ( n11106 & n11469 ) | ( n11106 & n11470 ) | ( n11469 & n11470 ) ;
  assign n11473 = ( n11106 & n11471 ) | ( n11106 & ~n11472 ) | ( n11471 & ~n11472 ) ;
  assign n11474 = ( ~n1802 & n11468 ) | ( ~n1802 & n11473 ) | ( n11468 & n11473 ) ;
  assign n11475 = ( n1802 & ~n11107 ) | ( n1802 & n11252 ) | ( ~n11107 & n11252 ) ;
  assign n11476 = n1802 & ~n11107 ;
  assign n11477 = ( n11112 & n11475 ) | ( n11112 & n11476 ) | ( n11475 & n11476 ) ;
  assign n11478 = ( ~n11112 & n11475 ) | ( ~n11112 & n11476 ) | ( n11475 & n11476 ) ;
  assign n11479 = ( n11112 & ~n11477 ) | ( n11112 & n11478 ) | ( ~n11477 & n11478 ) ;
  assign n11480 = ( ~n1661 & n11474 ) | ( ~n1661 & n11479 ) | ( n11474 & n11479 ) ;
  assign n11481 = ( n1661 & ~n11113 ) | ( n1661 & n11252 ) | ( ~n11113 & n11252 ) ;
  assign n11482 = n1661 & ~n11113 ;
  assign n11483 = ( n11118 & n11481 ) | ( n11118 & n11482 ) | ( n11481 & n11482 ) ;
  assign n11484 = ( ~n11118 & n11481 ) | ( ~n11118 & n11482 ) | ( n11481 & n11482 ) ;
  assign n11485 = ( n11118 & ~n11483 ) | ( n11118 & n11484 ) | ( ~n11483 & n11484 ) ;
  assign n11486 = ( ~n1523 & n11480 ) | ( ~n1523 & n11485 ) | ( n11480 & n11485 ) ;
  assign n11487 = ( n1523 & ~n11119 ) | ( n1523 & n11252 ) | ( ~n11119 & n11252 ) ;
  assign n11488 = n1523 & ~n11119 ;
  assign n11489 = ( n11124 & n11487 ) | ( n11124 & n11488 ) | ( n11487 & n11488 ) ;
  assign n11490 = ( ~n11124 & n11487 ) | ( ~n11124 & n11488 ) | ( n11487 & n11488 ) ;
  assign n11491 = ( n11124 & ~n11489 ) | ( n11124 & n11490 ) | ( ~n11489 & n11490 ) ;
  assign n11492 = ( ~n1393 & n11486 ) | ( ~n1393 & n11491 ) | ( n11486 & n11491 ) ;
  assign n11493 = ( n1393 & ~n11125 ) | ( n1393 & n11252 ) | ( ~n11125 & n11252 ) ;
  assign n11494 = n1393 & ~n11125 ;
  assign n11495 = ( n11130 & n11493 ) | ( n11130 & n11494 ) | ( n11493 & n11494 ) ;
  assign n11496 = ( ~n11130 & n11493 ) | ( ~n11130 & n11494 ) | ( n11493 & n11494 ) ;
  assign n11497 = ( n11130 & ~n11495 ) | ( n11130 & n11496 ) | ( ~n11495 & n11496 ) ;
  assign n11498 = ( ~n1266 & n11492 ) | ( ~n1266 & n11497 ) | ( n11492 & n11497 ) ;
  assign n11499 = ( n1266 & ~n11131 ) | ( n1266 & n11252 ) | ( ~n11131 & n11252 ) ;
  assign n11500 = n1266 & ~n11131 ;
  assign n11501 = ( n11136 & n11499 ) | ( n11136 & n11500 ) | ( n11499 & n11500 ) ;
  assign n11502 = ( ~n11136 & n11499 ) | ( ~n11136 & n11500 ) | ( n11499 & n11500 ) ;
  assign n11503 = ( n11136 & ~n11501 ) | ( n11136 & n11502 ) | ( ~n11501 & n11502 ) ;
  assign n11504 = ( ~n1150 & n11498 ) | ( ~n1150 & n11503 ) | ( n11498 & n11503 ) ;
  assign n11505 = ( n1150 & ~n11137 ) | ( n1150 & n11252 ) | ( ~n11137 & n11252 ) ;
  assign n11506 = n1150 & ~n11137 ;
  assign n11507 = ( n11142 & n11505 ) | ( n11142 & n11506 ) | ( n11505 & n11506 ) ;
  assign n11508 = ( ~n11142 & n11505 ) | ( ~n11142 & n11506 ) | ( n11505 & n11506 ) ;
  assign n11509 = ( n11142 & ~n11507 ) | ( n11142 & n11508 ) | ( ~n11507 & n11508 ) ;
  assign n11510 = ( ~n1038 & n11504 ) | ( ~n1038 & n11509 ) | ( n11504 & n11509 ) ;
  assign n11511 = ( n1038 & ~n11143 ) | ( n1038 & n11252 ) | ( ~n11143 & n11252 ) ;
  assign n11512 = n1038 & ~n11143 ;
  assign n11513 = ( n11148 & n11511 ) | ( n11148 & n11512 ) | ( n11511 & n11512 ) ;
  assign n11514 = ( ~n11148 & n11511 ) | ( ~n11148 & n11512 ) | ( n11511 & n11512 ) ;
  assign n11515 = ( n11148 & ~n11513 ) | ( n11148 & n11514 ) | ( ~n11513 & n11514 ) ;
  assign n11516 = ( ~n933 & n11510 ) | ( ~n933 & n11515 ) | ( n11510 & n11515 ) ;
  assign n11517 = ( n933 & ~n11149 ) | ( n933 & n11252 ) | ( ~n11149 & n11252 ) ;
  assign n11518 = n933 & ~n11149 ;
  assign n11519 = ( n11154 & n11517 ) | ( n11154 & n11518 ) | ( n11517 & n11518 ) ;
  assign n11520 = ( ~n11154 & n11517 ) | ( ~n11154 & n11518 ) | ( n11517 & n11518 ) ;
  assign n11521 = ( n11154 & ~n11519 ) | ( n11154 & n11520 ) | ( ~n11519 & n11520 ) ;
  assign n11522 = ( ~n839 & n11516 ) | ( ~n839 & n11521 ) | ( n11516 & n11521 ) ;
  assign n11523 = ~n839 & n11155 ;
  assign n11524 = ( ~n839 & n11155 ) | ( ~n839 & n11252 ) | ( n11155 & n11252 ) ;
  assign n11525 = ( n11160 & n11523 ) | ( n11160 & n11524 ) | ( n11523 & n11524 ) ;
  assign n11526 = ( ~n11160 & n11523 ) | ( ~n11160 & n11524 ) | ( n11523 & n11524 ) ;
  assign n11527 = ( n11160 & ~n11525 ) | ( n11160 & n11526 ) | ( ~n11525 & n11526 ) ;
  assign n11528 = ( ~n746 & n11522 ) | ( ~n746 & n11527 ) | ( n11522 & n11527 ) ;
  assign n11529 = ~n746 & n11161 ;
  assign n11530 = ( ~n746 & n11161 ) | ( ~n746 & n11252 ) | ( n11161 & n11252 ) ;
  assign n11531 = ( n11166 & n11529 ) | ( n11166 & n11530 ) | ( n11529 & n11530 ) ;
  assign n11532 = ( ~n11166 & n11529 ) | ( ~n11166 & n11530 ) | ( n11529 & n11530 ) ;
  assign n11533 = ( n11166 & ~n11531 ) | ( n11166 & n11532 ) | ( ~n11531 & n11532 ) ;
  assign n11534 = ( ~n664 & n11528 ) | ( ~n664 & n11533 ) | ( n11528 & n11533 ) ;
  assign n11535 = ~n664 & n11167 ;
  assign n11536 = ( ~n664 & n11167 ) | ( ~n664 & n11252 ) | ( n11167 & n11252 ) ;
  assign n11537 = ( ~n11172 & n11535 ) | ( ~n11172 & n11536 ) | ( n11535 & n11536 ) ;
  assign n11538 = ( n11172 & n11535 ) | ( n11172 & n11536 ) | ( n11535 & n11536 ) ;
  assign n11539 = ( n11172 & n11537 ) | ( n11172 & ~n11538 ) | ( n11537 & ~n11538 ) ;
  assign n11540 = ( ~n588 & n11534 ) | ( ~n588 & n11539 ) | ( n11534 & n11539 ) ;
  assign n11541 = ( n588 & ~n11173 ) | ( n588 & n11252 ) | ( ~n11173 & n11252 ) ;
  assign n11542 = n588 & ~n11173 ;
  assign n11543 = ( n11178 & n11541 ) | ( n11178 & n11542 ) | ( n11541 & n11542 ) ;
  assign n11544 = ( ~n11178 & n11541 ) | ( ~n11178 & n11542 ) | ( n11541 & n11542 ) ;
  assign n11545 = ( n11178 & ~n11543 ) | ( n11178 & n11544 ) | ( ~n11543 & n11544 ) ;
  assign n11546 = ( ~n518 & n11540 ) | ( ~n518 & n11545 ) | ( n11540 & n11545 ) ;
  assign n11547 = ( n518 & ~n11179 ) | ( n518 & n11252 ) | ( ~n11179 & n11252 ) ;
  assign n11548 = n518 & ~n11179 ;
  assign n11549 = ( n11184 & n11547 ) | ( n11184 & n11548 ) | ( n11547 & n11548 ) ;
  assign n11550 = ( ~n11184 & n11547 ) | ( ~n11184 & n11548 ) | ( n11547 & n11548 ) ;
  assign n11551 = ( n11184 & ~n11549 ) | ( n11184 & n11550 ) | ( ~n11549 & n11550 ) ;
  assign n11552 = ( ~n454 & n11546 ) | ( ~n454 & n11551 ) | ( n11546 & n11551 ) ;
  assign n11553 = n454 & ~n11185 ;
  assign n11554 = ( n454 & ~n11185 ) | ( n454 & n11252 ) | ( ~n11185 & n11252 ) ;
  assign n11555 = ( n11190 & n11553 ) | ( n11190 & n11554 ) | ( n11553 & n11554 ) ;
  assign n11556 = ( ~n11190 & n11553 ) | ( ~n11190 & n11554 ) | ( n11553 & n11554 ) ;
  assign n11557 = ( n11190 & ~n11555 ) | ( n11190 & n11556 ) | ( ~n11555 & n11556 ) ;
  assign n11558 = ( ~n396 & n11552 ) | ( ~n396 & n11557 ) | ( n11552 & n11557 ) ;
  assign n11559 = ( n396 & ~n11191 ) | ( n396 & n11252 ) | ( ~n11191 & n11252 ) ;
  assign n11560 = n396 & ~n11191 ;
  assign n11561 = ( n11196 & n11559 ) | ( n11196 & n11560 ) | ( n11559 & n11560 ) ;
  assign n11562 = ( ~n11196 & n11559 ) | ( ~n11196 & n11560 ) | ( n11559 & n11560 ) ;
  assign n11563 = ( n11196 & ~n11561 ) | ( n11196 & n11562 ) | ( ~n11561 & n11562 ) ;
  assign n11564 = ( ~n344 & n11558 ) | ( ~n344 & n11563 ) | ( n11558 & n11563 ) ;
  assign n11565 = ( n344 & ~n11197 ) | ( n344 & n11252 ) | ( ~n11197 & n11252 ) ;
  assign n11566 = n344 & ~n11197 ;
  assign n11567 = ( n11202 & n11565 ) | ( n11202 & n11566 ) | ( n11565 & n11566 ) ;
  assign n11568 = ( ~n11202 & n11565 ) | ( ~n11202 & n11566 ) | ( n11565 & n11566 ) ;
  assign n11569 = ( n11202 & ~n11567 ) | ( n11202 & n11568 ) | ( ~n11567 & n11568 ) ;
  assign n11570 = ( ~n298 & n11564 ) | ( ~n298 & n11569 ) | ( n11564 & n11569 ) ;
  assign n11571 = ( n298 & ~n11203 ) | ( n298 & n11252 ) | ( ~n11203 & n11252 ) ;
  assign n11572 = n298 & ~n11203 ;
  assign n11573 = ( n11208 & n11571 ) | ( n11208 & n11572 ) | ( n11571 & n11572 ) ;
  assign n11574 = ( ~n11208 & n11571 ) | ( ~n11208 & n11572 ) | ( n11571 & n11572 ) ;
  assign n11575 = ( n11208 & ~n11573 ) | ( n11208 & n11574 ) | ( ~n11573 & n11574 ) ;
  assign n11576 = ( ~n258 & n11570 ) | ( ~n258 & n11575 ) | ( n11570 & n11575 ) ;
  assign n11577 = ~n258 & n11209 ;
  assign n11578 = ( ~n258 & n11209 ) | ( ~n258 & n11252 ) | ( n11209 & n11252 ) ;
  assign n11579 = ( ~n11214 & n11577 ) | ( ~n11214 & n11578 ) | ( n11577 & n11578 ) ;
  assign n11580 = ( n11214 & n11577 ) | ( n11214 & n11578 ) | ( n11577 & n11578 ) ;
  assign n11581 = ( n11214 & n11579 ) | ( n11214 & ~n11580 ) | ( n11579 & ~n11580 ) ;
  assign n11582 = ( ~n225 & n11576 ) | ( ~n225 & n11581 ) | ( n11576 & n11581 ) ;
  assign n11583 = ( n225 & ~n11215 ) | ( n225 & n11252 ) | ( ~n11215 & n11252 ) ;
  assign n11584 = n225 & ~n11215 ;
  assign n11585 = ( n11220 & n11583 ) | ( n11220 & n11584 ) | ( n11583 & n11584 ) ;
  assign n11586 = ( ~n11220 & n11583 ) | ( ~n11220 & n11584 ) | ( n11583 & n11584 ) ;
  assign n11587 = ( n11220 & ~n11585 ) | ( n11220 & n11586 ) | ( ~n11585 & n11586 ) ;
  assign n11588 = ( ~n197 & n11582 ) | ( ~n197 & n11587 ) | ( n11582 & n11587 ) ;
  assign n11589 = ~n197 & n11221 ;
  assign n11590 = ( ~n197 & n11221 ) | ( ~n197 & n11252 ) | ( n11221 & n11252 ) ;
  assign n11591 = ( ~n11226 & n11589 ) | ( ~n11226 & n11590 ) | ( n11589 & n11590 ) ;
  assign n11592 = ( n11226 & n11589 ) | ( n11226 & n11590 ) | ( n11589 & n11590 ) ;
  assign n11593 = ( n11226 & n11591 ) | ( n11226 & ~n11592 ) | ( n11591 & ~n11592 ) ;
  assign n11594 = ( ~n170 & n11588 ) | ( ~n170 & n11593 ) | ( n11588 & n11593 ) ;
  assign n11595 = ( n170 & ~n11227 ) | ( n170 & n11252 ) | ( ~n11227 & n11252 ) ;
  assign n11596 = n170 & ~n11227 ;
  assign n11597 = ( n11232 & n11595 ) | ( n11232 & n11596 ) | ( n11595 & n11596 ) ;
  assign n11598 = ( ~n11232 & n11595 ) | ( ~n11232 & n11596 ) | ( n11595 & n11596 ) ;
  assign n11599 = ( n11232 & ~n11597 ) | ( n11232 & n11598 ) | ( ~n11597 & n11598 ) ;
  assign n11600 = ( ~n142 & n11594 ) | ( ~n142 & n11599 ) | ( n11594 & n11599 ) ;
  assign n11601 = ~n11245 & n11250 ;
  assign n11602 = n10892 & n11245 ;
  assign n11603 = ( ~n11251 & n11601 ) | ( ~n11251 & n11602 ) | ( n11601 & n11602 ) ;
  assign n11604 = ( n142 & ~n11233 ) | ( n142 & n11252 ) | ( ~n11233 & n11252 ) ;
  assign n11605 = n142 & ~n11233 ;
  assign n11606 = ( n11238 & n11604 ) | ( n11238 & n11605 ) | ( n11604 & n11605 ) ;
  assign n11607 = ( ~n11238 & n11604 ) | ( ~n11238 & n11605 ) | ( n11604 & n11605 ) ;
  assign n11608 = ( n11238 & ~n11606 ) | ( n11238 & n11607 ) | ( ~n11606 & n11607 ) ;
  assign n11609 = ( ~n132 & n11600 ) | ( ~n132 & n11608 ) | ( n11600 & n11608 ) ;
  assign n11610 = ( n132 & ~n11239 ) | ( n132 & n11252 ) | ( ~n11239 & n11252 ) ;
  assign n11611 = n132 & ~n11239 ;
  assign n11612 = ( n11244 & n11610 ) | ( n11244 & n11611 ) | ( n11610 & n11611 ) ;
  assign n11613 = ( ~n11244 & n11610 ) | ( ~n11244 & n11611 ) | ( n11610 & n11611 ) ;
  assign n11614 = ( n11244 & ~n11612 ) | ( n11244 & n11613 ) | ( ~n11612 & n11613 ) ;
  assign n11615 = ( n11245 & ~n11250 ) | ( n11245 & n11609 ) | ( ~n11250 & n11609 ) ;
  assign n11616 = ( n10897 & n11245 ) | ( n10897 & ~n11601 ) | ( n11245 & ~n11601 ) ;
  assign n11617 = n11614 | n11616 ;
  assign n11618 = ( n11614 & ~n11615 ) | ( n11614 & n11617 ) | ( ~n11615 & n11617 ) ;
  assign n11619 = ( ~n131 & n11609 ) | ( ~n131 & n11618 ) | ( n11609 & n11618 ) ;
  assign n11620 = n11603 | n11619 ;
  assign n11621 = ( n132 & ~n11600 ) | ( n132 & n11620 ) | ( ~n11600 & n11620 ) ;
  assign n11622 = n132 & ~n11600 ;
  assign n11623 = ( n11608 & n11621 ) | ( n11608 & n11622 ) | ( n11621 & n11622 ) ;
  assign n11624 = ( n11608 & ~n11621 ) | ( n11608 & n11622 ) | ( ~n11621 & n11622 ) ;
  assign n11625 = ( n11621 & ~n11623 ) | ( n11621 & n11624 ) | ( ~n11623 & n11624 ) ;
  assign n11626 = ~n11258 & n11620 ;
  assign n11627 = n11252 & ~n11620 ;
  assign n11628 = ( x6 & n11626 ) | ( x6 & n11627 ) | ( n11626 & n11627 ) ;
  assign n11629 = ( ~x6 & n11626 ) | ( ~x6 & n11627 ) | ( n11626 & n11627 ) ;
  assign n11630 = ( x6 & ~n11628 ) | ( x6 & n11629 ) | ( ~n11628 & n11629 ) ;
  assign n11631 = x2 | x3 ;
  assign n11632 = x4 | n11631 ;
  assign n11633 = n11252 & ~n11632 ;
  assign n11634 = ~n11252 & n11632 ;
  assign n11635 = ( x5 & ~n11620 ) | ( x5 & n11634 ) | ( ~n11620 & n11634 ) ;
  assign n11636 = ( n11626 & ~n11633 ) | ( n11626 & n11635 ) | ( ~n11633 & n11635 ) ;
  assign n11637 = ( ~n10888 & n11630 ) | ( ~n10888 & n11636 ) | ( n11630 & n11636 ) ;
  assign n11638 = ~n10888 & n11252 ;
  assign n11639 = ( n11253 & n11620 ) | ( n11253 & n11638 ) | ( n11620 & n11638 ) ;
  assign n11640 = ( ~x7 & n11629 ) | ( ~x7 & n11639 ) | ( n11629 & n11639 ) ;
  assign n11641 = ( x7 & n11629 ) | ( x7 & n11639 ) | ( n11629 & n11639 ) ;
  assign n11642 = ( x7 & n11640 ) | ( x7 & ~n11641 ) | ( n11640 & ~n11641 ) ;
  assign n11643 = ( ~n10533 & n11637 ) | ( ~n10533 & n11642 ) | ( n11637 & n11642 ) ;
  assign n11644 = n10533 & ~n11263 ;
  assign n11645 = ( n10533 & ~n11263 ) | ( n10533 & n11620 ) | ( ~n11263 & n11620 ) ;
  assign n11646 = ( n11257 & n11644 ) | ( n11257 & n11645 ) | ( n11644 & n11645 ) ;
  assign n11647 = ( ~n11257 & n11644 ) | ( ~n11257 & n11645 ) | ( n11644 & n11645 ) ;
  assign n11648 = ( n11257 & ~n11646 ) | ( n11257 & n11647 ) | ( ~n11646 & n11647 ) ;
  assign n11649 = ( ~n10180 & n11643 ) | ( ~n10180 & n11648 ) | ( n11643 & n11648 ) ;
  assign n11650 = n10180 & ~n11264 ;
  assign n11651 = ( n10180 & ~n11264 ) | ( n10180 & n11620 ) | ( ~n11264 & n11620 ) ;
  assign n11652 = ( n11269 & n11650 ) | ( n11269 & n11651 ) | ( n11650 & n11651 ) ;
  assign n11653 = ( ~n11269 & n11650 ) | ( ~n11269 & n11651 ) | ( n11650 & n11651 ) ;
  assign n11654 = ( n11269 & ~n11652 ) | ( n11269 & n11653 ) | ( ~n11652 & n11653 ) ;
  assign n11655 = ( ~n9834 & n11649 ) | ( ~n9834 & n11654 ) | ( n11649 & n11654 ) ;
  assign n11656 = ( n9834 & ~n11270 ) | ( n9834 & n11620 ) | ( ~n11270 & n11620 ) ;
  assign n11657 = n9834 & ~n11270 ;
  assign n11658 = ( n11275 & n11656 ) | ( n11275 & n11657 ) | ( n11656 & n11657 ) ;
  assign n11659 = ( ~n11275 & n11656 ) | ( ~n11275 & n11657 ) | ( n11656 & n11657 ) ;
  assign n11660 = ( n11275 & ~n11658 ) | ( n11275 & n11659 ) | ( ~n11658 & n11659 ) ;
  assign n11661 = ( ~n9497 & n11655 ) | ( ~n9497 & n11660 ) | ( n11655 & n11660 ) ;
  assign n11662 = ~n9497 & n11276 ;
  assign n11663 = ( ~n9497 & n11276 ) | ( ~n9497 & n11620 ) | ( n11276 & n11620 ) ;
  assign n11664 = ( n11281 & n11662 ) | ( n11281 & n11663 ) | ( n11662 & n11663 ) ;
  assign n11665 = ( ~n11281 & n11662 ) | ( ~n11281 & n11663 ) | ( n11662 & n11663 ) ;
  assign n11666 = ( n11281 & ~n11664 ) | ( n11281 & n11665 ) | ( ~n11664 & n11665 ) ;
  assign n11667 = ( ~n9167 & n11661 ) | ( ~n9167 & n11666 ) | ( n11661 & n11666 ) ;
  assign n11668 = ( n9167 & ~n11282 ) | ( n9167 & n11620 ) | ( ~n11282 & n11620 ) ;
  assign n11669 = n9167 & ~n11282 ;
  assign n11670 = ( n11287 & n11668 ) | ( n11287 & n11669 ) | ( n11668 & n11669 ) ;
  assign n11671 = ( ~n11287 & n11668 ) | ( ~n11287 & n11669 ) | ( n11668 & n11669 ) ;
  assign n11672 = ( n11287 & ~n11670 ) | ( n11287 & n11671 ) | ( ~n11670 & n11671 ) ;
  assign n11673 = ( ~n8838 & n11667 ) | ( ~n8838 & n11672 ) | ( n11667 & n11672 ) ;
  assign n11674 = ~n8838 & n11288 ;
  assign n11675 = ( ~n8838 & n11288 ) | ( ~n8838 & n11620 ) | ( n11288 & n11620 ) ;
  assign n11676 = ( ~n11293 & n11674 ) | ( ~n11293 & n11675 ) | ( n11674 & n11675 ) ;
  assign n11677 = ( n11293 & n11674 ) | ( n11293 & n11675 ) | ( n11674 & n11675 ) ;
  assign n11678 = ( n11293 & n11676 ) | ( n11293 & ~n11677 ) | ( n11676 & ~n11677 ) ;
  assign n11679 = ( ~n8517 & n11673 ) | ( ~n8517 & n11678 ) | ( n11673 & n11678 ) ;
  assign n11680 = n8517 & ~n11294 ;
  assign n11681 = ( n8517 & ~n11294 ) | ( n8517 & n11620 ) | ( ~n11294 & n11620 ) ;
  assign n11682 = ( n11299 & n11680 ) | ( n11299 & n11681 ) | ( n11680 & n11681 ) ;
  assign n11683 = ( ~n11299 & n11680 ) | ( ~n11299 & n11681 ) | ( n11680 & n11681 ) ;
  assign n11684 = ( n11299 & ~n11682 ) | ( n11299 & n11683 ) | ( ~n11682 & n11683 ) ;
  assign n11685 = ( ~n8201 & n11679 ) | ( ~n8201 & n11684 ) | ( n11679 & n11684 ) ;
  assign n11686 = ( n8201 & ~n11300 ) | ( n8201 & n11620 ) | ( ~n11300 & n11620 ) ;
  assign n11687 = n8201 & ~n11300 ;
  assign n11688 = ( n11305 & n11686 ) | ( n11305 & n11687 ) | ( n11686 & n11687 ) ;
  assign n11689 = ( ~n11305 & n11686 ) | ( ~n11305 & n11687 ) | ( n11686 & n11687 ) ;
  assign n11690 = ( n11305 & ~n11688 ) | ( n11305 & n11689 ) | ( ~n11688 & n11689 ) ;
  assign n11691 = ( ~n7897 & n11685 ) | ( ~n7897 & n11690 ) | ( n11685 & n11690 ) ;
  assign n11692 = ~n7897 & n11306 ;
  assign n11693 = ( ~n7897 & n11306 ) | ( ~n7897 & n11620 ) | ( n11306 & n11620 ) ;
  assign n11694 = ( ~n11311 & n11692 ) | ( ~n11311 & n11693 ) | ( n11692 & n11693 ) ;
  assign n11695 = ( n11311 & n11692 ) | ( n11311 & n11693 ) | ( n11692 & n11693 ) ;
  assign n11696 = ( n11311 & n11694 ) | ( n11311 & ~n11695 ) | ( n11694 & ~n11695 ) ;
  assign n11697 = ( ~n7594 & n11691 ) | ( ~n7594 & n11696 ) | ( n11691 & n11696 ) ;
  assign n11698 = ~n7594 & n11312 ;
  assign n11699 = ( ~n7594 & n11312 ) | ( ~n7594 & n11620 ) | ( n11312 & n11620 ) ;
  assign n11700 = ( ~n11317 & n11698 ) | ( ~n11317 & n11699 ) | ( n11698 & n11699 ) ;
  assign n11701 = ( n11317 & n11698 ) | ( n11317 & n11699 ) | ( n11698 & n11699 ) ;
  assign n11702 = ( n11317 & n11700 ) | ( n11317 & ~n11701 ) | ( n11700 & ~n11701 ) ;
  assign n11703 = ( ~n7296 & n11697 ) | ( ~n7296 & n11702 ) | ( n11697 & n11702 ) ;
  assign n11704 = ~n7296 & n11318 ;
  assign n11705 = ( ~n7296 & n11318 ) | ( ~n7296 & n11620 ) | ( n11318 & n11620 ) ;
  assign n11706 = ( n11323 & n11704 ) | ( n11323 & n11705 ) | ( n11704 & n11705 ) ;
  assign n11707 = ( ~n11323 & n11704 ) | ( ~n11323 & n11705 ) | ( n11704 & n11705 ) ;
  assign n11708 = ( n11323 & ~n11706 ) | ( n11323 & n11707 ) | ( ~n11706 & n11707 ) ;
  assign n11709 = ( ~n7006 & n11703 ) | ( ~n7006 & n11708 ) | ( n11703 & n11708 ) ;
  assign n11710 = ( n7006 & ~n11324 ) | ( n7006 & n11620 ) | ( ~n11324 & n11620 ) ;
  assign n11711 = n7006 & ~n11324 ;
  assign n11712 = ( n11329 & n11710 ) | ( n11329 & n11711 ) | ( n11710 & n11711 ) ;
  assign n11713 = ( ~n11329 & n11710 ) | ( ~n11329 & n11711 ) | ( n11710 & n11711 ) ;
  assign n11714 = ( n11329 & ~n11712 ) | ( n11329 & n11713 ) | ( ~n11712 & n11713 ) ;
  assign n11715 = ( ~n6723 & n11709 ) | ( ~n6723 & n11714 ) | ( n11709 & n11714 ) ;
  assign n11716 = ( n6723 & ~n11330 ) | ( n6723 & n11620 ) | ( ~n11330 & n11620 ) ;
  assign n11717 = n6723 & ~n11330 ;
  assign n11718 = ( n11335 & n11716 ) | ( n11335 & n11717 ) | ( n11716 & n11717 ) ;
  assign n11719 = ( ~n11335 & n11716 ) | ( ~n11335 & n11717 ) | ( n11716 & n11717 ) ;
  assign n11720 = ( n11335 & ~n11718 ) | ( n11335 & n11719 ) | ( ~n11718 & n11719 ) ;
  assign n11721 = ( ~n6442 & n11715 ) | ( ~n6442 & n11720 ) | ( n11715 & n11720 ) ;
  assign n11722 = ( n6442 & ~n11336 ) | ( n6442 & n11620 ) | ( ~n11336 & n11620 ) ;
  assign n11723 = n6442 & ~n11336 ;
  assign n11724 = ( n11341 & n11722 ) | ( n11341 & n11723 ) | ( n11722 & n11723 ) ;
  assign n11725 = ( ~n11341 & n11722 ) | ( ~n11341 & n11723 ) | ( n11722 & n11723 ) ;
  assign n11726 = ( n11341 & ~n11724 ) | ( n11341 & n11725 ) | ( ~n11724 & n11725 ) ;
  assign n11727 = ( ~n6172 & n11721 ) | ( ~n6172 & n11726 ) | ( n11721 & n11726 ) ;
  assign n11728 = ( n6172 & ~n11342 ) | ( n6172 & n11620 ) | ( ~n11342 & n11620 ) ;
  assign n11729 = n6172 & ~n11342 ;
  assign n11730 = ( n11347 & n11728 ) | ( n11347 & n11729 ) | ( n11728 & n11729 ) ;
  assign n11731 = ( ~n11347 & n11728 ) | ( ~n11347 & n11729 ) | ( n11728 & n11729 ) ;
  assign n11732 = ( n11347 & ~n11730 ) | ( n11347 & n11731 ) | ( ~n11730 & n11731 ) ;
  assign n11733 = ( ~n5905 & n11727 ) | ( ~n5905 & n11732 ) | ( n11727 & n11732 ) ;
  assign n11734 = ~n5905 & n11348 ;
  assign n11735 = ( ~n5905 & n11348 ) | ( ~n5905 & n11620 ) | ( n11348 & n11620 ) ;
  assign n11736 = ( n11353 & n11734 ) | ( n11353 & n11735 ) | ( n11734 & n11735 ) ;
  assign n11737 = ( ~n11353 & n11734 ) | ( ~n11353 & n11735 ) | ( n11734 & n11735 ) ;
  assign n11738 = ( n11353 & ~n11736 ) | ( n11353 & n11737 ) | ( ~n11736 & n11737 ) ;
  assign n11739 = ( ~n5642 & n11733 ) | ( ~n5642 & n11738 ) | ( n11733 & n11738 ) ;
  assign n11740 = ( n5642 & ~n11354 ) | ( n5642 & n11620 ) | ( ~n11354 & n11620 ) ;
  assign n11741 = n5642 & ~n11354 ;
  assign n11742 = ( n11359 & n11740 ) | ( n11359 & n11741 ) | ( n11740 & n11741 ) ;
  assign n11743 = ( ~n11359 & n11740 ) | ( ~n11359 & n11741 ) | ( n11740 & n11741 ) ;
  assign n11744 = ( n11359 & ~n11742 ) | ( n11359 & n11743 ) | ( ~n11742 & n11743 ) ;
  assign n11745 = ( ~n5386 & n11739 ) | ( ~n5386 & n11744 ) | ( n11739 & n11744 ) ;
  assign n11746 = n5386 & ~n11360 ;
  assign n11747 = ( n5386 & ~n11360 ) | ( n5386 & n11620 ) | ( ~n11360 & n11620 ) ;
  assign n11748 = ( n11365 & n11746 ) | ( n11365 & n11747 ) | ( n11746 & n11747 ) ;
  assign n11749 = ( ~n11365 & n11746 ) | ( ~n11365 & n11747 ) | ( n11746 & n11747 ) ;
  assign n11750 = ( n11365 & ~n11748 ) | ( n11365 & n11749 ) | ( ~n11748 & n11749 ) ;
  assign n11751 = ( ~n5139 & n11745 ) | ( ~n5139 & n11750 ) | ( n11745 & n11750 ) ;
  assign n11752 = ( n5139 & ~n11366 ) | ( n5139 & n11620 ) | ( ~n11366 & n11620 ) ;
  assign n11753 = n5139 & ~n11366 ;
  assign n11754 = ( n11371 & n11752 ) | ( n11371 & n11753 ) | ( n11752 & n11753 ) ;
  assign n11755 = ( ~n11371 & n11752 ) | ( ~n11371 & n11753 ) | ( n11752 & n11753 ) ;
  assign n11756 = ( n11371 & ~n11754 ) | ( n11371 & n11755 ) | ( ~n11754 & n11755 ) ;
  assign n11757 = ( ~n4898 & n11751 ) | ( ~n4898 & n11756 ) | ( n11751 & n11756 ) ;
  assign n11758 = ( n4898 & ~n11372 ) | ( n4898 & n11620 ) | ( ~n11372 & n11620 ) ;
  assign n11759 = n4898 & ~n11372 ;
  assign n11760 = ( n11377 & n11758 ) | ( n11377 & n11759 ) | ( n11758 & n11759 ) ;
  assign n11761 = ( ~n11377 & n11758 ) | ( ~n11377 & n11759 ) | ( n11758 & n11759 ) ;
  assign n11762 = ( n11377 & ~n11760 ) | ( n11377 & n11761 ) | ( ~n11760 & n11761 ) ;
  assign n11763 = ( ~n4661 & n11757 ) | ( ~n4661 & n11762 ) | ( n11757 & n11762 ) ;
  assign n11764 = ~n4661 & n11378 ;
  assign n11765 = ( ~n4661 & n11378 ) | ( ~n4661 & n11620 ) | ( n11378 & n11620 ) ;
  assign n11766 = ( ~n11383 & n11764 ) | ( ~n11383 & n11765 ) | ( n11764 & n11765 ) ;
  assign n11767 = ( n11383 & n11764 ) | ( n11383 & n11765 ) | ( n11764 & n11765 ) ;
  assign n11768 = ( n11383 & n11766 ) | ( n11383 & ~n11767 ) | ( n11766 & ~n11767 ) ;
  assign n11769 = ( ~n4432 & n11763 ) | ( ~n4432 & n11768 ) | ( n11763 & n11768 ) ;
  assign n11770 = ( n4432 & ~n11384 ) | ( n4432 & n11620 ) | ( ~n11384 & n11620 ) ;
  assign n11771 = n4432 & ~n11384 ;
  assign n11772 = ( n11389 & n11770 ) | ( n11389 & n11771 ) | ( n11770 & n11771 ) ;
  assign n11773 = ( ~n11389 & n11770 ) | ( ~n11389 & n11771 ) | ( n11770 & n11771 ) ;
  assign n11774 = ( n11389 & ~n11772 ) | ( n11389 & n11773 ) | ( ~n11772 & n11773 ) ;
  assign n11775 = ( ~n4203 & n11769 ) | ( ~n4203 & n11774 ) | ( n11769 & n11774 ) ;
  assign n11776 = ( n4203 & ~n11390 ) | ( n4203 & n11620 ) | ( ~n11390 & n11620 ) ;
  assign n11777 = n4203 & ~n11390 ;
  assign n11778 = ( n11395 & n11776 ) | ( n11395 & n11777 ) | ( n11776 & n11777 ) ;
  assign n11779 = ( ~n11395 & n11776 ) | ( ~n11395 & n11777 ) | ( n11776 & n11777 ) ;
  assign n11780 = ( n11395 & ~n11778 ) | ( n11395 & n11779 ) | ( ~n11778 & n11779 ) ;
  assign n11781 = ( ~n3985 & n11775 ) | ( ~n3985 & n11780 ) | ( n11775 & n11780 ) ;
  assign n11782 = ( n3985 & ~n11396 ) | ( n3985 & n11620 ) | ( ~n11396 & n11620 ) ;
  assign n11783 = n3985 & ~n11396 ;
  assign n11784 = ( n11401 & n11782 ) | ( n11401 & n11783 ) | ( n11782 & n11783 ) ;
  assign n11785 = ( ~n11401 & n11782 ) | ( ~n11401 & n11783 ) | ( n11782 & n11783 ) ;
  assign n11786 = ( n11401 & ~n11784 ) | ( n11401 & n11785 ) | ( ~n11784 & n11785 ) ;
  assign n11787 = ( ~n3772 & n11781 ) | ( ~n3772 & n11786 ) | ( n11781 & n11786 ) ;
  assign n11788 = ( n3772 & ~n11402 ) | ( n3772 & n11620 ) | ( ~n11402 & n11620 ) ;
  assign n11789 = n3772 & ~n11402 ;
  assign n11790 = ( n11407 & n11788 ) | ( n11407 & n11789 ) | ( n11788 & n11789 ) ;
  assign n11791 = ( ~n11407 & n11788 ) | ( ~n11407 & n11789 ) | ( n11788 & n11789 ) ;
  assign n11792 = ( n11407 & ~n11790 ) | ( n11407 & n11791 ) | ( ~n11790 & n11791 ) ;
  assign n11793 = ( ~n3567 & n11787 ) | ( ~n3567 & n11792 ) | ( n11787 & n11792 ) ;
  assign n11794 = ( n3567 & ~n11408 ) | ( n3567 & n11620 ) | ( ~n11408 & n11620 ) ;
  assign n11795 = n3567 & ~n11408 ;
  assign n11796 = ( n11413 & n11794 ) | ( n11413 & n11795 ) | ( n11794 & n11795 ) ;
  assign n11797 = ( ~n11413 & n11794 ) | ( ~n11413 & n11795 ) | ( n11794 & n11795 ) ;
  assign n11798 = ( n11413 & ~n11796 ) | ( n11413 & n11797 ) | ( ~n11796 & n11797 ) ;
  assign n11799 = ( ~n3362 & n11793 ) | ( ~n3362 & n11798 ) | ( n11793 & n11798 ) ;
  assign n11800 = ( n3362 & ~n11414 ) | ( n3362 & n11620 ) | ( ~n11414 & n11620 ) ;
  assign n11801 = n3362 & ~n11414 ;
  assign n11802 = ( n11419 & n11800 ) | ( n11419 & n11801 ) | ( n11800 & n11801 ) ;
  assign n11803 = ( ~n11419 & n11800 ) | ( ~n11419 & n11801 ) | ( n11800 & n11801 ) ;
  assign n11804 = ( n11419 & ~n11802 ) | ( n11419 & n11803 ) | ( ~n11802 & n11803 ) ;
  assign n11805 = ( ~n3169 & n11799 ) | ( ~n3169 & n11804 ) | ( n11799 & n11804 ) ;
  assign n11806 = ( n3169 & ~n11420 ) | ( n3169 & n11620 ) | ( ~n11420 & n11620 ) ;
  assign n11807 = n3169 & ~n11420 ;
  assign n11808 = ( n11425 & n11806 ) | ( n11425 & n11807 ) | ( n11806 & n11807 ) ;
  assign n11809 = ( ~n11425 & n11806 ) | ( ~n11425 & n11807 ) | ( n11806 & n11807 ) ;
  assign n11810 = ( n11425 & ~n11808 ) | ( n11425 & n11809 ) | ( ~n11808 & n11809 ) ;
  assign n11811 = ( ~n2979 & n11805 ) | ( ~n2979 & n11810 ) | ( n11805 & n11810 ) ;
  assign n11812 = ( n2979 & ~n11426 ) | ( n2979 & n11620 ) | ( ~n11426 & n11620 ) ;
  assign n11813 = n2979 & ~n11426 ;
  assign n11814 = ( n11431 & n11812 ) | ( n11431 & n11813 ) | ( n11812 & n11813 ) ;
  assign n11815 = ( ~n11431 & n11812 ) | ( ~n11431 & n11813 ) | ( n11812 & n11813 ) ;
  assign n11816 = ( n11431 & ~n11814 ) | ( n11431 & n11815 ) | ( ~n11814 & n11815 ) ;
  assign n11817 = ( ~n2791 & n11811 ) | ( ~n2791 & n11816 ) | ( n11811 & n11816 ) ;
  assign n11818 = ~n2791 & n11432 ;
  assign n11819 = ( ~n2791 & n11432 ) | ( ~n2791 & n11620 ) | ( n11432 & n11620 ) ;
  assign n11820 = ( n11437 & n11818 ) | ( n11437 & n11819 ) | ( n11818 & n11819 ) ;
  assign n11821 = ( ~n11437 & n11818 ) | ( ~n11437 & n11819 ) | ( n11818 & n11819 ) ;
  assign n11822 = ( n11437 & ~n11820 ) | ( n11437 & n11821 ) | ( ~n11820 & n11821 ) ;
  assign n11823 = ( ~n2615 & n11817 ) | ( ~n2615 & n11822 ) | ( n11817 & n11822 ) ;
  assign n11824 = ~n2615 & n11438 ;
  assign n11825 = ( ~n2615 & n11438 ) | ( ~n2615 & n11620 ) | ( n11438 & n11620 ) ;
  assign n11826 = ( ~n11443 & n11824 ) | ( ~n11443 & n11825 ) | ( n11824 & n11825 ) ;
  assign n11827 = ( n11443 & n11824 ) | ( n11443 & n11825 ) | ( n11824 & n11825 ) ;
  assign n11828 = ( n11443 & n11826 ) | ( n11443 & ~n11827 ) | ( n11826 & ~n11827 ) ;
  assign n11829 = ( ~n2443 & n11823 ) | ( ~n2443 & n11828 ) | ( n11823 & n11828 ) ;
  assign n11830 = ~n2443 & n11444 ;
  assign n11831 = ( ~n2443 & n11444 ) | ( ~n2443 & n11620 ) | ( n11444 & n11620 ) ;
  assign n11832 = ( ~n11449 & n11830 ) | ( ~n11449 & n11831 ) | ( n11830 & n11831 ) ;
  assign n11833 = ( n11449 & n11830 ) | ( n11449 & n11831 ) | ( n11830 & n11831 ) ;
  assign n11834 = ( n11449 & n11832 ) | ( n11449 & ~n11833 ) | ( n11832 & ~n11833 ) ;
  assign n11835 = ( ~n2277 & n11829 ) | ( ~n2277 & n11834 ) | ( n11829 & n11834 ) ;
  assign n11836 = ( n2277 & ~n11450 ) | ( n2277 & n11620 ) | ( ~n11450 & n11620 ) ;
  assign n11837 = n2277 & ~n11450 ;
  assign n11838 = ( n11455 & n11836 ) | ( n11455 & n11837 ) | ( n11836 & n11837 ) ;
  assign n11839 = ( ~n11455 & n11836 ) | ( ~n11455 & n11837 ) | ( n11836 & n11837 ) ;
  assign n11840 = ( n11455 & ~n11838 ) | ( n11455 & n11839 ) | ( ~n11838 & n11839 ) ;
  assign n11841 = ( ~n2111 & n11835 ) | ( ~n2111 & n11840 ) | ( n11835 & n11840 ) ;
  assign n11842 = ( n2111 & ~n11456 ) | ( n2111 & n11620 ) | ( ~n11456 & n11620 ) ;
  assign n11843 = n2111 & ~n11456 ;
  assign n11844 = ( n11461 & n11842 ) | ( n11461 & n11843 ) | ( n11842 & n11843 ) ;
  assign n11845 = ( ~n11461 & n11842 ) | ( ~n11461 & n11843 ) | ( n11842 & n11843 ) ;
  assign n11846 = ( n11461 & ~n11844 ) | ( n11461 & n11845 ) | ( ~n11844 & n11845 ) ;
  assign n11847 = ( ~n1949 & n11841 ) | ( ~n1949 & n11846 ) | ( n11841 & n11846 ) ;
  assign n11848 = ( n1949 & ~n11462 ) | ( n1949 & n11620 ) | ( ~n11462 & n11620 ) ;
  assign n11849 = n1949 & ~n11462 ;
  assign n11850 = ( n11467 & n11848 ) | ( n11467 & n11849 ) | ( n11848 & n11849 ) ;
  assign n11851 = ( ~n11467 & n11848 ) | ( ~n11467 & n11849 ) | ( n11848 & n11849 ) ;
  assign n11852 = ( n11467 & ~n11850 ) | ( n11467 & n11851 ) | ( ~n11850 & n11851 ) ;
  assign n11853 = ( ~n1802 & n11847 ) | ( ~n1802 & n11852 ) | ( n11847 & n11852 ) ;
  assign n11854 = ~n1802 & n11468 ;
  assign n11855 = ( ~n1802 & n11468 ) | ( ~n1802 & n11620 ) | ( n11468 & n11620 ) ;
  assign n11856 = ( ~n11473 & n11854 ) | ( ~n11473 & n11855 ) | ( n11854 & n11855 ) ;
  assign n11857 = ( n11473 & n11854 ) | ( n11473 & n11855 ) | ( n11854 & n11855 ) ;
  assign n11858 = ( n11473 & n11856 ) | ( n11473 & ~n11857 ) | ( n11856 & ~n11857 ) ;
  assign n11859 = ( ~n1661 & n11853 ) | ( ~n1661 & n11858 ) | ( n11853 & n11858 ) ;
  assign n11860 = n1661 & ~n11474 ;
  assign n11861 = ( n1661 & ~n11474 ) | ( n1661 & n11620 ) | ( ~n11474 & n11620 ) ;
  assign n11862 = ( n11479 & n11860 ) | ( n11479 & n11861 ) | ( n11860 & n11861 ) ;
  assign n11863 = ( ~n11479 & n11860 ) | ( ~n11479 & n11861 ) | ( n11860 & n11861 ) ;
  assign n11864 = ( n11479 & ~n11862 ) | ( n11479 & n11863 ) | ( ~n11862 & n11863 ) ;
  assign n11865 = ( ~n1523 & n11859 ) | ( ~n1523 & n11864 ) | ( n11859 & n11864 ) ;
  assign n11866 = ~n1523 & n11480 ;
  assign n11867 = ( ~n1523 & n11480 ) | ( ~n1523 & n11620 ) | ( n11480 & n11620 ) ;
  assign n11868 = ( n11485 & n11866 ) | ( n11485 & n11867 ) | ( n11866 & n11867 ) ;
  assign n11869 = ( ~n11485 & n11866 ) | ( ~n11485 & n11867 ) | ( n11866 & n11867 ) ;
  assign n11870 = ( n11485 & ~n11868 ) | ( n11485 & n11869 ) | ( ~n11868 & n11869 ) ;
  assign n11871 = ( ~n1393 & n11865 ) | ( ~n1393 & n11870 ) | ( n11865 & n11870 ) ;
  assign n11872 = ~n1393 & n11486 ;
  assign n11873 = ( ~n1393 & n11486 ) | ( ~n1393 & n11620 ) | ( n11486 & n11620 ) ;
  assign n11874 = ( n11491 & n11872 ) | ( n11491 & n11873 ) | ( n11872 & n11873 ) ;
  assign n11875 = ( ~n11491 & n11872 ) | ( ~n11491 & n11873 ) | ( n11872 & n11873 ) ;
  assign n11876 = ( n11491 & ~n11874 ) | ( n11491 & n11875 ) | ( ~n11874 & n11875 ) ;
  assign n11877 = ( ~n1266 & n11871 ) | ( ~n1266 & n11876 ) | ( n11871 & n11876 ) ;
  assign n11878 = ( n1266 & ~n11492 ) | ( n1266 & n11620 ) | ( ~n11492 & n11620 ) ;
  assign n11879 = n1266 & ~n11492 ;
  assign n11880 = ( n11497 & n11878 ) | ( n11497 & n11879 ) | ( n11878 & n11879 ) ;
  assign n11881 = ( ~n11497 & n11878 ) | ( ~n11497 & n11879 ) | ( n11878 & n11879 ) ;
  assign n11882 = ( n11497 & ~n11880 ) | ( n11497 & n11881 ) | ( ~n11880 & n11881 ) ;
  assign n11883 = ( ~n1150 & n11877 ) | ( ~n1150 & n11882 ) | ( n11877 & n11882 ) ;
  assign n11884 = ( n1150 & ~n11498 ) | ( n1150 & n11620 ) | ( ~n11498 & n11620 ) ;
  assign n11885 = n1150 & ~n11498 ;
  assign n11886 = ( n11503 & n11884 ) | ( n11503 & n11885 ) | ( n11884 & n11885 ) ;
  assign n11887 = ( ~n11503 & n11884 ) | ( ~n11503 & n11885 ) | ( n11884 & n11885 ) ;
  assign n11888 = ( n11503 & ~n11886 ) | ( n11503 & n11887 ) | ( ~n11886 & n11887 ) ;
  assign n11889 = ( ~n1038 & n11883 ) | ( ~n1038 & n11888 ) | ( n11883 & n11888 ) ;
  assign n11890 = ( n1038 & ~n11504 ) | ( n1038 & n11620 ) | ( ~n11504 & n11620 ) ;
  assign n11891 = n1038 & ~n11504 ;
  assign n11892 = ( n11509 & n11890 ) | ( n11509 & n11891 ) | ( n11890 & n11891 ) ;
  assign n11893 = ( ~n11509 & n11890 ) | ( ~n11509 & n11891 ) | ( n11890 & n11891 ) ;
  assign n11894 = ( n11509 & ~n11892 ) | ( n11509 & n11893 ) | ( ~n11892 & n11893 ) ;
  assign n11895 = ( ~n933 & n11889 ) | ( ~n933 & n11894 ) | ( n11889 & n11894 ) ;
  assign n11896 = ( n933 & ~n11510 ) | ( n933 & n11620 ) | ( ~n11510 & n11620 ) ;
  assign n11897 = n933 & ~n11510 ;
  assign n11898 = ( n11515 & n11896 ) | ( n11515 & n11897 ) | ( n11896 & n11897 ) ;
  assign n11899 = ( ~n11515 & n11896 ) | ( ~n11515 & n11897 ) | ( n11896 & n11897 ) ;
  assign n11900 = ( n11515 & ~n11898 ) | ( n11515 & n11899 ) | ( ~n11898 & n11899 ) ;
  assign n11901 = ( ~n839 & n11895 ) | ( ~n839 & n11900 ) | ( n11895 & n11900 ) ;
  assign n11902 = ( n839 & ~n11516 ) | ( n839 & n11620 ) | ( ~n11516 & n11620 ) ;
  assign n11903 = n839 & ~n11516 ;
  assign n11904 = ( n11521 & n11902 ) | ( n11521 & n11903 ) | ( n11902 & n11903 ) ;
  assign n11905 = ( ~n11521 & n11902 ) | ( ~n11521 & n11903 ) | ( n11902 & n11903 ) ;
  assign n11906 = ( n11521 & ~n11904 ) | ( n11521 & n11905 ) | ( ~n11904 & n11905 ) ;
  assign n11907 = ( ~n746 & n11901 ) | ( ~n746 & n11906 ) | ( n11901 & n11906 ) ;
  assign n11908 = ~n746 & n11522 ;
  assign n11909 = ( ~n746 & n11522 ) | ( ~n746 & n11620 ) | ( n11522 & n11620 ) ;
  assign n11910 = ( n11527 & n11908 ) | ( n11527 & n11909 ) | ( n11908 & n11909 ) ;
  assign n11911 = ( ~n11527 & n11908 ) | ( ~n11527 & n11909 ) | ( n11908 & n11909 ) ;
  assign n11912 = ( n11527 & ~n11910 ) | ( n11527 & n11911 ) | ( ~n11910 & n11911 ) ;
  assign n11913 = ( ~n664 & n11907 ) | ( ~n664 & n11912 ) | ( n11907 & n11912 ) ;
  assign n11914 = ~n664 & n11528 ;
  assign n11915 = ( ~n664 & n11528 ) | ( ~n664 & n11620 ) | ( n11528 & n11620 ) ;
  assign n11916 = ( n11533 & n11914 ) | ( n11533 & n11915 ) | ( n11914 & n11915 ) ;
  assign n11917 = ( ~n11533 & n11914 ) | ( ~n11533 & n11915 ) | ( n11914 & n11915 ) ;
  assign n11918 = ( n11533 & ~n11916 ) | ( n11533 & n11917 ) | ( ~n11916 & n11917 ) ;
  assign n11919 = ( ~n588 & n11913 ) | ( ~n588 & n11918 ) | ( n11913 & n11918 ) ;
  assign n11920 = n588 & ~n11534 ;
  assign n11921 = ( n588 & ~n11534 ) | ( n588 & n11620 ) | ( ~n11534 & n11620 ) ;
  assign n11922 = ( n11539 & n11920 ) | ( n11539 & n11921 ) | ( n11920 & n11921 ) ;
  assign n11923 = ( ~n11539 & n11920 ) | ( ~n11539 & n11921 ) | ( n11920 & n11921 ) ;
  assign n11924 = ( n11539 & ~n11922 ) | ( n11539 & n11923 ) | ( ~n11922 & n11923 ) ;
  assign n11925 = ( ~n518 & n11919 ) | ( ~n518 & n11924 ) | ( n11919 & n11924 ) ;
  assign n11926 = ( n518 & ~n11540 ) | ( n518 & n11620 ) | ( ~n11540 & n11620 ) ;
  assign n11927 = n518 & ~n11540 ;
  assign n11928 = ( n11545 & n11926 ) | ( n11545 & n11927 ) | ( n11926 & n11927 ) ;
  assign n11929 = ( ~n11545 & n11926 ) | ( ~n11545 & n11927 ) | ( n11926 & n11927 ) ;
  assign n11930 = ( n11545 & ~n11928 ) | ( n11545 & n11929 ) | ( ~n11928 & n11929 ) ;
  assign n11931 = ( ~n454 & n11925 ) | ( ~n454 & n11930 ) | ( n11925 & n11930 ) ;
  assign n11932 = ~n454 & n11546 ;
  assign n11933 = ( ~n454 & n11546 ) | ( ~n454 & n11620 ) | ( n11546 & n11620 ) ;
  assign n11934 = ( n11551 & n11932 ) | ( n11551 & n11933 ) | ( n11932 & n11933 ) ;
  assign n11935 = ( ~n11551 & n11932 ) | ( ~n11551 & n11933 ) | ( n11932 & n11933 ) ;
  assign n11936 = ( n11551 & ~n11934 ) | ( n11551 & n11935 ) | ( ~n11934 & n11935 ) ;
  assign n11937 = ( ~n396 & n11931 ) | ( ~n396 & n11936 ) | ( n11931 & n11936 ) ;
  assign n11938 = ( n396 & ~n11552 ) | ( n396 & n11620 ) | ( ~n11552 & n11620 ) ;
  assign n11939 = n396 & ~n11552 ;
  assign n11940 = ( n11557 & n11938 ) | ( n11557 & n11939 ) | ( n11938 & n11939 ) ;
  assign n11941 = ( ~n11557 & n11938 ) | ( ~n11557 & n11939 ) | ( n11938 & n11939 ) ;
  assign n11942 = ( n11557 & ~n11940 ) | ( n11557 & n11941 ) | ( ~n11940 & n11941 ) ;
  assign n11943 = ( ~n344 & n11937 ) | ( ~n344 & n11942 ) | ( n11937 & n11942 ) ;
  assign n11944 = n344 & ~n11558 ;
  assign n11945 = ( n344 & ~n11558 ) | ( n344 & n11620 ) | ( ~n11558 & n11620 ) ;
  assign n11946 = ( ~n11563 & n11944 ) | ( ~n11563 & n11945 ) | ( n11944 & n11945 ) ;
  assign n11947 = ( n11563 & n11944 ) | ( n11563 & n11945 ) | ( n11944 & n11945 ) ;
  assign n11948 = ( n11563 & n11946 ) | ( n11563 & ~n11947 ) | ( n11946 & ~n11947 ) ;
  assign n11949 = ( ~n298 & n11943 ) | ( ~n298 & n11948 ) | ( n11943 & n11948 ) ;
  assign n11950 = ( n298 & ~n11564 ) | ( n298 & n11620 ) | ( ~n11564 & n11620 ) ;
  assign n11951 = n298 & ~n11564 ;
  assign n11952 = ( n11569 & n11950 ) | ( n11569 & n11951 ) | ( n11950 & n11951 ) ;
  assign n11953 = ( ~n11569 & n11950 ) | ( ~n11569 & n11951 ) | ( n11950 & n11951 ) ;
  assign n11954 = ( n11569 & ~n11952 ) | ( n11569 & n11953 ) | ( ~n11952 & n11953 ) ;
  assign n11955 = ( ~n258 & n11949 ) | ( ~n258 & n11954 ) | ( n11949 & n11954 ) ;
  assign n11956 = ~n258 & n11570 ;
  assign n11957 = ( ~n258 & n11570 ) | ( ~n258 & n11620 ) | ( n11570 & n11620 ) ;
  assign n11958 = ( n11575 & n11956 ) | ( n11575 & n11957 ) | ( n11956 & n11957 ) ;
  assign n11959 = ( ~n11575 & n11956 ) | ( ~n11575 & n11957 ) | ( n11956 & n11957 ) ;
  assign n11960 = ( n11575 & ~n11958 ) | ( n11575 & n11959 ) | ( ~n11958 & n11959 ) ;
  assign n11961 = ( ~n225 & n11955 ) | ( ~n225 & n11960 ) | ( n11955 & n11960 ) ;
  assign n11962 = ( n225 & ~n11576 ) | ( n225 & n11620 ) | ( ~n11576 & n11620 ) ;
  assign n11963 = n225 & ~n11576 ;
  assign n11964 = ( n11581 & n11962 ) | ( n11581 & n11963 ) | ( n11962 & n11963 ) ;
  assign n11965 = ( ~n11581 & n11962 ) | ( ~n11581 & n11963 ) | ( n11962 & n11963 ) ;
  assign n11966 = ( n11581 & ~n11964 ) | ( n11581 & n11965 ) | ( ~n11964 & n11965 ) ;
  assign n11967 = ( ~n197 & n11961 ) | ( ~n197 & n11966 ) | ( n11961 & n11966 ) ;
  assign n11968 = ( n197 & ~n11582 ) | ( n197 & n11620 ) | ( ~n11582 & n11620 ) ;
  assign n11969 = n197 & ~n11582 ;
  assign n11970 = ( n11587 & n11968 ) | ( n11587 & n11969 ) | ( n11968 & n11969 ) ;
  assign n11971 = ( ~n11587 & n11968 ) | ( ~n11587 & n11969 ) | ( n11968 & n11969 ) ;
  assign n11972 = ( n11587 & ~n11970 ) | ( n11587 & n11971 ) | ( ~n11970 & n11971 ) ;
  assign n11973 = ( ~n170 & n11967 ) | ( ~n170 & n11972 ) | ( n11967 & n11972 ) ;
  assign n11974 = n170 & ~n11588 ;
  assign n11975 = ( n170 & ~n11588 ) | ( n170 & n11620 ) | ( ~n11588 & n11620 ) ;
  assign n11976 = ( n11593 & n11974 ) | ( n11593 & n11975 ) | ( n11974 & n11975 ) ;
  assign n11977 = ( ~n11593 & n11974 ) | ( ~n11593 & n11975 ) | ( n11974 & n11975 ) ;
  assign n11978 = ( n11593 & ~n11976 ) | ( n11593 & n11977 ) | ( ~n11976 & n11977 ) ;
  assign n11979 = ( ~n142 & n11973 ) | ( ~n142 & n11978 ) | ( n11973 & n11978 ) ;
  assign n11980 = ~n142 & n11594 ;
  assign n11981 = ( ~n142 & n11594 ) | ( ~n142 & n11620 ) | ( n11594 & n11620 ) ;
  assign n11982 = ( n11599 & n11980 ) | ( n11599 & n11981 ) | ( n11980 & n11981 ) ;
  assign n11983 = ( ~n11599 & n11980 ) | ( ~n11599 & n11981 ) | ( n11980 & n11981 ) ;
  assign n11984 = ( n11599 & ~n11982 ) | ( n11599 & n11983 ) | ( ~n11982 & n11983 ) ;
  assign n11985 = ( ~n132 & n11979 ) | ( ~n132 & n11984 ) | ( n11979 & n11984 ) ;
  assign n11986 = n11625 & ~n11985 ;
  assign n11987 = n11625 | n11985 ;
  assign n11988 = ~n11609 & n11614 ;
  assign n11989 = ( n131 & n11618 ) | ( n131 & ~n11988 ) | ( n11618 & ~n11988 ) ;
  assign n11990 = ( n131 & ~n11987 ) | ( n131 & n11989 ) | ( ~n11987 & n11989 ) ;
  assign n11991 = ( n11625 & ~n11986 ) | ( n11625 & n11990 ) | ( ~n11986 & n11990 ) ;
  assign n11992 = ( n11625 & ~n11985 ) | ( n11625 & n11989 ) | ( ~n11985 & n11989 ) ;
  assign n11993 = ( n11603 & ~n11609 ) | ( n11603 & n11614 ) | ( ~n11609 & n11614 ) ;
  assign n11994 = n11603 & ~n11993 ;
  assign n11995 = n11988 | n11994 ;
  assign n11996 = n131 & ~n11995 ;
  assign n11997 = ( n11985 & n11992 ) | ( n11985 & ~n11996 ) | ( n11992 & ~n11996 ) ;
  assign n11998 = ( n132 & ~n11979 ) | ( n132 & n11997 ) | ( ~n11979 & n11997 ) ;
  assign n11999 = n132 & ~n11979 ;
  assign n12000 = ( n11984 & ~n11998 ) | ( n11984 & n11999 ) | ( ~n11998 & n11999 ) ;
  assign n12001 = ( n11984 & n11998 ) | ( n11984 & n11999 ) | ( n11998 & n11999 ) ;
  assign n12002 = ( n11998 & n12000 ) | ( n11998 & ~n12001 ) | ( n12000 & ~n12001 ) ;
  assign n12003 = n11991 | n12002 ;
  assign n12004 = n131 & ~n12002 ;
  assign n12005 = n170 & ~n11967 ;
  assign n12006 = ( n170 & ~n11967 ) | ( n170 & n11997 ) | ( ~n11967 & n11997 ) ;
  assign n12007 = ( n11972 & n12005 ) | ( n11972 & n12006 ) | ( n12005 & n12006 ) ;
  assign n12008 = ( ~n11972 & n12005 ) | ( ~n11972 & n12006 ) | ( n12005 & n12006 ) ;
  assign n12009 = ( n11972 & ~n12007 ) | ( n11972 & n12008 ) | ( ~n12007 & n12008 ) ;
  assign n12010 = n197 & ~n11961 ;
  assign n12011 = ( n197 & ~n11961 ) | ( n197 & n11997 ) | ( ~n11961 & n11997 ) ;
  assign n12012 = ( n11966 & n12010 ) | ( n11966 & n12011 ) | ( n12010 & n12011 ) ;
  assign n12013 = ( ~n11966 & n12010 ) | ( ~n11966 & n12011 ) | ( n12010 & n12011 ) ;
  assign n12014 = ( n11966 & ~n12012 ) | ( n11966 & n12013 ) | ( ~n12012 & n12013 ) ;
  assign n12015 = ( n258 & ~n11949 ) | ( n258 & n11997 ) | ( ~n11949 & n11997 ) ;
  assign n12016 = n258 & ~n11949 ;
  assign n12017 = ( n11954 & n12015 ) | ( n11954 & n12016 ) | ( n12015 & n12016 ) ;
  assign n12018 = ( ~n11954 & n12015 ) | ( ~n11954 & n12016 ) | ( n12015 & n12016 ) ;
  assign n12019 = ( n11954 & ~n12017 ) | ( n11954 & n12018 ) | ( ~n12017 & n12018 ) ;
  assign n12020 = ( n344 & ~n11937 ) | ( n344 & n11997 ) | ( ~n11937 & n11997 ) ;
  assign n12021 = n344 & ~n11937 ;
  assign n12022 = ( n11942 & n12020 ) | ( n11942 & n12021 ) | ( n12020 & n12021 ) ;
  assign n12023 = ( ~n11942 & n12020 ) | ( ~n11942 & n12021 ) | ( n12020 & n12021 ) ;
  assign n12024 = ( n11942 & ~n12022 ) | ( n11942 & n12023 ) | ( ~n12022 & n12023 ) ;
  assign n12025 = n454 & ~n11925 ;
  assign n12026 = ( n454 & ~n11925 ) | ( n454 & n11997 ) | ( ~n11925 & n11997 ) ;
  assign n12027 = ( ~n11930 & n12025 ) | ( ~n11930 & n12026 ) | ( n12025 & n12026 ) ;
  assign n12028 = ( n11930 & n12025 ) | ( n11930 & n12026 ) | ( n12025 & n12026 ) ;
  assign n12029 = ( n11930 & n12027 ) | ( n11930 & ~n12028 ) | ( n12027 & ~n12028 ) ;
  assign n12030 = ( n518 & ~n11919 ) | ( n518 & n11997 ) | ( ~n11919 & n11997 ) ;
  assign n12031 = n518 & ~n11919 ;
  assign n12032 = ( n11924 & n12030 ) | ( n11924 & n12031 ) | ( n12030 & n12031 ) ;
  assign n12033 = ( ~n11924 & n12030 ) | ( ~n11924 & n12031 ) | ( n12030 & n12031 ) ;
  assign n12034 = ( n11924 & ~n12032 ) | ( n11924 & n12033 ) | ( ~n12032 & n12033 ) ;
  assign n12035 = ( n664 & ~n11907 ) | ( n664 & n11997 ) | ( ~n11907 & n11997 ) ;
  assign n12036 = n664 & ~n11907 ;
  assign n12037 = ( n11912 & n12035 ) | ( n11912 & n12036 ) | ( n12035 & n12036 ) ;
  assign n12038 = ( ~n11912 & n12035 ) | ( ~n11912 & n12036 ) | ( n12035 & n12036 ) ;
  assign n12039 = ( n11912 & ~n12037 ) | ( n11912 & n12038 ) | ( ~n12037 & n12038 ) ;
  assign n12040 = ( n933 & ~n11889 ) | ( n933 & n11997 ) | ( ~n11889 & n11997 ) ;
  assign n12041 = n933 & ~n11889 ;
  assign n12042 = ( n11894 & n12040 ) | ( n11894 & n12041 ) | ( n12040 & n12041 ) ;
  assign n12043 = ( ~n11894 & n12040 ) | ( ~n11894 & n12041 ) | ( n12040 & n12041 ) ;
  assign n12044 = ( n11894 & ~n12042 ) | ( n11894 & n12043 ) | ( ~n12042 & n12043 ) ;
  assign n12045 = ( n1150 & ~n11877 ) | ( n1150 & n11997 ) | ( ~n11877 & n11997 ) ;
  assign n12046 = n1150 & ~n11877 ;
  assign n12047 = ( n11882 & n12045 ) | ( n11882 & n12046 ) | ( n12045 & n12046 ) ;
  assign n12048 = ( ~n11882 & n12045 ) | ( ~n11882 & n12046 ) | ( n12045 & n12046 ) ;
  assign n12049 = ( n11882 & ~n12047 ) | ( n11882 & n12048 ) | ( ~n12047 & n12048 ) ;
  assign n12050 = ( n1266 & ~n11871 ) | ( n1266 & n11997 ) | ( ~n11871 & n11997 ) ;
  assign n12051 = n1266 & ~n11871 ;
  assign n12052 = ( n11876 & n12050 ) | ( n11876 & n12051 ) | ( n12050 & n12051 ) ;
  assign n12053 = ( ~n11876 & n12050 ) | ( ~n11876 & n12051 ) | ( n12050 & n12051 ) ;
  assign n12054 = ( n11876 & ~n12052 ) | ( n11876 & n12053 ) | ( ~n12052 & n12053 ) ;
  assign n12055 = ( n1949 & ~n11841 ) | ( n1949 & n11997 ) | ( ~n11841 & n11997 ) ;
  assign n12056 = n1949 & ~n11841 ;
  assign n12057 = ( n11846 & n12055 ) | ( n11846 & n12056 ) | ( n12055 & n12056 ) ;
  assign n12058 = ( ~n11846 & n12055 ) | ( ~n11846 & n12056 ) | ( n12055 & n12056 ) ;
  assign n12059 = ( n11846 & ~n12057 ) | ( n11846 & n12058 ) | ( ~n12057 & n12058 ) ;
  assign n12060 = ( n2277 & ~n11829 ) | ( n2277 & n11997 ) | ( ~n11829 & n11997 ) ;
  assign n12061 = n2277 & ~n11829 ;
  assign n12062 = ( n11834 & n12060 ) | ( n11834 & n12061 ) | ( n12060 & n12061 ) ;
  assign n12063 = ( ~n11834 & n12060 ) | ( ~n11834 & n12061 ) | ( n12060 & n12061 ) ;
  assign n12064 = ( n11834 & ~n12062 ) | ( n11834 & n12063 ) | ( ~n12062 & n12063 ) ;
  assign n12065 = ( n2443 & ~n11823 ) | ( n2443 & n11997 ) | ( ~n11823 & n11997 ) ;
  assign n12066 = n2443 & ~n11823 ;
  assign n12067 = ( n11828 & n12065 ) | ( n11828 & n12066 ) | ( n12065 & n12066 ) ;
  assign n12068 = ( ~n11828 & n12065 ) | ( ~n11828 & n12066 ) | ( n12065 & n12066 ) ;
  assign n12069 = ( n11828 & ~n12067 ) | ( n11828 & n12068 ) | ( ~n12067 & n12068 ) ;
  assign n12070 = ~n2615 & n11817 ;
  assign n12071 = ( ~n2615 & n11817 ) | ( ~n2615 & n11997 ) | ( n11817 & n11997 ) ;
  assign n12072 = ( ~n11822 & n12070 ) | ( ~n11822 & n12071 ) | ( n12070 & n12071 ) ;
  assign n12073 = ( n11822 & n12070 ) | ( n11822 & n12071 ) | ( n12070 & n12071 ) ;
  assign n12074 = ( n11822 & n12072 ) | ( n11822 & ~n12073 ) | ( n12072 & ~n12073 ) ;
  assign n12075 = ( n2979 & ~n11805 ) | ( n2979 & n11997 ) | ( ~n11805 & n11997 ) ;
  assign n12076 = n2979 & ~n11805 ;
  assign n12077 = ( n11810 & n12075 ) | ( n11810 & n12076 ) | ( n12075 & n12076 ) ;
  assign n12078 = ( ~n11810 & n12075 ) | ( ~n11810 & n12076 ) | ( n12075 & n12076 ) ;
  assign n12079 = ( n11810 & ~n12077 ) | ( n11810 & n12078 ) | ( ~n12077 & n12078 ) ;
  assign n12080 = ( n3362 & ~n11793 ) | ( n3362 & n11997 ) | ( ~n11793 & n11997 ) ;
  assign n12081 = n3362 & ~n11793 ;
  assign n12082 = ( n11798 & n12080 ) | ( n11798 & n12081 ) | ( n12080 & n12081 ) ;
  assign n12083 = ( ~n11798 & n12080 ) | ( ~n11798 & n12081 ) | ( n12080 & n12081 ) ;
  assign n12084 = ( n11798 & ~n12082 ) | ( n11798 & n12083 ) | ( ~n12082 & n12083 ) ;
  assign n12085 = ( n3567 & ~n11787 ) | ( n3567 & n11997 ) | ( ~n11787 & n11997 ) ;
  assign n12086 = n3567 & ~n11787 ;
  assign n12087 = ( n11792 & n12085 ) | ( n11792 & n12086 ) | ( n12085 & n12086 ) ;
  assign n12088 = ( ~n11792 & n12085 ) | ( ~n11792 & n12086 ) | ( n12085 & n12086 ) ;
  assign n12089 = ( n11792 & ~n12087 ) | ( n11792 & n12088 ) | ( ~n12087 & n12088 ) ;
  assign n12090 = ( n3772 & ~n11781 ) | ( n3772 & n11997 ) | ( ~n11781 & n11997 ) ;
  assign n12091 = n3772 & ~n11781 ;
  assign n12092 = ( n11786 & n12090 ) | ( n11786 & n12091 ) | ( n12090 & n12091 ) ;
  assign n12093 = ( ~n11786 & n12090 ) | ( ~n11786 & n12091 ) | ( n12090 & n12091 ) ;
  assign n12094 = ( n11786 & ~n12092 ) | ( n11786 & n12093 ) | ( ~n12092 & n12093 ) ;
  assign n12095 = n4203 & ~n11769 ;
  assign n12096 = ( n4203 & ~n11769 ) | ( n4203 & n11997 ) | ( ~n11769 & n11997 ) ;
  assign n12097 = ( n11774 & n12095 ) | ( n11774 & n12096 ) | ( n12095 & n12096 ) ;
  assign n12098 = ( ~n11774 & n12095 ) | ( ~n11774 & n12096 ) | ( n12095 & n12096 ) ;
  assign n12099 = ( n11774 & ~n12097 ) | ( n11774 & n12098 ) | ( ~n12097 & n12098 ) ;
  assign n12100 = n4432 & ~n11763 ;
  assign n12101 = ( n4432 & ~n11763 ) | ( n4432 & n11997 ) | ( ~n11763 & n11997 ) ;
  assign n12102 = ( n11768 & n12100 ) | ( n11768 & n12101 ) | ( n12100 & n12101 ) ;
  assign n12103 = ( ~n11768 & n12100 ) | ( ~n11768 & n12101 ) | ( n12100 & n12101 ) ;
  assign n12104 = ( n11768 & ~n12102 ) | ( n11768 & n12103 ) | ( ~n12102 & n12103 ) ;
  assign n12105 = ( n4661 & ~n11757 ) | ( n4661 & n11997 ) | ( ~n11757 & n11997 ) ;
  assign n12106 = n4661 & ~n11757 ;
  assign n12107 = ( n11762 & n12105 ) | ( n11762 & n12106 ) | ( n12105 & n12106 ) ;
  assign n12108 = ( ~n11762 & n12105 ) | ( ~n11762 & n12106 ) | ( n12105 & n12106 ) ;
  assign n12109 = ( n11762 & ~n12107 ) | ( n11762 & n12108 ) | ( ~n12107 & n12108 ) ;
  assign n12110 = ~n4898 & n11751 ;
  assign n12111 = ( ~n4898 & n11751 ) | ( ~n4898 & n11997 ) | ( n11751 & n11997 ) ;
  assign n12112 = ( ~n11756 & n12110 ) | ( ~n11756 & n12111 ) | ( n12110 & n12111 ) ;
  assign n12113 = ( n11756 & n12110 ) | ( n11756 & n12111 ) | ( n12110 & n12111 ) ;
  assign n12114 = ( n11756 & n12112 ) | ( n11756 & ~n12113 ) | ( n12112 & ~n12113 ) ;
  assign n12115 = ( n5139 & ~n11745 ) | ( n5139 & n11997 ) | ( ~n11745 & n11997 ) ;
  assign n12116 = n5139 & ~n11745 ;
  assign n12117 = ( n11750 & n12115 ) | ( n11750 & n12116 ) | ( n12115 & n12116 ) ;
  assign n12118 = ( ~n11750 & n12115 ) | ( ~n11750 & n12116 ) | ( n12115 & n12116 ) ;
  assign n12119 = ( n11750 & ~n12117 ) | ( n11750 & n12118 ) | ( ~n12117 & n12118 ) ;
  assign n12120 = ~n5386 & n11739 ;
  assign n12121 = ( ~n5386 & n11739 ) | ( ~n5386 & n11997 ) | ( n11739 & n11997 ) ;
  assign n12122 = ( ~n11744 & n12120 ) | ( ~n11744 & n12121 ) | ( n12120 & n12121 ) ;
  assign n12123 = ( n11744 & n12120 ) | ( n11744 & n12121 ) | ( n12120 & n12121 ) ;
  assign n12124 = ( n11744 & n12122 ) | ( n11744 & ~n12123 ) | ( n12122 & ~n12123 ) ;
  assign n12125 = ( n6172 & ~n11721 ) | ( n6172 & n11997 ) | ( ~n11721 & n11997 ) ;
  assign n12126 = n6172 & ~n11721 ;
  assign n12127 = ( n11726 & n12125 ) | ( n11726 & n12126 ) | ( n12125 & n12126 ) ;
  assign n12128 = ( ~n11726 & n12125 ) | ( ~n11726 & n12126 ) | ( n12125 & n12126 ) ;
  assign n12129 = ( n11726 & ~n12127 ) | ( n11726 & n12128 ) | ( ~n12127 & n12128 ) ;
  assign n12130 = ( n7006 & ~n11703 ) | ( n7006 & n11997 ) | ( ~n11703 & n11997 ) ;
  assign n12131 = n7006 & ~n11703 ;
  assign n12132 = ( n11708 & n12130 ) | ( n11708 & n12131 ) | ( n12130 & n12131 ) ;
  assign n12133 = ( ~n11708 & n12130 ) | ( ~n11708 & n12131 ) | ( n12130 & n12131 ) ;
  assign n12134 = ( n11708 & ~n12132 ) | ( n11708 & n12133 ) | ( ~n12132 & n12133 ) ;
  assign n12135 = ( n7296 & ~n11697 ) | ( n7296 & n11997 ) | ( ~n11697 & n11997 ) ;
  assign n12136 = n7296 & ~n11697 ;
  assign n12137 = ( n11702 & n12135 ) | ( n11702 & n12136 ) | ( n12135 & n12136 ) ;
  assign n12138 = ( ~n11702 & n12135 ) | ( ~n11702 & n12136 ) | ( n12135 & n12136 ) ;
  assign n12139 = ( n11702 & ~n12137 ) | ( n11702 & n12138 ) | ( ~n12137 & n12138 ) ;
  assign n12140 = ~n7897 & n11685 ;
  assign n12141 = ( ~n7897 & n11685 ) | ( ~n7897 & n11997 ) | ( n11685 & n11997 ) ;
  assign n12142 = ( n11690 & n12140 ) | ( n11690 & n12141 ) | ( n12140 & n12141 ) ;
  assign n12143 = ( ~n11690 & n12140 ) | ( ~n11690 & n12141 ) | ( n12140 & n12141 ) ;
  assign n12144 = ( n11690 & ~n12142 ) | ( n11690 & n12143 ) | ( ~n12142 & n12143 ) ;
  assign n12145 = ~n8201 & n11679 ;
  assign n12146 = ( ~n8201 & n11679 ) | ( ~n8201 & n11997 ) | ( n11679 & n11997 ) ;
  assign n12147 = ( n11684 & n12145 ) | ( n11684 & n12146 ) | ( n12145 & n12146 ) ;
  assign n12148 = ( ~n11684 & n12145 ) | ( ~n11684 & n12146 ) | ( n12145 & n12146 ) ;
  assign n12149 = ( n11684 & ~n12147 ) | ( n11684 & n12148 ) | ( ~n12147 & n12148 ) ;
  assign n12150 = ( n8517 & ~n11673 ) | ( n8517 & n11997 ) | ( ~n11673 & n11997 ) ;
  assign n12151 = n8517 & ~n11673 ;
  assign n12152 = ( n11678 & n12150 ) | ( n11678 & n12151 ) | ( n12150 & n12151 ) ;
  assign n12153 = ( ~n11678 & n12150 ) | ( ~n11678 & n12151 ) | ( n12150 & n12151 ) ;
  assign n12154 = ( n11678 & ~n12152 ) | ( n11678 & n12153 ) | ( ~n12152 & n12153 ) ;
  assign n12155 = n8838 & ~n11667 ;
  assign n12156 = ( n8838 & ~n11667 ) | ( n8838 & n11997 ) | ( ~n11667 & n11997 ) ;
  assign n12157 = ( ~n11672 & n12155 ) | ( ~n11672 & n12156 ) | ( n12155 & n12156 ) ;
  assign n12158 = ( n11672 & n12155 ) | ( n11672 & n12156 ) | ( n12155 & n12156 ) ;
  assign n12159 = ( n11672 & n12157 ) | ( n11672 & ~n12158 ) | ( n12157 & ~n12158 ) ;
  assign n12160 = n9167 & ~n11661 ;
  assign n12161 = ( n9167 & ~n11661 ) | ( n9167 & n11997 ) | ( ~n11661 & n11997 ) ;
  assign n12162 = ( n11666 & n12160 ) | ( n11666 & n12161 ) | ( n12160 & n12161 ) ;
  assign n12163 = ( ~n11666 & n12160 ) | ( ~n11666 & n12161 ) | ( n12160 & n12161 ) ;
  assign n12164 = ( n11666 & ~n12162 ) | ( n11666 & n12163 ) | ( ~n12162 & n12163 ) ;
  assign n12165 = ( n9497 & ~n11655 ) | ( n9497 & n11997 ) | ( ~n11655 & n11997 ) ;
  assign n12166 = n9497 & ~n11655 ;
  assign n12167 = ( n11660 & n12165 ) | ( n11660 & n12166 ) | ( n12165 & n12166 ) ;
  assign n12168 = ( ~n11660 & n12165 ) | ( ~n11660 & n12166 ) | ( n12165 & n12166 ) ;
  assign n12169 = ( n11660 & ~n12167 ) | ( n11660 & n12168 ) | ( ~n12167 & n12168 ) ;
  assign n12170 = ( n10533 & ~n11637 ) | ( n10533 & n11997 ) | ( ~n11637 & n11997 ) ;
  assign n12171 = n10533 & ~n11637 ;
  assign n12172 = ( n11642 & n12170 ) | ( n11642 & n12171 ) | ( n12170 & n12171 ) ;
  assign n12173 = ( ~n11642 & n12170 ) | ( ~n11642 & n12171 ) | ( n12170 & n12171 ) ;
  assign n12174 = ( n11642 & ~n12172 ) | ( n11642 & n12173 ) | ( ~n12172 & n12173 ) ;
  assign n12175 = n10888 & ~n11636 ;
  assign n12176 = ( n10888 & ~n11636 ) | ( n10888 & n11997 ) | ( ~n11636 & n11997 ) ;
  assign n12177 = ( ~n11630 & n12175 ) | ( ~n11630 & n12176 ) | ( n12175 & n12176 ) ;
  assign n12178 = ( n11630 & n12175 ) | ( n11630 & n12176 ) | ( n12175 & n12176 ) ;
  assign n12179 = ( n11630 & n12177 ) | ( n11630 & ~n12178 ) | ( n12177 & ~n12178 ) ;
  assign n12180 = n11620 & ~n11997 ;
  assign n12181 = ~n11631 & n11997 ;
  assign n12182 = ( x4 & n12180 ) | ( x4 & n12181 ) | ( n12180 & n12181 ) ;
  assign n12183 = ( ~x4 & n12180 ) | ( ~x4 & n12181 ) | ( n12180 & n12181 ) ;
  assign n12184 = ( x4 & ~n12182 ) | ( x4 & n12183 ) | ( ~n12182 & n12183 ) ;
  assign n12185 = x0 | x1 ;
  assign n12186 = x2 | n12185 ;
  assign n12187 = n11620 & ~n12186 ;
  assign n12188 = ~n11620 & n12186 ;
  assign n12189 = ( x3 & ~n11997 ) | ( x3 & n12188 ) | ( ~n11997 & n12188 ) ;
  assign n12190 = ( n12181 & ~n12187 ) | ( n12181 & n12189 ) | ( ~n12187 & n12189 ) ;
  assign n12191 = ( ~n11252 & n12184 ) | ( ~n11252 & n12190 ) | ( n12184 & n12190 ) ;
  assign n12192 = ~n11252 & n11620 ;
  assign n12193 = ( n11627 & n11997 ) | ( n11627 & n12192 ) | ( n11997 & n12192 ) ;
  assign n12194 = ( ~x5 & n12183 ) | ( ~x5 & n12193 ) | ( n12183 & n12193 ) ;
  assign n12195 = ( x5 & n12183 ) | ( x5 & n12193 ) | ( n12183 & n12193 ) ;
  assign n12196 = ( x5 & n12194 ) | ( x5 & ~n12195 ) | ( n12194 & ~n12195 ) ;
  assign n12197 = ( ~n10888 & n12191 ) | ( ~n10888 & n12196 ) | ( n12191 & n12196 ) ;
  assign n12198 = ( ~n10533 & n12179 ) | ( ~n10533 & n12197 ) | ( n12179 & n12197 ) ;
  assign n12199 = ( ~n10180 & n12174 ) | ( ~n10180 & n12198 ) | ( n12174 & n12198 ) ;
  assign n12200 = ( n10180 & ~n11643 ) | ( n10180 & n11997 ) | ( ~n11643 & n11997 ) ;
  assign n12201 = n10180 & ~n11643 ;
  assign n12202 = ( n11648 & n12200 ) | ( n11648 & n12201 ) | ( n12200 & n12201 ) ;
  assign n12203 = ( ~n11648 & n12200 ) | ( ~n11648 & n12201 ) | ( n12200 & n12201 ) ;
  assign n12204 = ( n11648 & ~n12202 ) | ( n11648 & n12203 ) | ( ~n12202 & n12203 ) ;
  assign n12205 = ( ~n9834 & n12199 ) | ( ~n9834 & n12204 ) | ( n12199 & n12204 ) ;
  assign n12206 = ~n9834 & n11649 ;
  assign n12207 = ( ~n9834 & n11649 ) | ( ~n9834 & n11997 ) | ( n11649 & n11997 ) ;
  assign n12208 = ( n11654 & n12206 ) | ( n11654 & n12207 ) | ( n12206 & n12207 ) ;
  assign n12209 = ( ~n11654 & n12206 ) | ( ~n11654 & n12207 ) | ( n12206 & n12207 ) ;
  assign n12210 = ( n11654 & ~n12208 ) | ( n11654 & n12209 ) | ( ~n12208 & n12209 ) ;
  assign n12211 = ( ~n9497 & n12205 ) | ( ~n9497 & n12210 ) | ( n12205 & n12210 ) ;
  assign n12212 = ( ~n9167 & n12169 ) | ( ~n9167 & n12211 ) | ( n12169 & n12211 ) ;
  assign n12213 = ( ~n8838 & n12164 ) | ( ~n8838 & n12212 ) | ( n12164 & n12212 ) ;
  assign n12214 = ( ~n8517 & n12159 ) | ( ~n8517 & n12213 ) | ( n12159 & n12213 ) ;
  assign n12215 = ( ~n8201 & n12154 ) | ( ~n8201 & n12214 ) | ( n12154 & n12214 ) ;
  assign n12216 = ( ~n7897 & n12149 ) | ( ~n7897 & n12215 ) | ( n12149 & n12215 ) ;
  assign n12217 = ( ~n7594 & n12144 ) | ( ~n7594 & n12216 ) | ( n12144 & n12216 ) ;
  assign n12218 = ( n7594 & ~n11691 ) | ( n7594 & n11997 ) | ( ~n11691 & n11997 ) ;
  assign n12219 = n7594 & ~n11691 ;
  assign n12220 = ( n11696 & n12218 ) | ( n11696 & n12219 ) | ( n12218 & n12219 ) ;
  assign n12221 = ( ~n11696 & n12218 ) | ( ~n11696 & n12219 ) | ( n12218 & n12219 ) ;
  assign n12222 = ( n11696 & ~n12220 ) | ( n11696 & n12221 ) | ( ~n12220 & n12221 ) ;
  assign n12223 = ( ~n7296 & n12217 ) | ( ~n7296 & n12222 ) | ( n12217 & n12222 ) ;
  assign n12224 = ( ~n7006 & n12139 ) | ( ~n7006 & n12223 ) | ( n12139 & n12223 ) ;
  assign n12225 = ( ~n6723 & n12134 ) | ( ~n6723 & n12224 ) | ( n12134 & n12224 ) ;
  assign n12226 = ( n6723 & ~n11709 ) | ( n6723 & n11997 ) | ( ~n11709 & n11997 ) ;
  assign n12227 = n6723 & ~n11709 ;
  assign n12228 = ( n11714 & n12226 ) | ( n11714 & n12227 ) | ( n12226 & n12227 ) ;
  assign n12229 = ( ~n11714 & n12226 ) | ( ~n11714 & n12227 ) | ( n12226 & n12227 ) ;
  assign n12230 = ( n11714 & ~n12228 ) | ( n11714 & n12229 ) | ( ~n12228 & n12229 ) ;
  assign n12231 = ( ~n6442 & n12225 ) | ( ~n6442 & n12230 ) | ( n12225 & n12230 ) ;
  assign n12232 = ( n6442 & ~n11715 ) | ( n6442 & n11997 ) | ( ~n11715 & n11997 ) ;
  assign n12233 = n6442 & ~n11715 ;
  assign n12234 = ( n11720 & n12232 ) | ( n11720 & n12233 ) | ( n12232 & n12233 ) ;
  assign n12235 = ( ~n11720 & n12232 ) | ( ~n11720 & n12233 ) | ( n12232 & n12233 ) ;
  assign n12236 = ( n11720 & ~n12234 ) | ( n11720 & n12235 ) | ( ~n12234 & n12235 ) ;
  assign n12237 = ( ~n6172 & n12231 ) | ( ~n6172 & n12236 ) | ( n12231 & n12236 ) ;
  assign n12238 = ( ~n5905 & n12129 ) | ( ~n5905 & n12237 ) | ( n12129 & n12237 ) ;
  assign n12239 = ~n5905 & n11727 ;
  assign n12240 = ( ~n5905 & n11727 ) | ( ~n5905 & n11997 ) | ( n11727 & n11997 ) ;
  assign n12241 = ( ~n11732 & n12239 ) | ( ~n11732 & n12240 ) | ( n12239 & n12240 ) ;
  assign n12242 = ( n11732 & n12239 ) | ( n11732 & n12240 ) | ( n12239 & n12240 ) ;
  assign n12243 = ( n11732 & n12241 ) | ( n11732 & ~n12242 ) | ( n12241 & ~n12242 ) ;
  assign n12244 = ( ~n5642 & n12238 ) | ( ~n5642 & n12243 ) | ( n12238 & n12243 ) ;
  assign n12245 = ( n5642 & ~n11733 ) | ( n5642 & n11997 ) | ( ~n11733 & n11997 ) ;
  assign n12246 = n5642 & ~n11733 ;
  assign n12247 = ( n11738 & n12245 ) | ( n11738 & n12246 ) | ( n12245 & n12246 ) ;
  assign n12248 = ( ~n11738 & n12245 ) | ( ~n11738 & n12246 ) | ( n12245 & n12246 ) ;
  assign n12249 = ( n11738 & ~n12247 ) | ( n11738 & n12248 ) | ( ~n12247 & n12248 ) ;
  assign n12250 = ( ~n5386 & n12244 ) | ( ~n5386 & n12249 ) | ( n12244 & n12249 ) ;
  assign n12251 = ( ~n5139 & n12124 ) | ( ~n5139 & n12250 ) | ( n12124 & n12250 ) ;
  assign n12252 = ( ~n4898 & n12119 ) | ( ~n4898 & n12251 ) | ( n12119 & n12251 ) ;
  assign n12253 = ( ~n4661 & n12114 ) | ( ~n4661 & n12252 ) | ( n12114 & n12252 ) ;
  assign n12254 = ( ~n4432 & n12109 ) | ( ~n4432 & n12253 ) | ( n12109 & n12253 ) ;
  assign n12255 = ( ~n4203 & n12104 ) | ( ~n4203 & n12254 ) | ( n12104 & n12254 ) ;
  assign n12256 = ( ~n3985 & n12099 ) | ( ~n3985 & n12255 ) | ( n12099 & n12255 ) ;
  assign n12257 = ( n3985 & ~n11775 ) | ( n3985 & n11997 ) | ( ~n11775 & n11997 ) ;
  assign n12258 = n3985 & ~n11775 ;
  assign n12259 = ( n11780 & n12257 ) | ( n11780 & n12258 ) | ( n12257 & n12258 ) ;
  assign n12260 = ( ~n11780 & n12257 ) | ( ~n11780 & n12258 ) | ( n12257 & n12258 ) ;
  assign n12261 = ( n11780 & ~n12259 ) | ( n11780 & n12260 ) | ( ~n12259 & n12260 ) ;
  assign n12262 = ( ~n3772 & n12256 ) | ( ~n3772 & n12261 ) | ( n12256 & n12261 ) ;
  assign n12263 = ( ~n3567 & n12094 ) | ( ~n3567 & n12262 ) | ( n12094 & n12262 ) ;
  assign n12264 = ( ~n3362 & n12089 ) | ( ~n3362 & n12263 ) | ( n12089 & n12263 ) ;
  assign n12265 = ( ~n3169 & n12084 ) | ( ~n3169 & n12264 ) | ( n12084 & n12264 ) ;
  assign n12266 = ( n3169 & ~n11799 ) | ( n3169 & n11997 ) | ( ~n11799 & n11997 ) ;
  assign n12267 = n3169 & ~n11799 ;
  assign n12268 = ( n11804 & n12266 ) | ( n11804 & n12267 ) | ( n12266 & n12267 ) ;
  assign n12269 = ( ~n11804 & n12266 ) | ( ~n11804 & n12267 ) | ( n12266 & n12267 ) ;
  assign n12270 = ( n11804 & ~n12268 ) | ( n11804 & n12269 ) | ( ~n12268 & n12269 ) ;
  assign n12271 = ( ~n2979 & n12265 ) | ( ~n2979 & n12270 ) | ( n12265 & n12270 ) ;
  assign n12272 = ( ~n2791 & n12079 ) | ( ~n2791 & n12271 ) | ( n12079 & n12271 ) ;
  assign n12273 = n2791 & ~n11811 ;
  assign n12274 = ( n2791 & ~n11811 ) | ( n2791 & n11997 ) | ( ~n11811 & n11997 ) ;
  assign n12275 = ( n11816 & n12273 ) | ( n11816 & n12274 ) | ( n12273 & n12274 ) ;
  assign n12276 = ( ~n11816 & n12273 ) | ( ~n11816 & n12274 ) | ( n12273 & n12274 ) ;
  assign n12277 = ( n11816 & ~n12275 ) | ( n11816 & n12276 ) | ( ~n12275 & n12276 ) ;
  assign n12278 = ( ~n2615 & n12272 ) | ( ~n2615 & n12277 ) | ( n12272 & n12277 ) ;
  assign n12279 = ( ~n2443 & n12074 ) | ( ~n2443 & n12278 ) | ( n12074 & n12278 ) ;
  assign n12280 = ( ~n2277 & n12069 ) | ( ~n2277 & n12279 ) | ( n12069 & n12279 ) ;
  assign n12281 = ( ~n2111 & n12064 ) | ( ~n2111 & n12280 ) | ( n12064 & n12280 ) ;
  assign n12282 = ( n2111 & ~n11835 ) | ( n2111 & n11997 ) | ( ~n11835 & n11997 ) ;
  assign n12283 = n2111 & ~n11835 ;
  assign n12284 = ( n11840 & n12282 ) | ( n11840 & n12283 ) | ( n12282 & n12283 ) ;
  assign n12285 = ( ~n11840 & n12282 ) | ( ~n11840 & n12283 ) | ( n12282 & n12283 ) ;
  assign n12286 = ( n11840 & ~n12284 ) | ( n11840 & n12285 ) | ( ~n12284 & n12285 ) ;
  assign n12287 = ( ~n1949 & n12281 ) | ( ~n1949 & n12286 ) | ( n12281 & n12286 ) ;
  assign n12288 = ( ~n1802 & n12059 ) | ( ~n1802 & n12287 ) | ( n12059 & n12287 ) ;
  assign n12289 = ~n1802 & n11847 ;
  assign n12290 = ( ~n1802 & n11847 ) | ( ~n1802 & n11997 ) | ( n11847 & n11997 ) ;
  assign n12291 = ( ~n11852 & n12289 ) | ( ~n11852 & n12290 ) | ( n12289 & n12290 ) ;
  assign n12292 = ( n11852 & n12289 ) | ( n11852 & n12290 ) | ( n12289 & n12290 ) ;
  assign n12293 = ( n11852 & n12291 ) | ( n11852 & ~n12292 ) | ( n12291 & ~n12292 ) ;
  assign n12294 = ( ~n1661 & n12288 ) | ( ~n1661 & n12293 ) | ( n12288 & n12293 ) ;
  assign n12295 = n1661 & ~n11853 ;
  assign n12296 = ( n1661 & ~n11853 ) | ( n1661 & n11997 ) | ( ~n11853 & n11997 ) ;
  assign n12297 = ( n11858 & n12295 ) | ( n11858 & n12296 ) | ( n12295 & n12296 ) ;
  assign n12298 = ( ~n11858 & n12295 ) | ( ~n11858 & n12296 ) | ( n12295 & n12296 ) ;
  assign n12299 = ( n11858 & ~n12297 ) | ( n11858 & n12298 ) | ( ~n12297 & n12298 ) ;
  assign n12300 = ( ~n1523 & n12294 ) | ( ~n1523 & n12299 ) | ( n12294 & n12299 ) ;
  assign n12301 = n1523 & ~n11859 ;
  assign n12302 = ( n1523 & ~n11859 ) | ( n1523 & n11997 ) | ( ~n11859 & n11997 ) ;
  assign n12303 = ( ~n11864 & n12301 ) | ( ~n11864 & n12302 ) | ( n12301 & n12302 ) ;
  assign n12304 = ( n11864 & n12301 ) | ( n11864 & n12302 ) | ( n12301 & n12302 ) ;
  assign n12305 = ( n11864 & n12303 ) | ( n11864 & ~n12304 ) | ( n12303 & ~n12304 ) ;
  assign n12306 = ( ~n1393 & n12300 ) | ( ~n1393 & n12305 ) | ( n12300 & n12305 ) ;
  assign n12307 = ( n1393 & ~n11865 ) | ( n1393 & n11997 ) | ( ~n11865 & n11997 ) ;
  assign n12308 = n1393 & ~n11865 ;
  assign n12309 = ( n11870 & n12307 ) | ( n11870 & n12308 ) | ( n12307 & n12308 ) ;
  assign n12310 = ( ~n11870 & n12307 ) | ( ~n11870 & n12308 ) | ( n12307 & n12308 ) ;
  assign n12311 = ( n11870 & ~n12309 ) | ( n11870 & n12310 ) | ( ~n12309 & n12310 ) ;
  assign n12312 = ( ~n1266 & n12306 ) | ( ~n1266 & n12311 ) | ( n12306 & n12311 ) ;
  assign n12313 = ( ~n1150 & n12054 ) | ( ~n1150 & n12312 ) | ( n12054 & n12312 ) ;
  assign n12314 = ( ~n1038 & n12049 ) | ( ~n1038 & n12313 ) | ( n12049 & n12313 ) ;
  assign n12315 = n1038 & ~n11883 ;
  assign n12316 = ( n1038 & ~n11883 ) | ( n1038 & n11997 ) | ( ~n11883 & n11997 ) ;
  assign n12317 = ( ~n11888 & n12315 ) | ( ~n11888 & n12316 ) | ( n12315 & n12316 ) ;
  assign n12318 = ( n11888 & n12315 ) | ( n11888 & n12316 ) | ( n12315 & n12316 ) ;
  assign n12319 = ( n11888 & n12317 ) | ( n11888 & ~n12318 ) | ( n12317 & ~n12318 ) ;
  assign n12320 = ( ~n933 & n12314 ) | ( ~n933 & n12319 ) | ( n12314 & n12319 ) ;
  assign n12321 = ( ~n839 & n12044 ) | ( ~n839 & n12320 ) | ( n12044 & n12320 ) ;
  assign n12322 = ( n839 & ~n11895 ) | ( n839 & n11997 ) | ( ~n11895 & n11997 ) ;
  assign n12323 = n839 & ~n11895 ;
  assign n12324 = ( n11900 & n12322 ) | ( n11900 & n12323 ) | ( n12322 & n12323 ) ;
  assign n12325 = ( ~n11900 & n12322 ) | ( ~n11900 & n12323 ) | ( n12322 & n12323 ) ;
  assign n12326 = ( n11900 & ~n12324 ) | ( n11900 & n12325 ) | ( ~n12324 & n12325 ) ;
  assign n12327 = ( ~n746 & n12321 ) | ( ~n746 & n12326 ) | ( n12321 & n12326 ) ;
  assign n12328 = n746 & ~n11901 ;
  assign n12329 = ( n746 & ~n11901 ) | ( n746 & n11997 ) | ( ~n11901 & n11997 ) ;
  assign n12330 = ( n11906 & n12328 ) | ( n11906 & n12329 ) | ( n12328 & n12329 ) ;
  assign n12331 = ( ~n11906 & n12328 ) | ( ~n11906 & n12329 ) | ( n12328 & n12329 ) ;
  assign n12332 = ( n11906 & ~n12330 ) | ( n11906 & n12331 ) | ( ~n12330 & n12331 ) ;
  assign n12333 = ( ~n664 & n12327 ) | ( ~n664 & n12332 ) | ( n12327 & n12332 ) ;
  assign n12334 = ( ~n588 & n12039 ) | ( ~n588 & n12333 ) | ( n12039 & n12333 ) ;
  assign n12335 = ~n588 & n11913 ;
  assign n12336 = ( ~n588 & n11913 ) | ( ~n588 & n11997 ) | ( n11913 & n11997 ) ;
  assign n12337 = ( ~n11918 & n12335 ) | ( ~n11918 & n12336 ) | ( n12335 & n12336 ) ;
  assign n12338 = ( n11918 & n12335 ) | ( n11918 & n12336 ) | ( n12335 & n12336 ) ;
  assign n12339 = ( n11918 & n12337 ) | ( n11918 & ~n12338 ) | ( n12337 & ~n12338 ) ;
  assign n12340 = ( ~n518 & n12334 ) | ( ~n518 & n12339 ) | ( n12334 & n12339 ) ;
  assign n12341 = ( ~n454 & n12034 ) | ( ~n454 & n12340 ) | ( n12034 & n12340 ) ;
  assign n12342 = ( ~n396 & n12029 ) | ( ~n396 & n12341 ) | ( n12029 & n12341 ) ;
  assign n12343 = ( n396 & ~n11931 ) | ( n396 & n11997 ) | ( ~n11931 & n11997 ) ;
  assign n12344 = n396 & ~n11931 ;
  assign n12345 = ( n11936 & n12343 ) | ( n11936 & n12344 ) | ( n12343 & n12344 ) ;
  assign n12346 = ( ~n11936 & n12343 ) | ( ~n11936 & n12344 ) | ( n12343 & n12344 ) ;
  assign n12347 = ( n11936 & ~n12345 ) | ( n11936 & n12346 ) | ( ~n12345 & n12346 ) ;
  assign n12348 = ( ~n344 & n12342 ) | ( ~n344 & n12347 ) | ( n12342 & n12347 ) ;
  assign n12349 = ( ~n298 & n12024 ) | ( ~n298 & n12348 ) | ( n12024 & n12348 ) ;
  assign n12350 = ( n298 & ~n11943 ) | ( n298 & n11997 ) | ( ~n11943 & n11997 ) ;
  assign n12351 = n298 & ~n11943 ;
  assign n12352 = ( n11948 & n12350 ) | ( n11948 & n12351 ) | ( n12350 & n12351 ) ;
  assign n12353 = ( ~n11948 & n12350 ) | ( ~n11948 & n12351 ) | ( n12350 & n12351 ) ;
  assign n12354 = ( n11948 & ~n12352 ) | ( n11948 & n12353 ) | ( ~n12352 & n12353 ) ;
  assign n12355 = ( ~n258 & n12349 ) | ( ~n258 & n12354 ) | ( n12349 & n12354 ) ;
  assign n12356 = ( ~n225 & n12019 ) | ( ~n225 & n12355 ) | ( n12019 & n12355 ) ;
  assign n12357 = ( n225 & ~n11955 ) | ( n225 & n11997 ) | ( ~n11955 & n11997 ) ;
  assign n12358 = n225 & ~n11955 ;
  assign n12359 = ( n11960 & n12357 ) | ( n11960 & n12358 ) | ( n12357 & n12358 ) ;
  assign n12360 = ( ~n11960 & n12357 ) | ( ~n11960 & n12358 ) | ( n12357 & n12358 ) ;
  assign n12361 = ( n11960 & ~n12359 ) | ( n11960 & n12360 ) | ( ~n12359 & n12360 ) ;
  assign n12362 = ( ~n197 & n12356 ) | ( ~n197 & n12361 ) | ( n12356 & n12361 ) ;
  assign n12363 = ( ~n170 & n12014 ) | ( ~n170 & n12362 ) | ( n12014 & n12362 ) ;
  assign n12364 = ( ~n142 & n12009 ) | ( ~n142 & n12363 ) | ( n12009 & n12363 ) ;
  assign n12365 = n142 & ~n11973 ;
  assign n12366 = ( n142 & ~n11973 ) | ( n142 & n11997 ) | ( ~n11973 & n11997 ) ;
  assign n12367 = ( n11978 & n12365 ) | ( n11978 & n12366 ) | ( n12365 & n12366 ) ;
  assign n12368 = ( ~n11978 & n12365 ) | ( ~n11978 & n12366 ) | ( n12365 & n12366 ) ;
  assign n12369 = ( n11978 & ~n12367 ) | ( n11978 & n12368 ) | ( ~n12367 & n12368 ) ;
  assign n12370 = ( ~n132 & n12364 ) | ( ~n132 & n12369 ) | ( n12364 & n12369 ) ;
  assign n12371 = ~n12004 & n12370 ;
  assign n12372 = ( n131 & n11625 ) | ( n131 & ~n11995 ) | ( n11625 & ~n11995 ) ;
  assign n12373 = ( n131 & ~n11625 ) | ( n131 & n11985 ) | ( ~n11625 & n11985 ) ;
  assign n12374 = ( ~n11987 & n12372 ) | ( ~n11987 & n12373 ) | ( n12372 & n12373 ) ;
  assign n12375 = ( n12003 & n12371 ) | ( n12003 & ~n12374 ) | ( n12371 & ~n12374 ) ;
  assign y0 = n12375 ;
  assign y1 = n11997 ;
  assign y2 = n11620 ;
  assign y3 = n11252 ;
  assign y4 = n10888 ;
  assign y5 = n10533 ;
  assign y6 = n10180 ;
  assign y7 = n9834 ;
  assign y8 = n9497 ;
  assign y9 = n9167 ;
  assign y10 = n8838 ;
  assign y11 = n8517 ;
  assign y12 = n8201 ;
  assign y13 = n7897 ;
  assign y14 = n7594 ;
  assign y15 = n7296 ;
  assign y16 = n7006 ;
  assign y17 = n6723 ;
  assign y18 = n6442 ;
  assign y19 = n6172 ;
  assign y20 = n5905 ;
  assign y21 = n5642 ;
  assign y22 = n5386 ;
  assign y23 = n5139 ;
  assign y24 = n4898 ;
  assign y25 = n4661 ;
  assign y26 = n4432 ;
  assign y27 = n4203 ;
  assign y28 = n3985 ;
  assign y29 = n3772 ;
  assign y30 = n3567 ;
  assign y31 = n3362 ;
  assign y32 = n3169 ;
  assign y33 = n2979 ;
  assign y34 = n2791 ;
  assign y35 = n2615 ;
  assign y36 = n2443 ;
  assign y37 = n2277 ;
  assign y38 = n2111 ;
  assign y39 = n1949 ;
  assign y40 = n1802 ;
  assign y41 = n1661 ;
  assign y42 = n1523 ;
  assign y43 = n1393 ;
  assign y44 = n1266 ;
  assign y45 = n1150 ;
  assign y46 = n1038 ;
  assign y47 = n933 ;
  assign y48 = n839 ;
  assign y49 = n746 ;
  assign y50 = n664 ;
  assign y51 = n588 ;
  assign y52 = n518 ;
  assign y53 = n454 ;
  assign y54 = n396 ;
  assign y55 = n344 ;
  assign y56 = n298 ;
  assign y57 = n258 ;
  assign y58 = n225 ;
  assign y59 = n197 ;
  assign y60 = n170 ;
  assign y61 = n142 ;
  assign y62 = n132 ;
  assign y63 = n131 ;
endmodule
