module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 ;
  assign n9 = x4 | x5 ;
  assign n10 = ~x6 & x7 ;
  assign n11 = ~n9 & n10 ;
  assign n12 = x0 | x2 ;
  assign n13 = x1 | x3 ;
  assign n14 = n12 | n13 ;
  assign n15 = n11 & ~n14 ;
  assign n16 = x0 & ~x2 ;
  assign n17 = ~n13 & n16 ;
  assign n18 = n11 & n17 ;
  assign n19 = x1 & ~x3 ;
  assign n20 = ~n12 & n19 ;
  assign n21 = n11 & n20 ;
  assign n22 = n16 & n19 ;
  assign n23 = n11 & n22 ;
  assign n24 = ~x0 & x2 ;
  assign n25 = ~n13 & n24 ;
  assign n26 = n11 & n25 ;
  assign n27 = x0 & x2 ;
  assign n28 = ~n13 & n27 ;
  assign n29 = n11 & n28 ;
  assign n30 = n19 & n24 ;
  assign n31 = n11 & n30 ;
  assign n32 = n19 & n27 ;
  assign n33 = n11 & n32 ;
  assign n34 = ~x1 & x3 ;
  assign n35 = ~n12 & n34 ;
  assign n36 = n11 & n35 ;
  assign n37 = n16 & n34 ;
  assign n38 = n11 & n37 ;
  assign n39 = x1 & x3 ;
  assign n40 = ~n12 & n39 ;
  assign n41 = n11 & n40 ;
  assign n42 = n16 & n39 ;
  assign n43 = n11 & n42 ;
  assign n44 = n24 & n34 ;
  assign n45 = n11 & n44 ;
  assign n46 = n27 & n34 ;
  assign n47 = n11 & n46 ;
  assign n48 = n24 & n39 ;
  assign n49 = n11 & n48 ;
  assign n50 = n27 & n39 ;
  assign n51 = n11 & n50 ;
  assign n52 = x4 & ~x5 ;
  assign n53 = n10 & n52 ;
  assign n54 = ~n14 & n53 ;
  assign n55 = n17 & n53 ;
  assign n56 = n20 & n53 ;
  assign n57 = n22 & n53 ;
  assign n58 = n25 & n53 ;
  assign n59 = n28 & n53 ;
  assign n60 = n30 & n53 ;
  assign n61 = n32 & n53 ;
  assign n62 = n35 & n53 ;
  assign n63 = n37 & n53 ;
  assign n64 = n40 & n53 ;
  assign n65 = n42 & n53 ;
  assign n66 = n44 & n53 ;
  assign n67 = n46 & n53 ;
  assign n68 = n48 & n53 ;
  assign n69 = n50 & n53 ;
  assign n70 = ~x4 & x5 ;
  assign n71 = n10 & n70 ;
  assign n72 = ~n14 & n71 ;
  assign n73 = n17 & n71 ;
  assign n74 = n20 & n71 ;
  assign n75 = n22 & n71 ;
  assign n76 = n25 & n71 ;
  assign n77 = n28 & n71 ;
  assign n78 = n30 & n71 ;
  assign n79 = n32 & n71 ;
  assign n80 = n35 & n71 ;
  assign n81 = n37 & n71 ;
  assign n82 = n40 & n71 ;
  assign n83 = n42 & n71 ;
  assign n84 = n44 & n71 ;
  assign n85 = n46 & n71 ;
  assign n86 = n48 & n71 ;
  assign n87 = n50 & n71 ;
  assign n88 = x4 & x5 ;
  assign n89 = n10 & n88 ;
  assign n90 = ~n14 & n89 ;
  assign n91 = n17 & n89 ;
  assign n92 = n20 & n89 ;
  assign n93 = n22 & n89 ;
  assign n94 = n25 & n89 ;
  assign n95 = n28 & n89 ;
  assign n96 = n30 & n89 ;
  assign n97 = n32 & n89 ;
  assign n98 = n35 & n89 ;
  assign n99 = n37 & n89 ;
  assign n100 = n40 & n89 ;
  assign n101 = n42 & n89 ;
  assign n102 = n44 & n89 ;
  assign n103 = n46 & n89 ;
  assign n104 = n48 & n89 ;
  assign n105 = n50 & n89 ;
  assign n106 = x6 & x7 ;
  assign n107 = ~n9 & n106 ;
  assign n108 = ~n14 & n107 ;
  assign n109 = n17 & n107 ;
  assign n110 = n20 & n107 ;
  assign n111 = n22 & n107 ;
  assign n112 = n25 & n107 ;
  assign n113 = n28 & n107 ;
  assign n114 = n30 & n107 ;
  assign n115 = n32 & n107 ;
  assign n116 = n35 & n107 ;
  assign n117 = n37 & n107 ;
  assign n118 = n40 & n107 ;
  assign n119 = n42 & n107 ;
  assign n120 = n44 & n107 ;
  assign n121 = n46 & n107 ;
  assign n122 = n48 & n107 ;
  assign n123 = n50 & n107 ;
  assign n124 = n52 & n106 ;
  assign n125 = ~n14 & n124 ;
  assign n126 = n17 & n124 ;
  assign n127 = n20 & n124 ;
  assign n128 = n22 & n124 ;
  assign n129 = n25 & n124 ;
  assign n130 = n28 & n124 ;
  assign n131 = n30 & n124 ;
  assign n132 = n32 & n124 ;
  assign n133 = n35 & n124 ;
  assign n134 = n37 & n124 ;
  assign n135 = n40 & n124 ;
  assign n136 = n42 & n124 ;
  assign n137 = n44 & n124 ;
  assign n138 = n46 & n124 ;
  assign n139 = n48 & n124 ;
  assign n140 = n50 & n124 ;
  assign n141 = n70 & n106 ;
  assign n142 = ~n14 & n141 ;
  assign n143 = n17 & n141 ;
  assign n144 = n20 & n141 ;
  assign n145 = n22 & n141 ;
  assign n146 = n25 & n141 ;
  assign n147 = n28 & n141 ;
  assign n148 = n30 & n141 ;
  assign n149 = n32 & n141 ;
  assign n150 = n35 & n141 ;
  assign n151 = n37 & n141 ;
  assign n152 = n40 & n141 ;
  assign n153 = n42 & n141 ;
  assign n154 = n44 & n141 ;
  assign n155 = n46 & n141 ;
  assign n156 = n48 & n141 ;
  assign n157 = n50 & n141 ;
  assign n158 = n88 & n106 ;
  assign n159 = ~n14 & n158 ;
  assign n160 = n17 & n158 ;
  assign n161 = n20 & n158 ;
  assign n162 = n22 & n158 ;
  assign n163 = n25 & n158 ;
  assign n164 = n28 & n158 ;
  assign n165 = n30 & n158 ;
  assign n166 = n32 & n158 ;
  assign n167 = n35 & n158 ;
  assign n168 = n37 & n158 ;
  assign n169 = n40 & n158 ;
  assign n170 = n42 & n158 ;
  assign n171 = n44 & n158 ;
  assign n172 = n46 & n158 ;
  assign n173 = n48 & n158 ;
  assign n174 = n50 & n158 ;
  assign n175 = x6 | x7 ;
  assign n176 = n9 | n175 ;
  assign n177 = n14 | n176 ;
  assign n178 = n17 & ~n176 ;
  assign n179 = n20 & ~n176 ;
  assign n180 = n22 & ~n176 ;
  assign n181 = n25 & ~n176 ;
  assign n182 = n28 & ~n176 ;
  assign n183 = n30 & ~n176 ;
  assign n184 = n32 & ~n176 ;
  assign n185 = n35 & ~n176 ;
  assign n186 = n37 & ~n176 ;
  assign n187 = n40 & ~n176 ;
  assign n188 = n42 & ~n176 ;
  assign n189 = n44 & ~n176 ;
  assign n190 = n46 & ~n176 ;
  assign n191 = n48 & ~n176 ;
  assign n192 = n50 & ~n176 ;
  assign n193 = n52 & ~n175 ;
  assign n194 = ~n14 & n193 ;
  assign n195 = n17 & n193 ;
  assign n196 = n20 & n193 ;
  assign n197 = n22 & n193 ;
  assign n198 = n25 & n193 ;
  assign n199 = n28 & n193 ;
  assign n200 = n30 & n193 ;
  assign n201 = n32 & n193 ;
  assign n202 = n35 & n193 ;
  assign n203 = n37 & n193 ;
  assign n204 = n40 & n193 ;
  assign n205 = n42 & n193 ;
  assign n206 = n44 & n193 ;
  assign n207 = n46 & n193 ;
  assign n208 = n48 & n193 ;
  assign n209 = n50 & n193 ;
  assign n210 = n70 & ~n175 ;
  assign n211 = ~n14 & n210 ;
  assign n212 = n17 & n210 ;
  assign n213 = n20 & n210 ;
  assign n214 = n22 & n210 ;
  assign n215 = n25 & n210 ;
  assign n216 = n28 & n210 ;
  assign n217 = n30 & n210 ;
  assign n218 = n32 & n210 ;
  assign n219 = n35 & n210 ;
  assign n220 = n37 & n210 ;
  assign n221 = n40 & n210 ;
  assign n222 = n42 & n210 ;
  assign n223 = n44 & n210 ;
  assign n224 = n46 & n210 ;
  assign n225 = n48 & n210 ;
  assign n226 = n50 & n210 ;
  assign n227 = n88 & ~n175 ;
  assign n228 = ~n14 & n227 ;
  assign n229 = n17 & n227 ;
  assign n230 = n20 & n227 ;
  assign n231 = n22 & n227 ;
  assign n232 = n25 & n227 ;
  assign n233 = n28 & n227 ;
  assign n234 = n30 & n227 ;
  assign n235 = n32 & n227 ;
  assign n236 = n35 & n227 ;
  assign n237 = n37 & n227 ;
  assign n238 = n40 & n227 ;
  assign n239 = n42 & n227 ;
  assign n240 = n44 & n227 ;
  assign n241 = n46 & n227 ;
  assign n242 = n48 & n227 ;
  assign n243 = n50 & n227 ;
  assign n244 = x6 & ~x7 ;
  assign n245 = ~n9 & n244 ;
  assign n246 = ~n14 & n245 ;
  assign n247 = n17 & n245 ;
  assign n248 = n20 & n245 ;
  assign n249 = n22 & n245 ;
  assign n250 = n25 & n245 ;
  assign n251 = n28 & n245 ;
  assign n252 = n30 & n245 ;
  assign n253 = n32 & n245 ;
  assign n254 = n35 & n245 ;
  assign n255 = n37 & n245 ;
  assign n256 = n40 & n245 ;
  assign n257 = n42 & n245 ;
  assign n258 = n44 & n245 ;
  assign n259 = n46 & n245 ;
  assign n260 = n48 & n245 ;
  assign n261 = n50 & n245 ;
  assign n262 = n52 & n244 ;
  assign n263 = ~n14 & n262 ;
  assign n264 = n17 & n262 ;
  assign n265 = n20 & n262 ;
  assign n266 = n22 & n262 ;
  assign n267 = n25 & n262 ;
  assign n268 = n28 & n262 ;
  assign n269 = n30 & n262 ;
  assign n270 = n32 & n262 ;
  assign n271 = n35 & n262 ;
  assign n272 = n37 & n262 ;
  assign n273 = n40 & n262 ;
  assign n274 = n42 & n262 ;
  assign n275 = n44 & n262 ;
  assign n276 = n46 & n262 ;
  assign n277 = n48 & n262 ;
  assign n278 = n50 & n262 ;
  assign n279 = n70 & n244 ;
  assign n280 = ~n14 & n279 ;
  assign n281 = n17 & n279 ;
  assign n282 = n20 & n279 ;
  assign n283 = n22 & n279 ;
  assign n284 = n25 & n279 ;
  assign n285 = n28 & n279 ;
  assign n286 = n30 & n279 ;
  assign n287 = n32 & n279 ;
  assign n288 = n35 & n279 ;
  assign n289 = n37 & n279 ;
  assign n290 = n40 & n279 ;
  assign n291 = n42 & n279 ;
  assign n292 = n44 & n279 ;
  assign n293 = n46 & n279 ;
  assign n294 = n48 & n279 ;
  assign n295 = n50 & n279 ;
  assign n296 = n88 & n244 ;
  assign n297 = ~n14 & n296 ;
  assign n298 = n17 & n296 ;
  assign n299 = n20 & n296 ;
  assign n300 = n22 & n296 ;
  assign n301 = n25 & n296 ;
  assign n302 = n28 & n296 ;
  assign n303 = n30 & n296 ;
  assign n304 = n32 & n296 ;
  assign n305 = n35 & n296 ;
  assign n306 = n37 & n296 ;
  assign n307 = n40 & n296 ;
  assign n308 = n42 & n296 ;
  assign n309 = n44 & n296 ;
  assign n310 = n46 & n296 ;
  assign n311 = n48 & n296 ;
  assign n312 = n50 & n296 ;
  assign y0 = n15 ;
  assign y1 = n18 ;
  assign y2 = n21 ;
  assign y3 = n23 ;
  assign y4 = n26 ;
  assign y5 = n29 ;
  assign y6 = n31 ;
  assign y7 = n33 ;
  assign y8 = n36 ;
  assign y9 = n38 ;
  assign y10 = n41 ;
  assign y11 = n43 ;
  assign y12 = n45 ;
  assign y13 = n47 ;
  assign y14 = n49 ;
  assign y15 = n51 ;
  assign y16 = n54 ;
  assign y17 = n55 ;
  assign y18 = n56 ;
  assign y19 = n57 ;
  assign y20 = n58 ;
  assign y21 = n59 ;
  assign y22 = n60 ;
  assign y23 = n61 ;
  assign y24 = n62 ;
  assign y25 = n63 ;
  assign y26 = n64 ;
  assign y27 = n65 ;
  assign y28 = n66 ;
  assign y29 = n67 ;
  assign y30 = n68 ;
  assign y31 = n69 ;
  assign y32 = n72 ;
  assign y33 = n73 ;
  assign y34 = n74 ;
  assign y35 = n75 ;
  assign y36 = n76 ;
  assign y37 = n77 ;
  assign y38 = n78 ;
  assign y39 = n79 ;
  assign y40 = n80 ;
  assign y41 = n81 ;
  assign y42 = n82 ;
  assign y43 = n83 ;
  assign y44 = n84 ;
  assign y45 = n85 ;
  assign y46 = n86 ;
  assign y47 = n87 ;
  assign y48 = n90 ;
  assign y49 = n91 ;
  assign y50 = n92 ;
  assign y51 = n93 ;
  assign y52 = n94 ;
  assign y53 = n95 ;
  assign y54 = n96 ;
  assign y55 = n97 ;
  assign y56 = n98 ;
  assign y57 = n99 ;
  assign y58 = n100 ;
  assign y59 = n101 ;
  assign y60 = n102 ;
  assign y61 = n103 ;
  assign y62 = n104 ;
  assign y63 = n105 ;
  assign y64 = n108 ;
  assign y65 = n109 ;
  assign y66 = n110 ;
  assign y67 = n111 ;
  assign y68 = n112 ;
  assign y69 = n113 ;
  assign y70 = n114 ;
  assign y71 = n115 ;
  assign y72 = n116 ;
  assign y73 = n117 ;
  assign y74 = n118 ;
  assign y75 = n119 ;
  assign y76 = n120 ;
  assign y77 = n121 ;
  assign y78 = n122 ;
  assign y79 = n123 ;
  assign y80 = n125 ;
  assign y81 = n126 ;
  assign y82 = n127 ;
  assign y83 = n128 ;
  assign y84 = n129 ;
  assign y85 = n130 ;
  assign y86 = n131 ;
  assign y87 = n132 ;
  assign y88 = n133 ;
  assign y89 = n134 ;
  assign y90 = n135 ;
  assign y91 = n136 ;
  assign y92 = n137 ;
  assign y93 = n138 ;
  assign y94 = n139 ;
  assign y95 = n140 ;
  assign y96 = n142 ;
  assign y97 = n143 ;
  assign y98 = n144 ;
  assign y99 = n145 ;
  assign y100 = n146 ;
  assign y101 = n147 ;
  assign y102 = n148 ;
  assign y103 = n149 ;
  assign y104 = n150 ;
  assign y105 = n151 ;
  assign y106 = n152 ;
  assign y107 = n153 ;
  assign y108 = n154 ;
  assign y109 = n155 ;
  assign y110 = n156 ;
  assign y111 = n157 ;
  assign y112 = n159 ;
  assign y113 = n160 ;
  assign y114 = n161 ;
  assign y115 = n162 ;
  assign y116 = n163 ;
  assign y117 = n164 ;
  assign y118 = n165 ;
  assign y119 = n166 ;
  assign y120 = n167 ;
  assign y121 = n168 ;
  assign y122 = n169 ;
  assign y123 = n170 ;
  assign y124 = n171 ;
  assign y125 = n172 ;
  assign y126 = n173 ;
  assign y127 = n174 ;
  assign y128 = ~n177 ;
  assign y129 = n178 ;
  assign y130 = n179 ;
  assign y131 = n180 ;
  assign y132 = n181 ;
  assign y133 = n182 ;
  assign y134 = n183 ;
  assign y135 = n184 ;
  assign y136 = n185 ;
  assign y137 = n186 ;
  assign y138 = n187 ;
  assign y139 = n188 ;
  assign y140 = n189 ;
  assign y141 = n190 ;
  assign y142 = n191 ;
  assign y143 = n192 ;
  assign y144 = n194 ;
  assign y145 = n195 ;
  assign y146 = n196 ;
  assign y147 = n197 ;
  assign y148 = n198 ;
  assign y149 = n199 ;
  assign y150 = n200 ;
  assign y151 = n201 ;
  assign y152 = n202 ;
  assign y153 = n203 ;
  assign y154 = n204 ;
  assign y155 = n205 ;
  assign y156 = n206 ;
  assign y157 = n207 ;
  assign y158 = n208 ;
  assign y159 = n209 ;
  assign y160 = n211 ;
  assign y161 = n212 ;
  assign y162 = n213 ;
  assign y163 = n214 ;
  assign y164 = n215 ;
  assign y165 = n216 ;
  assign y166 = n217 ;
  assign y167 = n218 ;
  assign y168 = n219 ;
  assign y169 = n220 ;
  assign y170 = n221 ;
  assign y171 = n222 ;
  assign y172 = n223 ;
  assign y173 = n224 ;
  assign y174 = n225 ;
  assign y175 = n226 ;
  assign y176 = n228 ;
  assign y177 = n229 ;
  assign y178 = n230 ;
  assign y179 = n231 ;
  assign y180 = n232 ;
  assign y181 = n233 ;
  assign y182 = n234 ;
  assign y183 = n235 ;
  assign y184 = n236 ;
  assign y185 = n237 ;
  assign y186 = n238 ;
  assign y187 = n239 ;
  assign y188 = n240 ;
  assign y189 = n241 ;
  assign y190 = n242 ;
  assign y191 = n243 ;
  assign y192 = n246 ;
  assign y193 = n247 ;
  assign y194 = n248 ;
  assign y195 = n249 ;
  assign y196 = n250 ;
  assign y197 = n251 ;
  assign y198 = n252 ;
  assign y199 = n253 ;
  assign y200 = n254 ;
  assign y201 = n255 ;
  assign y202 = n256 ;
  assign y203 = n257 ;
  assign y204 = n258 ;
  assign y205 = n259 ;
  assign y206 = n260 ;
  assign y207 = n261 ;
  assign y208 = n263 ;
  assign y209 = n264 ;
  assign y210 = n265 ;
  assign y211 = n266 ;
  assign y212 = n267 ;
  assign y213 = n268 ;
  assign y214 = n269 ;
  assign y215 = n270 ;
  assign y216 = n271 ;
  assign y217 = n272 ;
  assign y218 = n273 ;
  assign y219 = n274 ;
  assign y220 = n275 ;
  assign y221 = n276 ;
  assign y222 = n277 ;
  assign y223 = n278 ;
  assign y224 = n280 ;
  assign y225 = n281 ;
  assign y226 = n282 ;
  assign y227 = n283 ;
  assign y228 = n284 ;
  assign y229 = n285 ;
  assign y230 = n286 ;
  assign y231 = n287 ;
  assign y232 = n288 ;
  assign y233 = n289 ;
  assign y234 = n290 ;
  assign y235 = n291 ;
  assign y236 = n292 ;
  assign y237 = n293 ;
  assign y238 = n294 ;
  assign y239 = n295 ;
  assign y240 = n297 ;
  assign y241 = n298 ;
  assign y242 = n299 ;
  assign y243 = n300 ;
  assign y244 = n301 ;
  assign y245 = n302 ;
  assign y246 = n303 ;
  assign y247 = n304 ;
  assign y248 = n305 ;
  assign y249 = n306 ;
  assign y250 = n307 ;
  assign y251 = n308 ;
  assign y252 = n309 ;
  assign y253 = n310 ;
  assign y254 = n311 ;
  assign y255 = n312 ;
endmodule
