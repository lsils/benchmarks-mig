module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 ;
  assign n513 = x127 & x255 ;
  assign n514 = x368 & ~x496 ;
  assign n515 = ( x369 & ~x497 ) | ( x369 & n514 ) | ( ~x497 & n514 ) ;
  assign n516 = x342 & ~x470 ;
  assign n517 = ( x343 & ~x471 ) | ( x343 & n516 ) | ( ~x471 & n516 ) ;
  assign n518 = ( x344 & ~x472 ) | ( x344 & n517 ) | ( ~x472 & n517 ) ;
  assign n519 = ~x342 & x470 ;
  assign n520 = ~x341 & x469 ;
  assign n521 = ~x344 & x472 ;
  assign n522 = n520 | n521 ;
  assign n523 = n519 & ~n522 ;
  assign n524 = ~x343 & x471 ;
  assign n525 = ( n522 & ~n523 ) | ( n522 & n524 ) | ( ~n523 & n524 ) ;
  assign n526 = ( ~n518 & n523 ) | ( ~n518 & n525 ) | ( n523 & n525 ) ;
  assign n527 = x292 & ~x420 ;
  assign n528 = ( x293 & ~x421 ) | ( x293 & n527 ) | ( ~x421 & n527 ) ;
  assign n529 = ~x284 & x412 ;
  assign n530 = ~x290 & x418 ;
  assign n531 = ~x285 & x413 ;
  assign n532 = ( ~n529 & n530 ) | ( ~n529 & n531 ) | ( n530 & n531 ) ;
  assign n533 = n529 | n532 ;
  assign n534 = ~x287 & x415 ;
  assign n535 = ~x286 & x414 ;
  assign n536 = ~x288 & x416 ;
  assign n537 = ~x289 & x417 ;
  assign n538 = ( ~n534 & n536 ) | ( ~n534 & n537 ) | ( n536 & n537 ) ;
  assign n539 = ( ~n534 & n535 ) | ( ~n534 & n538 ) | ( n535 & n538 ) ;
  assign n540 = n534 | n539 ;
  assign n541 = n533 | n540 ;
  assign n542 = x256 & ~x384 ;
  assign n543 = ( x257 & ~x385 ) | ( x257 & n542 ) | ( ~x385 & n542 ) ;
  assign n544 = ( x258 & ~x386 ) | ( x258 & n543 ) | ( ~x386 & n543 ) ;
  assign n545 = ( x259 & ~x387 ) | ( x259 & n544 ) | ( ~x387 & n544 ) ;
  assign n546 = ( x260 & ~x388 ) | ( x260 & n545 ) | ( ~x388 & n545 ) ;
  assign n547 = ( x261 & ~x389 ) | ( x261 & n546 ) | ( ~x389 & n546 ) ;
  assign n548 = ( x262 & ~x390 ) | ( x262 & n547 ) | ( ~x390 & n547 ) ;
  assign n549 = ( x263 & ~x391 ) | ( x263 & n548 ) | ( ~x391 & n548 ) ;
  assign n550 = ( x264 & ~x392 ) | ( x264 & n549 ) | ( ~x392 & n549 ) ;
  assign n551 = ( x265 & ~x393 ) | ( x265 & n550 ) | ( ~x393 & n550 ) ;
  assign n552 = ( x266 & ~x394 ) | ( x266 & n551 ) | ( ~x394 & n551 ) ;
  assign n553 = ( x267 & ~x395 ) | ( x267 & n552 ) | ( ~x395 & n552 ) ;
  assign n554 = ( x268 & ~x396 ) | ( x268 & n553 ) | ( ~x396 & n553 ) ;
  assign n555 = ( x269 & ~x397 ) | ( x269 & n554 ) | ( ~x397 & n554 ) ;
  assign n556 = ( x270 & ~x398 ) | ( x270 & n555 ) | ( ~x398 & n555 ) ;
  assign n557 = ( x271 & ~x399 ) | ( x271 & n556 ) | ( ~x399 & n556 ) ;
  assign n558 = ( x272 & ~x400 ) | ( x272 & n557 ) | ( ~x400 & n557 ) ;
  assign n559 = ( x273 & ~x401 ) | ( x273 & n558 ) | ( ~x401 & n558 ) ;
  assign n560 = ( x274 & ~x402 ) | ( x274 & n559 ) | ( ~x402 & n559 ) ;
  assign n561 = ( x275 & ~x403 ) | ( x275 & n560 ) | ( ~x403 & n560 ) ;
  assign n562 = ( x276 & ~x404 ) | ( x276 & n561 ) | ( ~x404 & n561 ) ;
  assign n563 = ( x277 & ~x405 ) | ( x277 & n562 ) | ( ~x405 & n562 ) ;
  assign n564 = ( x278 & ~x406 ) | ( x278 & n563 ) | ( ~x406 & n563 ) ;
  assign n565 = ( x279 & ~x407 ) | ( x279 & n564 ) | ( ~x407 & n564 ) ;
  assign n566 = ( x280 & ~x408 ) | ( x280 & n565 ) | ( ~x408 & n565 ) ;
  assign n567 = ~x283 & x411 ;
  assign n568 = ~x282 & x410 ;
  assign n569 = ~x281 & x409 ;
  assign n570 = ( ~n567 & n568 ) | ( ~n567 & n569 ) | ( n568 & n569 ) ;
  assign n571 = n567 | n570 ;
  assign n572 = n566 & ~n571 ;
  assign n573 = x281 & ~x409 ;
  assign n574 = ( x282 & ~x410 ) | ( x282 & n573 ) | ( ~x410 & n573 ) ;
  assign n575 = ( x283 & ~x411 ) | ( x283 & n574 ) | ( ~x411 & n574 ) ;
  assign n576 = ( x284 & ~x412 ) | ( x284 & n575 ) | ( ~x412 & n575 ) ;
  assign n577 = ~n541 & n576 ;
  assign n578 = ( ~n541 & n572 ) | ( ~n541 & n577 ) | ( n572 & n577 ) ;
  assign n579 = x285 & ~x413 ;
  assign n580 = ( x286 & ~x414 ) | ( x286 & n579 ) | ( ~x414 & n579 ) ;
  assign n581 = ( x287 & ~x415 ) | ( x287 & n580 ) | ( ~x415 & n580 ) ;
  assign n582 = ( x288 & ~x416 ) | ( x288 & n581 ) | ( ~x416 & n581 ) ;
  assign n583 = ( x289 & ~x417 ) | ( x289 & n582 ) | ( ~x417 & n582 ) ;
  assign n584 = ( x290 & ~x418 ) | ( x290 & n583 ) | ( ~x418 & n583 ) ;
  assign n585 = n578 | n584 ;
  assign n586 = ( x291 & ~x419 ) | ( x291 & n585 ) | ( ~x419 & n585 ) ;
  assign n587 = ~x292 & x420 ;
  assign n588 = ( ~x293 & x421 ) | ( ~x293 & n587 ) | ( x421 & n587 ) ;
  assign n589 = ( n528 & n586 ) | ( n528 & ~n588 ) | ( n586 & ~n588 ) ;
  assign n590 = ( x294 & ~x422 ) | ( x294 & n589 ) | ( ~x422 & n589 ) ;
  assign n591 = ( x295 & ~x423 ) | ( x295 & n590 ) | ( ~x423 & n590 ) ;
  assign n592 = ( x296 & ~x424 ) | ( x296 & n591 ) | ( ~x424 & n591 ) ;
  assign n593 = ( x297 & ~x425 ) | ( x297 & n592 ) | ( ~x425 & n592 ) ;
  assign n594 = ( x298 & ~x426 ) | ( x298 & n593 ) | ( ~x426 & n593 ) ;
  assign n595 = ( x299 & ~x427 ) | ( x299 & n594 ) | ( ~x427 & n594 ) ;
  assign n596 = ( x300 & ~x428 ) | ( x300 & n595 ) | ( ~x428 & n595 ) ;
  assign n597 = ( x301 & ~x429 ) | ( x301 & n596 ) | ( ~x429 & n596 ) ;
  assign n598 = ~x307 & x435 ;
  assign n599 = ~x303 & x431 ;
  assign n600 = ~x309 & x437 ;
  assign n601 = ~x304 & x432 ;
  assign n602 = ( ~n598 & n600 ) | ( ~n598 & n601 ) | ( n600 & n601 ) ;
  assign n603 = ( ~n598 & n599 ) | ( ~n598 & n602 ) | ( n599 & n602 ) ;
  assign n604 = n598 | n603 ;
  assign n605 = x303 & ~x431 ;
  assign n606 = ~x302 & x430 ;
  assign n607 = ~n605 & n606 ;
  assign n608 = ~x308 & x436 ;
  assign n609 = ~x305 & x433 ;
  assign n610 = n608 | n609 ;
  assign n611 = n607 | n610 ;
  assign n612 = ~x311 & x439 ;
  assign n613 = ~x306 & x434 ;
  assign n614 = ~x310 & x438 ;
  assign n615 = ( ~n612 & n613 ) | ( ~n612 & n614 ) | ( n613 & n614 ) ;
  assign n616 = n612 | n615 ;
  assign n617 = n611 | n616 ;
  assign n618 = n604 | n617 ;
  assign n619 = x302 & ~x430 ;
  assign n620 = n605 | n619 ;
  assign n621 = ~n618 & n620 ;
  assign n622 = ( n597 & ~n618 ) | ( n597 & n621 ) | ( ~n618 & n621 ) ;
  assign n623 = x304 & ~x432 ;
  assign n624 = ( x305 & ~x433 ) | ( x305 & n623 ) | ( ~x433 & n623 ) ;
  assign n625 = ( x306 & ~x434 ) | ( x306 & n624 ) | ( ~x434 & n624 ) ;
  assign n626 = ( x307 & ~x435 ) | ( x307 & n625 ) | ( ~x435 & n625 ) ;
  assign n627 = ( x308 & ~x436 ) | ( x308 & n626 ) | ( ~x436 & n626 ) ;
  assign n628 = ( x309 & ~x437 ) | ( x309 & n627 ) | ( ~x437 & n627 ) ;
  assign n629 = ( x310 & ~x438 ) | ( x310 & n628 ) | ( ~x438 & n628 ) ;
  assign n630 = ( x311 & ~x439 ) | ( x311 & n629 ) | ( ~x439 & n629 ) ;
  assign n631 = n622 | n630 ;
  assign n632 = ( x312 & ~x440 ) | ( x312 & n631 ) | ( ~x440 & n631 ) ;
  assign n633 = ( x313 & ~x441 ) | ( x313 & n632 ) | ( ~x441 & n632 ) ;
  assign n634 = x315 & ~x443 ;
  assign n635 = x314 & ~x442 ;
  assign n636 = n634 | n635 ;
  assign n637 = n633 | n636 ;
  assign n638 = ~x323 & x451 ;
  assign n639 = ~x322 & x450 ;
  assign n640 = ~x315 & x443 ;
  assign n641 = ~x316 & x444 ;
  assign n642 = ( ~n638 & n640 ) | ( ~n638 & n641 ) | ( n640 & n641 ) ;
  assign n643 = ( ~n638 & n639 ) | ( ~n638 & n642 ) | ( n639 & n642 ) ;
  assign n644 = n638 | n643 ;
  assign n645 = ~x318 & x446 ;
  assign n646 = ~x317 & x445 ;
  assign n647 = ~x319 & x447 ;
  assign n648 = ( ~n645 & n646 ) | ( ~n645 & n647 ) | ( n646 & n647 ) ;
  assign n649 = n645 | n648 ;
  assign n650 = ~x314 & x442 ;
  assign n651 = n634 & n650 ;
  assign n652 = ( n649 & n650 ) | ( n649 & ~n651 ) | ( n650 & ~n651 ) ;
  assign n653 = n644 | n652 ;
  assign n654 = ~x320 & x448 ;
  assign n655 = ( ~x321 & x449 ) | ( ~x321 & n654 ) | ( x449 & n654 ) ;
  assign n656 = x322 & ~x450 ;
  assign n657 = n655 & n656 ;
  assign n658 = ( n653 & n655 ) | ( n653 & ~n657 ) | ( n655 & ~n657 ) ;
  assign n659 = n637 & ~n658 ;
  assign n660 = x316 & ~x444 ;
  assign n661 = ( x317 & ~x445 ) | ( x317 & n660 ) | ( ~x445 & n660 ) ;
  assign n662 = ( x318 & ~x446 ) | ( x318 & n661 ) | ( ~x446 & n661 ) ;
  assign n663 = ( x319 & ~x447 ) | ( x319 & n662 ) | ( ~x447 & n662 ) ;
  assign n664 = ( x320 & ~x448 ) | ( x320 & n663 ) | ( ~x448 & n663 ) ;
  assign n665 = ( x321 & ~x449 ) | ( x321 & n664 ) | ( ~x449 & n664 ) ;
  assign n666 = ( x322 & ~x450 ) | ( x322 & n665 ) | ( ~x450 & n665 ) ;
  assign n667 = ( x323 & ~x451 ) | ( x323 & n666 ) | ( ~x451 & n666 ) ;
  assign n668 = n659 | n667 ;
  assign n669 = ( x324 & ~x452 ) | ( x324 & n668 ) | ( ~x452 & n668 ) ;
  assign n670 = ( x325 & ~x453 ) | ( x325 & n669 ) | ( ~x453 & n669 ) ;
  assign n671 = ( x326 & ~x454 ) | ( x326 & n670 ) | ( ~x454 & n670 ) ;
  assign n672 = ( x327 & ~x455 ) | ( x327 & n671 ) | ( ~x455 & n671 ) ;
  assign n673 = ( x328 & ~x456 ) | ( x328 & n672 ) | ( ~x456 & n672 ) ;
  assign n674 = ( x329 & ~x457 ) | ( x329 & n673 ) | ( ~x457 & n673 ) ;
  assign n675 = ( x330 & ~x458 ) | ( x330 & n674 ) | ( ~x458 & n674 ) ;
  assign n676 = ( x331 & ~x459 ) | ( x331 & n675 ) | ( ~x459 & n675 ) ;
  assign n677 = ( x332 & ~x460 ) | ( x332 & n676 ) | ( ~x460 & n676 ) ;
  assign n678 = ( x333 & ~x461 ) | ( x333 & n677 ) | ( ~x461 & n677 ) ;
  assign n679 = ( x334 & ~x462 ) | ( x334 & n678 ) | ( ~x462 & n678 ) ;
  assign n680 = ( x335 & ~x463 ) | ( x335 & n679 ) | ( ~x463 & n679 ) ;
  assign n681 = ( x336 & ~x464 ) | ( x336 & n680 ) | ( ~x464 & n680 ) ;
  assign n682 = ( x337 & ~x465 ) | ( x337 & n681 ) | ( ~x465 & n681 ) ;
  assign n683 = ~x339 & x467 ;
  assign n684 = ~x340 & x468 ;
  assign n685 = ~x338 & x466 ;
  assign n686 = ( ~n683 & n684 ) | ( ~n683 & n685 ) | ( n684 & n685 ) ;
  assign n687 = n683 | n686 ;
  assign n688 = n682 & ~n687 ;
  assign n689 = x338 & ~x466 ;
  assign n690 = ( x339 & ~x467 ) | ( x339 & n689 ) | ( ~x467 & n689 ) ;
  assign n691 = ( x340 & ~x468 ) | ( x340 & n690 ) | ( ~x468 & n690 ) ;
  assign n692 = ( x341 & ~x469 ) | ( x341 & n691 ) | ( ~x469 & n691 ) ;
  assign n693 = ( ~n518 & n688 ) | ( ~n518 & n692 ) | ( n688 & n692 ) ;
  assign n694 = ( n518 & ~n526 ) | ( n518 & n693 ) | ( ~n526 & n693 ) ;
  assign n695 = ( x345 & ~x473 ) | ( x345 & n694 ) | ( ~x473 & n694 ) ;
  assign n696 = ( x346 & ~x474 ) | ( x346 & n695 ) | ( ~x474 & n695 ) ;
  assign n697 = ( x347 & ~x475 ) | ( x347 & n696 ) | ( ~x475 & n696 ) ;
  assign n698 = ( x348 & ~x476 ) | ( x348 & n697 ) | ( ~x476 & n697 ) ;
  assign n699 = ( x349 & ~x477 ) | ( x349 & n698 ) | ( ~x477 & n698 ) ;
  assign n700 = ( x350 & ~x478 ) | ( x350 & n699 ) | ( ~x478 & n699 ) ;
  assign n701 = ( x351 & ~x479 ) | ( x351 & n700 ) | ( ~x479 & n700 ) ;
  assign n702 = ( x352 & ~x480 ) | ( x352 & n701 ) | ( ~x480 & n701 ) ;
  assign n703 = ( x353 & ~x481 ) | ( x353 & n702 ) | ( ~x481 & n702 ) ;
  assign n704 = ( x354 & ~x482 ) | ( x354 & n703 ) | ( ~x482 & n703 ) ;
  assign n705 = ( x355 & ~x483 ) | ( x355 & n704 ) | ( ~x483 & n704 ) ;
  assign n706 = ( x356 & ~x484 ) | ( x356 & n705 ) | ( ~x484 & n705 ) ;
  assign n707 = ( x357 & ~x485 ) | ( x357 & n706 ) | ( ~x485 & n706 ) ;
  assign n708 = ( x358 & ~x486 ) | ( x358 & n707 ) | ( ~x486 & n707 ) ;
  assign n709 = ( x359 & ~x487 ) | ( x359 & n708 ) | ( ~x487 & n708 ) ;
  assign n710 = ( x360 & ~x488 ) | ( x360 & n709 ) | ( ~x488 & n709 ) ;
  assign n711 = ( x361 & ~x489 ) | ( x361 & n710 ) | ( ~x489 & n710 ) ;
  assign n712 = ( x362 & ~x490 ) | ( x362 & n711 ) | ( ~x490 & n711 ) ;
  assign n713 = ( x363 & ~x491 ) | ( x363 & n712 ) | ( ~x491 & n712 ) ;
  assign n714 = ( x364 & ~x492 ) | ( x364 & n713 ) | ( ~x492 & n713 ) ;
  assign n715 = ( x365 & ~x493 ) | ( x365 & n714 ) | ( ~x493 & n714 ) ;
  assign n716 = ( x366 & ~x494 ) | ( x366 & n715 ) | ( ~x494 & n715 ) ;
  assign n717 = ( x367 & ~x495 ) | ( x367 & n716 ) | ( ~x495 & n716 ) ;
  assign n718 = ~x368 & x496 ;
  assign n719 = ( ~x369 & x497 ) | ( ~x369 & n718 ) | ( x497 & n718 ) ;
  assign n720 = ( n515 & n717 ) | ( n515 & ~n719 ) | ( n717 & ~n719 ) ;
  assign n721 = ( x370 & ~x498 ) | ( x370 & n720 ) | ( ~x498 & n720 ) ;
  assign n722 = ( x371 & ~x499 ) | ( x371 & n721 ) | ( ~x499 & n721 ) ;
  assign n723 = ( x372 & ~x500 ) | ( x372 & n722 ) | ( ~x500 & n722 ) ;
  assign n724 = ( x373 & ~x501 ) | ( x373 & n723 ) | ( ~x501 & n723 ) ;
  assign n725 = ( x374 & ~x502 ) | ( x374 & n724 ) | ( ~x502 & n724 ) ;
  assign n726 = ( x375 & ~x503 ) | ( x375 & n725 ) | ( ~x503 & n725 ) ;
  assign n727 = ( x376 & ~x504 ) | ( x376 & n726 ) | ( ~x504 & n726 ) ;
  assign n728 = ( x377 & ~x505 ) | ( x377 & n727 ) | ( ~x505 & n727 ) ;
  assign n729 = ( x378 & ~x506 ) | ( x378 & n728 ) | ( ~x506 & n728 ) ;
  assign n730 = ( x379 & ~x507 ) | ( x379 & n729 ) | ( ~x507 & n729 ) ;
  assign n731 = ~x380 & x508 ;
  assign n732 = ( ~x381 & x509 ) | ( ~x381 & n731 ) | ( x509 & n731 ) ;
  assign n733 = x380 & ~x508 ;
  assign n734 = ( x381 & ~x509 ) | ( x381 & n733 ) | ( ~x509 & n733 ) ;
  assign n735 = ( n730 & ~n732 ) | ( n730 & n734 ) | ( ~n732 & n734 ) ;
  assign n736 = ( x382 & ~x510 ) | ( x382 & n735 ) | ( ~x510 & n735 ) ;
  assign n737 = ( ~x383 & x511 ) | ( ~x383 & n736 ) | ( x511 & n736 ) ;
  assign n738 = x370 & n737 ;
  assign n739 = x498 & ~n737 ;
  assign n740 = n738 | n739 ;
  assign n741 = x124 & ~x252 ;
  assign n742 = ( x125 & ~x253 ) | ( x125 & n741 ) | ( ~x253 & n741 ) ;
  assign n743 = ( x126 & ~x254 ) | ( x126 & n742 ) | ( ~x254 & n742 ) ;
  assign n744 = ( ~x127 & x255 ) | ( ~x127 & n743 ) | ( x255 & n743 ) ;
  assign n745 = ~x99 & x227 ;
  assign n746 = ~x103 & x231 ;
  assign n747 = ~x100 & x228 ;
  assign n748 = ( ~n745 & n746 ) | ( ~n745 & n747 ) | ( n746 & n747 ) ;
  assign n749 = n745 | n748 ;
  assign n750 = ~x101 & x229 ;
  assign n751 = ~x102 & x230 ;
  assign n752 = ( ~n749 & n750 ) | ( ~n749 & n751 ) | ( n750 & n751 ) ;
  assign n753 = n749 | n752 ;
  assign n754 = ~x105 & x233 ;
  assign n755 = ~x106 & x234 ;
  assign n756 = n754 | n755 ;
  assign n757 = ~x104 & x232 ;
  assign n758 = ( ~n753 & n756 ) | ( ~n753 & n757 ) | ( n756 & n757 ) ;
  assign n759 = n753 | n758 ;
  assign n760 = x66 & ~x194 ;
  assign n761 = ( x67 & ~x195 ) | ( x67 & n760 ) | ( ~x195 & n760 ) ;
  assign n762 = ( x68 & ~x196 ) | ( x68 & n761 ) | ( ~x196 & n761 ) ;
  assign n763 = ( x69 & ~x197 ) | ( x69 & n762 ) | ( ~x197 & n762 ) ;
  assign n764 = ( x70 & ~x198 ) | ( x70 & n763 ) | ( ~x198 & n763 ) ;
  assign n765 = ( x71 & ~x199 ) | ( x71 & n764 ) | ( ~x199 & n764 ) ;
  assign n766 = ( x72 & ~x200 ) | ( x72 & n765 ) | ( ~x200 & n765 ) ;
  assign n767 = ( x73 & ~x201 ) | ( x73 & n766 ) | ( ~x201 & n766 ) ;
  assign n768 = ( x74 & ~x202 ) | ( x74 & n767 ) | ( ~x202 & n767 ) ;
  assign n769 = ( x75 & ~x203 ) | ( x75 & n768 ) | ( ~x203 & n768 ) ;
  assign n770 = x65 & ~x193 ;
  assign n771 = x63 & ~x191 ;
  assign n772 = x64 & ~x192 ;
  assign n773 = ~x57 & x185 ;
  assign n774 = ( ~x58 & x186 ) | ( ~x58 & n773 ) | ( x186 & n773 ) ;
  assign n775 = x56 & ~x184 ;
  assign n776 = x57 & ~x185 ;
  assign n777 = ( x58 & ~x186 ) | ( x58 & n776 ) | ( ~x186 & n776 ) ;
  assign n778 = ( ~n774 & n775 ) | ( ~n774 & n777 ) | ( n775 & n777 ) ;
  assign n779 = ( x59 & ~x187 ) | ( x59 & n778 ) | ( ~x187 & n778 ) ;
  assign n780 = ( x60 & ~x188 ) | ( x60 & n779 ) | ( ~x188 & n779 ) ;
  assign n781 = ~x54 & x182 ;
  assign n782 = ~x53 & x181 ;
  assign n783 = ~x47 & x175 ;
  assign n784 = ~x48 & x176 ;
  assign n785 = ( ~n781 & n783 ) | ( ~n781 & n784 ) | ( n783 & n784 ) ;
  assign n786 = ( ~n781 & n782 ) | ( ~n781 & n785 ) | ( n782 & n785 ) ;
  assign n787 = n781 | n786 ;
  assign n788 = ~x50 & x178 ;
  assign n789 = ~x49 & x177 ;
  assign n790 = ~x52 & x180 ;
  assign n791 = ~x51 & x179 ;
  assign n792 = ( ~n788 & n790 ) | ( ~n788 & n791 ) | ( n790 & n791 ) ;
  assign n793 = ( ~n788 & n789 ) | ( ~n788 & n792 ) | ( n789 & n792 ) ;
  assign n794 = n788 | n793 ;
  assign n795 = n787 | n794 ;
  assign n796 = x0 & ~x128 ;
  assign n797 = ( x1 & ~x129 ) | ( x1 & n796 ) | ( ~x129 & n796 ) ;
  assign n798 = ( x2 & ~x130 ) | ( x2 & n797 ) | ( ~x130 & n797 ) ;
  assign n799 = ( x3 & ~x131 ) | ( x3 & n798 ) | ( ~x131 & n798 ) ;
  assign n800 = ( x4 & ~x132 ) | ( x4 & n799 ) | ( ~x132 & n799 ) ;
  assign n801 = ( x5 & ~x133 ) | ( x5 & n800 ) | ( ~x133 & n800 ) ;
  assign n802 = ( x6 & ~x134 ) | ( x6 & n801 ) | ( ~x134 & n801 ) ;
  assign n803 = ( x7 & ~x135 ) | ( x7 & n802 ) | ( ~x135 & n802 ) ;
  assign n804 = ( x8 & ~x136 ) | ( x8 & n803 ) | ( ~x136 & n803 ) ;
  assign n805 = ( x9 & ~x137 ) | ( x9 & n804 ) | ( ~x137 & n804 ) ;
  assign n806 = ( x10 & ~x138 ) | ( x10 & n805 ) | ( ~x138 & n805 ) ;
  assign n807 = ( x11 & ~x139 ) | ( x11 & n806 ) | ( ~x139 & n806 ) ;
  assign n808 = ( x12 & ~x140 ) | ( x12 & n807 ) | ( ~x140 & n807 ) ;
  assign n809 = ( x13 & ~x141 ) | ( x13 & n808 ) | ( ~x141 & n808 ) ;
  assign n810 = ( x14 & ~x142 ) | ( x14 & n809 ) | ( ~x142 & n809 ) ;
  assign n811 = ( x15 & ~x143 ) | ( x15 & n810 ) | ( ~x143 & n810 ) ;
  assign n812 = ( x16 & ~x144 ) | ( x16 & n811 ) | ( ~x144 & n811 ) ;
  assign n813 = ( x17 & ~x145 ) | ( x17 & n812 ) | ( ~x145 & n812 ) ;
  assign n814 = ( x18 & ~x146 ) | ( x18 & n813 ) | ( ~x146 & n813 ) ;
  assign n815 = ( x19 & ~x147 ) | ( x19 & n814 ) | ( ~x147 & n814 ) ;
  assign n816 = ( x20 & ~x148 ) | ( x20 & n815 ) | ( ~x148 & n815 ) ;
  assign n817 = ( x21 & ~x149 ) | ( x21 & n816 ) | ( ~x149 & n816 ) ;
  assign n818 = ( x22 & ~x150 ) | ( x22 & n817 ) | ( ~x150 & n817 ) ;
  assign n819 = ( x23 & ~x151 ) | ( x23 & n818 ) | ( ~x151 & n818 ) ;
  assign n820 = ( x24 & ~x152 ) | ( x24 & n819 ) | ( ~x152 & n819 ) ;
  assign n821 = ( x25 & ~x153 ) | ( x25 & n820 ) | ( ~x153 & n820 ) ;
  assign n822 = ( x26 & ~x154 ) | ( x26 & n821 ) | ( ~x154 & n821 ) ;
  assign n823 = ( x27 & ~x155 ) | ( x27 & n822 ) | ( ~x155 & n822 ) ;
  assign n824 = ( x28 & ~x156 ) | ( x28 & n823 ) | ( ~x156 & n823 ) ;
  assign n825 = ( x29 & ~x157 ) | ( x29 & n824 ) | ( ~x157 & n824 ) ;
  assign n826 = ( x30 & ~x158 ) | ( x30 & n825 ) | ( ~x158 & n825 ) ;
  assign n827 = ( x31 & ~x159 ) | ( x31 & n826 ) | ( ~x159 & n826 ) ;
  assign n828 = ( x32 & ~x160 ) | ( x32 & n827 ) | ( ~x160 & n827 ) ;
  assign n829 = ( x33 & ~x161 ) | ( x33 & n828 ) | ( ~x161 & n828 ) ;
  assign n830 = ( x34 & ~x162 ) | ( x34 & n829 ) | ( ~x162 & n829 ) ;
  assign n831 = ( x35 & ~x163 ) | ( x35 & n830 ) | ( ~x163 & n830 ) ;
  assign n832 = ( x36 & ~x164 ) | ( x36 & n831 ) | ( ~x164 & n831 ) ;
  assign n833 = ( x37 & ~x165 ) | ( x37 & n832 ) | ( ~x165 & n832 ) ;
  assign n834 = ( x38 & ~x166 ) | ( x38 & n833 ) | ( ~x166 & n833 ) ;
  assign n835 = ( x39 & ~x167 ) | ( x39 & n834 ) | ( ~x167 & n834 ) ;
  assign n836 = ( x40 & ~x168 ) | ( x40 & n835 ) | ( ~x168 & n835 ) ;
  assign n837 = ( x41 & ~x169 ) | ( x41 & n836 ) | ( ~x169 & n836 ) ;
  assign n838 = ( x42 & ~x170 ) | ( x42 & n837 ) | ( ~x170 & n837 ) ;
  assign n839 = ( x43 & ~x171 ) | ( x43 & n838 ) | ( ~x171 & n838 ) ;
  assign n840 = ( x44 & ~x172 ) | ( x44 & n839 ) | ( ~x172 & n839 ) ;
  assign n841 = ( x45 & ~x173 ) | ( x45 & n840 ) | ( ~x173 & n840 ) ;
  assign n842 = ( x46 & ~x174 ) | ( x46 & n841 ) | ( ~x174 & n841 ) ;
  assign n843 = ( x47 & ~x175 ) | ( x47 & n842 ) | ( ~x175 & n842 ) ;
  assign n844 = ~n795 & n843 ;
  assign n845 = x48 & ~x176 ;
  assign n846 = ( x49 & ~x177 ) | ( x49 & n845 ) | ( ~x177 & n845 ) ;
  assign n847 = ( x50 & ~x178 ) | ( x50 & n846 ) | ( ~x178 & n846 ) ;
  assign n848 = ( x51 & ~x179 ) | ( x51 & n847 ) | ( ~x179 & n847 ) ;
  assign n849 = ( x52 & ~x180 ) | ( x52 & n848 ) | ( ~x180 & n848 ) ;
  assign n850 = ( x53 & ~x181 ) | ( x53 & n849 ) | ( ~x181 & n849 ) ;
  assign n851 = ( x54 & ~x182 ) | ( x54 & n850 ) | ( ~x182 & n850 ) ;
  assign n852 = n844 | n851 ;
  assign n853 = ( x55 & ~x183 ) | ( x55 & n852 ) | ( ~x183 & n852 ) ;
  assign n854 = ~x60 & x188 ;
  assign n855 = ~x56 & x184 ;
  assign n856 = ~x59 & x187 ;
  assign n857 = ( ~n854 & n855 ) | ( ~n854 & n856 ) | ( n855 & n856 ) ;
  assign n858 = n854 | n857 ;
  assign n859 = n774 | n858 ;
  assign n860 = ~n780 & n859 ;
  assign n861 = ( n780 & n853 ) | ( n780 & ~n860 ) | ( n853 & ~n860 ) ;
  assign n862 = ( x61 & ~x189 ) | ( x61 & n861 ) | ( ~x189 & n861 ) ;
  assign n863 = ( x62 & ~x190 ) | ( x62 & n862 ) | ( ~x190 & n862 ) ;
  assign n864 = ( ~n771 & n772 ) | ( ~n771 & n863 ) | ( n772 & n863 ) ;
  assign n865 = ( ~n770 & n771 ) | ( ~n770 & n864 ) | ( n771 & n864 ) ;
  assign n866 = ~x63 & x191 ;
  assign n867 = ( ~x64 & x192 ) | ( ~x64 & n866 ) | ( x192 & n866 ) ;
  assign n868 = ~n770 & n867 ;
  assign n869 = ( n770 & n865 ) | ( n770 & ~n868 ) | ( n865 & ~n868 ) ;
  assign n870 = ~x72 & x200 ;
  assign n871 = ~x71 & x199 ;
  assign n872 = ~x74 & x202 ;
  assign n873 = ~x73 & x201 ;
  assign n874 = ( ~n870 & n872 ) | ( ~n870 & n873 ) | ( n872 & n873 ) ;
  assign n875 = ( ~n870 & n871 ) | ( ~n870 & n874 ) | ( n871 & n874 ) ;
  assign n876 = n870 | n875 ;
  assign n877 = ~x68 & x196 ;
  assign n878 = ~x67 & x195 ;
  assign n879 = ~x70 & x198 ;
  assign n880 = ~x69 & x197 ;
  assign n881 = ( ~n877 & n879 ) | ( ~n877 & n880 ) | ( n879 & n880 ) ;
  assign n882 = ( ~n877 & n878 ) | ( ~n877 & n881 ) | ( n878 & n881 ) ;
  assign n883 = n877 | n882 ;
  assign n884 = ~x75 & x203 ;
  assign n885 = ~x65 & x193 ;
  assign n886 = ~x66 & x194 ;
  assign n887 = ( ~n884 & n885 ) | ( ~n884 & n886 ) | ( n885 & n886 ) ;
  assign n888 = n884 | n887 ;
  assign n889 = ( ~n876 & n883 ) | ( ~n876 & n888 ) | ( n883 & n888 ) ;
  assign n890 = n876 | n889 ;
  assign n891 = n869 & ~n890 ;
  assign n892 = n769 | n891 ;
  assign n893 = ( x76 & ~x204 ) | ( x76 & n892 ) | ( ~x204 & n892 ) ;
  assign n894 = ( x77 & ~x205 ) | ( x77 & n893 ) | ( ~x205 & n893 ) ;
  assign n895 = ( x78 & ~x206 ) | ( x78 & n894 ) | ( ~x206 & n894 ) ;
  assign n896 = ( x79 & ~x207 ) | ( x79 & n895 ) | ( ~x207 & n895 ) ;
  assign n897 = ( x80 & ~x208 ) | ( x80 & n896 ) | ( ~x208 & n896 ) ;
  assign n898 = ( x81 & ~x209 ) | ( x81 & n897 ) | ( ~x209 & n897 ) ;
  assign n899 = ( x82 & ~x210 ) | ( x82 & n898 ) | ( ~x210 & n898 ) ;
  assign n900 = ( x83 & ~x211 ) | ( x83 & n899 ) | ( ~x211 & n899 ) ;
  assign n901 = ( x84 & ~x212 ) | ( x84 & n900 ) | ( ~x212 & n900 ) ;
  assign n902 = ( x85 & ~x213 ) | ( x85 & n901 ) | ( ~x213 & n901 ) ;
  assign n903 = ( x86 & ~x214 ) | ( x86 & n902 ) | ( ~x214 & n902 ) ;
  assign n904 = ( x87 & ~x215 ) | ( x87 & n903 ) | ( ~x215 & n903 ) ;
  assign n905 = ( x88 & ~x216 ) | ( x88 & n904 ) | ( ~x216 & n904 ) ;
  assign n906 = ( x89 & ~x217 ) | ( x89 & n905 ) | ( ~x217 & n905 ) ;
  assign n907 = ( x90 & ~x218 ) | ( x90 & n906 ) | ( ~x218 & n906 ) ;
  assign n908 = ( x91 & ~x219 ) | ( x91 & n907 ) | ( ~x219 & n907 ) ;
  assign n909 = ~x91 & x219 ;
  assign n910 = ~x95 & x223 ;
  assign n911 = ~x97 & x225 ;
  assign n912 = ~x92 & x220 ;
  assign n913 = ( ~n910 & n911 ) | ( ~n910 & n912 ) | ( n911 & n912 ) ;
  assign n914 = ( ~n909 & n910 ) | ( ~n909 & n913 ) | ( n910 & n913 ) ;
  assign n915 = ~x94 & x222 ;
  assign n916 = ~x93 & x221 ;
  assign n917 = ~x98 & x226 ;
  assign n918 = ~x96 & x224 ;
  assign n919 = ( ~n915 & n917 ) | ( ~n915 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ( ~n915 & n916 ) | ( ~n915 & n919 ) | ( n916 & n919 ) ;
  assign n921 = n915 | n920 ;
  assign n922 = n914 | n921 ;
  assign n923 = n908 & ~n922 ;
  assign n924 = x92 & ~x220 ;
  assign n925 = ( x93 & ~x221 ) | ( x93 & n924 ) | ( ~x221 & n924 ) ;
  assign n926 = ( x94 & ~x222 ) | ( x94 & n925 ) | ( ~x222 & n925 ) ;
  assign n927 = ( x95 & ~x223 ) | ( x95 & n926 ) | ( ~x223 & n926 ) ;
  assign n928 = ( x96 & ~x224 ) | ( x96 & n927 ) | ( ~x224 & n927 ) ;
  assign n929 = ( x97 & ~x225 ) | ( x97 & n928 ) | ( ~x225 & n928 ) ;
  assign n930 = ( x98 & ~x226 ) | ( x98 & n929 ) | ( ~x226 & n929 ) ;
  assign n931 = ( x99 & ~x227 ) | ( x99 & n930 ) | ( ~x227 & n930 ) ;
  assign n932 = ~n759 & n931 ;
  assign n933 = ( ~n759 & n923 ) | ( ~n759 & n932 ) | ( n923 & n932 ) ;
  assign n934 = x100 & ~x228 ;
  assign n935 = ( x101 & ~x229 ) | ( x101 & n934 ) | ( ~x229 & n934 ) ;
  assign n936 = ( x102 & ~x230 ) | ( x102 & n935 ) | ( ~x230 & n935 ) ;
  assign n937 = ( x103 & ~x231 ) | ( x103 & n936 ) | ( ~x231 & n936 ) ;
  assign n938 = ~n756 & n937 ;
  assign n939 = ( x104 & ~x232 ) | ( x104 & n938 ) | ( ~x232 & n938 ) ;
  assign n940 = ( x105 & ~x233 ) | ( x105 & n939 ) | ( ~x233 & n939 ) ;
  assign n941 = ( x106 & ~x234 ) | ( x106 & n940 ) | ( ~x234 & n940 ) ;
  assign n942 = n933 | n941 ;
  assign n943 = ( x107 & ~x235 ) | ( x107 & n942 ) | ( ~x235 & n942 ) ;
  assign n944 = ( x108 & ~x236 ) | ( x108 & n943 ) | ( ~x236 & n943 ) ;
  assign n945 = ( x109 & ~x237 ) | ( x109 & n944 ) | ( ~x237 & n944 ) ;
  assign n946 = ( x110 & ~x238 ) | ( x110 & n945 ) | ( ~x238 & n945 ) ;
  assign n947 = ( x111 & ~x239 ) | ( x111 & n946 ) | ( ~x239 & n946 ) ;
  assign n948 = ~x112 & x240 ;
  assign n949 = ( ~x113 & x241 ) | ( ~x113 & n948 ) | ( x241 & n948 ) ;
  assign n950 = x112 & ~x240 ;
  assign n951 = ( x113 & ~x241 ) | ( x113 & n950 ) | ( ~x241 & n950 ) ;
  assign n952 = ( n947 & ~n949 ) | ( n947 & n951 ) | ( ~n949 & n951 ) ;
  assign n953 = ( x114 & ~x242 ) | ( x114 & n952 ) | ( ~x242 & n952 ) ;
  assign n954 = ( x115 & ~x243 ) | ( x115 & n953 ) | ( ~x243 & n953 ) ;
  assign n955 = ( x116 & ~x244 ) | ( x116 & n954 ) | ( ~x244 & n954 ) ;
  assign n956 = ( x117 & ~x245 ) | ( x117 & n955 ) | ( ~x245 & n955 ) ;
  assign n957 = ( x118 & ~x246 ) | ( x118 & n956 ) | ( ~x246 & n956 ) ;
  assign n958 = ( x119 & ~x247 ) | ( x119 & n957 ) | ( ~x247 & n957 ) ;
  assign n959 = ( x120 & ~x248 ) | ( x120 & n958 ) | ( ~x248 & n958 ) ;
  assign n960 = ( x121 & ~x249 ) | ( x121 & n959 ) | ( ~x249 & n959 ) ;
  assign n961 = ( x122 & ~x250 ) | ( x122 & n960 ) | ( ~x250 & n960 ) ;
  assign n962 = ( x123 & ~x251 ) | ( x123 & n961 ) | ( ~x251 & n961 ) ;
  assign n963 = ~x125 & x253 ;
  assign n964 = ~x124 & x252 ;
  assign n965 = ~x126 & x254 ;
  assign n966 = ( ~n963 & n964 ) | ( ~n963 & n965 ) | ( n964 & n965 ) ;
  assign n967 = ( ~n743 & n963 ) | ( ~n743 & n966 ) | ( n963 & n966 ) ;
  assign n968 = ( x127 & ~x255 ) | ( x127 & n967 ) | ( ~x255 & n967 ) ;
  assign n969 = ( n744 & n962 ) | ( n744 & ~n968 ) | ( n962 & ~n968 ) ;
  assign n970 = ~x114 & n969 ;
  assign n971 = x242 & ~n969 ;
  assign n972 = ( n969 & ~n970 ) | ( n969 & n971 ) | ( ~n970 & n971 ) ;
  assign n973 = x369 & n737 ;
  assign n974 = x497 & ~n737 ;
  assign n975 = n973 | n974 ;
  assign n976 = x241 | n969 ;
  assign n977 = ~x113 & n969 ;
  assign n978 = n976 & ~n977 ;
  assign n979 = x368 & n737 ;
  assign n980 = x496 & ~n737 ;
  assign n981 = n979 | n980 ;
  assign n982 = x240 | n969 ;
  assign n983 = ~x112 & n969 ;
  assign n984 = n982 & ~n983 ;
  assign n985 = ~n981 & n984 ;
  assign n986 = ( ~n975 & n978 ) | ( ~n975 & n985 ) | ( n978 & n985 ) ;
  assign n987 = ( ~n740 & n972 ) | ( ~n740 & n986 ) | ( n972 & n986 ) ;
  assign n988 = x371 & n737 ;
  assign n989 = x499 & ~n737 ;
  assign n990 = n988 | n989 ;
  assign n991 = x243 | n969 ;
  assign n992 = ~x115 & n969 ;
  assign n993 = n991 & ~n992 ;
  assign n994 = ~n990 & n993 ;
  assign n995 = n987 | n994 ;
  assign n996 = x366 & n737 ;
  assign n997 = x494 & ~n737 ;
  assign n998 = x238 | n969 ;
  assign n999 = ~x110 & n969 ;
  assign n1000 = n998 & ~n999 ;
  assign n1001 = ( n996 & n997 ) | ( n996 & ~n1000 ) | ( n997 & ~n1000 ) ;
  assign n1002 = ~x365 & n737 ;
  assign n1003 = x493 | n737 ;
  assign n1004 = x237 | n969 ;
  assign n1005 = ~x109 & n969 ;
  assign n1006 = n1004 & ~n1005 ;
  assign n1007 = ( n1002 & n1003 ) | ( n1002 & ~n1006 ) | ( n1003 & ~n1006 ) ;
  assign n1008 = ( n1001 & ~n1002 ) | ( n1001 & n1007 ) | ( ~n1002 & n1007 ) ;
  assign n1009 = x489 & ~n737 ;
  assign n1010 = x361 & n737 ;
  assign n1011 = x233 | n969 ;
  assign n1012 = ~x105 & n969 ;
  assign n1013 = n1011 & ~n1012 ;
  assign n1014 = ( n1009 & n1010 ) | ( n1009 & ~n1013 ) | ( n1010 & ~n1013 ) ;
  assign n1015 = x488 & ~n737 ;
  assign n1016 = x360 & n737 ;
  assign n1017 = x232 | n969 ;
  assign n1018 = ~x104 & n969 ;
  assign n1019 = n1017 & ~n1018 ;
  assign n1020 = ( n1015 & n1016 ) | ( n1015 & ~n1019 ) | ( n1016 & ~n1019 ) ;
  assign n1021 = n1014 | n1020 ;
  assign n1022 = x490 & ~n737 ;
  assign n1023 = x362 & n737 ;
  assign n1024 = x234 | n969 ;
  assign n1025 = ~x106 & n969 ;
  assign n1026 = n1024 & ~n1025 ;
  assign n1027 = ( n1022 & n1023 ) | ( n1022 & ~n1026 ) | ( n1023 & ~n1026 ) ;
  assign n1028 = n1021 | n1027 ;
  assign n1029 = x364 & n737 ;
  assign n1030 = x492 & ~n737 ;
  assign n1031 = x236 | n969 ;
  assign n1032 = ~x108 & n969 ;
  assign n1033 = n1031 & ~n1032 ;
  assign n1034 = ( n1029 & n1030 ) | ( n1029 & ~n1033 ) | ( n1030 & ~n1033 ) ;
  assign n1035 = x363 & n737 ;
  assign n1036 = x491 & ~n737 ;
  assign n1037 = x235 | n969 ;
  assign n1038 = ~x107 & n969 ;
  assign n1039 = n1037 & ~n1038 ;
  assign n1040 = ( n1035 & n1036 ) | ( n1035 & ~n1039 ) | ( n1036 & ~n1039 ) ;
  assign n1041 = n1034 | n1040 ;
  assign n1042 = x358 & n737 ;
  assign n1043 = x486 & ~n737 ;
  assign n1044 = x230 | n969 ;
  assign n1045 = ~x102 & n969 ;
  assign n1046 = n1044 & ~n1045 ;
  assign n1047 = ( n1042 & n1043 ) | ( n1042 & ~n1046 ) | ( n1043 & ~n1046 ) ;
  assign n1048 = x487 & ~n737 ;
  assign n1049 = x359 & n737 ;
  assign n1050 = x231 | n969 ;
  assign n1051 = ~x103 & n969 ;
  assign n1052 = n1050 & ~n1051 ;
  assign n1053 = ( n1048 & n1049 ) | ( n1048 & ~n1052 ) | ( n1049 & ~n1052 ) ;
  assign n1054 = ( ~n1028 & n1047 ) | ( ~n1028 & n1053 ) | ( n1047 & n1053 ) ;
  assign n1055 = ( ~n1028 & n1041 ) | ( ~n1028 & n1054 ) | ( n1041 & n1054 ) ;
  assign n1056 = n1028 | n1055 ;
  assign n1057 = x485 | n737 ;
  assign n1058 = ~x357 & n737 ;
  assign n1059 = n1057 & ~n1058 ;
  assign n1060 = x229 | n969 ;
  assign n1061 = ~x101 & n969 ;
  assign n1062 = n1060 & ~n1061 ;
  assign n1063 = x219 | n969 ;
  assign n1064 = ~x91 & n969 ;
  assign n1065 = n1063 & ~n1064 ;
  assign n1066 = x347 & n737 ;
  assign n1067 = x475 & ~n737 ;
  assign n1068 = n1066 | n1067 ;
  assign n1069 = x218 | n969 ;
  assign n1070 = ~x90 & n969 ;
  assign n1071 = n1069 & ~n1070 ;
  assign n1072 = x474 & ~n737 ;
  assign n1073 = x346 & n737 ;
  assign n1074 = n1072 | n1073 ;
  assign n1075 = x217 | n969 ;
  assign n1076 = ~x89 & n969 ;
  assign n1077 = n1075 & ~n1076 ;
  assign n1078 = x473 & ~n737 ;
  assign n1079 = x345 & n737 ;
  assign n1080 = n1078 | n1079 ;
  assign n1081 = x216 | n969 ;
  assign n1082 = ~x88 & n969 ;
  assign n1083 = n1081 & ~n1082 ;
  assign n1084 = x472 & ~n737 ;
  assign n1085 = x344 & n737 ;
  assign n1086 = n1084 | n1085 ;
  assign n1087 = n1083 & ~n1086 ;
  assign n1088 = ( n1077 & ~n1080 ) | ( n1077 & n1087 ) | ( ~n1080 & n1087 ) ;
  assign n1089 = ( n1071 & ~n1074 ) | ( n1071 & n1088 ) | ( ~n1074 & n1088 ) ;
  assign n1090 = ( n1065 & ~n1068 ) | ( n1065 & n1089 ) | ( ~n1068 & n1089 ) ;
  assign n1091 = ( ~n1071 & n1072 ) | ( ~n1071 & n1073 ) | ( n1072 & n1073 ) ;
  assign n1092 = ( ~n1077 & n1078 ) | ( ~n1077 & n1079 ) | ( n1078 & n1079 ) ;
  assign n1093 = n1091 | n1092 ;
  assign n1094 = x471 & ~n737 ;
  assign n1095 = x342 & n737 ;
  assign n1096 = x470 & ~n737 ;
  assign n1097 = x214 | n969 ;
  assign n1098 = ~x86 & n969 ;
  assign n1099 = n1097 & ~n1098 ;
  assign n1100 = ( n1095 & n1096 ) | ( n1095 & ~n1099 ) | ( n1096 & ~n1099 ) ;
  assign n1101 = x343 & n737 ;
  assign n1102 = x215 | n969 ;
  assign n1103 = ~x87 & n969 ;
  assign n1104 = n1102 & ~n1103 ;
  assign n1105 = ( n1094 & ~n1101 ) | ( n1094 & n1104 ) | ( ~n1101 & n1104 ) ;
  assign n1106 = ( n1094 & n1100 ) | ( n1094 & ~n1105 ) | ( n1100 & ~n1105 ) ;
  assign n1107 = ~n1090 & n1106 ;
  assign n1108 = ( ~n1090 & n1093 ) | ( ~n1090 & n1107 ) | ( n1093 & n1107 ) ;
  assign n1109 = n1094 | n1101 ;
  assign n1110 = x341 & n737 ;
  assign n1111 = x469 & ~n737 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = x213 | n969 ;
  assign n1114 = ~x85 & n969 ;
  assign n1115 = n1113 & ~n1114 ;
  assign n1116 = ~n1112 & n1115 ;
  assign n1117 = n1095 | n1096 ;
  assign n1118 = n1099 | n1117 ;
  assign n1119 = ( n1116 & ~n1117 ) | ( n1116 & n1118 ) | ( ~n1117 & n1118 ) ;
  assign n1120 = ( n1104 & ~n1109 ) | ( n1104 & n1119 ) | ( ~n1109 & n1119 ) ;
  assign n1121 = n1112 & ~n1115 ;
  assign n1122 = x468 | n737 ;
  assign n1123 = ~x340 & n737 ;
  assign n1124 = n1122 & ~n1123 ;
  assign n1125 = x212 | n969 ;
  assign n1126 = ~x84 & n969 ;
  assign n1127 = n1125 & ~n1126 ;
  assign n1128 = x467 | n737 ;
  assign n1129 = ~x339 & n737 ;
  assign n1130 = n1128 & ~n1129 ;
  assign n1131 = x211 | n969 ;
  assign n1132 = ~x83 & n969 ;
  assign n1133 = n1131 & ~n1132 ;
  assign n1134 = x465 | n737 ;
  assign n1135 = ~x337 & n737 ;
  assign n1136 = n1134 & ~n1135 ;
  assign n1137 = x209 | n969 ;
  assign n1138 = ~x81 & n969 ;
  assign n1139 = n1137 & ~n1138 ;
  assign n1140 = x464 | n737 ;
  assign n1141 = ~x336 & n737 ;
  assign n1142 = n1140 & ~n1141 ;
  assign n1143 = x208 | n969 ;
  assign n1144 = ~x80 & n969 ;
  assign n1145 = n1143 & ~n1144 ;
  assign n1146 = x463 | n737 ;
  assign n1147 = ~x335 & n737 ;
  assign n1148 = n1146 & ~n1147 ;
  assign n1149 = x462 | n737 ;
  assign n1150 = ~x334 & n737 ;
  assign n1151 = n1149 & ~n1150 ;
  assign n1152 = x206 | n969 ;
  assign n1153 = ~x78 & n969 ;
  assign n1154 = n1152 & ~n1153 ;
  assign n1155 = x461 | n737 ;
  assign n1156 = ~x333 & n737 ;
  assign n1157 = n1155 & ~n1156 ;
  assign n1158 = x460 | n737 ;
  assign n1159 = ~x332 & n737 ;
  assign n1160 = n1158 & ~n1159 ;
  assign n1161 = x204 | n969 ;
  assign n1162 = ~x76 & n969 ;
  assign n1163 = n1161 & ~n1162 ;
  assign n1164 = x456 & ~n737 ;
  assign n1165 = x328 & n737 ;
  assign n1166 = x200 | n969 ;
  assign n1167 = ~x72 & n969 ;
  assign n1168 = n1166 & ~n1167 ;
  assign n1169 = ( n1164 & n1165 ) | ( n1164 & ~n1168 ) | ( n1165 & ~n1168 ) ;
  assign n1170 = x451 & ~n737 ;
  assign n1171 = x323 & n737 ;
  assign n1172 = x195 | n969 ;
  assign n1173 = ~x67 & n969 ;
  assign n1174 = n1172 & ~n1173 ;
  assign n1175 = ( n1170 & n1171 ) | ( n1170 & ~n1174 ) | ( n1171 & ~n1174 ) ;
  assign n1176 = n1169 | n1175 ;
  assign n1177 = x325 & n737 ;
  assign n1178 = x453 & ~n737 ;
  assign n1179 = x197 | n969 ;
  assign n1180 = ~x69 & n969 ;
  assign n1181 = n1179 & ~n1180 ;
  assign n1182 = ( n1177 & n1178 ) | ( n1177 & ~n1181 ) | ( n1178 & ~n1181 ) ;
  assign n1183 = x326 & n737 ;
  assign n1184 = x454 & ~n737 ;
  assign n1185 = x198 | n969 ;
  assign n1186 = ~x70 & n969 ;
  assign n1187 = n1185 & ~n1186 ;
  assign n1188 = ( n1183 & n1184 ) | ( n1183 & ~n1187 ) | ( n1184 & ~n1187 ) ;
  assign n1189 = n1182 | n1188 ;
  assign n1190 = x455 | n737 ;
  assign n1191 = x324 & n737 ;
  assign n1192 = x452 & ~n737 ;
  assign n1193 = x196 | n969 ;
  assign n1194 = ~x68 & n969 ;
  assign n1195 = n1193 & ~n1194 ;
  assign n1196 = ( n1191 & n1192 ) | ( n1191 & ~n1195 ) | ( n1192 & ~n1195 ) ;
  assign n1197 = ~x327 & n737 ;
  assign n1198 = ~x71 & n969 ;
  assign n1199 = x199 | n969 ;
  assign n1200 = ~n1198 & n1199 ;
  assign n1201 = ( n1190 & n1197 ) | ( n1190 & n1200 ) | ( n1197 & n1200 ) ;
  assign n1202 = ( n1190 & n1196 ) | ( n1190 & ~n1201 ) | ( n1196 & ~n1201 ) ;
  assign n1203 = x329 & n737 ;
  assign n1204 = x457 & ~n737 ;
  assign n1205 = x201 | n969 ;
  assign n1206 = ~x73 & n969 ;
  assign n1207 = n1205 & ~n1206 ;
  assign n1208 = ( n1203 & n1204 ) | ( n1203 & ~n1207 ) | ( n1204 & ~n1207 ) ;
  assign n1209 = ( ~n1176 & n1202 ) | ( ~n1176 & n1208 ) | ( n1202 & n1208 ) ;
  assign n1210 = ( ~n1176 & n1189 ) | ( ~n1176 & n1209 ) | ( n1189 & n1209 ) ;
  assign n1211 = n1176 | n1210 ;
  assign n1212 = x446 & ~n737 ;
  assign n1213 = x190 | n969 ;
  assign n1214 = ~x62 & n969 ;
  assign n1215 = n1213 & ~n1214 ;
  assign n1216 = x318 & n737 ;
  assign n1217 = x445 & ~n737 ;
  assign n1218 = x317 & n737 ;
  assign n1219 = n1217 | n1218 ;
  assign n1220 = x189 | n969 ;
  assign n1221 = ~x61 & n969 ;
  assign n1222 = n1220 & ~n1221 ;
  assign n1223 = x316 & n737 ;
  assign n1224 = x444 & ~n737 ;
  assign n1225 = n1223 | n1224 ;
  assign n1226 = x188 | n969 ;
  assign n1227 = ~x60 & n969 ;
  assign n1228 = n1226 & ~n1227 ;
  assign n1229 = x443 & ~n737 ;
  assign n1230 = x315 & n737 ;
  assign n1231 = n1229 | n1230 ;
  assign n1232 = x187 | n969 ;
  assign n1233 = ~x59 & n969 ;
  assign n1234 = n1232 & ~n1233 ;
  assign n1235 = x314 & n737 ;
  assign n1236 = x442 & ~n737 ;
  assign n1237 = n1235 | n1236 ;
  assign n1238 = x186 | n969 ;
  assign n1239 = ~x58 & n969 ;
  assign n1240 = n1238 & ~n1239 ;
  assign n1241 = x441 & ~n737 ;
  assign n1242 = x313 & n737 ;
  assign n1243 = n1241 | n1242 ;
  assign n1244 = x185 | n969 ;
  assign n1245 = ~x57 & n969 ;
  assign n1246 = n1244 & ~n1245 ;
  assign n1247 = x440 & ~n737 ;
  assign n1248 = x312 & n737 ;
  assign n1249 = n1247 | n1248 ;
  assign n1250 = x184 | n969 ;
  assign n1251 = ~x56 & n969 ;
  assign n1252 = n1250 & ~n1251 ;
  assign n1253 = ~n1249 & n1252 ;
  assign n1254 = ( ~n1243 & n1246 ) | ( ~n1243 & n1253 ) | ( n1246 & n1253 ) ;
  assign n1255 = ( ~n1237 & n1240 ) | ( ~n1237 & n1254 ) | ( n1240 & n1254 ) ;
  assign n1256 = ( ~n1231 & n1234 ) | ( ~n1231 & n1255 ) | ( n1234 & n1255 ) ;
  assign n1257 = ( ~n1225 & n1228 ) | ( ~n1225 & n1256 ) | ( n1228 & n1256 ) ;
  assign n1258 = ( ~n1219 & n1222 ) | ( ~n1219 & n1257 ) | ( n1222 & n1257 ) ;
  assign n1259 = ~n1216 & n1258 ;
  assign n1260 = ( ~n1212 & n1215 ) | ( ~n1212 & n1259 ) | ( n1215 & n1259 ) ;
  assign n1261 = x446 | n737 ;
  assign n1262 = ( n1215 & n1258 ) | ( n1215 & ~n1261 ) | ( n1258 & ~n1261 ) ;
  assign n1263 = ( ~x318 & n1260 ) | ( ~x318 & n1262 ) | ( n1260 & n1262 ) ;
  assign n1264 = x319 & n737 ;
  assign n1265 = x447 & ~n737 ;
  assign n1266 = n1264 | n1265 ;
  assign n1267 = x191 | n969 ;
  assign n1268 = ~x63 & n969 ;
  assign n1269 = n1267 & ~n1268 ;
  assign n1270 = ( n1263 & ~n1266 ) | ( n1263 & n1269 ) | ( ~n1266 & n1269 ) ;
  assign n1271 = x175 | n969 ;
  assign n1272 = ~x47 & n969 ;
  assign n1273 = n1271 & ~n1272 ;
  assign n1274 = x303 & n737 ;
  assign n1275 = x431 & ~n737 ;
  assign n1276 = n1274 | n1275 ;
  assign n1277 = x430 & ~n737 ;
  assign n1278 = x302 & n737 ;
  assign n1279 = n1277 | n1278 ;
  assign n1280 = x174 | n969 ;
  assign n1281 = ~x46 & n969 ;
  assign n1282 = n1280 & ~n1281 ;
  assign n1283 = x429 | n737 ;
  assign n1284 = ~x301 & n737 ;
  assign n1285 = n1283 & ~n1284 ;
  assign n1286 = x173 | n969 ;
  assign n1287 = ~x45 & n969 ;
  assign n1288 = n1286 & ~n1287 ;
  assign n1289 = x426 & ~n737 ;
  assign n1290 = x298 & n737 ;
  assign n1291 = n1289 | n1290 ;
  assign n1292 = x170 | n969 ;
  assign n1293 = ~x42 & n969 ;
  assign n1294 = n1292 & ~n1293 ;
  assign n1295 = x425 & ~n737 ;
  assign n1296 = x297 & n737 ;
  assign n1297 = n1295 | n1296 ;
  assign n1298 = x169 | n969 ;
  assign n1299 = ~x41 & n969 ;
  assign n1300 = n1298 & ~n1299 ;
  assign n1301 = x424 & ~n737 ;
  assign n1302 = x296 & n737 ;
  assign n1303 = n1301 | n1302 ;
  assign n1304 = x168 | n969 ;
  assign n1305 = ~x40 & n969 ;
  assign n1306 = n1304 & ~n1305 ;
  assign n1307 = x418 | n737 ;
  assign n1308 = ~x290 & n737 ;
  assign n1309 = n1307 & ~n1308 ;
  assign n1310 = x162 | n969 ;
  assign n1311 = ~x34 & n969 ;
  assign n1312 = n1310 & ~n1311 ;
  assign n1313 = x415 | n737 ;
  assign n1314 = ~x287 & n737 ;
  assign n1315 = n1313 & ~n1314 ;
  assign n1316 = x159 | n969 ;
  assign n1317 = ~x31 & n969 ;
  assign n1318 = n1316 & ~n1317 ;
  assign n1319 = n1315 & ~n1318 ;
  assign n1320 = x414 | n737 ;
  assign n1321 = ~x286 & n737 ;
  assign n1322 = n1320 & ~n1321 ;
  assign n1323 = x158 | n969 ;
  assign n1324 = ~x30 & n969 ;
  assign n1325 = n1323 & ~n1324 ;
  assign n1326 = x413 | n737 ;
  assign n1327 = ~x285 & n737 ;
  assign n1328 = n1326 & ~n1327 ;
  assign n1329 = x157 | n969 ;
  assign n1330 = ~x29 & n969 ;
  assign n1331 = n1329 & ~n1330 ;
  assign n1332 = x412 & ~n737 ;
  assign n1333 = x284 & n737 ;
  assign n1334 = x156 | n969 ;
  assign n1335 = ~x28 & n969 ;
  assign n1336 = n1334 & ~n1335 ;
  assign n1337 = ( n1332 & n1333 ) | ( n1332 & ~n1336 ) | ( n1333 & ~n1336 ) ;
  assign n1338 = ( n1328 & ~n1331 ) | ( n1328 & n1337 ) | ( ~n1331 & n1337 ) ;
  assign n1339 = x411 | n737 ;
  assign n1340 = ~x283 & n737 ;
  assign n1341 = n1339 & ~n1340 ;
  assign n1342 = x155 | n969 ;
  assign n1343 = ~x27 & n969 ;
  assign n1344 = n1342 & ~n1343 ;
  assign n1345 = x408 | n737 ;
  assign n1346 = ~x280 & n737 ;
  assign n1347 = n1345 & ~n1346 ;
  assign n1348 = x152 | n969 ;
  assign n1349 = ~x24 & n969 ;
  assign n1350 = n1348 & ~n1349 ;
  assign n1351 = x407 | n737 ;
  assign n1352 = ~x279 & n737 ;
  assign n1353 = n1351 & ~n1352 ;
  assign n1354 = x151 | n969 ;
  assign n1355 = ~x23 & n969 ;
  assign n1356 = n1354 & ~n1355 ;
  assign n1357 = x406 | n737 ;
  assign n1358 = ~x278 & n737 ;
  assign n1359 = x150 | n969 ;
  assign n1360 = ~x22 & n969 ;
  assign n1361 = n1359 & ~n1360 ;
  assign n1362 = ( ~n1357 & n1358 ) | ( ~n1357 & n1361 ) | ( n1358 & n1361 ) ;
  assign n1363 = ( ~n1351 & n1352 ) | ( ~n1351 & n1356 ) | ( n1352 & n1356 ) ;
  assign n1364 = n1362 | n1363 ;
  assign n1365 = x272 & n737 ;
  assign n1366 = x400 & ~n737 ;
  assign n1367 = x144 | n969 ;
  assign n1368 = ~x16 & n969 ;
  assign n1369 = n1367 & ~n1368 ;
  assign n1370 = ( n1365 & n1366 ) | ( n1365 & ~n1369 ) | ( n1366 & ~n1369 ) ;
  assign n1371 = x398 & ~n737 ;
  assign n1372 = x270 & n737 ;
  assign n1373 = x142 | n969 ;
  assign n1374 = ~x14 & n969 ;
  assign n1375 = n1373 & ~n1374 ;
  assign n1376 = ( n1371 & n1372 ) | ( n1371 & ~n1375 ) | ( n1372 & ~n1375 ) ;
  assign n1377 = x403 & ~n737 ;
  assign n1378 = x275 & n737 ;
  assign n1379 = x147 | n969 ;
  assign n1380 = ~x19 & n969 ;
  assign n1381 = n1379 & ~n1380 ;
  assign n1382 = ( n1377 & n1378 ) | ( n1377 & ~n1381 ) | ( n1378 & ~n1381 ) ;
  assign n1383 = x399 & ~n737 ;
  assign n1384 = x271 & n737 ;
  assign n1385 = x143 | n969 ;
  assign n1386 = ~x15 & n969 ;
  assign n1387 = n1385 & ~n1386 ;
  assign n1388 = ( n1383 & n1384 ) | ( n1383 & ~n1387 ) | ( n1384 & ~n1387 ) ;
  assign n1389 = ( ~n1370 & n1382 ) | ( ~n1370 & n1388 ) | ( n1382 & n1388 ) ;
  assign n1390 = ( ~n1370 & n1376 ) | ( ~n1370 & n1389 ) | ( n1376 & n1389 ) ;
  assign n1391 = n1370 | n1390 ;
  assign n1392 = x274 & n737 ;
  assign n1393 = x402 & ~n737 ;
  assign n1394 = x146 | n969 ;
  assign n1395 = ~x18 & n969 ;
  assign n1396 = n1394 & ~n1395 ;
  assign n1397 = ( n1392 & n1393 ) | ( n1392 & ~n1396 ) | ( n1393 & ~n1396 ) ;
  assign n1398 = x145 | n969 ;
  assign n1399 = ~x17 & n969 ;
  assign n1400 = n1398 & ~n1399 ;
  assign n1401 = x273 & n737 ;
  assign n1402 = x401 & ~n737 ;
  assign n1403 = ( ~n1400 & n1401 ) | ( ~n1400 & n1402 ) | ( n1401 & n1402 ) ;
  assign n1404 = n1397 | n1403 ;
  assign n1405 = n1391 | n1404 ;
  assign n1406 = x390 | n737 ;
  assign n1407 = ~x262 & n737 ;
  assign n1408 = n1406 & ~n1407 ;
  assign n1409 = x134 | n969 ;
  assign n1410 = ~x6 & n969 ;
  assign n1411 = n1409 & ~n1410 ;
  assign n1412 = x389 | n737 ;
  assign n1413 = ~x261 & n737 ;
  assign n1414 = n1412 & ~n1413 ;
  assign n1415 = x133 | n969 ;
  assign n1416 = ~x5 & n969 ;
  assign n1417 = n1415 & ~n1416 ;
  assign n1418 = x388 | n737 ;
  assign n1419 = ~x260 & n737 ;
  assign n1420 = n1418 & ~n1419 ;
  assign n1421 = x132 | n969 ;
  assign n1422 = ~x4 & n969 ;
  assign n1423 = n1421 & ~n1422 ;
  assign n1424 = x385 | n737 ;
  assign n1425 = ~x257 & n737 ;
  assign n1426 = n1424 & ~n1425 ;
  assign n1427 = x129 | n969 ;
  assign n1428 = ~x1 & n969 ;
  assign n1429 = n1427 & ~n1428 ;
  assign n1430 = x128 & ~n969 ;
  assign n1431 = ~x0 & n969 ;
  assign n1432 = ( n969 & n1430 ) | ( n969 & ~n1431 ) | ( n1430 & ~n1431 ) ;
  assign n1433 = x384 & ~n737 ;
  assign n1434 = x256 & n737 ;
  assign n1435 = n1433 | n1434 ;
  assign n1436 = n1432 & ~n1435 ;
  assign n1437 = ( ~n1426 & n1429 ) | ( ~n1426 & n1436 ) | ( n1429 & n1436 ) ;
  assign n1438 = ~x258 & n737 ;
  assign n1439 = x386 | n737 ;
  assign n1440 = ~n1438 & n1439 ;
  assign n1441 = x130 | n969 ;
  assign n1442 = ~x2 & n969 ;
  assign n1443 = n1441 & ~n1442 ;
  assign n1444 = ( n1437 & ~n1440 ) | ( n1437 & n1443 ) | ( ~n1440 & n1443 ) ;
  assign n1445 = x387 | n737 ;
  assign n1446 = ~x259 & n737 ;
  assign n1447 = n1445 & ~n1446 ;
  assign n1448 = x131 | n969 ;
  assign n1449 = ~x3 & n969 ;
  assign n1450 = n1448 & ~n1449 ;
  assign n1451 = ( n1444 & ~n1447 ) | ( n1444 & n1450 ) | ( ~n1447 & n1450 ) ;
  assign n1452 = ( ~n1420 & n1423 ) | ( ~n1420 & n1451 ) | ( n1423 & n1451 ) ;
  assign n1453 = ( ~n1414 & n1417 ) | ( ~n1414 & n1452 ) | ( n1417 & n1452 ) ;
  assign n1454 = ( ~n1408 & n1411 ) | ( ~n1408 & n1453 ) | ( n1411 & n1453 ) ;
  assign n1455 = x391 | n737 ;
  assign n1456 = ~x263 & n737 ;
  assign n1457 = n1455 & ~n1456 ;
  assign n1458 = x135 | n969 ;
  assign n1459 = ~x7 & n969 ;
  assign n1460 = n1458 & ~n1459 ;
  assign n1461 = ( n1454 & ~n1457 ) | ( n1454 & n1460 ) | ( ~n1457 & n1460 ) ;
  assign n1462 = x392 | n737 ;
  assign n1463 = ~x264 & n737 ;
  assign n1464 = n1462 & ~n1463 ;
  assign n1465 = x136 | n969 ;
  assign n1466 = ~x8 & n969 ;
  assign n1467 = n1465 & ~n1466 ;
  assign n1468 = ( n1461 & ~n1464 ) | ( n1461 & n1467 ) | ( ~n1464 & n1467 ) ;
  assign n1469 = x393 | n737 ;
  assign n1470 = ~x265 & n737 ;
  assign n1471 = n1469 & ~n1470 ;
  assign n1472 = x137 | n969 ;
  assign n1473 = ~x9 & n969 ;
  assign n1474 = n1472 & ~n1473 ;
  assign n1475 = ( n1468 & ~n1471 ) | ( n1468 & n1474 ) | ( ~n1471 & n1474 ) ;
  assign n1476 = x394 | n737 ;
  assign n1477 = ~x266 & n737 ;
  assign n1478 = n1476 & ~n1477 ;
  assign n1479 = x138 | n969 ;
  assign n1480 = ~x10 & n969 ;
  assign n1481 = n1479 & ~n1480 ;
  assign n1482 = ( n1475 & ~n1478 ) | ( n1475 & n1481 ) | ( ~n1478 & n1481 ) ;
  assign n1483 = x269 & n737 ;
  assign n1484 = x397 & ~n737 ;
  assign n1485 = x141 | n969 ;
  assign n1486 = ~x13 & n969 ;
  assign n1487 = n1485 & ~n1486 ;
  assign n1488 = ( n1483 & n1484 ) | ( n1483 & ~n1487 ) | ( n1484 & ~n1487 ) ;
  assign n1489 = x268 & n737 ;
  assign n1490 = x396 & ~n737 ;
  assign n1491 = x140 | n969 ;
  assign n1492 = ~x12 & n969 ;
  assign n1493 = n1491 & ~n1492 ;
  assign n1494 = ( n1489 & n1490 ) | ( n1489 & ~n1493 ) | ( n1490 & ~n1493 ) ;
  assign n1495 = n1488 | n1494 ;
  assign n1496 = x267 & n737 ;
  assign n1497 = x395 & ~n737 ;
  assign n1498 = x139 | n969 ;
  assign n1499 = ~x11 & n969 ;
  assign n1500 = n1498 & ~n1499 ;
  assign n1501 = ( n1496 & n1497 ) | ( n1496 & ~n1500 ) | ( n1497 & ~n1500 ) ;
  assign n1502 = n1495 | n1501 ;
  assign n1503 = n1482 & ~n1502 ;
  assign n1504 = n1483 | n1484 ;
  assign n1505 = n1489 | n1490 ;
  assign n1506 = n1496 | n1497 ;
  assign n1507 = n1500 & ~n1506 ;
  assign n1508 = ( n1493 & ~n1505 ) | ( n1493 & n1507 ) | ( ~n1505 & n1507 ) ;
  assign n1509 = ( n1487 & ~n1504 ) | ( n1487 & n1508 ) | ( ~n1504 & n1508 ) ;
  assign n1510 = n1371 | n1372 ;
  assign n1511 = n1375 & ~n1510 ;
  assign n1512 = n1509 | n1511 ;
  assign n1513 = ~n1405 & n1512 ;
  assign n1514 = ( ~n1405 & n1503 ) | ( ~n1405 & n1513 ) | ( n1503 & n1513 ) ;
  assign n1515 = n1377 | n1378 ;
  assign n1516 = n1392 | n1393 ;
  assign n1517 = n1401 | n1402 ;
  assign n1518 = n1365 | n1366 ;
  assign n1519 = n1383 | n1384 ;
  assign n1520 = n1387 & ~n1519 ;
  assign n1521 = ( n1369 & ~n1518 ) | ( n1369 & n1520 ) | ( ~n1518 & n1520 ) ;
  assign n1522 = ( n1400 & ~n1517 ) | ( n1400 & n1521 ) | ( ~n1517 & n1521 ) ;
  assign n1523 = ( n1396 & ~n1516 ) | ( n1396 & n1522 ) | ( ~n1516 & n1522 ) ;
  assign n1524 = ( n1381 & ~n1515 ) | ( n1381 & n1523 ) | ( ~n1515 & n1523 ) ;
  assign n1525 = x405 | n737 ;
  assign n1526 = ~x277 & n737 ;
  assign n1527 = n1525 & ~n1526 ;
  assign n1528 = x149 | n969 ;
  assign n1529 = ~x21 & n969 ;
  assign n1530 = n1528 & ~n1529 ;
  assign n1531 = x404 & ~n737 ;
  assign n1532 = x276 & n737 ;
  assign n1533 = n1531 | n1532 ;
  assign n1534 = x148 | n969 ;
  assign n1535 = ~x20 & n969 ;
  assign n1536 = n1534 & ~n1535 ;
  assign n1537 = ~n1533 & n1536 ;
  assign n1538 = ( ~n1527 & n1530 ) | ( ~n1527 & n1537 ) | ( n1530 & n1537 ) ;
  assign n1539 = n1524 | n1538 ;
  assign n1540 = n1514 | n1539 ;
  assign n1541 = ( n1531 & n1532 ) | ( n1531 & ~n1536 ) | ( n1532 & ~n1536 ) ;
  assign n1542 = ( n1527 & ~n1530 ) | ( n1527 & n1541 ) | ( ~n1530 & n1541 ) ;
  assign n1543 = n1357 & ~n1358 ;
  assign n1544 = ( ~n1361 & n1542 ) | ( ~n1361 & n1543 ) | ( n1542 & n1543 ) ;
  assign n1545 = ~n1364 & n1544 ;
  assign n1546 = ( n1364 & n1540 ) | ( n1364 & ~n1545 ) | ( n1540 & ~n1545 ) ;
  assign n1547 = ( ~n1353 & n1356 ) | ( ~n1353 & n1546 ) | ( n1356 & n1546 ) ;
  assign n1548 = ( ~n1347 & n1350 ) | ( ~n1347 & n1547 ) | ( n1350 & n1547 ) ;
  assign n1549 = x409 | n737 ;
  assign n1550 = ~x281 & n737 ;
  assign n1551 = n1549 & ~n1550 ;
  assign n1552 = x153 | n969 ;
  assign n1553 = ~x25 & n969 ;
  assign n1554 = n1552 & ~n1553 ;
  assign n1555 = ( n1548 & ~n1551 ) | ( n1548 & n1554 ) | ( ~n1551 & n1554 ) ;
  assign n1556 = x410 | n737 ;
  assign n1557 = ~x282 & n737 ;
  assign n1558 = n1556 & ~n1557 ;
  assign n1559 = x154 | n969 ;
  assign n1560 = ~x26 & n969 ;
  assign n1561 = n1559 & ~n1560 ;
  assign n1562 = ( n1555 & ~n1558 ) | ( n1555 & n1561 ) | ( ~n1558 & n1561 ) ;
  assign n1563 = ( ~n1341 & n1344 ) | ( ~n1341 & n1562 ) | ( n1344 & n1562 ) ;
  assign n1564 = ~n1338 & n1563 ;
  assign n1565 = n1332 | n1333 ;
  assign n1566 = n1336 & ~n1565 ;
  assign n1567 = ( ~n1328 & n1331 ) | ( ~n1328 & n1566 ) | ( n1331 & n1566 ) ;
  assign n1568 = n1564 | n1567 ;
  assign n1569 = ( ~n1322 & n1325 ) | ( ~n1322 & n1568 ) | ( n1325 & n1568 ) ;
  assign n1570 = ~n1319 & n1569 ;
  assign n1571 = x417 | n737 ;
  assign n1572 = ~x289 & n737 ;
  assign n1573 = n1571 & ~n1572 ;
  assign n1574 = x161 | n969 ;
  assign n1575 = ~x33 & n969 ;
  assign n1576 = n1574 & ~n1575 ;
  assign n1577 = x288 & n737 ;
  assign n1578 = x416 & ~n737 ;
  assign n1579 = x160 | n969 ;
  assign n1580 = ~x32 & n969 ;
  assign n1581 = n1579 & ~n1580 ;
  assign n1582 = ( n1577 & n1578 ) | ( n1577 & ~n1581 ) | ( n1578 & ~n1581 ) ;
  assign n1583 = ( n1573 & ~n1576 ) | ( n1573 & n1582 ) | ( ~n1576 & n1582 ) ;
  assign n1584 = n1577 | n1578 ;
  assign n1585 = n1581 & ~n1584 ;
  assign n1586 = ( ~n1573 & n1576 ) | ( ~n1573 & n1585 ) | ( n1576 & n1585 ) ;
  assign n1587 = ( ~n1313 & n1314 ) | ( ~n1313 & n1318 ) | ( n1314 & n1318 ) ;
  assign n1588 = ( ~n1570 & n1586 ) | ( ~n1570 & n1587 ) | ( n1586 & n1587 ) ;
  assign n1589 = ( n1570 & ~n1583 ) | ( n1570 & n1588 ) | ( ~n1583 & n1588 ) ;
  assign n1590 = ( ~n1309 & n1312 ) | ( ~n1309 & n1589 ) | ( n1312 & n1589 ) ;
  assign n1591 = x419 | n737 ;
  assign n1592 = ~x291 & n737 ;
  assign n1593 = n1591 & ~n1592 ;
  assign n1594 = x163 | n969 ;
  assign n1595 = ~x35 & n969 ;
  assign n1596 = n1594 & ~n1595 ;
  assign n1597 = ( n1590 & ~n1593 ) | ( n1590 & n1596 ) | ( ~n1593 & n1596 ) ;
  assign n1598 = x421 | n737 ;
  assign n1599 = ~x293 & n737 ;
  assign n1600 = n1598 & ~n1599 ;
  assign n1601 = x165 | n969 ;
  assign n1602 = ~x37 & n969 ;
  assign n1603 = n1601 & ~n1602 ;
  assign n1604 = x420 & ~n737 ;
  assign n1605 = x292 & n737 ;
  assign n1606 = x164 | n969 ;
  assign n1607 = ~x36 & n969 ;
  assign n1608 = n1606 & ~n1607 ;
  assign n1609 = ( n1604 & n1605 ) | ( n1604 & ~n1608 ) | ( n1605 & ~n1608 ) ;
  assign n1610 = ( n1600 & ~n1603 ) | ( n1600 & n1609 ) | ( ~n1603 & n1609 ) ;
  assign n1611 = n1604 | n1605 ;
  assign n1612 = n1608 & ~n1611 ;
  assign n1613 = ( ~n1600 & n1603 ) | ( ~n1600 & n1612 ) | ( n1603 & n1612 ) ;
  assign n1614 = ( n1597 & ~n1610 ) | ( n1597 & n1613 ) | ( ~n1610 & n1613 ) ;
  assign n1615 = x422 | n737 ;
  assign n1616 = ~x294 & n737 ;
  assign n1617 = n1615 & ~n1616 ;
  assign n1618 = x166 | n969 ;
  assign n1619 = ~x38 & n969 ;
  assign n1620 = n1618 & ~n1619 ;
  assign n1621 = ( n1614 & ~n1617 ) | ( n1614 & n1620 ) | ( ~n1617 & n1620 ) ;
  assign n1622 = x423 | n737 ;
  assign n1623 = ~x295 & n737 ;
  assign n1624 = n1622 & ~n1623 ;
  assign n1625 = x167 | n969 ;
  assign n1626 = ~x39 & n969 ;
  assign n1627 = n1625 & ~n1626 ;
  assign n1628 = ( n1621 & ~n1624 ) | ( n1621 & n1627 ) | ( ~n1624 & n1627 ) ;
  assign n1629 = ( ~n1303 & n1306 ) | ( ~n1303 & n1628 ) | ( n1306 & n1628 ) ;
  assign n1630 = ( ~n1297 & n1300 ) | ( ~n1297 & n1629 ) | ( n1300 & n1629 ) ;
  assign n1631 = ( ~n1291 & n1294 ) | ( ~n1291 & n1630 ) | ( n1294 & n1630 ) ;
  assign n1632 = x427 | n737 ;
  assign n1633 = ~x299 & n737 ;
  assign n1634 = n1632 & ~n1633 ;
  assign n1635 = x171 | n969 ;
  assign n1636 = ~x43 & n969 ;
  assign n1637 = n1635 & ~n1636 ;
  assign n1638 = ( n1631 & ~n1634 ) | ( n1631 & n1637 ) | ( ~n1634 & n1637 ) ;
  assign n1639 = x428 | n737 ;
  assign n1640 = ~x300 & n737 ;
  assign n1641 = n1639 & ~n1640 ;
  assign n1642 = x172 | n969 ;
  assign n1643 = ~x44 & n969 ;
  assign n1644 = n1642 & ~n1643 ;
  assign n1645 = ( n1638 & ~n1641 ) | ( n1638 & n1644 ) | ( ~n1641 & n1644 ) ;
  assign n1646 = ( ~n1285 & n1288 ) | ( ~n1285 & n1645 ) | ( n1288 & n1645 ) ;
  assign n1647 = ( ~n1279 & n1282 ) | ( ~n1279 & n1646 ) | ( n1282 & n1646 ) ;
  assign n1648 = ( n1273 & ~n1276 ) | ( n1273 & n1647 ) | ( ~n1276 & n1647 ) ;
  assign n1649 = x182 | n969 ;
  assign n1650 = ~x54 & n969 ;
  assign n1651 = n1649 & ~n1650 ;
  assign n1652 = x438 | n737 ;
  assign n1653 = x181 | n969 ;
  assign n1654 = ~x53 & n969 ;
  assign n1655 = n1653 & ~n1654 ;
  assign n1656 = x437 & ~n737 ;
  assign n1657 = x309 & n737 ;
  assign n1658 = n1656 | n1657 ;
  assign n1659 = x180 | n969 ;
  assign n1660 = ~x52 & n969 ;
  assign n1661 = n1659 & ~n1660 ;
  assign n1662 = x436 & ~n737 ;
  assign n1663 = x308 & n737 ;
  assign n1664 = n1662 | n1663 ;
  assign n1665 = x179 | n969 ;
  assign n1666 = ~x51 & n969 ;
  assign n1667 = n1665 & ~n1666 ;
  assign n1668 = x435 & ~n737 ;
  assign n1669 = x307 & n737 ;
  assign n1670 = n1668 | n1669 ;
  assign n1671 = x178 | n969 ;
  assign n1672 = ~x50 & n969 ;
  assign n1673 = n1671 & ~n1672 ;
  assign n1674 = x434 & ~n737 ;
  assign n1675 = x306 & n737 ;
  assign n1676 = n1674 | n1675 ;
  assign n1677 = x177 | n969 ;
  assign n1678 = ~x49 & n969 ;
  assign n1679 = n1677 & ~n1678 ;
  assign n1680 = x433 & ~n737 ;
  assign n1681 = x305 & n737 ;
  assign n1682 = n1680 | n1681 ;
  assign n1683 = x176 | n969 ;
  assign n1684 = ~x48 & n969 ;
  assign n1685 = n1683 & ~n1684 ;
  assign n1686 = x304 & n737 ;
  assign n1687 = x432 & ~n737 ;
  assign n1688 = n1686 | n1687 ;
  assign n1689 = n1685 & ~n1688 ;
  assign n1690 = ( n1679 & ~n1682 ) | ( n1679 & n1689 ) | ( ~n1682 & n1689 ) ;
  assign n1691 = ( n1673 & ~n1676 ) | ( n1673 & n1690 ) | ( ~n1676 & n1690 ) ;
  assign n1692 = ( n1667 & ~n1670 ) | ( n1667 & n1691 ) | ( ~n1670 & n1691 ) ;
  assign n1693 = ( n1661 & ~n1664 ) | ( n1661 & n1692 ) | ( ~n1664 & n1692 ) ;
  assign n1694 = ( n1655 & ~n1658 ) | ( n1655 & n1693 ) | ( ~n1658 & n1693 ) ;
  assign n1695 = ( n1651 & ~n1652 ) | ( n1651 & n1694 ) | ( ~n1652 & n1694 ) ;
  assign n1696 = x438 & ~n737 ;
  assign n1697 = x310 & n737 ;
  assign n1698 = n1694 & ~n1697 ;
  assign n1699 = ( n1651 & ~n1696 ) | ( n1651 & n1698 ) | ( ~n1696 & n1698 ) ;
  assign n1700 = ( ~x310 & n1695 ) | ( ~x310 & n1699 ) | ( n1695 & n1699 ) ;
  assign n1701 = x311 & n737 ;
  assign n1702 = x439 & ~n737 ;
  assign n1703 = n1701 | n1702 ;
  assign n1704 = x183 | n969 ;
  assign n1705 = ~x55 & n969 ;
  assign n1706 = n1704 & ~n1705 ;
  assign n1707 = ~n1703 & n1706 ;
  assign n1708 = n1700 | n1707 ;
  assign n1709 = ( ~n1661 & n1662 ) | ( ~n1661 & n1663 ) | ( n1662 & n1663 ) ;
  assign n1710 = ( ~n1273 & n1274 ) | ( ~n1273 & n1275 ) | ( n1274 & n1275 ) ;
  assign n1711 = ( ~n1679 & n1680 ) | ( ~n1679 & n1681 ) | ( n1680 & n1681 ) ;
  assign n1712 = ( ~n1651 & n1696 ) | ( ~n1651 & n1697 ) | ( n1696 & n1697 ) ;
  assign n1713 = ( ~n1709 & n1711 ) | ( ~n1709 & n1712 ) | ( n1711 & n1712 ) ;
  assign n1714 = ( ~n1709 & n1710 ) | ( ~n1709 & n1713 ) | ( n1710 & n1713 ) ;
  assign n1715 = n1709 | n1714 ;
  assign n1716 = ( ~n1667 & n1668 ) | ( ~n1667 & n1669 ) | ( n1668 & n1669 ) ;
  assign n1717 = ( ~n1673 & n1674 ) | ( ~n1673 & n1675 ) | ( n1674 & n1675 ) ;
  assign n1718 = ( ~n1655 & n1656 ) | ( ~n1655 & n1657 ) | ( n1656 & n1657 ) ;
  assign n1719 = ( ~n1685 & n1686 ) | ( ~n1685 & n1687 ) | ( n1686 & n1687 ) ;
  assign n1720 = ( ~n1716 & n1718 ) | ( ~n1716 & n1719 ) | ( n1718 & n1719 ) ;
  assign n1721 = ( ~n1716 & n1717 ) | ( ~n1716 & n1720 ) | ( n1717 & n1720 ) ;
  assign n1722 = n1716 | n1721 ;
  assign n1723 = n1715 | n1722 ;
  assign n1724 = ~n1708 & n1723 ;
  assign n1725 = ( n1648 & n1708 ) | ( n1648 & ~n1724 ) | ( n1708 & ~n1724 ) ;
  assign n1726 = ( n1241 & n1242 ) | ( n1241 & ~n1246 ) | ( n1242 & ~n1246 ) ;
  assign n1727 = ( n1247 & n1248 ) | ( n1247 & ~n1252 ) | ( n1248 & ~n1252 ) ;
  assign n1728 = ( n1701 & n1702 ) | ( n1701 & ~n1706 ) | ( n1702 & ~n1706 ) ;
  assign n1729 = ( n1235 & n1236 ) | ( n1235 & ~n1240 ) | ( n1236 & ~n1240 ) ;
  assign n1730 = ( ~n1726 & n1728 ) | ( ~n1726 & n1729 ) | ( n1728 & n1729 ) ;
  assign n1731 = ( ~n1726 & n1727 ) | ( ~n1726 & n1730 ) | ( n1727 & n1730 ) ;
  assign n1732 = n1726 | n1731 ;
  assign n1733 = ( n1229 & n1230 ) | ( n1229 & ~n1234 ) | ( n1230 & ~n1234 ) ;
  assign n1734 = ( n1223 & n1224 ) | ( n1223 & n1228 ) | ( n1224 & n1228 ) ;
  assign n1735 = ( n1225 & n1733 ) | ( n1225 & ~n1734 ) | ( n1733 & ~n1734 ) ;
  assign n1736 = ( n1212 & ~n1215 ) | ( n1212 & n1216 ) | ( ~n1215 & n1216 ) ;
  assign n1737 = ( n1217 & n1218 ) | ( n1217 & ~n1222 ) | ( n1218 & ~n1222 ) ;
  assign n1738 = n1736 | n1737 ;
  assign n1739 = n1735 | n1738 ;
  assign n1740 = n1732 | n1739 ;
  assign n1741 = ~n1270 & n1740 ;
  assign n1742 = ( n1270 & n1725 ) | ( n1270 & ~n1741 ) | ( n1725 & ~n1741 ) ;
  assign n1743 = ( n1264 & n1265 ) | ( n1264 & ~n1269 ) | ( n1265 & ~n1269 ) ;
  assign n1744 = x449 & ~n737 ;
  assign n1745 = x321 & n737 ;
  assign n1746 = x193 | n969 ;
  assign n1747 = ~x65 & n969 ;
  assign n1748 = n1746 & ~n1747 ;
  assign n1749 = ( n1744 & n1745 ) | ( n1744 & ~n1748 ) | ( n1745 & ~n1748 ) ;
  assign n1750 = x450 & ~n737 ;
  assign n1751 = x322 & n737 ;
  assign n1752 = x194 | n969 ;
  assign n1753 = ~x66 & n969 ;
  assign n1754 = n1752 & ~n1753 ;
  assign n1755 = ( n1750 & n1751 ) | ( n1750 & ~n1754 ) | ( n1751 & ~n1754 ) ;
  assign n1756 = x448 & ~n737 ;
  assign n1757 = x320 & n737 ;
  assign n1758 = x192 | n969 ;
  assign n1759 = ~x64 & n969 ;
  assign n1760 = n1758 & ~n1759 ;
  assign n1761 = ( n1756 & n1757 ) | ( n1756 & ~n1760 ) | ( n1757 & ~n1760 ) ;
  assign n1762 = ( ~n1743 & n1755 ) | ( ~n1743 & n1761 ) | ( n1755 & n1761 ) ;
  assign n1763 = ( ~n1743 & n1749 ) | ( ~n1743 & n1762 ) | ( n1749 & n1762 ) ;
  assign n1764 = n1743 | n1763 ;
  assign n1765 = n1742 & ~n1764 ;
  assign n1766 = n1170 | n1171 ;
  assign n1767 = n1174 & ~n1766 ;
  assign n1768 = n1750 | n1751 ;
  assign n1769 = n1744 | n1745 ;
  assign n1770 = n1756 | n1757 ;
  assign n1771 = n1760 & ~n1770 ;
  assign n1772 = ( n1748 & ~n1769 ) | ( n1748 & n1771 ) | ( ~n1769 & n1771 ) ;
  assign n1773 = ( n1754 & ~n1768 ) | ( n1754 & n1772 ) | ( ~n1768 & n1772 ) ;
  assign n1774 = n1767 | n1773 ;
  assign n1775 = ~n1211 & n1774 ;
  assign n1776 = ( ~n1211 & n1765 ) | ( ~n1211 & n1775 ) | ( n1765 & n1775 ) ;
  assign n1777 = n1203 | n1204 ;
  assign n1778 = n1164 | n1165 ;
  assign n1779 = n1190 & ~n1197 ;
  assign n1780 = n1183 | n1184 ;
  assign n1781 = n1177 | n1178 ;
  assign n1782 = n1191 | n1192 ;
  assign n1783 = n1195 & ~n1782 ;
  assign n1784 = ( n1181 & ~n1781 ) | ( n1181 & n1783 ) | ( ~n1781 & n1783 ) ;
  assign n1785 = ( n1187 & ~n1780 ) | ( n1187 & n1784 ) | ( ~n1780 & n1784 ) ;
  assign n1786 = ( n1200 & ~n1779 ) | ( n1200 & n1785 ) | ( ~n1779 & n1785 ) ;
  assign n1787 = ( n1168 & ~n1778 ) | ( n1168 & n1786 ) | ( ~n1778 & n1786 ) ;
  assign n1788 = ( n1207 & ~n1777 ) | ( n1207 & n1787 ) | ( ~n1777 & n1787 ) ;
  assign n1789 = n1776 | n1788 ;
  assign n1790 = x458 | n737 ;
  assign n1791 = ~x330 & n737 ;
  assign n1792 = n1790 & ~n1791 ;
  assign n1793 = x202 | n969 ;
  assign n1794 = ~x74 & n969 ;
  assign n1795 = n1793 & ~n1794 ;
  assign n1796 = ( n1789 & ~n1792 ) | ( n1789 & n1795 ) | ( ~n1792 & n1795 ) ;
  assign n1797 = x459 | n737 ;
  assign n1798 = ~x331 & n737 ;
  assign n1799 = n1797 & ~n1798 ;
  assign n1800 = x203 | n969 ;
  assign n1801 = ~x75 & n969 ;
  assign n1802 = n1800 & ~n1801 ;
  assign n1803 = ( n1796 & ~n1799 ) | ( n1796 & n1802 ) | ( ~n1799 & n1802 ) ;
  assign n1804 = ( ~n1160 & n1163 ) | ( ~n1160 & n1803 ) | ( n1163 & n1803 ) ;
  assign n1805 = x205 | n969 ;
  assign n1806 = ~x77 & n969 ;
  assign n1807 = n1805 & ~n1806 ;
  assign n1808 = ( ~n1157 & n1804 ) | ( ~n1157 & n1807 ) | ( n1804 & n1807 ) ;
  assign n1809 = ( ~n1151 & n1154 ) | ( ~n1151 & n1808 ) | ( n1154 & n1808 ) ;
  assign n1810 = x207 | n969 ;
  assign n1811 = ~x79 & n969 ;
  assign n1812 = n1810 & ~n1811 ;
  assign n1813 = ( ~n1148 & n1809 ) | ( ~n1148 & n1812 ) | ( n1809 & n1812 ) ;
  assign n1814 = ( ~n1142 & n1145 ) | ( ~n1142 & n1813 ) | ( n1145 & n1813 ) ;
  assign n1815 = ( ~n1136 & n1139 ) | ( ~n1136 & n1814 ) | ( n1139 & n1814 ) ;
  assign n1816 = x466 | n737 ;
  assign n1817 = ~x338 & n737 ;
  assign n1818 = n1816 & ~n1817 ;
  assign n1819 = x210 | n969 ;
  assign n1820 = ~x82 & n969 ;
  assign n1821 = n1819 & ~n1820 ;
  assign n1822 = ( n1815 & ~n1818 ) | ( n1815 & n1821 ) | ( ~n1818 & n1821 ) ;
  assign n1823 = ( ~n1130 & n1133 ) | ( ~n1130 & n1822 ) | ( n1133 & n1822 ) ;
  assign n1824 = ( ~n1124 & n1127 ) | ( ~n1124 & n1823 ) | ( n1127 & n1823 ) ;
  assign n1825 = n1120 | n1824 ;
  assign n1826 = ( n1120 & ~n1121 ) | ( n1120 & n1825 ) | ( ~n1121 & n1825 ) ;
  assign n1827 = ( ~n1083 & n1084 ) | ( ~n1083 & n1085 ) | ( n1084 & n1085 ) ;
  assign n1828 = ( n1094 & n1101 ) | ( n1094 & ~n1104 ) | ( n1101 & ~n1104 ) ;
  assign n1829 = ( ~n1065 & n1066 ) | ( ~n1065 & n1067 ) | ( n1066 & n1067 ) ;
  assign n1830 = ( ~n1827 & n1828 ) | ( ~n1827 & n1829 ) | ( n1828 & n1829 ) ;
  assign n1831 = n1827 | n1830 ;
  assign n1832 = n1826 & ~n1831 ;
  assign n1833 = ( n1090 & ~n1108 ) | ( n1090 & n1832 ) | ( ~n1108 & n1832 ) ;
  assign n1834 = x227 | n969 ;
  assign n1835 = ~x99 & n969 ;
  assign n1836 = n1834 & ~n1835 ;
  assign n1837 = x355 & n737 ;
  assign n1838 = x483 & ~n737 ;
  assign n1839 = n1837 | n1838 ;
  assign n1840 = x226 | n969 ;
  assign n1841 = ~x98 & n969 ;
  assign n1842 = n1840 & ~n1841 ;
  assign n1843 = x482 & ~n737 ;
  assign n1844 = x354 & n737 ;
  assign n1845 = n1843 | n1844 ;
  assign n1846 = x225 | n969 ;
  assign n1847 = ~x97 & n969 ;
  assign n1848 = n1846 & ~n1847 ;
  assign n1849 = x353 & n737 ;
  assign n1850 = x481 & ~n737 ;
  assign n1851 = n1849 | n1850 ;
  assign n1852 = x224 | n969 ;
  assign n1853 = ~x96 & n969 ;
  assign n1854 = n1852 & ~n1853 ;
  assign n1855 = x480 & ~n737 ;
  assign n1856 = x352 & n737 ;
  assign n1857 = n1855 | n1856 ;
  assign n1858 = x223 | n969 ;
  assign n1859 = ~x95 & n969 ;
  assign n1860 = n1858 & ~n1859 ;
  assign n1861 = x479 & ~n737 ;
  assign n1862 = x351 & n737 ;
  assign n1863 = n1861 | n1862 ;
  assign n1864 = x222 | n969 ;
  assign n1865 = ~x94 & n969 ;
  assign n1866 = n1864 & ~n1865 ;
  assign n1867 = x478 & ~n737 ;
  assign n1868 = x350 & n737 ;
  assign n1869 = n1867 | n1868 ;
  assign n1870 = x221 | n969 ;
  assign n1871 = ~x93 & n969 ;
  assign n1872 = n1870 & ~n1871 ;
  assign n1873 = x349 & n737 ;
  assign n1874 = x477 & ~n737 ;
  assign n1875 = n1873 | n1874 ;
  assign n1876 = x220 | n969 ;
  assign n1877 = ~x92 & n969 ;
  assign n1878 = n1876 & ~n1877 ;
  assign n1879 = x476 & ~n737 ;
  assign n1880 = x348 & n737 ;
  assign n1881 = n1879 | n1880 ;
  assign n1882 = n1878 & ~n1881 ;
  assign n1883 = ( n1872 & ~n1875 ) | ( n1872 & n1882 ) | ( ~n1875 & n1882 ) ;
  assign n1884 = ( n1866 & ~n1869 ) | ( n1866 & n1883 ) | ( ~n1869 & n1883 ) ;
  assign n1885 = ( n1860 & ~n1863 ) | ( n1860 & n1884 ) | ( ~n1863 & n1884 ) ;
  assign n1886 = ( n1854 & ~n1857 ) | ( n1854 & n1885 ) | ( ~n1857 & n1885 ) ;
  assign n1887 = ( n1848 & ~n1851 ) | ( n1848 & n1886 ) | ( ~n1851 & n1886 ) ;
  assign n1888 = ( n1842 & ~n1845 ) | ( n1842 & n1887 ) | ( ~n1845 & n1887 ) ;
  assign n1889 = ( n1836 & ~n1839 ) | ( n1836 & n1888 ) | ( ~n1839 & n1888 ) ;
  assign n1890 = ( ~n1842 & n1843 ) | ( ~n1842 & n1844 ) | ( n1843 & n1844 ) ;
  assign n1891 = ( ~n1860 & n1861 ) | ( ~n1860 & n1862 ) | ( n1861 & n1862 ) ;
  assign n1892 = ( ~n1878 & n1879 ) | ( ~n1878 & n1880 ) | ( n1879 & n1880 ) ;
  assign n1893 = ( ~n1836 & n1837 ) | ( ~n1836 & n1838 ) | ( n1837 & n1838 ) ;
  assign n1894 = ( ~n1890 & n1892 ) | ( ~n1890 & n1893 ) | ( n1892 & n1893 ) ;
  assign n1895 = ( ~n1890 & n1891 ) | ( ~n1890 & n1894 ) | ( n1891 & n1894 ) ;
  assign n1896 = n1890 | n1895 ;
  assign n1897 = ( ~n1854 & n1855 ) | ( ~n1854 & n1856 ) | ( n1855 & n1856 ) ;
  assign n1898 = ( ~n1848 & n1849 ) | ( ~n1848 & n1850 ) | ( n1849 & n1850 ) ;
  assign n1899 = ( ~n1866 & n1867 ) | ( ~n1866 & n1868 ) | ( n1867 & n1868 ) ;
  assign n1900 = ( ~n1872 & n1873 ) | ( ~n1872 & n1874 ) | ( n1873 & n1874 ) ;
  assign n1901 = ( ~n1897 & n1899 ) | ( ~n1897 & n1900 ) | ( n1899 & n1900 ) ;
  assign n1902 = ( ~n1897 & n1898 ) | ( ~n1897 & n1901 ) | ( n1898 & n1901 ) ;
  assign n1903 = n1897 | n1902 ;
  assign n1904 = n1896 | n1903 ;
  assign n1905 = ~n1889 & n1904 ;
  assign n1906 = ( n1833 & n1889 ) | ( n1833 & ~n1905 ) | ( n1889 & ~n1905 ) ;
  assign n1907 = x484 | n737 ;
  assign n1908 = ~x356 & n737 ;
  assign n1909 = n1907 & ~n1908 ;
  assign n1910 = x228 | n969 ;
  assign n1911 = ~x100 & n969 ;
  assign n1912 = n1910 & ~n1911 ;
  assign n1913 = ( n1906 & ~n1909 ) | ( n1906 & n1912 ) | ( ~n1909 & n1912 ) ;
  assign n1914 = ( ~n1059 & n1062 ) | ( ~n1059 & n1913 ) | ( n1062 & n1913 ) ;
  assign n1915 = ~n1056 & n1914 ;
  assign n1916 = n1035 | n1036 ;
  assign n1917 = n1022 | n1023 ;
  assign n1918 = n1015 | n1016 ;
  assign n1919 = n1048 | n1049 ;
  assign n1920 = n1052 & ~n1919 ;
  assign n1921 = ( n1019 & ~n1918 ) | ( n1019 & n1920 ) | ( ~n1918 & n1920 ) ;
  assign n1922 = x489 | n737 ;
  assign n1923 = ( x361 & n1009 ) | ( x361 & n1922 ) | ( n1009 & n1922 ) ;
  assign n1924 = ( n1013 & n1921 ) | ( n1013 & ~n1923 ) | ( n1921 & ~n1923 ) ;
  assign n1925 = ( n1026 & ~n1917 ) | ( n1026 & n1924 ) | ( ~n1917 & n1924 ) ;
  assign n1926 = ( n1039 & ~n1916 ) | ( n1039 & n1925 ) | ( ~n1916 & n1925 ) ;
  assign n1927 = ~n1041 & n1926 ;
  assign n1928 = n1042 | n1043 ;
  assign n1929 = ( n1046 & ~n1056 ) | ( n1046 & n1928 ) | ( ~n1056 & n1928 ) ;
  assign n1930 = ~n1928 & n1929 ;
  assign n1931 = ( n1002 & ~n1003 ) | ( n1002 & n1006 ) | ( ~n1003 & n1006 ) ;
  assign n1932 = ( ~n1029 & n1030 ) | ( ~n1029 & n1033 ) | ( n1030 & n1033 ) ;
  assign n1933 = ( ~n1030 & n1931 ) | ( ~n1030 & n1932 ) | ( n1931 & n1932 ) ;
  assign n1934 = ~n1008 & n1933 ;
  assign n1935 = ( ~n1008 & n1930 ) | ( ~n1008 & n1934 ) | ( n1930 & n1934 ) ;
  assign n1936 = ( ~n1008 & n1927 ) | ( ~n1008 & n1935 ) | ( n1927 & n1935 ) ;
  assign n1937 = ( ~n1008 & n1915 ) | ( ~n1008 & n1936 ) | ( n1915 & n1936 ) ;
  assign n1938 = n996 | n997 ;
  assign n1939 = n1000 & ~n1938 ;
  assign n1940 = x239 | n969 ;
  assign n1941 = ~x111 & n969 ;
  assign n1942 = n1940 & ~n1941 ;
  assign n1943 = x495 & ~n737 ;
  assign n1944 = x367 & n737 ;
  assign n1945 = n1943 | n1944 ;
  assign n1946 = ( n1939 & n1942 ) | ( n1939 & ~n1945 ) | ( n1942 & ~n1945 ) ;
  assign n1947 = n1937 | n1946 ;
  assign n1948 = ( n738 & n739 ) | ( n738 & ~n972 ) | ( n739 & ~n972 ) ;
  assign n1949 = ( ~n1942 & n1943 ) | ( ~n1942 & n1944 ) | ( n1943 & n1944 ) ;
  assign n1950 = ( n973 & n974 ) | ( n973 & ~n978 ) | ( n974 & ~n978 ) ;
  assign n1951 = ( n979 & n980 ) | ( n979 & ~n984 ) | ( n980 & ~n984 ) ;
  assign n1952 = ( ~n1948 & n1950 ) | ( ~n1948 & n1951 ) | ( n1950 & n1951 ) ;
  assign n1953 = ( ~n1948 & n1949 ) | ( ~n1948 & n1952 ) | ( n1949 & n1952 ) ;
  assign n1954 = n1948 | n1953 ;
  assign n1955 = ~n995 & n1954 ;
  assign n1956 = ( n995 & n1947 ) | ( n995 & ~n1955 ) | ( n1947 & ~n1955 ) ;
  assign n1957 = x506 & ~n737 ;
  assign n1958 = x378 & n737 ;
  assign n1959 = x250 & ~n969 ;
  assign n1960 = x122 & n969 ;
  assign n1961 = n1959 | n1960 ;
  assign n1962 = ( n1957 & n1958 ) | ( n1957 & ~n1961 ) | ( n1958 & ~n1961 ) ;
  assign n1963 = x375 & n737 ;
  assign n1964 = x503 & ~n737 ;
  assign n1965 = x247 | n969 ;
  assign n1966 = ~x119 & n969 ;
  assign n1967 = n1965 & ~n1966 ;
  assign n1968 = ( n1963 & n1964 ) | ( n1963 & ~n1967 ) | ( n1964 & ~n1967 ) ;
  assign n1969 = x381 & n737 ;
  assign n1970 = x509 & ~n737 ;
  assign n1971 = x253 & ~n744 ;
  assign n1972 = x125 & n744 ;
  assign n1973 = n1971 | n1972 ;
  assign n1974 = ( n1969 & n1970 ) | ( n1969 & ~n1973 ) | ( n1970 & ~n1973 ) ;
  assign n1975 = x374 & n737 ;
  assign n1976 = x502 & ~n737 ;
  assign n1977 = x246 | n969 ;
  assign n1978 = ~x118 & n969 ;
  assign n1979 = n1977 & ~n1978 ;
  assign n1980 = ( n1975 & n1976 ) | ( n1975 & ~n1979 ) | ( n1976 & ~n1979 ) ;
  assign n1981 = ( ~n1962 & n1974 ) | ( ~n1962 & n1980 ) | ( n1974 & n1980 ) ;
  assign n1982 = ( ~n1962 & n1968 ) | ( ~n1962 & n1981 ) | ( n1968 & n1981 ) ;
  assign n1983 = n1962 | n1982 ;
  assign n1984 = x380 & n737 ;
  assign n1985 = x508 & ~n737 ;
  assign n1986 = x252 | n744 ;
  assign n1987 = ~x124 & n744 ;
  assign n1988 = n1986 & ~n1987 ;
  assign n1989 = ( n1984 & n1985 ) | ( n1984 & ~n1988 ) | ( n1985 & ~n1988 ) ;
  assign n1990 = x507 & ~n737 ;
  assign n1991 = x379 & n737 ;
  assign n1992 = x123 & ~n968 ;
  assign n1993 = x251 & ~n744 ;
  assign n1994 = n1992 | n1993 ;
  assign n1995 = ( n1990 & n1991 ) | ( n1990 & ~n1994 ) | ( n1991 & ~n1994 ) ;
  assign n1996 = n1989 | n1995 ;
  assign n1997 = x377 & n737 ;
  assign n1998 = x505 & ~n737 ;
  assign n1999 = x249 | n969 ;
  assign n2000 = ~x121 & n969 ;
  assign n2001 = n1999 & ~n2000 ;
  assign n2002 = ( n1997 & n1998 ) | ( n1997 & ~n2001 ) | ( n1998 & ~n2001 ) ;
  assign n2003 = x504 & ~n737 ;
  assign n2004 = x376 & n737 ;
  assign n2005 = x248 | n969 ;
  assign n2006 = ~x120 & n969 ;
  assign n2007 = n2005 & ~n2006 ;
  assign n2008 = ( n2003 & n2004 ) | ( n2003 & ~n2007 ) | ( n2004 & ~n2007 ) ;
  assign n2009 = n2002 | n2008 ;
  assign n2010 = n1996 | n2009 ;
  assign n2011 = x373 & n737 ;
  assign n2012 = x501 & ~n737 ;
  assign n2013 = x245 | n969 ;
  assign n2014 = ~x117 & n969 ;
  assign n2015 = n2013 & ~n2014 ;
  assign n2016 = ( n2011 & n2012 ) | ( n2011 & ~n2015 ) | ( n2012 & ~n2015 ) ;
  assign n2017 = x510 & ~n737 ;
  assign n2018 = x382 & n737 ;
  assign n2019 = ( x127 & x254 ) | ( x127 & ~x255 ) | ( x254 & ~x255 ) ;
  assign n2020 = x126 & ~n2019 ;
  assign n2021 = ~x254 & n2019 ;
  assign n2022 = ( n2019 & n2020 ) | ( n2019 & ~n2021 ) | ( n2020 & ~n2021 ) ;
  assign n2023 = ( n2017 & n2018 ) | ( n2017 & ~n2022 ) | ( n2018 & ~n2022 ) ;
  assign n2024 = n2016 | n2023 ;
  assign n2025 = ( n988 & n989 ) | ( n988 & ~n993 ) | ( n989 & ~n993 ) ;
  assign n2026 = x372 & n737 ;
  assign n2027 = x500 & ~n737 ;
  assign n2028 = x244 | n969 ;
  assign n2029 = ~x116 & n969 ;
  assign n2030 = n2028 & ~n2029 ;
  assign n2031 = ( n2026 & n2027 ) | ( n2026 & ~n2030 ) | ( n2027 & ~n2030 ) ;
  assign n2032 = n2025 | n2031 ;
  assign n2033 = n2024 | n2032 ;
  assign n2034 = n2010 | n2033 ;
  assign n2035 = n1983 | n2034 ;
  assign n2036 = n1956 & ~n2035 ;
  assign n2037 = x510 | n737 ;
  assign n2038 = n1969 | n1970 ;
  assign n2039 = n1957 | n1958 ;
  assign n2040 = n1997 | n1998 ;
  assign n2041 = n2003 | n2004 ;
  assign n2042 = n1963 | n1964 ;
  assign n2043 = n1975 | n1976 ;
  assign n2044 = n2011 | n2012 ;
  assign n2045 = n2026 | n2027 ;
  assign n2046 = n2030 & ~n2045 ;
  assign n2047 = ( n2015 & ~n2044 ) | ( n2015 & n2046 ) | ( ~n2044 & n2046 ) ;
  assign n2048 = ( n1979 & ~n2043 ) | ( n1979 & n2047 ) | ( ~n2043 & n2047 ) ;
  assign n2049 = ( n1967 & ~n2042 ) | ( n1967 & n2048 ) | ( ~n2042 & n2048 ) ;
  assign n2050 = ( n2007 & ~n2041 ) | ( n2007 & n2049 ) | ( ~n2041 & n2049 ) ;
  assign n2051 = ( n2001 & ~n2040 ) | ( n2001 & n2050 ) | ( ~n2040 & n2050 ) ;
  assign n2052 = ( n1961 & ~n2039 ) | ( n1961 & n2051 ) | ( ~n2039 & n2051 ) ;
  assign n2053 = n1984 | n1985 ;
  assign n2054 = n1990 | n1991 ;
  assign n2055 = n1994 & ~n2054 ;
  assign n2056 = ( n1988 & ~n2053 ) | ( n1988 & n2055 ) | ( ~n2053 & n2055 ) ;
  assign n2057 = n1996 & ~n2056 ;
  assign n2058 = ( n2052 & n2056 ) | ( n2052 & ~n2057 ) | ( n2056 & ~n2057 ) ;
  assign n2059 = ( n1973 & ~n2038 ) | ( n1973 & n2058 ) | ( ~n2038 & n2058 ) ;
  assign n2060 = ( n2022 & ~n2037 ) | ( n2022 & n2059 ) | ( ~n2037 & n2059 ) ;
  assign n2061 = ~n2018 & n2059 ;
  assign n2062 = ( ~n2017 & n2022 ) | ( ~n2017 & n2061 ) | ( n2022 & n2061 ) ;
  assign n2063 = ( ~x382 & n2060 ) | ( ~x382 & n2062 ) | ( n2060 & n2062 ) ;
  assign n2064 = n2036 | n2063 ;
  assign n2065 = x383 & x511 ;
  assign n2066 = ( ~n513 & n2064 ) | ( ~n513 & n2065 ) | ( n2064 & n2065 ) ;
  assign n2067 = ~n1432 & n2066 ;
  assign n2068 = n1435 & ~n2066 ;
  assign n2069 = ( n2066 & ~n2067 ) | ( n2066 & n2068 ) | ( ~n2067 & n2068 ) ;
  assign n2070 = ~n1429 & n2066 ;
  assign n2071 = n1426 | n2066 ;
  assign n2072 = ~n2070 & n2071 ;
  assign n2073 = ~n1443 & n2066 ;
  assign n2074 = n1440 | n2066 ;
  assign n2075 = ~n2073 & n2074 ;
  assign n2076 = ~n1450 & n2066 ;
  assign n2077 = n1447 | n2066 ;
  assign n2078 = ~n2076 & n2077 ;
  assign n2079 = ~n1423 & n2066 ;
  assign n2080 = n1420 | n2066 ;
  assign n2081 = ~n2079 & n2080 ;
  assign n2082 = ~n1417 & n2066 ;
  assign n2083 = ( n1412 & ~n1413 ) | ( n1412 & n2066 ) | ( ~n1413 & n2066 ) ;
  assign n2084 = ~n2082 & n2083 ;
  assign n2085 = ~n1411 & n2066 ;
  assign n2086 = n1408 | n2066 ;
  assign n2087 = ~n2085 & n2086 ;
  assign n2088 = ~n1460 & n2066 ;
  assign n2089 = n1457 | n2066 ;
  assign n2090 = ~n2088 & n2089 ;
  assign n2091 = ~n1467 & n2066 ;
  assign n2092 = n1464 | n2066 ;
  assign n2093 = ~n2091 & n2092 ;
  assign n2094 = ~n1474 & n2066 ;
  assign n2095 = n1471 | n2066 ;
  assign n2096 = ~n2094 & n2095 ;
  assign n2097 = ~n1481 & n2066 ;
  assign n2098 = n1478 | n2066 ;
  assign n2099 = ~n2097 & n2098 ;
  assign n2100 = ~n1500 & n2066 ;
  assign n2101 = n1506 | n2066 ;
  assign n2102 = ~n2100 & n2101 ;
  assign n2103 = ~n1493 & n2066 ;
  assign n2104 = n1505 | n2066 ;
  assign n2105 = ~n2103 & n2104 ;
  assign n2106 = ~n1487 & n2066 ;
  assign n2107 = n1504 | n2066 ;
  assign n2108 = ~n2106 & n2107 ;
  assign n2109 = ~n1375 & n2066 ;
  assign n2110 = n1510 | n2066 ;
  assign n2111 = ~n2109 & n2110 ;
  assign n2112 = ~n1387 & n2066 ;
  assign n2113 = n1519 | n2066 ;
  assign n2114 = ~n2112 & n2113 ;
  assign n2115 = ~n1369 & n2066 ;
  assign n2116 = n1518 | n2066 ;
  assign n2117 = ~n2115 & n2116 ;
  assign n2118 = ~n1400 & n2066 ;
  assign n2119 = n1517 | n2066 ;
  assign n2120 = ~n2118 & n2119 ;
  assign n2121 = ~n1396 & n2066 ;
  assign n2122 = n1516 | n2066 ;
  assign n2123 = ~n2121 & n2122 ;
  assign n2124 = ~n1381 & n2066 ;
  assign n2125 = n1515 | n2066 ;
  assign n2126 = ~n2124 & n2125 ;
  assign n2127 = ~n1536 & n2066 ;
  assign n2128 = n1533 | n2066 ;
  assign n2129 = ~n2127 & n2128 ;
  assign n2130 = ~n1530 & n2066 ;
  assign n2131 = n1527 | n2066 ;
  assign n2132 = ~n2130 & n2131 ;
  assign n2133 = ~n1361 & n2066 ;
  assign n2134 = n1543 | n2066 ;
  assign n2135 = ~n2133 & n2134 ;
  assign n2136 = ~n1356 & n2066 ;
  assign n2137 = n1353 | n2066 ;
  assign n2138 = ~n2136 & n2137 ;
  assign n2139 = ~n1350 & n2066 ;
  assign n2140 = n1347 | n2066 ;
  assign n2141 = ~n2139 & n2140 ;
  assign n2142 = ~n1554 & n2066 ;
  assign n2143 = n1551 | n2066 ;
  assign n2144 = ~n2142 & n2143 ;
  assign n2145 = ~n1561 & n2066 ;
  assign n2146 = n1558 | n2066 ;
  assign n2147 = ~n2145 & n2146 ;
  assign n2148 = ~n1344 & n2066 ;
  assign n2149 = n1341 | n2066 ;
  assign n2150 = ~n2148 & n2149 ;
  assign n2151 = ~n1336 & n2066 ;
  assign n2152 = n1565 | n2066 ;
  assign n2153 = ~n2151 & n2152 ;
  assign n2154 = ~n1331 & n2066 ;
  assign n2155 = n1328 | n2066 ;
  assign n2156 = ~n2154 & n2155 ;
  assign n2157 = ~n1325 & n2066 ;
  assign n2158 = n1322 | n2066 ;
  assign n2159 = ~n2157 & n2158 ;
  assign n2160 = ~n1318 & n2066 ;
  assign n2161 = n1315 | n2066 ;
  assign n2162 = ~n2160 & n2161 ;
  assign n2163 = ~n1581 & n2066 ;
  assign n2164 = n1584 | n2066 ;
  assign n2165 = ~n2163 & n2164 ;
  assign n2166 = ~n1576 & n2066 ;
  assign n2167 = n1573 | n2066 ;
  assign n2168 = ~n2166 & n2167 ;
  assign n2169 = ~n1312 & n2066 ;
  assign n2170 = n1309 | n2066 ;
  assign n2171 = ~n2169 & n2170 ;
  assign n2172 = ~n1596 & n2066 ;
  assign n2173 = n1593 | n2066 ;
  assign n2174 = ~n2172 & n2173 ;
  assign n2175 = ~n1608 & n2066 ;
  assign n2176 = n1611 | n2066 ;
  assign n2177 = ~n2175 & n2176 ;
  assign n2178 = ~n1603 & n2066 ;
  assign n2179 = n1600 | n2066 ;
  assign n2180 = ~n2178 & n2179 ;
  assign n2181 = ~n1620 & n2066 ;
  assign n2182 = n1617 | n2066 ;
  assign n2183 = ~n2181 & n2182 ;
  assign n2184 = ~n1627 & n2066 ;
  assign n2185 = n1624 | n2066 ;
  assign n2186 = ~n2184 & n2185 ;
  assign n2187 = ~n1306 & n2066 ;
  assign n2188 = n1303 | n2066 ;
  assign n2189 = ~n2187 & n2188 ;
  assign n2190 = ~n1300 & n2066 ;
  assign n2191 = n1297 | n2066 ;
  assign n2192 = ~n2190 & n2191 ;
  assign n2193 = ~n1294 & n2066 ;
  assign n2194 = n1291 | n2066 ;
  assign n2195 = ~n2193 & n2194 ;
  assign n2196 = ~n1637 & n2066 ;
  assign n2197 = n1634 | n2066 ;
  assign n2198 = ~n2196 & n2197 ;
  assign n2199 = ~n1644 & n2066 ;
  assign n2200 = n1641 | n2066 ;
  assign n2201 = ~n2199 & n2200 ;
  assign n2202 = ~n1288 & n2066 ;
  assign n2203 = n1285 | n2066 ;
  assign n2204 = ~n2202 & n2203 ;
  assign n2205 = ~n1282 & n2066 ;
  assign n2206 = n1279 | n2066 ;
  assign n2207 = ~n2205 & n2206 ;
  assign n2208 = ~n1273 & n2066 ;
  assign n2209 = n1276 | n2066 ;
  assign n2210 = ~n2208 & n2209 ;
  assign n2211 = ~n1685 & n2066 ;
  assign n2212 = n1688 | n2066 ;
  assign n2213 = ~n2211 & n2212 ;
  assign n2214 = ~n1679 & n2066 ;
  assign n2215 = n1682 | n2066 ;
  assign n2216 = ~n2214 & n2215 ;
  assign n2217 = ~n1673 & n2066 ;
  assign n2218 = n1676 | n2066 ;
  assign n2219 = ~n2217 & n2218 ;
  assign n2220 = ~n1667 & n2066 ;
  assign n2221 = n1670 | n2066 ;
  assign n2222 = ~n2220 & n2221 ;
  assign n2223 = ~n1661 & n2066 ;
  assign n2224 = n1664 | n2066 ;
  assign n2225 = ~n2223 & n2224 ;
  assign n2226 = ~n1655 & n2066 ;
  assign n2227 = n1658 | n2066 ;
  assign n2228 = ~n2226 & n2227 ;
  assign n2229 = ~n1651 & n2066 ;
  assign n2230 = ( ~n1696 & n1697 ) | ( ~n1696 & n2066 ) | ( n1697 & n2066 ) ;
  assign n2231 = ( n1696 & ~n2229 ) | ( n1696 & n2230 ) | ( ~n2229 & n2230 ) ;
  assign n2232 = ~n1706 & n2066 ;
  assign n2233 = n1703 | n2066 ;
  assign n2234 = ~n2232 & n2233 ;
  assign n2235 = ~n1252 & n2066 ;
  assign n2236 = n1249 | n2066 ;
  assign n2237 = ~n2235 & n2236 ;
  assign n2238 = ~n1246 & n2066 ;
  assign n2239 = n1243 | n2066 ;
  assign n2240 = ~n2238 & n2239 ;
  assign n2241 = ~n1240 & n2066 ;
  assign n2242 = n1237 | n2066 ;
  assign n2243 = ~n2241 & n2242 ;
  assign n2244 = ~n1234 & n2066 ;
  assign n2245 = n1231 | n2066 ;
  assign n2246 = ~n2244 & n2245 ;
  assign n2247 = ~n1228 & n2066 ;
  assign n2248 = n1225 | n2066 ;
  assign n2249 = ~n2247 & n2248 ;
  assign n2250 = ~n1222 & n2066 ;
  assign n2251 = n1219 | n2066 ;
  assign n2252 = ~n2250 & n2251 ;
  assign n2253 = ~n1215 & n2066 ;
  assign n2254 = ( n1212 & ~n1216 ) | ( n1212 & n2066 ) | ( ~n1216 & n2066 ) ;
  assign n2255 = ( n1216 & ~n2253 ) | ( n1216 & n2254 ) | ( ~n2253 & n2254 ) ;
  assign n2256 = ~n1269 & n2066 ;
  assign n2257 = n1266 | n2066 ;
  assign n2258 = ~n2256 & n2257 ;
  assign n2259 = ~n1760 & n2066 ;
  assign n2260 = n1770 | n2066 ;
  assign n2261 = ~n2259 & n2260 ;
  assign n2262 = ~n1748 & n2066 ;
  assign n2263 = n1769 | n2066 ;
  assign n2264 = ~n2262 & n2263 ;
  assign n2265 = ~n1754 & n2066 ;
  assign n2266 = n1768 | n2066 ;
  assign n2267 = ~n2265 & n2266 ;
  assign n2268 = ~n1174 & n2066 ;
  assign n2269 = n1766 | n2066 ;
  assign n2270 = ~n2268 & n2269 ;
  assign n2271 = ~n1195 & n2066 ;
  assign n2272 = n1782 | n2066 ;
  assign n2273 = ~n2271 & n2272 ;
  assign n2274 = ~n1181 & n2066 ;
  assign n2275 = n1781 | n2066 ;
  assign n2276 = ~n2274 & n2275 ;
  assign n2277 = ~n1187 & n2066 ;
  assign n2278 = n1780 | n2066 ;
  assign n2279 = ~n2277 & n2278 ;
  assign n2280 = ~n1200 & n2066 ;
  assign n2281 = n1779 | n2066 ;
  assign n2282 = ~n2280 & n2281 ;
  assign n2283 = ~n1168 & n2066 ;
  assign n2284 = n1778 | n2066 ;
  assign n2285 = ~n2283 & n2284 ;
  assign n2286 = ~n1207 & n2066 ;
  assign n2287 = n1777 | n2066 ;
  assign n2288 = ~n2286 & n2287 ;
  assign n2289 = ~n1795 & n2066 ;
  assign n2290 = n1792 | n2066 ;
  assign n2291 = ~n2289 & n2290 ;
  assign n2292 = ~n1802 & n2066 ;
  assign n2293 = n1799 | n2066 ;
  assign n2294 = ~n2292 & n2293 ;
  assign n2295 = ~n1163 & n2066 ;
  assign n2296 = n1160 | n2066 ;
  assign n2297 = ~n2295 & n2296 ;
  assign n2298 = ~n1807 & n2066 ;
  assign n2299 = n1157 | n2066 ;
  assign n2300 = ~n2298 & n2299 ;
  assign n2301 = ~n1154 & n2066 ;
  assign n2302 = n1151 | n2066 ;
  assign n2303 = ~n2301 & n2302 ;
  assign n2304 = ~n1812 & n2066 ;
  assign n2305 = n1148 | n2066 ;
  assign n2306 = ~n2304 & n2305 ;
  assign n2307 = ~n1145 & n2066 ;
  assign n2308 = n1142 | n2066 ;
  assign n2309 = ~n2307 & n2308 ;
  assign n2310 = ~n1139 & n2066 ;
  assign n2311 = n1136 | n2066 ;
  assign n2312 = ~n2310 & n2311 ;
  assign n2313 = ~n1821 & n2066 ;
  assign n2314 = n1818 | n2066 ;
  assign n2315 = ~n2313 & n2314 ;
  assign n2316 = ~n1133 & n2066 ;
  assign n2317 = n1130 | n2066 ;
  assign n2318 = ~n2316 & n2317 ;
  assign n2319 = ~n1127 & n2066 ;
  assign n2320 = n1124 | n2066 ;
  assign n2321 = ~n2319 & n2320 ;
  assign n2322 = ~n1115 & n2066 ;
  assign n2323 = n1112 | n2066 ;
  assign n2324 = ~n2322 & n2323 ;
  assign n2325 = ~n1099 & n2066 ;
  assign n2326 = n1117 | n2066 ;
  assign n2327 = ~n2325 & n2326 ;
  assign n2328 = ~n1104 & n2066 ;
  assign n2329 = n1109 | n2066 ;
  assign n2330 = ~n2328 & n2329 ;
  assign n2331 = ~n1083 & n2066 ;
  assign n2332 = n1086 | n2066 ;
  assign n2333 = ~n2331 & n2332 ;
  assign n2334 = ~n1077 & n2066 ;
  assign n2335 = n1080 | n2066 ;
  assign n2336 = ~n2334 & n2335 ;
  assign n2337 = ~n1071 & n2066 ;
  assign n2338 = n1074 | n2066 ;
  assign n2339 = ~n2337 & n2338 ;
  assign n2340 = ~n1065 & n2066 ;
  assign n2341 = n1068 | n2066 ;
  assign n2342 = ~n2340 & n2341 ;
  assign n2343 = ~n1878 & n2066 ;
  assign n2344 = n1881 | n2066 ;
  assign n2345 = ~n2343 & n2344 ;
  assign n2346 = ~n1872 & n2066 ;
  assign n2347 = n1875 | n2066 ;
  assign n2348 = ~n2346 & n2347 ;
  assign n2349 = ~n1866 & n2066 ;
  assign n2350 = n1869 | n2066 ;
  assign n2351 = ~n2349 & n2350 ;
  assign n2352 = ~n1860 & n2066 ;
  assign n2353 = n1863 | n2066 ;
  assign n2354 = ~n2352 & n2353 ;
  assign n2355 = ~n1854 & n2066 ;
  assign n2356 = n1857 | n2066 ;
  assign n2357 = ~n2355 & n2356 ;
  assign n2358 = ~n1848 & n2066 ;
  assign n2359 = n1851 | n2066 ;
  assign n2360 = ~n2358 & n2359 ;
  assign n2361 = ~n1842 & n2066 ;
  assign n2362 = n1845 | n2066 ;
  assign n2363 = ~n2361 & n2362 ;
  assign n2364 = ~n1836 & n2066 ;
  assign n2365 = n1839 | n2066 ;
  assign n2366 = ~n2364 & n2365 ;
  assign n2367 = ~n1912 & n2066 ;
  assign n2368 = n1909 | n2066 ;
  assign n2369 = ~n2367 & n2368 ;
  assign n2370 = ~n1062 & n2066 ;
  assign n2371 = n1059 | n2066 ;
  assign n2372 = ~n2370 & n2371 ;
  assign n2373 = ~n1046 & n2066 ;
  assign n2374 = n1928 | n2066 ;
  assign n2375 = ~n2373 & n2374 ;
  assign n2376 = ~n1052 & n2066 ;
  assign n2377 = n1919 | n2066 ;
  assign n2378 = ~n2376 & n2377 ;
  assign n2379 = ~n1019 & n2066 ;
  assign n2380 = n1918 | n2066 ;
  assign n2381 = ~n2379 & n2380 ;
  assign n2382 = ~n1013 & n2066 ;
  assign n2383 = ( n1009 & ~n1010 ) | ( n1009 & n2066 ) | ( ~n1010 & n2066 ) ;
  assign n2384 = ( n1010 & ~n2382 ) | ( n1010 & n2383 ) | ( ~n2382 & n2383 ) ;
  assign n2385 = ~n1026 & n2066 ;
  assign n2386 = n1917 | n2066 ;
  assign n2387 = ~n2385 & n2386 ;
  assign n2388 = ~n1039 & n2066 ;
  assign n2389 = n1916 | n2066 ;
  assign n2390 = ~n2388 & n2389 ;
  assign n2391 = ~n1033 & n2066 ;
  assign n2392 = ( n1029 & ~n1030 ) | ( n1029 & n2066 ) | ( ~n1030 & n2066 ) ;
  assign n2393 = ( n1030 & ~n2391 ) | ( n1030 & n2392 ) | ( ~n2391 & n2392 ) ;
  assign n2394 = ~n1006 & n2066 ;
  assign n2395 = ( ~n1002 & n1003 ) | ( ~n1002 & n2066 ) | ( n1003 & n2066 ) ;
  assign n2396 = ~n2394 & n2395 ;
  assign n2397 = ~n1000 & n2066 ;
  assign n2398 = n1938 | n2066 ;
  assign n2399 = ~n2397 & n2398 ;
  assign n2400 = ~n1942 & n2066 ;
  assign n2401 = n1945 | n2066 ;
  assign n2402 = ~n2400 & n2401 ;
  assign n2403 = ~n984 & n2066 ;
  assign n2404 = n981 | n2066 ;
  assign n2405 = ~n2403 & n2404 ;
  assign n2406 = ~n978 & n2066 ;
  assign n2407 = n975 | n2066 ;
  assign n2408 = ~n2406 & n2407 ;
  assign n2409 = ~n972 & n2066 ;
  assign n2410 = n740 | n2066 ;
  assign n2411 = ~n2409 & n2410 ;
  assign n2412 = ~n993 & n2066 ;
  assign n2413 = n990 | n2066 ;
  assign n2414 = ~n2412 & n2413 ;
  assign n2415 = ~n2030 & n2066 ;
  assign n2416 = n2045 | n2066 ;
  assign n2417 = ~n2415 & n2416 ;
  assign n2418 = ~n2015 & n2066 ;
  assign n2419 = n2044 | n2066 ;
  assign n2420 = ~n2418 & n2419 ;
  assign n2421 = ~n1979 & n2066 ;
  assign n2422 = n2043 | n2066 ;
  assign n2423 = ~n2421 & n2422 ;
  assign n2424 = ~n1967 & n2066 ;
  assign n2425 = n2042 | n2066 ;
  assign n2426 = ~n2424 & n2425 ;
  assign n2427 = ~n2007 & n2066 ;
  assign n2428 = n2041 | n2066 ;
  assign n2429 = ~n2427 & n2428 ;
  assign n2430 = ~n2001 & n2066 ;
  assign n2431 = n2040 | n2066 ;
  assign n2432 = ~n2430 & n2431 ;
  assign n2433 = ~n1961 & n2066 ;
  assign n2434 = n2039 | n2066 ;
  assign n2435 = ~n2433 & n2434 ;
  assign n2436 = ~n1994 & n2066 ;
  assign n2437 = n2054 | n2066 ;
  assign n2438 = ~n2436 & n2437 ;
  assign n2439 = ~n1988 & n2066 ;
  assign n2440 = n2053 | n2066 ;
  assign n2441 = ~n2439 & n2440 ;
  assign n2442 = ~n1973 & n2066 ;
  assign n2443 = n2038 | n2066 ;
  assign n2444 = ~n2442 & n2443 ;
  assign n2445 = ~n2022 & n2066 ;
  assign n2446 = ( n2017 & ~n2018 ) | ( n2017 & n2066 ) | ( ~n2018 & n2066 ) ;
  assign n2447 = ( n2018 & ~n2445 ) | ( n2018 & n2446 ) | ( ~n2445 & n2446 ) ;
  assign n2448 = n513 & n2065 ;
  assign n2449 = ~n969 & n2066 ;
  assign n2450 = n737 | n2066 ;
  assign n2451 = ~n2449 & n2450 ;
  assign y0 = n2069 ;
  assign y1 = n2072 ;
  assign y2 = n2075 ;
  assign y3 = n2078 ;
  assign y4 = n2081 ;
  assign y5 = n2084 ;
  assign y6 = n2087 ;
  assign y7 = n2090 ;
  assign y8 = n2093 ;
  assign y9 = n2096 ;
  assign y10 = n2099 ;
  assign y11 = n2102 ;
  assign y12 = n2105 ;
  assign y13 = n2108 ;
  assign y14 = n2111 ;
  assign y15 = n2114 ;
  assign y16 = n2117 ;
  assign y17 = n2120 ;
  assign y18 = n2123 ;
  assign y19 = n2126 ;
  assign y20 = n2129 ;
  assign y21 = n2132 ;
  assign y22 = n2135 ;
  assign y23 = n2138 ;
  assign y24 = n2141 ;
  assign y25 = n2144 ;
  assign y26 = n2147 ;
  assign y27 = n2150 ;
  assign y28 = n2153 ;
  assign y29 = n2156 ;
  assign y30 = n2159 ;
  assign y31 = n2162 ;
  assign y32 = n2165 ;
  assign y33 = n2168 ;
  assign y34 = n2171 ;
  assign y35 = n2174 ;
  assign y36 = n2177 ;
  assign y37 = n2180 ;
  assign y38 = n2183 ;
  assign y39 = n2186 ;
  assign y40 = n2189 ;
  assign y41 = n2192 ;
  assign y42 = n2195 ;
  assign y43 = n2198 ;
  assign y44 = n2201 ;
  assign y45 = n2204 ;
  assign y46 = n2207 ;
  assign y47 = n2210 ;
  assign y48 = n2213 ;
  assign y49 = n2216 ;
  assign y50 = n2219 ;
  assign y51 = n2222 ;
  assign y52 = n2225 ;
  assign y53 = n2228 ;
  assign y54 = n2231 ;
  assign y55 = n2234 ;
  assign y56 = n2237 ;
  assign y57 = n2240 ;
  assign y58 = n2243 ;
  assign y59 = n2246 ;
  assign y60 = n2249 ;
  assign y61 = n2252 ;
  assign y62 = n2255 ;
  assign y63 = n2258 ;
  assign y64 = n2261 ;
  assign y65 = n2264 ;
  assign y66 = n2267 ;
  assign y67 = n2270 ;
  assign y68 = n2273 ;
  assign y69 = n2276 ;
  assign y70 = n2279 ;
  assign y71 = n2282 ;
  assign y72 = n2285 ;
  assign y73 = n2288 ;
  assign y74 = n2291 ;
  assign y75 = n2294 ;
  assign y76 = n2297 ;
  assign y77 = n2300 ;
  assign y78 = n2303 ;
  assign y79 = n2306 ;
  assign y80 = n2309 ;
  assign y81 = n2312 ;
  assign y82 = n2315 ;
  assign y83 = n2318 ;
  assign y84 = n2321 ;
  assign y85 = n2324 ;
  assign y86 = n2327 ;
  assign y87 = n2330 ;
  assign y88 = n2333 ;
  assign y89 = n2336 ;
  assign y90 = n2339 ;
  assign y91 = n2342 ;
  assign y92 = n2345 ;
  assign y93 = n2348 ;
  assign y94 = n2351 ;
  assign y95 = n2354 ;
  assign y96 = n2357 ;
  assign y97 = n2360 ;
  assign y98 = n2363 ;
  assign y99 = n2366 ;
  assign y100 = n2369 ;
  assign y101 = n2372 ;
  assign y102 = n2375 ;
  assign y103 = n2378 ;
  assign y104 = n2381 ;
  assign y105 = n2384 ;
  assign y106 = n2387 ;
  assign y107 = n2390 ;
  assign y108 = n2393 ;
  assign y109 = n2396 ;
  assign y110 = n2399 ;
  assign y111 = n2402 ;
  assign y112 = n2405 ;
  assign y113 = n2408 ;
  assign y114 = n2411 ;
  assign y115 = n2414 ;
  assign y116 = n2417 ;
  assign y117 = n2420 ;
  assign y118 = n2423 ;
  assign y119 = n2426 ;
  assign y120 = n2429 ;
  assign y121 = n2432 ;
  assign y122 = n2435 ;
  assign y123 = n2438 ;
  assign y124 = n2441 ;
  assign y125 = n2444 ;
  assign y126 = n2447 ;
  assign y127 = n2448 ;
  assign y128 = ~n2451 ;
  assign y129 = ~n2066 ;
endmodule
