module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 ;
  assign n25 = x0 | x1 ;
  assign n26 = ( x2 & x3 ) | ( x2 & ~n25 ) | ( x3 & ~n25 ) ;
  assign n27 = n25 | n26 ;
  assign n28 = x4 | n27 ;
  assign n29 = ( x5 & x6 ) | ( x5 & ~n28 ) | ( x6 & ~n28 ) ;
  assign n30 = n28 | n29 ;
  assign n31 = ( x7 & x8 ) | ( x7 & ~n30 ) | ( x8 & ~n30 ) ;
  assign n32 = n30 | n31 ;
  assign n33 = ( x9 & x10 ) | ( x9 & ~n32 ) | ( x10 & ~n32 ) ;
  assign n34 = n32 | n33 ;
  assign n35 = x11 | n34 ;
  assign n36 = x12 | n35 ;
  assign n37 = x13 | n36 ;
  assign n38 = ( x14 & x15 ) | ( x14 & ~n37 ) | ( x15 & ~n37 ) ;
  assign n39 = n37 | n38 ;
  assign n40 = x16 | n39 ;
  assign n41 = ( x17 & x18 ) | ( x17 & ~n40 ) | ( x18 & ~n40 ) ;
  assign n42 = n40 | n41 ;
  assign n43 = x19 | n42 ;
  assign n44 = x20 | n43 ;
  assign n45 = ( x21 & ~x22 ) | ( x21 & n44 ) | ( ~x22 & n44 ) ;
  assign n46 = x21 & ~x22 ;
  assign n47 = x22 | n43 ;
  assign n48 = ( x20 & x22 ) | ( x20 & n47 ) | ( x22 & n47 ) ;
  assign n49 = ( x20 & x22 ) | ( x20 & ~n47 ) | ( x22 & ~n47 ) ;
  assign n50 = ( n47 & ~n48 ) | ( n47 & n49 ) | ( ~n48 & n49 ) ;
  assign n51 = ( ~n45 & n46 ) | ( ~n45 & n50 ) | ( n46 & n50 ) ;
  assign n52 = ( ~x22 & n37 ) | ( ~x22 & n38 ) | ( n37 & n38 ) ;
  assign n53 = x15 & x22 ;
  assign n54 = ( x14 & ~x22 ) | ( x14 & n37 ) | ( ~x22 & n37 ) ;
  assign n55 = x15 & n54 ;
  assign n56 = ( n52 & n53 ) | ( n52 & ~n55 ) | ( n53 & ~n55 ) ;
  assign n57 = n51 & n56 ;
  assign n58 = ( x17 & ~x22 ) | ( x17 & n40 ) | ( ~x22 & n40 ) ;
  assign n59 = x17 & ~x22 ;
  assign n60 = x16 & x22 ;
  assign n61 = ( x16 & x22 ) | ( x16 & n39 ) | ( x22 & n39 ) ;
  assign n62 = ( n40 & n60 ) | ( n40 & ~n61 ) | ( n60 & ~n61 ) ;
  assign n63 = ( ~n58 & n59 ) | ( ~n58 & n62 ) | ( n59 & n62 ) ;
  assign n64 = ( ~x22 & n40 ) | ( ~x22 & n41 ) | ( n40 & n41 ) ;
  assign n65 = x18 & x22 ;
  assign n66 = x18 & n58 ;
  assign n67 = ( n64 & n65 ) | ( n64 & ~n66 ) | ( n65 & ~n66 ) ;
  assign n68 = ( x19 & ~x22 ) | ( x19 & n42 ) | ( ~x22 & n42 ) ;
  assign n69 = x19 & ~x22 ;
  assign n70 = x19 & ~n42 ;
  assign n71 = ( n68 & ~n69 ) | ( n68 & n70 ) | ( ~n69 & n70 ) ;
  assign n72 = ~n67 & n71 ;
  assign n73 = n63 & n72 ;
  assign n74 = ( n67 & ~n68 ) | ( n67 & n69 ) | ( ~n68 & n69 ) ;
  assign n75 = x17 & ~n40 ;
  assign n76 = ( n58 & ~n59 ) | ( n58 & n75 ) | ( ~n59 & n75 ) ;
  assign n77 = ~n62 & n76 ;
  assign n78 = n74 & n77 ;
  assign n79 = n62 | n76 ;
  assign n80 = n72 & ~n79 ;
  assign n81 = n78 | n80 ;
  assign n82 = ( n57 & n73 ) | ( n57 & n81 ) | ( n73 & n81 ) ;
  assign n83 = n51 & ~n56 ;
  assign n84 = n72 & n77 ;
  assign n85 = n83 & n84 ;
  assign n86 = n62 & n76 ;
  assign n87 = n74 & n86 ;
  assign n88 = n57 & n87 ;
  assign n89 = n85 | n88 ;
  assign n90 = ( n73 & n80 ) | ( n73 & n83 ) | ( n80 & n83 ) ;
  assign n91 = n63 & n74 ;
  assign n92 = n57 & n91 ;
  assign n93 = ( n78 & n83 ) | ( n78 & n87 ) | ( n83 & n87 ) ;
  assign n94 = n92 | n93 ;
  assign n95 = ( ~n89 & n90 ) | ( ~n89 & n94 ) | ( n90 & n94 ) ;
  assign n96 = ( ~n82 & n89 ) | ( ~n82 & n95 ) | ( n89 & n95 ) ;
  assign n97 = n82 | n96 ;
  assign n98 = n74 & ~n79 ;
  assign n99 = x21 & ~n44 ;
  assign n100 = ( n45 & ~n46 ) | ( n45 & n99 ) | ( ~n46 & n99 ) ;
  assign n101 = ~n50 & n100 ;
  assign n102 = ( n91 & n98 ) | ( n91 & n101 ) | ( n98 & n101 ) ;
  assign n103 = n67 | n71 ;
  assign n104 = n63 & ~n103 ;
  assign n105 = n86 & ~n103 ;
  assign n106 = n101 & n105 ;
  assign n107 = ~n56 & n101 ;
  assign n108 = ( n104 & n106 ) | ( n104 & n107 ) | ( n106 & n107 ) ;
  assign n109 = n57 & n84 ;
  assign n110 = n67 & n71 ;
  assign n111 = n77 & n110 ;
  assign n112 = n83 & n111 ;
  assign n113 = n109 | n112 ;
  assign n114 = n67 & n86 ;
  assign n115 = n71 & n114 ;
  assign n116 = n57 & n115 ;
  assign n117 = ( ~n108 & n113 ) | ( ~n108 & n116 ) | ( n113 & n116 ) ;
  assign n118 = n108 | n117 ;
  assign n119 = n79 | n103 ;
  assign n120 = n107 & ~n119 ;
  assign n121 = n78 & n107 ;
  assign n122 = n83 & n115 ;
  assign n123 = n121 | n122 ;
  assign n124 = ( ~n118 & n120 ) | ( ~n118 & n123 ) | ( n120 & n123 ) ;
  assign n125 = n118 | n124 ;
  assign n126 = n77 & ~n103 ;
  assign n127 = n107 & n126 ;
  assign n128 = ~n56 & n106 ;
  assign n129 = ( n106 & n127 ) | ( n106 & ~n128 ) | ( n127 & ~n128 ) ;
  assign n130 = n125 | n129 ;
  assign n131 = n72 & n86 ;
  assign n132 = n51 & n131 ;
  assign n133 = n57 & n111 ;
  assign n134 = n63 & n110 ;
  assign n135 = ~n76 & n110 ;
  assign n136 = ~n62 & n135 ;
  assign n137 = n57 & n136 ;
  assign n138 = ( n51 & n134 ) | ( n51 & n137 ) | ( n134 & n137 ) ;
  assign n139 = ( ~n132 & n133 ) | ( ~n132 & n138 ) | ( n133 & n138 ) ;
  assign n140 = n132 | n139 ;
  assign n141 = n56 & n101 ;
  assign n142 = ~n119 & n141 ;
  assign n143 = n83 & n136 ;
  assign n144 = n142 | n143 ;
  assign n145 = ( n104 & n126 ) | ( n104 & n141 ) | ( n126 & n141 ) ;
  assign n146 = n144 | n145 ;
  assign n147 = ( ~n130 & n140 ) | ( ~n130 & n146 ) | ( n140 & n146 ) ;
  assign n148 = n130 | n147 ;
  assign n149 = ( ~n97 & n102 ) | ( ~n97 & n148 ) | ( n102 & n148 ) ;
  assign n150 = n83 & n91 ;
  assign n151 = n83 & n98 ;
  assign n152 = ( n57 & n105 ) | ( n57 & n126 ) | ( n105 & n126 ) ;
  assign n153 = ( n83 & n105 ) | ( n83 & n126 ) | ( n105 & n126 ) ;
  assign n154 = n57 & n98 ;
  assign n155 = ( n51 & n104 ) | ( n51 & n154 ) | ( n104 & n154 ) ;
  assign n156 = n153 | n155 ;
  assign n157 = ( ~n151 & n152 ) | ( ~n151 & n156 ) | ( n152 & n156 ) ;
  assign n158 = n151 | n157 ;
  assign n159 = n150 | n158 ;
  assign n160 = n97 | n149 ;
  assign n161 = n159 | n160 ;
  assign n162 = n50 | n100 ;
  assign n163 = n56 & ~n162 ;
  assign n164 = n111 & n163 ;
  assign n165 = n83 & ~n119 ;
  assign n166 = n164 | n165 ;
  assign n167 = ( n91 & n98 ) | ( n91 & n107 ) | ( n98 & n107 ) ;
  assign n168 = n166 | n167 ;
  assign n169 = ( n134 & n136 ) | ( n134 & n163 ) | ( n136 & n163 ) ;
  assign n170 = n57 & ~n119 ;
  assign n171 = ( n91 & n98 ) | ( n91 & n141 ) | ( n98 & n141 ) ;
  assign n172 = n170 | n171 ;
  assign n173 = n115 & ~n162 ;
  assign n174 = n56 | n162 ;
  assign n175 = ( n111 & n134 ) | ( n111 & ~n174 ) | ( n134 & ~n174 ) ;
  assign n176 = ( ~n172 & n173 ) | ( ~n172 & n175 ) | ( n173 & n175 ) ;
  assign n177 = n172 | n176 ;
  assign n178 = ( ~n168 & n169 ) | ( ~n168 & n177 ) | ( n169 & n177 ) ;
  assign n179 = n168 | n178 ;
  assign n180 = ( n131 & n136 ) | ( n131 & ~n174 ) | ( n136 & ~n174 ) ;
  assign n181 = ( n84 & n131 ) | ( n84 & n163 ) | ( n131 & n163 ) ;
  assign n182 = ( ~n179 & n180 ) | ( ~n179 & n181 ) | ( n180 & n181 ) ;
  assign n183 = n179 | n182 ;
  assign n184 = n84 & ~n174 ;
  assign n185 = n148 | n184 ;
  assign n186 = n73 & ~n174 ;
  assign n187 = n80 & n163 ;
  assign n188 = n186 | n187 ;
  assign n189 = n73 & n163 ;
  assign n190 = ( ~n184 & n188 ) | ( ~n184 & n189 ) | ( n188 & n189 ) ;
  assign n191 = ( ~n183 & n185 ) | ( ~n183 & n190 ) | ( n185 & n190 ) ;
  assign n192 = n183 | n191 ;
  assign n193 = n161 | n192 ;
  assign n194 = ~n149 & n193 ;
  assign n195 = ( ~x22 & n25 ) | ( ~x22 & n26 ) | ( n25 & n26 ) ;
  assign n196 = x3 & x22 ;
  assign n197 = ( x2 & ~x22 ) | ( x2 & n25 ) | ( ~x22 & n25 ) ;
  assign n198 = x3 & n197 ;
  assign n199 = ( n195 & n196 ) | ( n195 & ~n198 ) | ( n196 & ~n198 ) ;
  assign n200 = n194 & n199 ;
  assign n201 = n50 & n100 ;
  assign n202 = n56 & n201 ;
  assign n203 = n126 & n202 ;
  assign n204 = n80 & n101 ;
  assign n205 = ( n56 & n203 ) | ( n56 & n204 ) | ( n203 & n204 ) ;
  assign n206 = ~n56 & n201 ;
  assign n207 = n78 & n206 ;
  assign n208 = n98 & n202 ;
  assign n209 = n207 | n208 ;
  assign n210 = n205 | n209 ;
  assign n211 = n98 & ~n174 ;
  assign n212 = n189 | n211 ;
  assign n213 = ( n57 & n84 ) | ( n57 & n98 ) | ( n84 & n98 ) ;
  assign n214 = n84 & n101 ;
  assign n215 = n164 | n214 ;
  assign n216 = ( n132 & ~n213 ) | ( n132 & n215 ) | ( ~n213 & n215 ) ;
  assign n217 = n213 | n216 ;
  assign n218 = ( ~n210 & n212 ) | ( ~n210 & n217 ) | ( n212 & n217 ) ;
  assign n219 = n210 | n218 ;
  assign n220 = n73 & n141 ;
  assign n221 = n119 | n174 ;
  assign n222 = ~n220 & n221 ;
  assign n223 = n87 & ~n174 ;
  assign n224 = n105 & n201 ;
  assign n225 = ( ~n56 & n223 ) | ( ~n56 & n224 ) | ( n223 & n224 ) ;
  assign n226 = ~n56 & n173 ;
  assign n227 = n91 & n201 ;
  assign n228 = n126 & n163 ;
  assign n229 = n78 & ~n174 ;
  assign n230 = n228 | n229 ;
  assign n231 = n227 | n230 ;
  assign n232 = n226 | n231 ;
  assign n233 = ( n222 & n225 ) | ( n222 & n232 ) | ( n225 & n232 ) ;
  assign n234 = n83 & n134 ;
  assign n235 = n222 & ~n234 ;
  assign n236 = n57 & n126 ;
  assign n237 = n101 & n111 ;
  assign n238 = n56 & n237 ;
  assign n239 = ( n235 & n236 ) | ( n235 & n238 ) | ( n236 & n238 ) ;
  assign n240 = n235 & ~n239 ;
  assign n241 = ( n219 & ~n233 ) | ( n219 & n240 ) | ( ~n233 & n240 ) ;
  assign n242 = ~n219 & n241 ;
  assign n243 = n136 & n201 ;
  assign n244 = n98 & n107 ;
  assign n245 = ( ~n202 & n243 ) | ( ~n202 & n244 ) | ( n243 & n244 ) ;
  assign n246 = n91 & n163 ;
  assign n247 = n126 & n141 ;
  assign n248 = n246 | n247 ;
  assign n249 = n245 | n248 ;
  assign n250 = n57 & n78 ;
  assign n251 = n143 | n250 ;
  assign n252 = n57 & n80 ;
  assign n253 = n98 & n141 ;
  assign n254 = n252 | n253 ;
  assign n255 = n131 & n163 ;
  assign n256 = n87 & n202 ;
  assign n257 = n73 & n107 ;
  assign n258 = ( ~n137 & n256 ) | ( ~n137 & n257 ) | ( n256 & n257 ) ;
  assign n259 = ( n137 & ~n255 ) | ( n137 & n258 ) | ( ~n255 & n258 ) ;
  assign n260 = n255 | n259 ;
  assign n261 = ( ~n248 & n254 ) | ( ~n248 & n260 ) | ( n254 & n260 ) ;
  assign n262 = ( ~n249 & n251 ) | ( ~n249 & n261 ) | ( n251 & n261 ) ;
  assign n263 = n249 | n262 ;
  assign n264 = ( n57 & n115 ) | ( n57 & n206 ) | ( n115 & n206 ) ;
  assign n265 = n87 & n107 ;
  assign n266 = n84 & n163 ;
  assign n267 = ( ~n264 & n265 ) | ( ~n264 & n266 ) | ( n265 & n266 ) ;
  assign n268 = n264 | n267 ;
  assign n269 = n133 | n150 ;
  assign n270 = n126 & ~n174 ;
  assign n271 = ~n56 & n237 ;
  assign n272 = ( n142 & n174 ) | ( n142 & n271 ) | ( n174 & n271 ) ;
  assign n273 = n270 | n272 ;
  assign n274 = n269 | n273 ;
  assign n275 = n56 & n243 ;
  assign n276 = n73 & n83 ;
  assign n277 = ( ~n56 & n106 ) | ( ~n56 & n276 ) | ( n106 & n276 ) ;
  assign n278 = n134 & ~n174 ;
  assign n279 = ( ~n275 & n277 ) | ( ~n275 & n278 ) | ( n277 & n278 ) ;
  assign n280 = n275 | n279 ;
  assign n281 = n51 & n104 ;
  assign n282 = n121 | n281 ;
  assign n283 = n101 & n134 ;
  assign n284 = ~n56 & n283 ;
  assign n285 = ( n80 & n115 ) | ( n80 & n202 ) | ( n115 & n202 ) ;
  assign n286 = ( n98 & n104 ) | ( n98 & n206 ) | ( n104 & n206 ) ;
  assign n287 = ( ~n284 & n285 ) | ( ~n284 & n286 ) | ( n285 & n286 ) ;
  assign n288 = n284 | n287 ;
  assign n289 = ( ~n280 & n282 ) | ( ~n280 & n288 ) | ( n282 & n288 ) ;
  assign n290 = ( ~n274 & n280 ) | ( ~n274 & n289 ) | ( n280 & n289 ) ;
  assign n291 = ( ~n268 & n274 ) | ( ~n268 & n290 ) | ( n274 & n290 ) ;
  assign n292 = n268 | n291 ;
  assign n293 = n263 | n292 ;
  assign n294 = n107 & n136 ;
  assign n295 = n88 | n294 ;
  assign n296 = ( ~n119 & n134 ) | ( ~n119 & n202 ) | ( n134 & n202 ) ;
  assign n297 = n83 & n126 ;
  assign n298 = ( n80 & ~n119 ) | ( n80 & n163 ) | ( ~n119 & n163 ) ;
  assign n299 = n297 | n298 ;
  assign n300 = n129 | n299 ;
  assign n301 = ( ~n295 & n296 ) | ( ~n295 & n300 ) | ( n296 & n300 ) ;
  assign n302 = n295 | n301 ;
  assign n303 = ( n242 & n293 ) | ( n242 & n302 ) | ( n293 & n302 ) ;
  assign n304 = n242 & ~n303 ;
  assign n305 = n80 & ~n174 ;
  assign n306 = ( n98 & n111 ) | ( n98 & n202 ) | ( n111 & n202 ) ;
  assign n307 = n305 | n306 ;
  assign n308 = n87 & n141 ;
  assign n309 = ( n56 & n227 ) | ( n56 & n308 ) | ( n227 & n308 ) ;
  assign n310 = n115 & n206 ;
  assign n311 = n57 & n73 ;
  assign n312 = n310 | n311 ;
  assign n313 = n217 | n312 ;
  assign n314 = n111 & n206 ;
  assign n315 = n83 & n105 ;
  assign n316 = ( ~n312 & n314 ) | ( ~n312 & n315 ) | ( n314 & n315 ) ;
  assign n317 = ( ~n309 & n313 ) | ( ~n309 & n316 ) | ( n313 & n316 ) ;
  assign n318 = n309 | n317 ;
  assign n319 = n307 | n318 ;
  assign n320 = ( n78 & n115 ) | ( n78 & n202 ) | ( n115 & n202 ) ;
  assign n321 = ( ~n206 & n220 ) | ( ~n206 & n243 ) | ( n220 & n243 ) ;
  assign n322 = n320 | n321 ;
  assign n323 = ( n145 & n212 ) | ( n145 & ~n322 ) | ( n212 & ~n322 ) ;
  assign n324 = n322 | n323 ;
  assign n325 = n91 & ~n174 ;
  assign n326 = n84 & n206 ;
  assign n327 = n325 | n326 ;
  assign n328 = n87 & n206 ;
  assign n329 = n80 & n202 ;
  assign n330 = n328 | n329 ;
  assign n331 = n134 & n163 ;
  assign n332 = n330 | n331 ;
  assign n333 = ( n120 & ~n327 ) | ( n120 & n332 ) | ( ~n327 & n332 ) ;
  assign n334 = n327 | n333 ;
  assign n335 = ( ~n319 & n324 ) | ( ~n319 & n334 ) | ( n324 & n334 ) ;
  assign n336 = n319 | n335 ;
  assign n337 = ~n56 & n281 ;
  assign n338 = ~n119 & n206 ;
  assign n339 = n107 & n115 ;
  assign n340 = n338 | n339 ;
  assign n341 = n136 & ~n174 ;
  assign n342 = n107 & n131 ;
  assign n343 = n341 | n342 ;
  assign n344 = n340 | n343 ;
  assign n345 = n223 | n257 ;
  assign n346 = ( n104 & ~n119 ) | ( n104 & n202 ) | ( ~n119 & n202 ) ;
  assign n347 = n104 & n163 ;
  assign n348 = ( n121 & ~n346 ) | ( n121 & n347 ) | ( ~n346 & n347 ) ;
  assign n349 = n346 | n348 ;
  assign n350 = ( ~n344 & n345 ) | ( ~n344 & n349 ) | ( n345 & n349 ) ;
  assign n351 = n344 | n350 ;
  assign n352 = ~n56 & n204 ;
  assign n353 = ( n237 & ~n271 ) | ( n237 & n352 ) | ( ~n271 & n352 ) ;
  assign n354 = n184 | n353 ;
  assign n355 = ( n87 & ~n119 ) | ( n87 & n163 ) | ( ~n119 & n163 ) ;
  assign n356 = n56 & n204 ;
  assign n357 = ( ~n354 & n355 ) | ( ~n354 & n356 ) | ( n355 & n356 ) ;
  assign n358 = n354 | n357 ;
  assign n359 = n255 | n283 ;
  assign n360 = ( ~n104 & n119 ) | ( ~n104 & n174 ) | ( n119 & n174 ) ;
  assign n361 = ( n358 & ~n359 ) | ( n358 & n360 ) | ( ~n359 & n360 ) ;
  assign n362 = ~n358 & n361 ;
  assign n363 = n131 & n141 ;
  assign n364 = n98 & n163 ;
  assign n365 = ( n171 & ~n363 ) | ( n171 & n364 ) | ( ~n363 & n364 ) ;
  assign n366 = n363 | n365 ;
  assign n367 = ( n351 & n362 ) | ( n351 & ~n366 ) | ( n362 & ~n366 ) ;
  assign n368 = ~n351 & n367 ;
  assign n369 = ~n337 & n368 ;
  assign n370 = ( ~n56 & n143 ) | ( ~n56 & n227 ) | ( n143 & n227 ) ;
  assign n371 = n98 & n206 ;
  assign n372 = ( n112 & ~n370 ) | ( n112 & n371 ) | ( ~n370 & n371 ) ;
  assign n373 = n370 | n372 ;
  assign n374 = n116 | n278 ;
  assign n375 = n138 | n374 ;
  assign n376 = ( n369 & n373 ) | ( n369 & n375 ) | ( n373 & n375 ) ;
  assign n377 = n369 & ~n376 ;
  assign n378 = n131 & n201 ;
  assign n379 = ~n56 & n378 ;
  assign n380 = n83 & n87 ;
  assign n381 = ( n83 & ~n119 ) | ( n83 & n380 ) | ( ~n119 & n380 ) ;
  assign n382 = ( n56 & n92 ) | ( n56 & n106 ) | ( n92 & n106 ) ;
  assign n383 = ( n83 & n98 ) | ( n83 & n126 ) | ( n98 & n126 ) ;
  assign n384 = n382 | n383 ;
  assign n385 = n381 | n384 ;
  assign n386 = n56 & n224 ;
  assign n387 = ( n73 & n78 ) | ( n73 & n206 ) | ( n78 & n206 ) ;
  assign n388 = ( ~n379 & n386 ) | ( ~n379 & n387 ) | ( n386 & n387 ) ;
  assign n389 = ( n379 & ~n385 ) | ( n379 & n388 ) | ( ~n385 & n388 ) ;
  assign n390 = ( n89 & n385 ) | ( n89 & ~n389 ) | ( n385 & ~n389 ) ;
  assign n391 = n389 | n390 ;
  assign n392 = ( n336 & n377 ) | ( n336 & ~n391 ) | ( n377 & ~n391 ) ;
  assign n393 = ~n336 & n392 ;
  assign n394 = n304 | n393 ;
  assign n395 = n57 & n105 ;
  assign n396 = ( n56 & ~n162 ) | ( n56 & n395 ) | ( ~n162 & n395 ) ;
  assign n397 = ( n105 & n173 ) | ( n105 & n396 ) | ( n173 & n396 ) ;
  assign n398 = ( n122 & n127 ) | ( n122 & ~n188 ) | ( n127 & ~n188 ) ;
  assign n399 = n188 | n398 ;
  assign n400 = n397 | n399 ;
  assign n401 = ( n83 & n84 ) | ( n83 & n202 ) | ( n84 & n202 ) ;
  assign n402 = n204 | n256 ;
  assign n403 = ( n105 & n173 ) | ( n105 & ~n174 ) | ( n173 & ~n174 ) ;
  assign n404 = ( ~n401 & n402 ) | ( ~n401 & n403 ) | ( n402 & n403 ) ;
  assign n405 = n401 | n404 ;
  assign n406 = n150 | n257 ;
  assign n407 = n386 | n406 ;
  assign n408 = n73 & n201 ;
  assign n409 = ( ~n56 & n265 ) | ( ~n56 & n408 ) | ( n265 & n408 ) ;
  assign n410 = n134 & n202 ;
  assign n411 = n276 | n410 ;
  assign n412 = ( ~n407 & n409 ) | ( ~n407 & n411 ) | ( n409 & n411 ) ;
  assign n413 = n407 | n412 ;
  assign n414 = ( ~n400 & n405 ) | ( ~n400 & n413 ) | ( n405 & n413 ) ;
  assign n415 = n400 | n414 ;
  assign n416 = ( n126 & n141 ) | ( n126 & ~n174 ) | ( n141 & ~n174 ) ;
  assign n417 = n222 & ~n416 ;
  assign n418 = ( n79 & n103 ) | ( n79 & ~n347 ) | ( n103 & ~n347 ) ;
  assign n419 = ( n202 & n347 ) | ( n202 & ~n418 ) | ( n347 & ~n418 ) ;
  assign n420 = ( n98 & n107 ) | ( n98 & n136 ) | ( n107 & n136 ) ;
  assign n421 = n419 | n420 ;
  assign n422 = n136 & n163 ;
  assign n423 = ( n56 & n214 ) | ( n56 & n237 ) | ( n214 & n237 ) ;
  assign n424 = ( ~n421 & n422 ) | ( ~n421 & n423 ) | ( n422 & n423 ) ;
  assign n425 = n421 | n424 ;
  assign n426 = n56 & n281 ;
  assign n427 = n104 & ~n174 ;
  assign n428 = n115 & n141 ;
  assign n429 = n427 | n428 ;
  assign n430 = ( n155 & ~n426 ) | ( n155 & n429 ) | ( ~n426 & n429 ) ;
  assign n431 = ( n417 & n425 ) | ( n417 & ~n430 ) | ( n425 & ~n430 ) ;
  assign n432 = n134 & n206 ;
  assign n433 = n112 | n432 ;
  assign n434 = ( n126 & n131 ) | ( n126 & n163 ) | ( n131 & n163 ) ;
  assign n435 = n223 | n434 ;
  assign n436 = n142 | n234 ;
  assign n437 = ( ~n433 & n435 ) | ( ~n433 & n436 ) | ( n435 & n436 ) ;
  assign n438 = n433 | n437 ;
  assign n439 = n104 & n206 ;
  assign n440 = ~n119 & n163 ;
  assign n441 = n439 | n440 ;
  assign n442 = ~n56 & n214 ;
  assign n443 = ( n343 & ~n441 ) | ( n343 & n442 ) | ( ~n441 & n442 ) ;
  assign n444 = n441 | n443 ;
  assign n445 = ( n57 & n87 ) | ( n57 & n104 ) | ( n87 & n104 ) ;
  assign n446 = n251 | n445 ;
  assign n447 = n87 & n163 ;
  assign n448 = n446 | n447 ;
  assign n449 = n136 & n141 ;
  assign n450 = ( n115 & n206 ) | ( n115 & n378 ) | ( n206 & n378 ) ;
  assign n451 = ( ~n448 & n449 ) | ( ~n448 & n450 ) | ( n449 & n450 ) ;
  assign n452 = n448 | n451 ;
  assign n453 = ( n438 & ~n444 ) | ( n438 & n452 ) | ( ~n444 & n452 ) ;
  assign n454 = n308 | n339 ;
  assign n455 = ( n80 & n83 ) | ( n80 & n105 ) | ( n83 & n105 ) ;
  assign n456 = ( n56 & n116 ) | ( n56 & n227 ) | ( n116 & n227 ) ;
  assign n457 = ( n454 & ~n455 ) | ( n454 & n456 ) | ( ~n455 & n456 ) ;
  assign n458 = n78 & n141 ;
  assign n459 = ( ~n202 & n314 ) | ( ~n202 & n458 ) | ( n314 & n458 ) ;
  assign n460 = n203 | n459 ;
  assign n461 = ( n455 & ~n457 ) | ( n455 & n460 ) | ( ~n457 & n460 ) ;
  assign n462 = n457 | n461 ;
  assign n463 = ( n444 & ~n453 ) | ( n444 & n462 ) | ( ~n453 & n462 ) ;
  assign n464 = n453 | n463 ;
  assign n465 = ( n425 & n431 ) | ( n425 & n464 ) | ( n431 & n464 ) ;
  assign n466 = n431 & ~n465 ;
  assign n467 = n115 & n202 ;
  assign n468 = n56 & n132 ;
  assign n469 = ( n132 & n467 ) | ( n132 & ~n468 ) | ( n467 & ~n468 ) ;
  assign n470 = n164 | n469 ;
  assign n471 = n78 & n202 ;
  assign n472 = ( n98 & n131 ) | ( n98 & n141 ) | ( n131 & n141 ) ;
  assign n473 = n471 | n472 ;
  assign n474 = ( n307 & ~n470 ) | ( n307 & n473 ) | ( ~n470 & n473 ) ;
  assign n475 = n470 | n474 ;
  assign n476 = ( n415 & n466 ) | ( n415 & ~n475 ) | ( n466 & ~n475 ) ;
  assign n477 = ~n415 & n476 ;
  assign n478 = ( n304 & n393 ) | ( n304 & n477 ) | ( n393 & n477 ) ;
  assign n479 = ( ~x22 & n32 ) | ( ~x22 & n33 ) | ( n32 & n33 ) ;
  assign n480 = x10 & x22 ;
  assign n481 = ( x9 & ~x22 ) | ( x9 & n32 ) | ( ~x22 & n32 ) ;
  assign n482 = x10 & n481 ;
  assign n483 = ( n479 & n480 ) | ( n479 & ~n482 ) | ( n480 & ~n482 ) ;
  assign n484 = ( ~n394 & n478 ) | ( ~n394 & n483 ) | ( n478 & n483 ) ;
  assign n485 = n304 & n393 ;
  assign n486 = ( n478 & n483 ) | ( n478 & ~n485 ) | ( n483 & ~n485 ) ;
  assign n487 = x9 & ~x22 ;
  assign n488 = x9 & ~n32 ;
  assign n489 = ( n481 & ~n487 ) | ( n481 & n488 ) | ( ~n487 & n488 ) ;
  assign n490 = n394 & ~n477 ;
  assign n491 = ( n477 & ~n485 ) | ( n477 & n490 ) | ( ~n485 & n490 ) ;
  assign n492 = n489 & ~n491 ;
  assign n493 = ( n394 & ~n485 ) | ( n394 & n490 ) | ( ~n485 & n490 ) ;
  assign n494 = ~n489 & n493 ;
  assign n495 = ( n489 & ~n492 ) | ( n489 & n494 ) | ( ~n492 & n494 ) ;
  assign n496 = ( n484 & ~n486 ) | ( n484 & n495 ) | ( ~n486 & n495 ) ;
  assign n497 = ( x5 & ~x22 ) | ( x5 & n28 ) | ( ~x22 & n28 ) ;
  assign n498 = x5 & ~n28 ;
  assign n499 = x5 & ~x22 ;
  assign n500 = ( n497 & n498 ) | ( n497 & ~n499 ) | ( n498 & ~n499 ) ;
  assign n501 = ( n57 & n126 ) | ( n57 & n136 ) | ( n126 & n136 ) ;
  assign n502 = ~n56 & n408 ;
  assign n503 = n111 & ~n174 ;
  assign n504 = n228 | n503 ;
  assign n505 = ( n88 & ~n502 ) | ( n88 & n504 ) | ( ~n502 & n504 ) ;
  assign n506 = n502 | n505 ;
  assign n507 = ( n172 & ~n501 ) | ( n172 & n506 ) | ( ~n501 & n506 ) ;
  assign n508 = n501 | n507 ;
  assign n509 = n80 & n206 ;
  assign n510 = ( n73 & n78 ) | ( n73 & n83 ) | ( n78 & n83 ) ;
  assign n511 = ( n426 & ~n509 ) | ( n426 & n510 ) | ( ~n509 & n510 ) ;
  assign n512 = n509 | n511 ;
  assign n513 = ( n164 & n305 ) | ( n164 & ~n512 ) | ( n305 & ~n512 ) ;
  assign n514 = n512 | n513 ;
  assign n515 = ( n73 & n141 ) | ( n73 & n363 ) | ( n141 & n363 ) ;
  assign n516 = ( n85 & n347 ) | ( n85 & ~n515 ) | ( n347 & ~n515 ) ;
  assign n517 = n515 | n516 ;
  assign n518 = ( ~n508 & n514 ) | ( ~n508 & n517 ) | ( n514 & n517 ) ;
  assign n519 = n508 | n518 ;
  assign n520 = n104 & n107 ;
  assign n521 = ( n126 & n141 ) | ( n126 & n283 ) | ( n141 & n283 ) ;
  assign n522 = n520 | n521 ;
  assign n523 = ( n98 & ~n119 ) | ( n98 & n202 ) | ( ~n119 & n202 ) ;
  assign n524 = n250 | n523 ;
  assign n525 = n522 | n524 ;
  assign n526 = n56 & n173 ;
  assign n527 = ( n308 & n315 ) | ( n308 & ~n526 ) | ( n315 & ~n526 ) ;
  assign n528 = n526 | n527 ;
  assign n529 = n131 & ~n174 ;
  assign n530 = n256 | n529 ;
  assign n531 = ( n468 & ~n528 ) | ( n468 & n530 ) | ( ~n528 & n530 ) ;
  assign n532 = n528 | n531 ;
  assign n533 = n105 & n163 ;
  assign n534 = n237 | n371 ;
  assign n535 = n533 | n534 ;
  assign n536 = ( n525 & ~n532 ) | ( n525 & n535 ) | ( ~n532 & n535 ) ;
  assign n537 = ( n224 & n352 ) | ( n224 & ~n386 ) | ( n352 & ~n386 ) ;
  assign n538 = n78 & n163 ;
  assign n539 = n252 | n538 ;
  assign n540 = ( n374 & ~n537 ) | ( n374 & n539 ) | ( ~n537 & n539 ) ;
  assign n541 = n537 | n540 ;
  assign n542 = ( n78 & n107 ) | ( n78 & n214 ) | ( n107 & n214 ) ;
  assign n543 = n150 | n294 ;
  assign n544 = ( n330 & ~n542 ) | ( n330 & n543 ) | ( ~n542 & n543 ) ;
  assign n545 = n542 | n544 ;
  assign n546 = ( n98 & n107 ) | ( n98 & n163 ) | ( n107 & n163 ) ;
  assign n547 = n246 | n546 ;
  assign n548 = ( n73 & n87 ) | ( n73 & ~n174 ) | ( n87 & ~n174 ) ;
  assign n549 = ( n112 & ~n547 ) | ( n112 & n548 ) | ( ~n547 & n548 ) ;
  assign n550 = n547 | n549 ;
  assign n551 = ( ~n541 & n545 ) | ( ~n541 & n550 ) | ( n545 & n550 ) ;
  assign n552 = n541 | n551 ;
  assign n553 = ( n100 & n338 ) | ( n100 & n386 ) | ( n338 & n386 ) ;
  assign n554 = ( n83 & n98 ) | ( n83 & n234 ) | ( n98 & n234 ) ;
  assign n555 = n441 | n554 ;
  assign n556 = ( n136 & ~n174 ) | ( n136 & n184 ) | ( ~n174 & n184 ) ;
  assign n557 = ( ~n553 & n555 ) | ( ~n553 & n556 ) | ( n555 & n556 ) ;
  assign n558 = n553 | n557 ;
  assign n559 = ( ~n532 & n552 ) | ( ~n532 & n558 ) | ( n552 & n558 ) ;
  assign n560 = n532 | n559 ;
  assign n561 = ( ~n519 & n536 ) | ( ~n519 & n560 ) | ( n536 & n560 ) ;
  assign n562 = n519 | n561 ;
  assign n563 = n89 | n371 ;
  assign n564 = ( n105 & n111 ) | ( n105 & n206 ) | ( n111 & n206 ) ;
  assign n565 = n91 & n141 ;
  assign n566 = ( ~n563 & n564 ) | ( ~n563 & n565 ) | ( n564 & n565 ) ;
  assign n567 = n563 | n566 ;
  assign n568 = ( n104 & n111 ) | ( n104 & n202 ) | ( n111 & n202 ) ;
  assign n569 = n56 & n378 ;
  assign n570 = ( n378 & n568 ) | ( n378 & ~n569 ) | ( n568 & ~n569 ) ;
  assign n571 = ( n327 & n380 ) | ( n327 & ~n570 ) | ( n380 & ~n570 ) ;
  assign n572 = n570 | n571 ;
  assign n573 = ( n78 & n91 ) | ( n78 & n107 ) | ( n91 & n107 ) ;
  assign n574 = ( n98 & n126 ) | ( n98 & n202 ) | ( n126 & n202 ) ;
  assign n575 = ( n56 & n378 ) | ( n56 & n447 ) | ( n378 & n447 ) ;
  assign n576 = ( n166 & ~n574 ) | ( n166 & n575 ) | ( ~n574 & n575 ) ;
  assign n577 = ( ~n573 & n574 ) | ( ~n573 & n576 ) | ( n574 & n576 ) ;
  assign n578 = n573 | n577 ;
  assign n579 = ( ~n567 & n572 ) | ( ~n567 & n578 ) | ( n572 & n578 ) ;
  assign n580 = n567 | n579 ;
  assign n581 = ( n305 & n467 ) | ( n305 & ~n580 ) | ( n467 & ~n580 ) ;
  assign n582 = n580 | n581 ;
  assign n583 = ( ~n56 & n234 ) | ( ~n56 & n237 ) | ( n234 & n237 ) ;
  assign n584 = ( n105 & n134 ) | ( n105 & n163 ) | ( n134 & n163 ) ;
  assign n585 = n583 | n584 ;
  assign n586 = ( n204 & ~n352 ) | ( n204 & n432 ) | ( ~n352 & n432 ) ;
  assign n587 = n154 | n310 ;
  assign n588 = ( n257 & n283 ) | ( n257 & ~n284 ) | ( n283 & ~n284 ) ;
  assign n589 = ( ~n321 & n587 ) | ( ~n321 & n588 ) | ( n587 & n588 ) ;
  assign n590 = ( n321 & ~n586 ) | ( n321 & n589 ) | ( ~n586 & n589 ) ;
  assign n591 = n586 | n590 ;
  assign n592 = n170 | n255 ;
  assign n593 = ( n297 & n347 ) | ( n297 & ~n592 ) | ( n347 & ~n592 ) ;
  assign n594 = n592 | n593 ;
  assign n595 = ( ~n585 & n591 ) | ( ~n585 & n594 ) | ( n591 & n594 ) ;
  assign n596 = ( n57 & n73 ) | ( n57 & n163 ) | ( n73 & n163 ) ;
  assign n597 = n122 | n449 ;
  assign n598 = n596 | n597 ;
  assign n599 = ( n111 & n141 ) | ( n111 & ~n174 ) | ( n141 & ~n174 ) ;
  assign n600 = ( ~n284 & n386 ) | ( ~n284 & n599 ) | ( n386 & n599 ) ;
  assign n601 = ( ~n56 & n214 ) | ( ~n56 & n315 ) | ( n214 & n315 ) ;
  assign n602 = n56 & n283 ;
  assign n603 = ( n283 & n601 ) | ( n283 & ~n602 ) | ( n601 & ~n602 ) ;
  assign n604 = ( n56 & n116 ) | ( n56 & n408 ) | ( n116 & n408 ) ;
  assign n605 = ( n243 & ~n275 ) | ( n243 & n604 ) | ( ~n275 & n604 ) ;
  assign n606 = ( n600 & ~n603 ) | ( n600 & n605 ) | ( ~n603 & n605 ) ;
  assign n607 = ( n83 & n136 ) | ( n83 & ~n174 ) | ( n136 & ~n174 ) ;
  assign n608 = n410 | n607 ;
  assign n609 = n126 & n206 ;
  assign n610 = n84 & n202 ;
  assign n611 = n127 | n610 ;
  assign n612 = n609 | n611 ;
  assign n613 = ( ~n603 & n608 ) | ( ~n603 & n612 ) | ( n608 & n612 ) ;
  assign n614 = n603 | n613 ;
  assign n615 = ( ~n598 & n606 ) | ( ~n598 & n614 ) | ( n606 & n614 ) ;
  assign n616 = n598 | n615 ;
  assign n617 = n104 & n141 ;
  assign n618 = n105 & ~n174 ;
  assign n619 = n617 | n618 ;
  assign n620 = ( n84 & n104 ) | ( n84 & ~n174 ) | ( n104 & ~n174 ) ;
  assign n621 = n269 | n620 ;
  assign n622 = ( n248 & ~n619 ) | ( n248 & n621 ) | ( ~n619 & n621 ) ;
  assign n623 = n619 | n622 ;
  assign n624 = n501 | n623 ;
  assign n625 = ( n585 & ~n616 ) | ( n585 & n624 ) | ( ~n616 & n624 ) ;
  assign n626 = n616 | n625 ;
  assign n627 = ( ~n582 & n595 ) | ( ~n582 & n626 ) | ( n595 & n626 ) ;
  assign n628 = n582 | n627 ;
  assign n629 = n562 & n628 ;
  assign n630 = n562 | n628 ;
  assign n631 = ~n629 & n630 ;
  assign n632 = n270 | n314 ;
  assign n633 = n121 | n359 ;
  assign n634 = ( n84 & n115 ) | ( n84 & n202 ) | ( n115 & n202 ) ;
  assign n635 = ( n378 & ~n379 ) | ( n378 & n634 ) | ( ~n379 & n634 ) ;
  assign n636 = ( ~n632 & n633 ) | ( ~n632 & n635 ) | ( n633 & n635 ) ;
  assign n637 = n632 | n636 ;
  assign n638 = n232 | n397 ;
  assign n639 = n311 | n529 ;
  assign n640 = ( ~n275 & n342 ) | ( ~n275 & n639 ) | ( n342 & n639 ) ;
  assign n641 = n275 | n640 ;
  assign n642 = n170 | n410 ;
  assign n643 = ( n245 & ~n641 ) | ( n245 & n642 ) | ( ~n641 & n642 ) ;
  assign n644 = n641 | n643 ;
  assign n645 = ( ~n637 & n638 ) | ( ~n637 & n644 ) | ( n638 & n644 ) ;
  assign n646 = n637 | n645 ;
  assign n647 = n85 | n565 ;
  assign n648 = ( ~n56 & n237 ) | ( ~n56 & n305 ) | ( n237 & n305 ) ;
  assign n649 = n56 & n214 ;
  assign n650 = n648 | n649 ;
  assign n651 = n647 | n650 ;
  assign n652 = ( n83 & n115 ) | ( n83 & ~n119 ) | ( n115 & ~n119 ) ;
  assign n653 = n252 | n652 ;
  assign n654 = n449 | n618 ;
  assign n655 = ( n91 & n107 ) | ( n91 & n136 ) | ( n107 & n136 ) ;
  assign n656 = n57 & n134 ;
  assign n657 = ( n128 & ~n655 ) | ( n128 & n656 ) | ( ~n655 & n656 ) ;
  assign n658 = n655 | n657 ;
  assign n659 = ( ~n653 & n654 ) | ( ~n653 & n658 ) | ( n654 & n658 ) ;
  assign n660 = ( ~n223 & n653 ) | ( ~n223 & n659 ) | ( n653 & n659 ) ;
  assign n661 = n56 & n106 ;
  assign n662 = n116 | n661 ;
  assign n663 = n341 | n473 ;
  assign n664 = ( n509 & ~n662 ) | ( n509 & n663 ) | ( ~n662 & n663 ) ;
  assign n665 = n662 | n664 ;
  assign n666 = ( n223 & ~n651 ) | ( n223 & n665 ) | ( ~n651 & n665 ) ;
  assign n667 = ( n651 & ~n660 ) | ( n651 & n666 ) | ( ~n660 & n666 ) ;
  assign n668 = ( n84 & n206 ) | ( n84 & n378 ) | ( n206 & n378 ) ;
  assign n669 = n111 & n202 ;
  assign n670 = n447 | n669 ;
  assign n671 = ( n269 & ~n668 ) | ( n269 & n670 ) | ( ~n668 & n670 ) ;
  assign n672 = n668 | n671 ;
  assign n673 = n328 | n538 ;
  assign n674 = ( n237 & ~n271 ) | ( n237 & n387 ) | ( ~n271 & n387 ) ;
  assign n675 = ( n73 & n87 ) | ( n73 & n202 ) | ( n87 & n202 ) ;
  assign n676 = n433 | n675 ;
  assign n677 = n674 | n676 ;
  assign n678 = ( ~n672 & n673 ) | ( ~n672 & n677 ) | ( n673 & n677 ) ;
  assign n679 = n672 | n678 ;
  assign n680 = ( n151 & n329 ) | ( n151 & ~n679 ) | ( n329 & ~n679 ) ;
  assign n681 = n679 | n680 ;
  assign n682 = n266 | n587 ;
  assign n683 = n90 | n682 ;
  assign n684 = ( ~n660 & n681 ) | ( ~n660 & n683 ) | ( n681 & n683 ) ;
  assign n685 = ( n660 & ~n667 ) | ( n660 & n684 ) | ( ~n667 & n684 ) ;
  assign n686 = ( ~n646 & n667 ) | ( ~n646 & n685 ) | ( n667 & n685 ) ;
  assign n687 = n646 | n686 ;
  assign n688 = ( ~x22 & n28 ) | ( ~x22 & n29 ) | ( n28 & n29 ) ;
  assign n689 = x6 & x22 ;
  assign n690 = x6 & n497 ;
  assign n691 = ( n688 & n689 ) | ( n688 & ~n690 ) | ( n689 & ~n690 ) ;
  assign n692 = ( n631 & n687 ) | ( n631 & ~n691 ) | ( n687 & ~n691 ) ;
  assign n693 = ( n631 & ~n687 ) | ( n631 & n691 ) | ( ~n687 & n691 ) ;
  assign n694 = n692 & n693 ;
  assign n695 = ~n629 & n687 ;
  assign n696 = ( ~n629 & n630 ) | ( ~n629 & n695 ) | ( n630 & n695 ) ;
  assign n697 = ( n500 & ~n694 ) | ( n500 & n696 ) | ( ~n694 & n696 ) ;
  assign n698 = ( n630 & n631 ) | ( n630 & ~n687 ) | ( n631 & ~n687 ) ;
  assign n699 = ( n500 & n694 ) | ( n500 & ~n698 ) | ( n694 & ~n698 ) ;
  assign n700 = n697 & ~n699 ;
  assign n701 = ( ~x22 & n30 ) | ( ~x22 & n31 ) | ( n30 & n31 ) ;
  assign n702 = x8 & x22 ;
  assign n703 = ( x7 & ~x22 ) | ( x7 & n30 ) | ( ~x22 & n30 ) ;
  assign n704 = x8 & n703 ;
  assign n705 = ( n701 & n702 ) | ( n701 & ~n704 ) | ( n702 & ~n704 ) ;
  assign n706 = n562 & ~n705 ;
  assign n707 = n275 | n509 ;
  assign n708 = ( n80 & n87 ) | ( n80 & ~n174 ) | ( n87 & ~n174 ) ;
  assign n709 = n428 | n520 ;
  assign n710 = n642 | n709 ;
  assign n711 = ( ~n288 & n583 ) | ( ~n288 & n710 ) | ( n583 & n710 ) ;
  assign n712 = n471 | n609 ;
  assign n713 = n189 | n712 ;
  assign n714 = ( n115 & n206 ) | ( n115 & n314 ) | ( n206 & n314 ) ;
  assign n715 = ~n56 & n243 ;
  assign n716 = n656 | n715 ;
  assign n717 = n714 | n716 ;
  assign n718 = ( n399 & ~n713 ) | ( n399 & n717 ) | ( ~n713 & n717 ) ;
  assign n719 = n713 | n718 ;
  assign n720 = ( n288 & ~n711 ) | ( n288 & n719 ) | ( ~n711 & n719 ) ;
  assign n721 = n711 | n720 ;
  assign n722 = ( ~n707 & n708 ) | ( ~n707 & n721 ) | ( n708 & n721 ) ;
  assign n723 = n707 | n722 ;
  assign n724 = n315 | n432 ;
  assign n725 = n142 | n265 ;
  assign n726 = ( n84 & n163 ) | ( n84 & n173 ) | ( n163 & n173 ) ;
  assign n727 = ( n724 & n725 ) | ( n724 & ~n726 ) | ( n725 & ~n726 ) ;
  assign n728 = ( n354 & n726 ) | ( n354 & ~n727 ) | ( n726 & ~n727 ) ;
  assign n729 = n727 | n728 ;
  assign n730 = n723 | n729 ;
  assign n731 = ( n73 & n107 ) | ( n73 & n276 ) | ( n107 & n276 ) ;
  assign n732 = n226 | n387 ;
  assign n733 = n731 | n732 ;
  assign n734 = ( n57 & n73 ) | ( n57 & n132 ) | ( n73 & n132 ) ;
  assign n735 = ( n106 & ~n128 ) | ( n106 & n734 ) | ( ~n128 & n734 ) ;
  assign n736 = n380 | n395 ;
  assign n737 = ( n151 & n214 ) | ( n151 & ~n649 ) | ( n214 & ~n649 ) ;
  assign n738 = ( n294 & n669 ) | ( n294 & ~n737 ) | ( n669 & ~n737 ) ;
  assign n739 = n737 | n738 ;
  assign n740 = ( ~n735 & n736 ) | ( ~n735 & n739 ) | ( n736 & n739 ) ;
  assign n741 = n735 | n740 ;
  assign n742 = ( n132 & n250 ) | ( n132 & ~n468 ) | ( n250 & ~n468 ) ;
  assign n743 = n342 | n742 ;
  assign n744 = ( n253 & n529 ) | ( n253 & ~n743 ) | ( n529 & ~n743 ) ;
  assign n745 = n743 | n744 ;
  assign n746 = ( ~n578 & n741 ) | ( ~n578 & n745 ) | ( n741 & n745 ) ;
  assign n747 = ( n578 & ~n733 ) | ( n578 & n746 ) | ( ~n733 & n746 ) ;
  assign n748 = ( ~n730 & n733 ) | ( ~n730 & n747 ) | ( n733 & n747 ) ;
  assign n749 = n730 | n748 ;
  assign n750 = n477 & ~n749 ;
  assign n751 = ~n477 & n749 ;
  assign n752 = n750 | n751 ;
  assign n753 = ( ~n562 & n705 ) | ( ~n562 & n752 ) | ( n705 & n752 ) ;
  assign n754 = x7 & x22 ;
  assign n755 = x7 & n30 ;
  assign n756 = ( n703 & n754 ) | ( n703 & ~n755 ) | ( n754 & ~n755 ) ;
  assign n757 = n562 & ~n756 ;
  assign n758 = n562 & ~n751 ;
  assign n759 = ( n562 & n750 ) | ( n562 & ~n758 ) | ( n750 & ~n758 ) ;
  assign n760 = n751 & ~n756 ;
  assign n761 = ( ~n757 & n759 ) | ( ~n757 & n760 ) | ( n759 & n760 ) ;
  assign n762 = ( n706 & n753 ) | ( n706 & ~n761 ) | ( n753 & ~n761 ) ;
  assign n763 = ( n496 & n700 ) | ( n496 & n762 ) | ( n700 & n762 ) ;
  assign n764 = ( n78 & n163 ) | ( n78 & n173 ) | ( n163 & n173 ) ;
  assign n765 = ~n56 & n227 ;
  assign n766 = ( n227 & n432 ) | ( n227 & ~n765 ) | ( n432 & ~n765 ) ;
  assign n767 = ( ~n709 & n764 ) | ( ~n709 & n766 ) | ( n764 & n766 ) ;
  assign n768 = ( n612 & n709 ) | ( n612 & ~n767 ) | ( n709 & ~n767 ) ;
  assign n769 = n767 | n768 ;
  assign n770 = ( ~n386 & n617 ) | ( ~n386 & n769 ) | ( n617 & n769 ) ;
  assign n771 = n386 | n770 ;
  assign n772 = n120 | n278 ;
  assign n773 = ( n87 & n173 ) | ( n87 & ~n174 ) | ( n173 & ~n174 ) ;
  assign n774 = n382 | n773 ;
  assign n775 = ( n245 & ~n772 ) | ( n245 & n774 ) | ( ~n772 & n774 ) ;
  assign n776 = n772 | n775 ;
  assign n777 = n247 | n250 ;
  assign n778 = ( n275 & n310 ) | ( n275 & ~n777 ) | ( n310 & ~n777 ) ;
  assign n779 = n777 | n778 ;
  assign n780 = ( n340 & n411 ) | ( n340 & ~n779 ) | ( n411 & ~n779 ) ;
  assign n781 = n779 | n780 ;
  assign n782 = ( n332 & ~n776 ) | ( n332 & n781 ) | ( ~n776 & n781 ) ;
  assign n783 = n776 | n782 ;
  assign n784 = ( n51 & ~n57 ) | ( n51 & n104 ) | ( ~n57 & n104 ) ;
  assign n785 = ( n80 & n206 ) | ( n80 & n784 ) | ( n206 & n784 ) ;
  assign n786 = ~n119 & n202 ;
  assign n787 = n765 | n786 ;
  assign n788 = ( n256 & n311 ) | ( n256 & ~n786 ) | ( n311 & ~n786 ) ;
  assign n789 = n787 | n788 ;
  assign n790 = n128 | n253 ;
  assign n791 = n142 | n422 ;
  assign n792 = n211 | n246 ;
  assign n793 = ( ~n790 & n791 ) | ( ~n790 & n792 ) | ( n791 & n792 ) ;
  assign n794 = n790 | n793 ;
  assign n795 = ( ~n785 & n789 ) | ( ~n785 & n794 ) | ( n789 & n794 ) ;
  assign n796 = n78 & n83 ;
  assign n797 = n252 | n796 ;
  assign n798 = ( n170 & ~n502 ) | ( n170 & n797 ) | ( ~n502 & n797 ) ;
  assign n799 = n502 | n798 ;
  assign n800 = n364 | n503 ;
  assign n801 = ( ~n206 & n229 ) | ( ~n206 & n408 ) | ( n229 & n408 ) ;
  assign n802 = ( n78 & n201 ) | ( n78 & n801 ) | ( n201 & n801 ) ;
  assign n803 = ( ~n799 & n800 ) | ( ~n799 & n802 ) | ( n800 & n802 ) ;
  assign n804 = n799 | n803 ;
  assign n805 = ( n785 & n795 ) | ( n785 & ~n804 ) | ( n795 & ~n804 ) ;
  assign n806 = ( n582 & n804 ) | ( n582 & ~n805 ) | ( n804 & ~n805 ) ;
  assign n807 = n805 | n806 ;
  assign n808 = ( ~n771 & n783 ) | ( ~n771 & n807 ) | ( n783 & n807 ) ;
  assign n809 = n771 | n808 ;
  assign n810 = n687 & n809 ;
  assign n811 = n192 & ~n810 ;
  assign n812 = n687 | n809 ;
  assign n813 = ~n810 & n812 ;
  assign n814 = n199 & n813 ;
  assign n815 = n811 & ~n814 ;
  assign n816 = x22 | n35 ;
  assign n817 = ( x12 & x22 ) | ( x12 & n816 ) | ( x22 & n816 ) ;
  assign n818 = ( x12 & x22 ) | ( x12 & ~n816 ) | ( x22 & ~n816 ) ;
  assign n819 = ( n816 & ~n817 ) | ( n816 & n818 ) | ( ~n817 & n818 ) ;
  assign n820 = ( n224 & ~n386 ) | ( n224 & n449 ) | ( ~n386 & n449 ) ;
  assign n821 = ( n84 & n201 ) | ( n84 & n379 ) | ( n201 & n379 ) ;
  assign n822 = ( n283 & ~n284 ) | ( n283 & n386 ) | ( ~n284 & n386 ) ;
  assign n823 = ( ~n820 & n821 ) | ( ~n820 & n822 ) | ( n821 & n822 ) ;
  assign n824 = n820 | n823 ;
  assign n825 = n92 | n427 ;
  assign n826 = n792 | n800 ;
  assign n827 = n825 | n826 ;
  assign n828 = ( n154 & ~n715 ) | ( n154 & n765 ) | ( ~n715 & n765 ) ;
  assign n829 = n715 | n828 ;
  assign n830 = ( ~n824 & n827 ) | ( ~n824 & n829 ) | ( n827 & n829 ) ;
  assign n831 = n824 | n830 ;
  assign n832 = ( n56 & n106 ) | ( n56 & n447 ) | ( n106 & n447 ) ;
  assign n833 = n221 & ~n832 ;
  assign n834 = ~n791 & n833 ;
  assign n835 = n85 | n170 ;
  assign n836 = ( n73 & n83 ) | ( n73 & ~n119 ) | ( n83 & ~n119 ) ;
  assign n837 = ( n834 & n835 ) | ( n834 & n836 ) | ( n835 & n836 ) ;
  assign n838 = n834 & ~n837 ;
  assign n839 = ~n831 & n838 ;
  assign n840 = ( ~n56 & n173 ) | ( ~n56 & n283 ) | ( n173 & n283 ) ;
  assign n841 = ( n395 & ~n658 ) | ( n395 & n840 ) | ( ~n658 & n840 ) ;
  assign n842 = n471 | n601 ;
  assign n843 = ( n509 & n568 ) | ( n509 & ~n786 ) | ( n568 & ~n786 ) ;
  assign n844 = n786 | n843 ;
  assign n845 = ( n353 & n772 ) | ( n353 & ~n844 ) | ( n772 & ~n844 ) ;
  assign n846 = n844 | n845 ;
  assign n847 = ( n658 & ~n842 ) | ( n658 & n846 ) | ( ~n842 & n846 ) ;
  assign n848 = ( ~n841 & n842 ) | ( ~n841 & n847 ) | ( n842 & n847 ) ;
  assign n849 = n841 | n848 ;
  assign n850 = ( n122 & n227 ) | ( n122 & ~n765 ) | ( n227 & ~n765 ) ;
  assign n851 = n116 | n220 ;
  assign n852 = ( n223 & n342 ) | ( n223 & ~n851 ) | ( n342 & ~n851 ) ;
  assign n853 = n851 | n852 ;
  assign n854 = ( n619 & ~n850 ) | ( n619 & n853 ) | ( ~n850 & n853 ) ;
  assign n855 = ( n416 & n850 ) | ( n416 & ~n854 ) | ( n850 & ~n854 ) ;
  assign n856 = n854 | n855 ;
  assign n857 = ( n839 & n849 ) | ( n839 & n856 ) | ( n849 & n856 ) ;
  assign n858 = n839 & ~n857 ;
  assign n859 = ( ~n304 & n819 ) | ( ~n304 & n858 ) | ( n819 & n858 ) ;
  assign n860 = ( x11 & ~x22 ) | ( x11 & n34 ) | ( ~x22 & n34 ) ;
  assign n861 = x11 & ~n34 ;
  assign n862 = x11 & ~x22 ;
  assign n863 = ( n860 & n861 ) | ( n860 & ~n862 ) | ( n861 & ~n862 ) ;
  assign n864 = n858 | n863 ;
  assign n865 = ( n859 & n863 ) | ( n859 & ~n864 ) | ( n863 & ~n864 ) ;
  assign n866 = n819 & n858 ;
  assign n867 = ( n304 & ~n819 ) | ( n304 & n866 ) | ( ~n819 & n866 ) ;
  assign n868 = n865 | n867 ;
  assign n869 = n815 & ~n868 ;
  assign n870 = ~n489 & n562 ;
  assign n871 = ( n489 & ~n562 ) | ( n489 & n752 ) | ( ~n562 & n752 ) ;
  assign n872 = ~n705 & n751 ;
  assign n873 = ( ~n706 & n759 ) | ( ~n706 & n872 ) | ( n759 & n872 ) ;
  assign n874 = ( n870 & n871 ) | ( n870 & ~n873 ) | ( n871 & ~n873 ) ;
  assign n875 = ( n631 & n687 ) | ( n631 & ~n756 ) | ( n687 & ~n756 ) ;
  assign n876 = ( n631 & ~n687 ) | ( n631 & n756 ) | ( ~n687 & n756 ) ;
  assign n877 = n875 & n876 ;
  assign n878 = ( n691 & n696 ) | ( n691 & ~n877 ) | ( n696 & ~n877 ) ;
  assign n879 = ( n691 & ~n698 ) | ( n691 & n877 ) | ( ~n698 & n877 ) ;
  assign n880 = n878 & ~n879 ;
  assign n881 = ( n869 & n874 ) | ( n869 & n880 ) | ( n874 & n880 ) ;
  assign n882 = ( ~n869 & n874 ) | ( ~n869 & n880 ) | ( n874 & n880 ) ;
  assign n883 = ( n869 & ~n881 ) | ( n869 & n882 ) | ( ~n881 & n882 ) ;
  assign n884 = ( n200 & n763 ) | ( n200 & n883 ) | ( n763 & n883 ) ;
  assign n885 = n115 | n126 ;
  assign n886 = ( n201 & n568 ) | ( n201 & n885 ) | ( n568 & n885 ) ;
  assign n887 = n339 | n569 ;
  assign n888 = n237 | n243 ;
  assign n889 = n887 | n888 ;
  assign n890 = n265 | n458 ;
  assign n891 = n207 | n890 ;
  assign n892 = n363 | n891 ;
  assign n893 = ( n73 & n206 ) | ( n73 & n227 ) | ( n206 & n227 ) ;
  assign n894 = n214 | n309 ;
  assign n895 = n342 | n509 ;
  assign n896 = ( n329 & ~n894 ) | ( n329 & n895 ) | ( ~n894 & n895 ) ;
  assign n897 = n894 | n896 ;
  assign n898 = ( ~n892 & n893 ) | ( ~n892 & n897 ) | ( n893 & n897 ) ;
  assign n899 = n892 | n898 ;
  assign n900 = ( n886 & n889 ) | ( n886 & ~n899 ) | ( n889 & ~n899 ) ;
  assign n901 = n338 | n428 ;
  assign n902 = n208 | n220 ;
  assign n903 = ( n87 & n98 ) | ( n87 & n206 ) | ( n98 & n206 ) ;
  assign n904 = ( n257 & n471 ) | ( n257 & ~n903 ) | ( n471 & ~n903 ) ;
  assign n905 = n903 | n904 ;
  assign n906 = ( n402 & ~n902 ) | ( n402 & n905 ) | ( ~n902 & n905 ) ;
  assign n907 = n902 | n906 ;
  assign n908 = ( n111 & n134 ) | ( n111 & n206 ) | ( n134 & n206 ) ;
  assign n909 = ( n408 & n439 ) | ( n408 & ~n502 ) | ( n439 & ~n502 ) ;
  assign n910 = n908 | n909 ;
  assign n911 = ( n296 & ~n901 ) | ( n296 & n910 ) | ( ~n901 & n910 ) ;
  assign n912 = ( ~n901 & n907 ) | ( ~n901 & n911 ) | ( n907 & n911 ) ;
  assign n913 = ( n107 & n136 ) | ( n107 & n283 ) | ( n136 & n283 ) ;
  assign n914 = n824 | n913 ;
  assign n915 = ( n901 & ~n912 ) | ( n901 & n914 ) | ( ~n912 & n914 ) ;
  assign n916 = n912 | n915 ;
  assign n917 = ( n899 & ~n900 ) | ( n899 & n916 ) | ( ~n900 & n916 ) ;
  assign n918 = n900 | n917 ;
  assign n919 = ( x4 & ~x22 ) | ( x4 & n27 ) | ( ~x22 & n27 ) ;
  assign n920 = x4 & ~n27 ;
  assign n921 = x4 & ~x22 ;
  assign n922 = ( n919 & n920 ) | ( n919 & ~n921 ) | ( n920 & ~n921 ) ;
  assign n923 = n918 & n922 ;
  assign n924 = ( n194 & n918 ) | ( n194 & ~n922 ) | ( n918 & ~n922 ) ;
  assign n925 = ( ~n918 & n923 ) | ( ~n918 & n924 ) | ( n923 & n924 ) ;
  assign n926 = ( ~n193 & n199 ) | ( ~n193 & n925 ) | ( n199 & n925 ) ;
  assign n927 = ( ~n149 & n194 ) | ( ~n149 & n918 ) | ( n194 & n918 ) ;
  assign n928 = ( n199 & ~n925 ) | ( n199 & n927 ) | ( ~n925 & n927 ) ;
  assign n929 = ~n926 & n928 ;
  assign n930 = ( ~n394 & n478 ) | ( ~n394 & n819 ) | ( n478 & n819 ) ;
  assign n931 = ( n478 & ~n485 ) | ( n478 & n819 ) | ( ~n485 & n819 ) ;
  assign n932 = ~n491 & n863 ;
  assign n933 = n493 & ~n863 ;
  assign n934 = ( n863 & ~n932 ) | ( n863 & n933 ) | ( ~n932 & n933 ) ;
  assign n935 = ( n930 & ~n931 ) | ( n930 & n934 ) | ( ~n931 & n934 ) ;
  assign n936 = ( x13 & ~x22 ) | ( x13 & n36 ) | ( ~x22 & n36 ) ;
  assign n937 = x13 & ~x22 ;
  assign n938 = x13 & ~n36 ;
  assign n939 = ( n936 & ~n937 ) | ( n936 & n938 ) | ( ~n937 & n938 ) ;
  assign n940 = n858 & n939 ;
  assign n941 = x14 & ~x22 ;
  assign n942 = x14 & ~n37 ;
  assign n943 = ( n54 & ~n941 ) | ( n54 & n942 ) | ( ~n941 & n942 ) ;
  assign n944 = ~n858 & n943 ;
  assign n945 = n304 & n944 ;
  assign n946 = ( n304 & ~n940 ) | ( n304 & n944 ) | ( ~n940 & n944 ) ;
  assign n947 = ( n940 & ~n945 ) | ( n940 & n946 ) | ( ~n945 & n946 ) ;
  assign n948 = n918 & ~n947 ;
  assign n949 = n918 & n947 ;
  assign n950 = ( n947 & n948 ) | ( n947 & ~n949 ) | ( n948 & ~n949 ) ;
  assign n951 = ( n929 & n935 ) | ( n929 & ~n950 ) | ( n935 & ~n950 ) ;
  assign n952 = ( n929 & ~n935 ) | ( n929 & n950 ) | ( ~n935 & n950 ) ;
  assign n953 = ( ~n929 & n951 ) | ( ~n929 & n952 ) | ( n951 & n952 ) ;
  assign n954 = ( ~n394 & n478 ) | ( ~n394 & n863 ) | ( n478 & n863 ) ;
  assign n955 = ( n478 & ~n485 ) | ( n478 & n863 ) | ( ~n485 & n863 ) ;
  assign n956 = n483 & ~n491 ;
  assign n957 = ~n483 & n493 ;
  assign n958 = ( n483 & ~n956 ) | ( n483 & n957 ) | ( ~n956 & n957 ) ;
  assign n959 = ( n954 & ~n955 ) | ( n954 & n958 ) | ( ~n955 & n958 ) ;
  assign n960 = ( n304 & n858 ) | ( n304 & n939 ) | ( n858 & n939 ) ;
  assign n961 = ~n858 & n960 ;
  assign n962 = ( n866 & n939 ) | ( n866 & ~n960 ) | ( n939 & ~n960 ) ;
  assign n963 = ( n304 & ~n961 ) | ( n304 & n962 ) | ( ~n961 & n962 ) ;
  assign n964 = ( ~n192 & n500 ) | ( ~n192 & n813 ) | ( n500 & n813 ) ;
  assign n965 = ( n192 & ~n500 ) | ( n192 & n813 ) | ( ~n500 & n813 ) ;
  assign n966 = n964 & n965 ;
  assign n967 = ( ~n810 & n811 ) | ( ~n810 & n812 ) | ( n811 & n812 ) ;
  assign n968 = ( n922 & ~n966 ) | ( n922 & n967 ) | ( ~n966 & n967 ) ;
  assign n969 = ( ~n192 & n812 ) | ( ~n192 & n813 ) | ( n812 & n813 ) ;
  assign n970 = ( n922 & n966 ) | ( n922 & ~n969 ) | ( n966 & ~n969 ) ;
  assign n971 = n968 & ~n970 ;
  assign n972 = ( n959 & ~n963 ) | ( n959 & n971 ) | ( ~n963 & n971 ) ;
  assign n973 = ( n192 & ~n691 ) | ( n192 & n813 ) | ( ~n691 & n813 ) ;
  assign n974 = ( ~n192 & n691 ) | ( ~n192 & n813 ) | ( n691 & n813 ) ;
  assign n975 = n973 & n974 ;
  assign n976 = ( n500 & n967 ) | ( n500 & ~n975 ) | ( n967 & ~n975 ) ;
  assign n977 = ( n500 & ~n969 ) | ( n500 & n975 ) | ( ~n969 & n975 ) ;
  assign n978 = n976 & ~n977 ;
  assign n979 = ( n631 & n687 ) | ( n631 & ~n705 ) | ( n687 & ~n705 ) ;
  assign n980 = ( n631 & ~n687 ) | ( n631 & n705 ) | ( ~n687 & n705 ) ;
  assign n981 = n979 & n980 ;
  assign n982 = ( n696 & n756 ) | ( n696 & ~n981 ) | ( n756 & ~n981 ) ;
  assign n983 = ( ~n698 & n756 ) | ( ~n698 & n981 ) | ( n756 & n981 ) ;
  assign n984 = n982 & ~n983 ;
  assign n985 = ( n483 & ~n562 ) | ( n483 & n752 ) | ( ~n562 & n752 ) ;
  assign n986 = ~n483 & n562 ;
  assign n987 = ~n489 & n751 ;
  assign n988 = ( n759 & ~n870 ) | ( n759 & n987 ) | ( ~n870 & n987 ) ;
  assign n989 = ( n985 & n986 ) | ( n985 & ~n988 ) | ( n986 & ~n988 ) ;
  assign n990 = ( n978 & n984 ) | ( n978 & n989 ) | ( n984 & n989 ) ;
  assign n991 = ( ~n978 & n984 ) | ( ~n978 & n989 ) | ( n984 & n989 ) ;
  assign n992 = ( n978 & ~n990 ) | ( n978 & n991 ) | ( ~n990 & n991 ) ;
  assign n993 = ( n881 & n972 ) | ( n881 & n992 ) | ( n972 & n992 ) ;
  assign n994 = ( n881 & ~n972 ) | ( n881 & n992 ) | ( ~n972 & n992 ) ;
  assign n995 = ( n972 & ~n993 ) | ( n972 & n994 ) | ( ~n993 & n994 ) ;
  assign n996 = ( n884 & ~n953 ) | ( n884 & n995 ) | ( ~n953 & n995 ) ;
  assign n997 = ( ~n394 & n478 ) | ( ~n394 & n489 ) | ( n478 & n489 ) ;
  assign n998 = ( n478 & ~n485 ) | ( n478 & n489 ) | ( ~n485 & n489 ) ;
  assign n999 = ~n491 & n705 ;
  assign n1000 = n493 & ~n705 ;
  assign n1001 = ( n705 & ~n999 ) | ( n705 & n1000 ) | ( ~n999 & n1000 ) ;
  assign n1002 = ( n997 & ~n998 ) | ( n997 & n1001 ) | ( ~n998 & n1001 ) ;
  assign n1003 = ~n483 & n858 ;
  assign n1004 = ( n304 & n858 ) | ( n304 & ~n864 ) | ( n858 & ~n864 ) ;
  assign n1005 = ( ~n304 & n858 ) | ( ~n304 & n864 ) | ( n858 & n864 ) ;
  assign n1006 = ( ~n1003 & n1004 ) | ( ~n1003 & n1005 ) | ( n1004 & n1005 ) ;
  assign n1007 = ( ~n562 & n752 ) | ( ~n562 & n756 ) | ( n752 & n756 ) ;
  assign n1008 = n562 & ~n691 ;
  assign n1009 = ~n691 & n751 ;
  assign n1010 = ( n759 & ~n1008 ) | ( n759 & n1009 ) | ( ~n1008 & n1009 ) ;
  assign n1011 = ( n757 & n1007 ) | ( n757 & ~n1010 ) | ( n1007 & ~n1010 ) ;
  assign n1012 = ( n1002 & ~n1006 ) | ( n1002 & n1011 ) | ( ~n1006 & n1011 ) ;
  assign n1013 = n815 & n868 ;
  assign n1014 = ( n868 & n869 ) | ( n868 & ~n1013 ) | ( n869 & ~n1013 ) ;
  assign n1015 = ( ~n192 & n813 ) | ( ~n192 & n922 ) | ( n813 & n922 ) ;
  assign n1016 = ( n192 & n813 ) | ( n192 & ~n922 ) | ( n813 & ~n922 ) ;
  assign n1017 = n1015 & n1016 ;
  assign n1018 = ( n199 & n967 ) | ( n199 & ~n1017 ) | ( n967 & ~n1017 ) ;
  assign n1019 = ( n199 & ~n969 ) | ( n199 & n1017 ) | ( ~n969 & n1017 ) ;
  assign n1020 = n1018 & ~n1019 ;
  assign n1021 = ( n1012 & ~n1014 ) | ( n1012 & n1020 ) | ( ~n1014 & n1020 ) ;
  assign n1022 = ( ~n959 & n963 ) | ( ~n959 & n971 ) | ( n963 & n971 ) ;
  assign n1023 = ( ~n971 & n972 ) | ( ~n971 & n1022 ) | ( n972 & n1022 ) ;
  assign n1024 = ( n200 & ~n763 ) | ( n200 & n883 ) | ( ~n763 & n883 ) ;
  assign n1025 = ( n763 & ~n884 ) | ( n763 & n1024 ) | ( ~n884 & n1024 ) ;
  assign n1026 = ( n1021 & ~n1023 ) | ( n1021 & n1025 ) | ( ~n1023 & n1025 ) ;
  assign n1027 = n199 & n631 ;
  assign n1028 = n695 & ~n1027 ;
  assign n1029 = ( ~n304 & n483 ) | ( ~n304 & n858 ) | ( n483 & n858 ) ;
  assign n1030 = n483 & ~n1029 ;
  assign n1031 = n489 | n858 ;
  assign n1032 = ( n489 & n1029 ) | ( n489 & ~n1031 ) | ( n1029 & ~n1031 ) ;
  assign n1033 = ( n304 & ~n1030 ) | ( n304 & n1032 ) | ( ~n1030 & n1032 ) ;
  assign n1034 = n1028 & ~n1033 ;
  assign n1035 = ( n500 & n631 ) | ( n500 & ~n687 ) | ( n631 & ~n687 ) ;
  assign n1036 = ( ~n500 & n631 ) | ( ~n500 & n687 ) | ( n631 & n687 ) ;
  assign n1037 = n1035 & n1036 ;
  assign n1038 = ( n696 & n922 ) | ( n696 & ~n1037 ) | ( n922 & ~n1037 ) ;
  assign n1039 = ( ~n698 & n922 ) | ( ~n698 & n1037 ) | ( n922 & n1037 ) ;
  assign n1040 = n1038 & ~n1039 ;
  assign n1041 = ( n814 & n1034 ) | ( n814 & n1040 ) | ( n1034 & n1040 ) ;
  assign n1042 = ( n496 & ~n700 ) | ( n496 & n762 ) | ( ~n700 & n762 ) ;
  assign n1043 = ( n700 & ~n763 ) | ( n700 & n1042 ) | ( ~n763 & n1042 ) ;
  assign n1044 = ( ~n1012 & n1014 ) | ( ~n1012 & n1020 ) | ( n1014 & n1020 ) ;
  assign n1045 = ( ~n1020 & n1021 ) | ( ~n1020 & n1044 ) | ( n1021 & n1044 ) ;
  assign n1046 = ( n1041 & n1043 ) | ( n1041 & ~n1045 ) | ( n1043 & ~n1045 ) ;
  assign n1047 = ( ~n394 & n478 ) | ( ~n394 & n705 ) | ( n478 & n705 ) ;
  assign n1048 = ( n478 & ~n485 ) | ( n478 & n705 ) | ( ~n485 & n705 ) ;
  assign n1049 = ~n491 & n756 ;
  assign n1050 = n493 & ~n756 ;
  assign n1051 = ( n756 & ~n1049 ) | ( n756 & n1050 ) | ( ~n1049 & n1050 ) ;
  assign n1052 = ( n1047 & ~n1048 ) | ( n1047 & n1051 ) | ( ~n1048 & n1051 ) ;
  assign n1053 = ( ~n562 & n691 ) | ( ~n562 & n752 ) | ( n691 & n752 ) ;
  assign n1054 = ( ~n500 & n562 ) | ( ~n500 & n752 ) | ( n562 & n752 ) ;
  assign n1055 = n500 & n750 ;
  assign n1056 = ( ~n758 & n1054 ) | ( ~n758 & n1055 ) | ( n1054 & n1055 ) ;
  assign n1057 = ( n1008 & n1053 ) | ( n1008 & ~n1056 ) | ( n1053 & ~n1056 ) ;
  assign n1058 = ( n631 & ~n687 ) | ( n631 & n922 ) | ( ~n687 & n922 ) ;
  assign n1059 = ( n631 & n687 ) | ( n631 & ~n922 ) | ( n687 & ~n922 ) ;
  assign n1060 = n1058 & n1059 ;
  assign n1061 = ( n199 & n696 ) | ( n199 & ~n1060 ) | ( n696 & ~n1060 ) ;
  assign n1062 = ( n199 & ~n698 ) | ( n199 & n1060 ) | ( ~n698 & n1060 ) ;
  assign n1063 = n1061 & ~n1062 ;
  assign n1064 = ( n1052 & n1057 ) | ( n1052 & n1063 ) | ( n1057 & n1063 ) ;
  assign n1065 = ( ~n1002 & n1006 ) | ( ~n1002 & n1011 ) | ( n1006 & n1011 ) ;
  assign n1066 = ( ~n1011 & n1012 ) | ( ~n1011 & n1065 ) | ( n1012 & n1065 ) ;
  assign n1067 = ( ~n814 & n1034 ) | ( ~n814 & n1040 ) | ( n1034 & n1040 ) ;
  assign n1068 = ( n814 & ~n1041 ) | ( n814 & n1067 ) | ( ~n1041 & n1067 ) ;
  assign n1069 = ( n1064 & ~n1066 ) | ( n1064 & n1068 ) | ( ~n1066 & n1068 ) ;
  assign n1070 = ( ~n394 & n478 ) | ( ~n394 & n756 ) | ( n478 & n756 ) ;
  assign n1071 = ( n478 & ~n485 ) | ( n478 & n756 ) | ( ~n485 & n756 ) ;
  assign n1072 = ~n491 & n691 ;
  assign n1073 = n493 & ~n691 ;
  assign n1074 = ( n691 & ~n1072 ) | ( n691 & n1073 ) | ( ~n1072 & n1073 ) ;
  assign n1075 = ( n1070 & ~n1071 ) | ( n1070 & n1074 ) | ( ~n1071 & n1074 ) ;
  assign n1076 = ~n705 & n858 ;
  assign n1077 = ( n304 & n858 ) | ( n304 & ~n1031 ) | ( n858 & ~n1031 ) ;
  assign n1078 = ( ~n304 & n858 ) | ( ~n304 & n1031 ) | ( n858 & n1031 ) ;
  assign n1079 = ( ~n1076 & n1077 ) | ( ~n1076 & n1078 ) | ( n1077 & n1078 ) ;
  assign n1080 = n500 & ~n562 ;
  assign n1081 = ( ~n562 & n752 ) | ( ~n562 & n922 ) | ( n752 & n922 ) ;
  assign n1082 = n751 & ~n922 ;
  assign n1083 = ( n759 & n1081 ) | ( n759 & n1082 ) | ( n1081 & n1082 ) ;
  assign n1084 = ( n1054 & n1080 ) | ( n1054 & ~n1083 ) | ( n1080 & ~n1083 ) ;
  assign n1085 = ( n1075 & ~n1079 ) | ( n1075 & n1084 ) | ( ~n1079 & n1084 ) ;
  assign n1086 = n1028 & n1033 ;
  assign n1087 = ( n1033 & n1034 ) | ( n1033 & ~n1086 ) | ( n1034 & ~n1086 ) ;
  assign n1088 = ( n1052 & ~n1057 ) | ( n1052 & n1063 ) | ( ~n1057 & n1063 ) ;
  assign n1089 = ( n1057 & ~n1064 ) | ( n1057 & n1088 ) | ( ~n1064 & n1088 ) ;
  assign n1090 = ( n1085 & ~n1087 ) | ( n1085 & n1089 ) | ( ~n1087 & n1089 ) ;
  assign n1091 = n199 & ~n752 ;
  assign n1092 = n758 & ~n1091 ;
  assign n1093 = ( ~n304 & n705 ) | ( ~n304 & n858 ) | ( n705 & n858 ) ;
  assign n1094 = n705 & ~n1093 ;
  assign n1095 = n756 | n858 ;
  assign n1096 = ( n756 & n1093 ) | ( n756 & ~n1095 ) | ( n1093 & ~n1095 ) ;
  assign n1097 = ( n304 & ~n1094 ) | ( n304 & n1096 ) | ( ~n1094 & n1096 ) ;
  assign n1098 = n1092 & ~n1097 ;
  assign n1099 = ( ~n394 & n478 ) | ( ~n394 & n691 ) | ( n478 & n691 ) ;
  assign n1100 = ( n478 & ~n485 ) | ( n478 & n691 ) | ( ~n485 & n691 ) ;
  assign n1101 = ~n491 & n500 ;
  assign n1102 = n493 & ~n500 ;
  assign n1103 = ( n500 & ~n1101 ) | ( n500 & n1102 ) | ( ~n1101 & n1102 ) ;
  assign n1104 = ( n1099 & ~n1100 ) | ( n1099 & n1103 ) | ( ~n1100 & n1103 ) ;
  assign n1105 = n199 & ~n759 ;
  assign n1106 = ( ~n562 & n751 ) | ( ~n562 & n752 ) | ( n751 & n752 ) ;
  assign n1107 = ~n199 & n1106 ;
  assign n1108 = ( n199 & ~n1105 ) | ( n199 & n1107 ) | ( ~n1105 & n1107 ) ;
  assign n1109 = n562 & ~n922 ;
  assign n1110 = ( n1081 & ~n1108 ) | ( n1081 & n1109 ) | ( ~n1108 & n1109 ) ;
  assign n1111 = n1092 & n1097 ;
  assign n1112 = ( n1097 & n1098 ) | ( n1097 & ~n1111 ) | ( n1098 & ~n1111 ) ;
  assign n1113 = ( n1104 & n1110 ) | ( n1104 & ~n1112 ) | ( n1110 & ~n1112 ) ;
  assign n1114 = ( n1027 & n1098 ) | ( n1027 & n1113 ) | ( n1098 & n1113 ) ;
  assign n1115 = ( ~n394 & n478 ) | ( ~n394 & n500 ) | ( n478 & n500 ) ;
  assign n1116 = ( n478 & ~n485 ) | ( n478 & n500 ) | ( ~n485 & n500 ) ;
  assign n1117 = ~n491 & n922 ;
  assign n1118 = n493 & ~n922 ;
  assign n1119 = ( n922 & ~n1117 ) | ( n922 & n1118 ) | ( ~n1117 & n1118 ) ;
  assign n1120 = ( n1115 & ~n1116 ) | ( n1115 & n1119 ) | ( ~n1116 & n1119 ) ;
  assign n1121 = ( ~n304 & n691 ) | ( ~n304 & n858 ) | ( n691 & n858 ) ;
  assign n1122 = n691 & ~n1121 ;
  assign n1123 = n500 | n858 ;
  assign n1124 = ( n500 & n1121 ) | ( n500 & ~n1123 ) | ( n1121 & ~n1123 ) ;
  assign n1125 = ( n304 & ~n1122 ) | ( n304 & n1124 ) | ( ~n1122 & n1124 ) ;
  assign n1126 = ( ~n199 & n304 ) | ( ~n199 & n393 ) | ( n304 & n393 ) ;
  assign n1127 = ~n477 & n1126 ;
  assign n1128 = ~n1125 & n1127 ;
  assign n1129 = ~n691 & n858 ;
  assign n1130 = ( n304 & n858 ) | ( n304 & ~n1095 ) | ( n858 & ~n1095 ) ;
  assign n1131 = ( ~n304 & n858 ) | ( ~n304 & n1095 ) | ( n858 & n1095 ) ;
  assign n1132 = ( ~n1129 & n1130 ) | ( ~n1129 & n1131 ) | ( n1130 & n1131 ) ;
  assign n1133 = ( n1120 & n1128 ) | ( n1120 & ~n1132 ) | ( n1128 & ~n1132 ) ;
  assign n1134 = n199 | n922 ;
  assign n1135 = ( n199 & ~n858 ) | ( n199 & n1134 ) | ( ~n858 & n1134 ) ;
  assign n1136 = n304 | n1135 ;
  assign n1137 = n394 & ~n1126 ;
  assign n1138 = n858 & ~n922 ;
  assign n1139 = ( n304 & n858 ) | ( n304 & ~n1123 ) | ( n858 & ~n1123 ) ;
  assign n1140 = ( ~n304 & n858 ) | ( ~n304 & n1123 ) | ( n858 & n1123 ) ;
  assign n1141 = ( ~n1138 & n1139 ) | ( ~n1138 & n1140 ) | ( n1139 & n1140 ) ;
  assign n1142 = ( n1136 & ~n1137 ) | ( n1136 & n1141 ) | ( ~n1137 & n1141 ) ;
  assign n1143 = ( ~n394 & n478 ) | ( ~n394 & n922 ) | ( n478 & n922 ) ;
  assign n1144 = ( n478 & ~n485 ) | ( n478 & n922 ) | ( ~n485 & n922 ) ;
  assign n1145 = n199 & ~n491 ;
  assign n1146 = ~n199 & n493 ;
  assign n1147 = ( n199 & ~n1145 ) | ( n199 & n1146 ) | ( ~n1145 & n1146 ) ;
  assign n1148 = ( n1143 & ~n1144 ) | ( n1143 & n1147 ) | ( ~n1144 & n1147 ) ;
  assign n1149 = n1125 | n1127 ;
  assign n1150 = ( ~n1127 & n1128 ) | ( ~n1127 & n1149 ) | ( n1128 & n1149 ) ;
  assign n1151 = ( n1142 & ~n1148 ) | ( n1142 & n1150 ) | ( ~n1148 & n1150 ) ;
  assign n1152 = ( n1120 & ~n1128 ) | ( n1120 & n1132 ) | ( ~n1128 & n1132 ) ;
  assign n1153 = ( ~n1120 & n1133 ) | ( ~n1120 & n1152 ) | ( n1133 & n1152 ) ;
  assign n1154 = ( ~n1091 & n1151 ) | ( ~n1091 & n1153 ) | ( n1151 & n1153 ) ;
  assign n1155 = ( n1104 & ~n1110 ) | ( n1104 & n1112 ) | ( ~n1110 & n1112 ) ;
  assign n1156 = ( ~n1104 & n1113 ) | ( ~n1104 & n1155 ) | ( n1113 & n1155 ) ;
  assign n1157 = ( ~n1133 & n1154 ) | ( ~n1133 & n1156 ) | ( n1154 & n1156 ) ;
  assign n1158 = ( n1027 & ~n1098 ) | ( n1027 & n1113 ) | ( ~n1098 & n1113 ) ;
  assign n1159 = ( n1098 & ~n1114 ) | ( n1098 & n1158 ) | ( ~n1114 & n1158 ) ;
  assign n1160 = ( ~n1075 & n1079 ) | ( ~n1075 & n1084 ) | ( n1079 & n1084 ) ;
  assign n1161 = ( ~n1084 & n1085 ) | ( ~n1084 & n1160 ) | ( n1085 & n1160 ) ;
  assign n1162 = ( n1157 & ~n1159 ) | ( n1157 & n1161 ) | ( ~n1159 & n1161 ) ;
  assign n1163 = ( ~n1085 & n1087 ) | ( ~n1085 & n1089 ) | ( n1087 & n1089 ) ;
  assign n1164 = ( ~n1089 & n1090 ) | ( ~n1089 & n1163 ) | ( n1090 & n1163 ) ;
  assign n1165 = ( ~n1114 & n1162 ) | ( ~n1114 & n1164 ) | ( n1162 & n1164 ) ;
  assign n1166 = ( n1064 & n1066 ) | ( n1064 & n1068 ) | ( n1066 & n1068 ) ;
  assign n1167 = ( n1066 & n1069 ) | ( n1066 & ~n1166 ) | ( n1069 & ~n1166 ) ;
  assign n1168 = ( ~n1090 & n1165 ) | ( ~n1090 & n1167 ) | ( n1165 & n1167 ) ;
  assign n1169 = ( n1041 & n1043 ) | ( n1041 & n1045 ) | ( n1043 & n1045 ) ;
  assign n1170 = ( n1045 & n1046 ) | ( n1045 & ~n1169 ) | ( n1046 & ~n1169 ) ;
  assign n1171 = ( ~n1069 & n1168 ) | ( ~n1069 & n1170 ) | ( n1168 & n1170 ) ;
  assign n1172 = ( n1021 & n1023 ) | ( n1021 & n1025 ) | ( n1023 & n1025 ) ;
  assign n1173 = ( n1023 & n1026 ) | ( n1023 & ~n1172 ) | ( n1026 & ~n1172 ) ;
  assign n1174 = ( ~n1046 & n1171 ) | ( ~n1046 & n1173 ) | ( n1171 & n1173 ) ;
  assign n1175 = ( n884 & n953 ) | ( n884 & n995 ) | ( n953 & n995 ) ;
  assign n1176 = ( n953 & n996 ) | ( n953 & ~n1175 ) | ( n996 & ~n1175 ) ;
  assign n1177 = ( ~n1026 & n1174 ) | ( ~n1026 & n1176 ) | ( n1174 & n1176 ) ;
  assign n1178 = ( ~n562 & n752 ) | ( ~n562 & n863 ) | ( n752 & n863 ) ;
  assign n1179 = n562 & ~n863 ;
  assign n1180 = ~n483 & n751 ;
  assign n1181 = ( n759 & n985 ) | ( n759 & n1180 ) | ( n985 & n1180 ) ;
  assign n1182 = ( n1178 & n1179 ) | ( n1178 & ~n1181 ) | ( n1179 & ~n1181 ) ;
  assign n1183 = ( n489 & n631 ) | ( n489 & ~n687 ) | ( n631 & ~n687 ) ;
  assign n1184 = ( ~n489 & n631 ) | ( ~n489 & n687 ) | ( n631 & n687 ) ;
  assign n1185 = n1183 & n1184 ;
  assign n1186 = ( n696 & n705 ) | ( n696 & ~n1185 ) | ( n705 & ~n1185 ) ;
  assign n1187 = ( ~n698 & n705 ) | ( ~n698 & n1185 ) | ( n705 & n1185 ) ;
  assign n1188 = n1186 & ~n1187 ;
  assign n1189 = ( n192 & ~n756 ) | ( n192 & n813 ) | ( ~n756 & n813 ) ;
  assign n1190 = ( ~n192 & n756 ) | ( ~n192 & n813 ) | ( n756 & n813 ) ;
  assign n1191 = n1189 & n1190 ;
  assign n1192 = ( n691 & n967 ) | ( n691 & ~n1191 ) | ( n967 & ~n1191 ) ;
  assign n1193 = ( n691 & ~n969 ) | ( n691 & n1191 ) | ( ~n969 & n1191 ) ;
  assign n1194 = n1192 & ~n1193 ;
  assign n1195 = ( n1182 & n1188 ) | ( n1182 & n1194 ) | ( n1188 & n1194 ) ;
  assign n1196 = ( ~n1182 & n1188 ) | ( ~n1182 & n1194 ) | ( n1188 & n1194 ) ;
  assign n1197 = ( n1182 & ~n1195 ) | ( n1182 & n1196 ) | ( ~n1195 & n1196 ) ;
  assign n1198 = ( n304 & n943 ) | ( n304 & ~n944 ) | ( n943 & ~n944 ) ;
  assign n1199 = n199 & n918 ;
  assign n1200 = ( ~n394 & n478 ) | ( ~n394 & n939 ) | ( n478 & n939 ) ;
  assign n1201 = ( n478 & ~n485 ) | ( n478 & n939 ) | ( ~n485 & n939 ) ;
  assign n1202 = ~n491 & n819 ;
  assign n1203 = n493 & ~n819 ;
  assign n1204 = ( n819 & ~n1202 ) | ( n819 & n1203 ) | ( ~n1202 & n1203 ) ;
  assign n1205 = ( n1200 & ~n1201 ) | ( n1200 & n1204 ) | ( ~n1201 & n1204 ) ;
  assign n1206 = ( ~n1198 & n1199 ) | ( ~n1198 & n1205 ) | ( n1199 & n1205 ) ;
  assign n1207 = ( n1199 & n1205 ) | ( n1199 & ~n1206 ) | ( n1205 & ~n1206 ) ;
  assign n1208 = ( n1198 & n1206 ) | ( n1198 & ~n1207 ) | ( n1206 & ~n1207 ) ;
  assign n1209 = ( n951 & n1197 ) | ( n951 & ~n1208 ) | ( n1197 & ~n1208 ) ;
  assign n1210 = ( ~n951 & n1197 ) | ( ~n951 & n1208 ) | ( n1197 & n1208 ) ;
  assign n1211 = ( ~n1197 & n1209 ) | ( ~n1197 & n1210 ) | ( n1209 & n1210 ) ;
  assign n1212 = n194 & ~n500 ;
  assign n1213 = ( n922 & n927 ) | ( n922 & ~n1212 ) | ( n927 & ~n1212 ) ;
  assign n1214 = ( ~n193 & n922 ) | ( ~n193 & n1212 ) | ( n922 & n1212 ) ;
  assign n1215 = n1213 & ~n1214 ;
  assign n1216 = ( n948 & n990 ) | ( n948 & n1215 ) | ( n990 & n1215 ) ;
  assign n1217 = ( n948 & ~n990 ) | ( n948 & n1215 ) | ( ~n990 & n1215 ) ;
  assign n1218 = ( n990 & ~n1216 ) | ( n990 & n1217 ) | ( ~n1216 & n1217 ) ;
  assign n1219 = ( n993 & ~n1211 ) | ( n993 & n1218 ) | ( ~n1211 & n1218 ) ;
  assign n1220 = ( n993 & n1211 ) | ( n993 & n1218 ) | ( n1211 & n1218 ) ;
  assign n1221 = ( n1211 & n1219 ) | ( n1211 & ~n1220 ) | ( n1219 & ~n1220 ) ;
  assign n1222 = ( ~n996 & n1177 ) | ( ~n996 & n1221 ) | ( n1177 & n1221 ) ;
  assign n1223 = ( n1177 & n1221 ) | ( n1177 & ~n1222 ) | ( n1221 & ~n1222 ) ;
  assign n1224 = ( n996 & n1222 ) | ( n996 & ~n1223 ) | ( n1222 & ~n1223 ) ;
  assign n1225 = ( n50 & ~n56 ) | ( n50 & n119 ) | ( ~n56 & n119 ) ;
  assign n1226 = ( ~n119 & n137 ) | ( ~n119 & n1225 ) | ( n137 & n1225 ) ;
  assign n1227 = n787 | n1226 ;
  assign n1228 = n539 | n1227 ;
  assign n1229 = n172 | n282 ;
  assign n1230 = ( n92 & n112 ) | ( n92 & ~n352 ) | ( n112 & ~n352 ) ;
  assign n1231 = n353 | n1230 ;
  assign n1232 = ( n717 & ~n1229 ) | ( n717 & n1231 ) | ( ~n1229 & n1231 ) ;
  assign n1233 = n1229 | n1232 ;
  assign n1234 = n230 | n447 ;
  assign n1235 = ( ~n1228 & n1233 ) | ( ~n1228 & n1234 ) | ( n1233 & n1234 ) ;
  assign n1236 = n1228 | n1235 ;
  assign n1237 = n297 | n800 ;
  assign n1238 = n280 | n1237 ;
  assign n1239 = n80 & n83 ;
  assign n1240 = ( n106 & ~n128 ) | ( n106 & n1239 ) | ( ~n128 & n1239 ) ;
  assign n1241 = ( n189 & n325 ) | ( n189 & ~n1240 ) | ( n325 & ~n1240 ) ;
  assign n1242 = n1240 | n1241 ;
  assign n1243 = n186 | n308 ;
  assign n1244 = n250 | n1243 ;
  assign n1245 = ( n436 & ~n635 ) | ( n436 & n1244 ) | ( ~n635 & n1244 ) ;
  assign n1246 = n635 | n1245 ;
  assign n1247 = ( n905 & ~n1242 ) | ( n905 & n1246 ) | ( ~n1242 & n1246 ) ;
  assign n1248 = n1242 | n1247 ;
  assign n1249 = ( n517 & ~n1238 ) | ( n517 & n1248 ) | ( ~n1238 & n1248 ) ;
  assign n1250 = n1238 | n1249 ;
  assign n1251 = n283 | n522 ;
  assign n1252 = n211 | n444 ;
  assign n1253 = ( n132 & ~n468 ) | ( n132 & n649 ) | ( ~n468 & n649 ) ;
  assign n1254 = ( ~n1251 & n1252 ) | ( ~n1251 & n1253 ) | ( n1252 & n1253 ) ;
  assign n1255 = n1251 | n1254 ;
  assign n1256 = ( ~n1236 & n1250 ) | ( ~n1236 & n1255 ) | ( n1250 & n1255 ) ;
  assign n1257 = n1236 | n1256 ;
  assign n1258 = n1224 & ~n1257 ;
  assign n1259 = ~n1224 & n1257 ;
  assign n1260 = x2 & ~n25 ;
  assign n1261 = x2 & ~x22 ;
  assign n1262 = ( n197 & n1260 ) | ( n197 & ~n1261 ) | ( n1260 & ~n1261 ) ;
  assign n1263 = n199 | n1262 ;
  assign n1264 = ( n199 & n1262 ) | ( n199 & ~n1263 ) | ( n1262 & ~n1263 ) ;
  assign n1265 = n1263 & ~n1264 ;
  assign n1266 = ( n1258 & n1259 ) | ( n1258 & n1265 ) | ( n1259 & n1265 ) ;
  assign n1267 = ( n1224 & ~n1257 ) | ( n1224 & n1262 ) | ( ~n1257 & n1262 ) ;
  assign n1268 = ~n1258 & n1267 ;
  assign n1269 = n251 | n547 ;
  assign n1270 = n266 | n325 ;
  assign n1271 = ( n311 & n409 ) | ( n311 & ~n1239 ) | ( n409 & ~n1239 ) ;
  assign n1272 = n1239 | n1271 ;
  assign n1273 = ( ~n1269 & n1270 ) | ( ~n1269 & n1272 ) | ( n1270 & n1272 ) ;
  assign n1274 = n1269 | n1273 ;
  assign n1275 = ( n107 & n115 ) | ( n107 & n127 ) | ( n115 & n127 ) ;
  assign n1276 = ( ~n92 & n538 ) | ( ~n92 & n1275 ) | ( n538 & n1275 ) ;
  assign n1277 = ( n92 & n410 ) | ( n92 & ~n1276 ) | ( n410 & ~n1276 ) ;
  assign n1278 = n1276 | n1277 ;
  assign n1279 = n87 & ~n162 ;
  assign n1280 = ( ~n56 & n106 ) | ( ~n56 & n151 ) | ( n106 & n151 ) ;
  assign n1281 = n122 | n229 ;
  assign n1282 = ( n204 & n207 ) | ( n204 & ~n352 ) | ( n207 & ~n352 ) ;
  assign n1283 = ( n378 & ~n1281 ) | ( n378 & n1282 ) | ( ~n1281 & n1282 ) ;
  assign n1284 = n1281 | n1283 ;
  assign n1285 = ( n617 & ~n1280 ) | ( n617 & n1284 ) | ( ~n1280 & n1284 ) ;
  assign n1286 = ( ~n1279 & n1280 ) | ( ~n1279 & n1285 ) | ( n1280 & n1285 ) ;
  assign n1287 = ( ~n1278 & n1279 ) | ( ~n1278 & n1286 ) | ( n1279 & n1286 ) ;
  assign n1288 = n1278 | n1287 ;
  assign n1289 = ( n408 & ~n502 ) | ( n408 & n765 ) | ( ~n502 & n765 ) ;
  assign n1290 = ( ~n1274 & n1288 ) | ( ~n1274 & n1289 ) | ( n1288 & n1289 ) ;
  assign n1291 = n255 | n656 ;
  assign n1292 = n709 | n1291 ;
  assign n1293 = n166 | n585 ;
  assign n1294 = ( n73 & n141 ) | ( n73 & ~n174 ) | ( n141 & ~n174 ) ;
  assign n1295 = ( n56 & n109 ) | ( n56 & n214 ) | ( n109 & n214 ) ;
  assign n1296 = ( n380 & n509 ) | ( n380 & ~n1295 ) | ( n509 & ~n1295 ) ;
  assign n1297 = n1295 | n1296 ;
  assign n1298 = ( ~n1293 & n1294 ) | ( ~n1293 & n1297 ) | ( n1294 & n1297 ) ;
  assign n1299 = n1293 | n1298 ;
  assign n1300 = ( ~n1289 & n1292 ) | ( ~n1289 & n1299 ) | ( n1292 & n1299 ) ;
  assign n1301 = ( ~n1274 & n1290 ) | ( ~n1274 & n1300 ) | ( n1290 & n1300 ) ;
  assign n1302 = n1274 | n1301 ;
  assign n1303 = n562 & ~n819 ;
  assign n1304 = ( ~n562 & n752 ) | ( ~n562 & n819 ) | ( n752 & n819 ) ;
  assign n1305 = n751 & ~n863 ;
  assign n1306 = ( n759 & n1178 ) | ( n759 & n1305 ) | ( n1178 & n1305 ) ;
  assign n1307 = ( n1303 & n1304 ) | ( n1303 & ~n1306 ) | ( n1304 & ~n1306 ) ;
  assign n1308 = ( n483 & n631 ) | ( n483 & ~n687 ) | ( n631 & ~n687 ) ;
  assign n1309 = ( ~n483 & n631 ) | ( ~n483 & n687 ) | ( n631 & n687 ) ;
  assign n1310 = n1308 & n1309 ;
  assign n1311 = ( n489 & n696 ) | ( n489 & ~n1310 ) | ( n696 & ~n1310 ) ;
  assign n1312 = ( n489 & ~n698 ) | ( n489 & n1310 ) | ( ~n698 & n1310 ) ;
  assign n1313 = n1311 & ~n1312 ;
  assign n1314 = ( n192 & ~n705 ) | ( n192 & n813 ) | ( ~n705 & n813 ) ;
  assign n1315 = ( ~n192 & n705 ) | ( ~n192 & n813 ) | ( n705 & n813 ) ;
  assign n1316 = n1314 & n1315 ;
  assign n1317 = ( n756 & n967 ) | ( n756 & ~n1316 ) | ( n967 & ~n1316 ) ;
  assign n1318 = ( n756 & ~n969 ) | ( n756 & n1316 ) | ( ~n969 & n1316 ) ;
  assign n1319 = n1317 & ~n1318 ;
  assign n1320 = ( n1307 & n1313 ) | ( n1307 & n1319 ) | ( n1313 & n1319 ) ;
  assign n1321 = ( ~n1307 & n1313 ) | ( ~n1307 & n1319 ) | ( n1313 & n1319 ) ;
  assign n1322 = ( n1307 & ~n1320 ) | ( n1307 & n1321 ) | ( ~n1320 & n1321 ) ;
  assign n1323 = ( n478 & ~n485 ) | ( n478 & n943 ) | ( ~n485 & n943 ) ;
  assign n1324 = ( ~n394 & n478 ) | ( ~n394 & n943 ) | ( n478 & n943 ) ;
  assign n1325 = ~n491 & n939 ;
  assign n1326 = ~n493 & n939 ;
  assign n1327 = ( n493 & ~n1325 ) | ( n493 & n1326 ) | ( ~n1325 & n1326 ) ;
  assign n1328 = ( ~n1323 & n1324 ) | ( ~n1323 & n1327 ) | ( n1324 & n1327 ) ;
  assign n1329 = ( ~n304 & n923 ) | ( ~n304 & n1328 ) | ( n923 & n1328 ) ;
  assign n1330 = ( n304 & n923 ) | ( n304 & ~n1328 ) | ( n923 & ~n1328 ) ;
  assign n1331 = ( ~n923 & n1329 ) | ( ~n923 & n1330 ) | ( n1329 & n1330 ) ;
  assign n1332 = ( n1216 & n1322 ) | ( n1216 & ~n1331 ) | ( n1322 & ~n1331 ) ;
  assign n1333 = ( ~n1216 & n1322 ) | ( ~n1216 & n1331 ) | ( n1322 & n1331 ) ;
  assign n1334 = ( ~n1322 & n1332 ) | ( ~n1322 & n1333 ) | ( n1332 & n1333 ) ;
  assign n1335 = n194 & ~n691 ;
  assign n1336 = ( n500 & n927 ) | ( n500 & ~n1335 ) | ( n927 & ~n1335 ) ;
  assign n1337 = ( ~n193 & n500 ) | ( ~n193 & n1335 ) | ( n500 & n1335 ) ;
  assign n1338 = n1336 & ~n1337 ;
  assign n1339 = ( n1195 & n1206 ) | ( n1195 & n1338 ) | ( n1206 & n1338 ) ;
  assign n1340 = ( ~n1195 & n1206 ) | ( ~n1195 & n1338 ) | ( n1206 & n1338 ) ;
  assign n1341 = ( n1195 & ~n1339 ) | ( n1195 & n1340 ) | ( ~n1339 & n1340 ) ;
  assign n1342 = ( n1209 & ~n1334 ) | ( n1209 & n1341 ) | ( ~n1334 & n1341 ) ;
  assign n1343 = ( n1209 & n1334 ) | ( n1209 & n1341 ) | ( n1334 & n1341 ) ;
  assign n1344 = ( n1334 & n1342 ) | ( n1334 & ~n1343 ) | ( n1342 & ~n1343 ) ;
  assign n1345 = ( ~n1219 & n1222 ) | ( ~n1219 & n1344 ) | ( n1222 & n1344 ) ;
  assign n1346 = ( n1222 & n1344 ) | ( n1222 & ~n1345 ) | ( n1344 & ~n1345 ) ;
  assign n1347 = ( n1219 & n1345 ) | ( n1219 & ~n1346 ) | ( n1345 & ~n1346 ) ;
  assign n1348 = ( n1258 & ~n1302 ) | ( n1258 & n1347 ) | ( ~n1302 & n1347 ) ;
  assign n1349 = ( n631 & ~n687 ) | ( n631 & n863 ) | ( ~n687 & n863 ) ;
  assign n1350 = ( n631 & n687 ) | ( n631 & ~n863 ) | ( n687 & ~n863 ) ;
  assign n1351 = n1349 & n1350 ;
  assign n1352 = ( n483 & n696 ) | ( n483 & ~n1351 ) | ( n696 & ~n1351 ) ;
  assign n1353 = ( n483 & ~n698 ) | ( n483 & n1351 ) | ( ~n698 & n1351 ) ;
  assign n1354 = n1352 & ~n1353 ;
  assign n1355 = ( ~n562 & n752 ) | ( ~n562 & n939 ) | ( n752 & n939 ) ;
  assign n1356 = n562 & ~n939 ;
  assign n1357 = n751 & ~n819 ;
  assign n1358 = ( n759 & ~n1303 ) | ( n759 & n1357 ) | ( ~n1303 & n1357 ) ;
  assign n1359 = ( n1355 & n1356 ) | ( n1355 & ~n1358 ) | ( n1356 & ~n1358 ) ;
  assign n1360 = ( ~n192 & n489 ) | ( ~n192 & n813 ) | ( n489 & n813 ) ;
  assign n1361 = ( n192 & ~n489 ) | ( n192 & n813 ) | ( ~n489 & n813 ) ;
  assign n1362 = n1360 & n1361 ;
  assign n1363 = ( n705 & n967 ) | ( n705 & ~n1362 ) | ( n967 & ~n1362 ) ;
  assign n1364 = ( n705 & ~n969 ) | ( n705 & n1362 ) | ( ~n969 & n1362 ) ;
  assign n1365 = n1363 & ~n1364 ;
  assign n1366 = ( n1354 & n1359 ) | ( n1354 & n1365 ) | ( n1359 & n1365 ) ;
  assign n1367 = ( ~n1354 & n1359 ) | ( ~n1354 & n1365 ) | ( n1359 & n1365 ) ;
  assign n1368 = ( n1354 & ~n1366 ) | ( n1354 & n1367 ) | ( ~n1366 & n1367 ) ;
  assign n1369 = n478 & n943 ;
  assign n1370 = n477 & n943 ;
  assign n1371 = ( n490 & ~n1369 ) | ( n490 & n1370 ) | ( ~n1369 & n1370 ) ;
  assign n1372 = n500 & n918 ;
  assign n1373 = ( ~n304 & n1371 ) | ( ~n304 & n1372 ) | ( n1371 & n1372 ) ;
  assign n1374 = ( n304 & n1371 ) | ( n304 & ~n1372 ) | ( n1371 & ~n1372 ) ;
  assign n1375 = ( ~n1371 & n1373 ) | ( ~n1371 & n1374 ) | ( n1373 & n1374 ) ;
  assign n1376 = ( n1339 & n1368 ) | ( n1339 & ~n1375 ) | ( n1368 & ~n1375 ) ;
  assign n1377 = ( ~n1339 & n1368 ) | ( ~n1339 & n1375 ) | ( n1368 & n1375 ) ;
  assign n1378 = ( ~n1368 & n1376 ) | ( ~n1368 & n1377 ) | ( n1376 & n1377 ) ;
  assign n1379 = n756 & n918 ;
  assign n1380 = ( n194 & ~n756 ) | ( n194 & n918 ) | ( ~n756 & n918 ) ;
  assign n1381 = ( ~n918 & n1379 ) | ( ~n918 & n1380 ) | ( n1379 & n1380 ) ;
  assign n1382 = ( ~n193 & n691 ) | ( ~n193 & n1381 ) | ( n691 & n1381 ) ;
  assign n1383 = ( n691 & n927 ) | ( n691 & ~n1381 ) | ( n927 & ~n1381 ) ;
  assign n1384 = ~n1382 & n1383 ;
  assign n1385 = ( n1320 & n1329 ) | ( n1320 & n1384 ) | ( n1329 & n1384 ) ;
  assign n1386 = ( ~n1320 & n1329 ) | ( ~n1320 & n1384 ) | ( n1329 & n1384 ) ;
  assign n1387 = ( n1320 & ~n1385 ) | ( n1320 & n1386 ) | ( ~n1385 & n1386 ) ;
  assign n1388 = ( n1332 & ~n1378 ) | ( n1332 & n1387 ) | ( ~n1378 & n1387 ) ;
  assign n1389 = ( n1332 & n1378 ) | ( n1332 & n1387 ) | ( n1378 & n1387 ) ;
  assign n1390 = ( n1378 & n1388 ) | ( n1378 & ~n1389 ) | ( n1388 & ~n1389 ) ;
  assign n1391 = ( ~n1342 & n1345 ) | ( ~n1342 & n1390 ) | ( n1345 & n1390 ) ;
  assign n1392 = ( n1345 & n1390 ) | ( n1345 & ~n1391 ) | ( n1390 & ~n1391 ) ;
  assign n1393 = ( n1342 & n1391 ) | ( n1342 & ~n1392 ) | ( n1391 & ~n1392 ) ;
  assign n1394 = ( n83 & n104 ) | ( n83 & n136 ) | ( n104 & n136 ) ;
  assign n1395 = ( n98 & n126 ) | ( n98 & ~n174 ) | ( n126 & ~n174 ) ;
  assign n1396 = ( n331 & ~n1394 ) | ( n331 & n1395 ) | ( ~n1394 & n1395 ) ;
  assign n1397 = n1394 | n1396 ;
  assign n1398 = ( n107 & n163 ) | ( n107 & ~n418 ) | ( n163 & ~n418 ) ;
  assign n1399 = n94 | n1398 ;
  assign n1400 = n1291 | n1399 ;
  assign n1401 = n151 | n278 ;
  assign n1402 = n189 | n726 ;
  assign n1403 = ( ~n1400 & n1401 ) | ( ~n1400 & n1402 ) | ( n1401 & n1402 ) ;
  assign n1404 = n1400 | n1403 ;
  assign n1405 = ( n223 & ~n468 ) | ( n223 & n533 ) | ( ~n468 & n533 ) ;
  assign n1406 = n468 | n1405 ;
  assign n1407 = ( n399 & n1237 ) | ( n399 & ~n1406 ) | ( n1237 & ~n1406 ) ;
  assign n1408 = n1406 | n1407 ;
  assign n1409 = ( ~n1397 & n1404 ) | ( ~n1397 & n1408 ) | ( n1404 & n1408 ) ;
  assign n1410 = n1397 | n1409 ;
  assign n1411 = n288 | n462 ;
  assign n1412 = ( ~n226 & n252 ) | ( ~n226 & n901 ) | ( n252 & n901 ) ;
  assign n1413 = n226 | n1412 ;
  assign n1414 = ( n167 & n213 ) | ( n167 & ~n1413 ) | ( n213 & ~n1413 ) ;
  assign n1415 = n1413 | n1414 ;
  assign n1416 = ( n679 & ~n1411 ) | ( n679 & n1415 ) | ( ~n1411 & n1415 ) ;
  assign n1417 = n88 | n305 ;
  assign n1418 = ( n204 & n228 ) | ( n204 & ~n356 ) | ( n228 & ~n356 ) ;
  assign n1419 = n588 | n786 ;
  assign n1420 = ( ~n202 & n609 ) | ( ~n202 & n661 ) | ( n609 & n661 ) ;
  assign n1421 = ( ~n1418 & n1419 ) | ( ~n1418 & n1420 ) | ( n1419 & n1420 ) ;
  assign n1422 = n1418 | n1421 ;
  assign n1423 = n222 & ~n895 ;
  assign n1424 = ( n1417 & n1422 ) | ( n1417 & n1423 ) | ( n1422 & n1423 ) ;
  assign n1425 = ( ~n1411 & n1423 ) | ( ~n1411 & n1424 ) | ( n1423 & n1424 ) ;
  assign n1426 = ~n1424 & n1425 ;
  assign n1427 = ( n1410 & ~n1416 ) | ( n1410 & n1426 ) | ( ~n1416 & n1426 ) ;
  assign n1428 = ~n1410 & n1427 ;
  assign n1429 = ( n1348 & n1393 ) | ( n1348 & n1428 ) | ( n1393 & n1428 ) ;
  assign n1430 = ( ~n1348 & n1393 ) | ( ~n1348 & n1428 ) | ( n1393 & n1428 ) ;
  assign n1431 = ( n1348 & ~n1429 ) | ( n1348 & n1430 ) | ( ~n1429 & n1430 ) ;
  assign n1432 = ( n1258 & n1302 ) | ( n1258 & n1347 ) | ( n1302 & n1347 ) ;
  assign n1433 = ( ~n1259 & n1302 ) | ( ~n1259 & n1347 ) | ( n1302 & n1347 ) ;
  assign n1434 = ~n1432 & n1433 ;
  assign n1435 = x0 & ~x22 ;
  assign n1436 = ( ~x1 & n1262 ) | ( ~x1 & n1435 ) | ( n1262 & n1435 ) ;
  assign n1437 = ( n1262 & n1435 ) | ( n1262 & ~n1436 ) | ( n1435 & ~n1436 ) ;
  assign n1438 = ( x1 & n1436 ) | ( x1 & ~n1437 ) | ( n1436 & ~n1437 ) ;
  assign n1439 = x0 & n1438 ;
  assign n1440 = ( n1302 & n1348 ) | ( n1302 & ~n1432 ) | ( n1348 & ~n1432 ) ;
  assign n1441 = ( n1258 & n1259 ) | ( n1258 & ~n1440 ) | ( n1259 & ~n1440 ) ;
  assign n1442 = n1439 & ~n1441 ;
  assign n1443 = ( n1431 & n1434 ) | ( n1431 & ~n1442 ) | ( n1434 & ~n1442 ) ;
  assign n1444 = n1431 & ~n1443 ;
  assign n1445 = ( x0 & ~n1431 ) | ( x0 & n1439 ) | ( ~n1431 & n1439 ) ;
  assign n1446 = ( n25 & n1440 ) | ( n25 & n1445 ) | ( n1440 & n1445 ) ;
  assign n1447 = ( n1268 & n1444 ) | ( n1268 & ~n1446 ) | ( n1444 & ~n1446 ) ;
  assign n1448 = n1260 & n1440 ;
  assign n1449 = x0 & ~n1438 ;
  assign n1450 = ~x0 & x1 ;
  assign n1451 = ~n1431 & n1450 ;
  assign n1452 = ( n631 & n687 ) | ( n631 & ~n819 ) | ( n687 & ~n819 ) ;
  assign n1453 = ( n631 & ~n687 ) | ( n631 & n819 ) | ( ~n687 & n819 ) ;
  assign n1454 = n1452 & n1453 ;
  assign n1455 = ( n696 & n863 ) | ( n696 & ~n1454 ) | ( n863 & ~n1454 ) ;
  assign n1456 = ( ~n698 & n863 ) | ( ~n698 & n1454 ) | ( n863 & n1454 ) ;
  assign n1457 = n1455 & ~n1456 ;
  assign n1458 = n691 & n918 ;
  assign n1459 = ( n304 & ~n490 ) | ( n304 & n1458 ) | ( ~n490 & n1458 ) ;
  assign n1460 = ( n304 & n1458 ) | ( n304 & ~n1459 ) | ( n1458 & ~n1459 ) ;
  assign n1461 = ( n490 & n1459 ) | ( n490 & ~n1460 ) | ( n1459 & ~n1460 ) ;
  assign n1462 = ( n1373 & n1457 ) | ( n1373 & ~n1461 ) | ( n1457 & ~n1461 ) ;
  assign n1463 = ( ~n1373 & n1457 ) | ( ~n1373 & n1461 ) | ( n1457 & n1461 ) ;
  assign n1464 = ( ~n1457 & n1462 ) | ( ~n1457 & n1463 ) | ( n1462 & n1463 ) ;
  assign n1465 = ~n562 & n943 ;
  assign n1466 = ( n562 & n752 ) | ( n562 & ~n943 ) | ( n752 & ~n943 ) ;
  assign n1467 = n751 & ~n939 ;
  assign n1468 = ( n759 & n1355 ) | ( n759 & n1467 ) | ( n1355 & n1467 ) ;
  assign n1469 = ( n1465 & n1466 ) | ( n1465 & ~n1468 ) | ( n1466 & ~n1468 ) ;
  assign n1470 = n705 & n918 ;
  assign n1471 = ( n194 & ~n705 ) | ( n194 & n918 ) | ( ~n705 & n918 ) ;
  assign n1472 = ( ~n918 & n1470 ) | ( ~n918 & n1471 ) | ( n1470 & n1471 ) ;
  assign n1473 = ( ~n193 & n756 ) | ( ~n193 & n1472 ) | ( n756 & n1472 ) ;
  assign n1474 = ( n756 & n927 ) | ( n756 & ~n1472 ) | ( n927 & ~n1472 ) ;
  assign n1475 = ~n1473 & n1474 ;
  assign n1476 = ( n192 & ~n483 ) | ( n192 & n813 ) | ( ~n483 & n813 ) ;
  assign n1477 = ( ~n192 & n483 ) | ( ~n192 & n813 ) | ( n483 & n813 ) ;
  assign n1478 = n1476 & n1477 ;
  assign n1479 = ( n489 & n967 ) | ( n489 & ~n1478 ) | ( n967 & ~n1478 ) ;
  assign n1480 = ( n489 & ~n969 ) | ( n489 & n1478 ) | ( ~n969 & n1478 ) ;
  assign n1481 = n1479 & ~n1480 ;
  assign n1482 = ( n1469 & n1475 ) | ( n1469 & n1481 ) | ( n1475 & n1481 ) ;
  assign n1483 = ( ~n1469 & n1475 ) | ( ~n1469 & n1481 ) | ( n1475 & n1481 ) ;
  assign n1484 = ( n1469 & ~n1482 ) | ( n1469 & n1483 ) | ( ~n1482 & n1483 ) ;
  assign n1485 = ( n1366 & n1385 ) | ( n1366 & n1484 ) | ( n1385 & n1484 ) ;
  assign n1486 = ( n1366 & ~n1385 ) | ( n1366 & n1484 ) | ( ~n1385 & n1484 ) ;
  assign n1487 = ( n1385 & ~n1485 ) | ( n1385 & n1486 ) | ( ~n1485 & n1486 ) ;
  assign n1488 = ( n1376 & ~n1464 ) | ( n1376 & n1487 ) | ( ~n1464 & n1487 ) ;
  assign n1489 = ( n1376 & n1464 ) | ( n1376 & n1487 ) | ( n1464 & n1487 ) ;
  assign n1490 = ( n1464 & n1488 ) | ( n1464 & ~n1489 ) | ( n1488 & ~n1489 ) ;
  assign n1491 = ( ~n1388 & n1391 ) | ( ~n1388 & n1490 ) | ( n1391 & n1490 ) ;
  assign n1492 = ( n1391 & n1490 ) | ( n1391 & ~n1491 ) | ( n1490 & ~n1491 ) ;
  assign n1493 = ( n1388 & n1491 ) | ( n1388 & ~n1492 ) | ( n1491 & ~n1492 ) ;
  assign n1494 = ( n237 & ~n238 ) | ( n237 & n329 ) | ( ~n238 & n329 ) ;
  assign n1495 = n269 | n654 ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = ( n56 & n224 ) | ( n56 & n255 ) | ( n224 & n255 ) ;
  assign n1498 = ( ~n356 & n427 ) | ( ~n356 & n1497 ) | ( n427 & n1497 ) ;
  assign n1499 = n356 | n1498 ;
  assign n1500 = n229 | n422 ;
  assign n1501 = n395 | n1500 ;
  assign n1502 = ( n717 & ~n1499 ) | ( n717 & n1501 ) | ( ~n1499 & n1501 ) ;
  assign n1503 = n1499 | n1502 ;
  assign n1504 = ( ~n519 & n1496 ) | ( ~n519 & n1503 ) | ( n1496 & n1503 ) ;
  assign n1505 = ( n519 & ~n1415 ) | ( n519 & n1504 ) | ( ~n1415 & n1504 ) ;
  assign n1506 = ( n1248 & n1415 ) | ( n1248 & ~n1505 ) | ( n1415 & ~n1505 ) ;
  assign n1507 = n1505 | n1506 ;
  assign n1508 = ( n1429 & n1493 ) | ( n1429 & ~n1507 ) | ( n1493 & ~n1507 ) ;
  assign n1509 = ( ~n1429 & n1493 ) | ( ~n1429 & n1507 ) | ( n1493 & n1507 ) ;
  assign n1510 = ( ~n1493 & n1508 ) | ( ~n1493 & n1509 ) | ( n1508 & n1509 ) ;
  assign n1511 = n1449 & n1510 ;
  assign n1512 = n1451 | n1511 ;
  assign n1513 = n1431 & n1434 ;
  assign n1514 = n1440 & ~n1513 ;
  assign n1515 = ( ~n1431 & n1510 ) | ( ~n1431 & n1514 ) | ( n1510 & n1514 ) ;
  assign n1516 = ( n1431 & n1510 ) | ( n1431 & n1514 ) | ( n1510 & n1514 ) ;
  assign n1517 = ( n1431 & n1515 ) | ( n1431 & ~n1516 ) | ( n1515 & ~n1516 ) ;
  assign n1518 = ( x0 & n1449 ) | ( x0 & ~n1517 ) | ( n1449 & ~n1517 ) ;
  assign n1519 = ( ~n1449 & n1512 ) | ( ~n1449 & n1518 ) | ( n1512 & n1518 ) ;
  assign n1520 = ~n1262 & n1519 ;
  assign n1521 = n1262 & ~n1519 ;
  assign n1522 = ( ~n1448 & n1520 ) | ( ~n1448 & n1521 ) | ( n1520 & n1521 ) ;
  assign n1523 = ( n1266 & n1447 ) | ( n1266 & n1522 ) | ( n1447 & n1522 ) ;
  assign n1524 = ( ~n497 & n499 ) | ( ~n497 & n922 ) | ( n499 & n922 ) ;
  assign n1525 = n500 & ~n922 ;
  assign n1526 = n1524 | n1525 ;
  assign n1527 = n1265 & n1526 ;
  assign n1528 = ( n1434 & n1441 ) | ( n1434 & n1527 ) | ( n1441 & n1527 ) ;
  assign n1529 = n500 & n1266 ;
  assign n1530 = ( ~n919 & n921 ) | ( ~n919 & n1262 ) | ( n921 & n1262 ) ;
  assign n1531 = ( n1134 & ~n1263 ) | ( n1134 & n1530 ) | ( ~n1263 & n1530 ) ;
  assign n1532 = ( n1258 & n1259 ) | ( n1258 & n1531 ) | ( n1259 & n1531 ) ;
  assign n1533 = ( ~n1265 & n1440 ) | ( ~n1265 & n1527 ) | ( n1440 & n1527 ) ;
  assign n1534 = ( n1440 & n1532 ) | ( n1440 & ~n1533 ) | ( n1532 & ~n1533 ) ;
  assign n1535 = ( ~n1528 & n1529 ) | ( ~n1528 & n1534 ) | ( n1529 & n1534 ) ;
  assign n1536 = ( n1528 & n1529 ) | ( n1528 & n1534 ) | ( n1529 & n1534 ) ;
  assign n1537 = n1528 & ~n1529 ;
  assign n1538 = ( n1535 & ~n1536 ) | ( n1535 & n1537 ) | ( ~n1536 & n1537 ) ;
  assign n1539 = n489 & n918 ;
  assign n1540 = ( n194 & ~n489 ) | ( n194 & n918 ) | ( ~n489 & n918 ) ;
  assign n1541 = ( ~n918 & n1539 ) | ( ~n918 & n1540 ) | ( n1539 & n1540 ) ;
  assign n1542 = ( ~n193 & n705 ) | ( ~n193 & n1541 ) | ( n705 & n1541 ) ;
  assign n1543 = ( n705 & n927 ) | ( n705 & ~n1541 ) | ( n927 & ~n1541 ) ;
  assign n1544 = ~n1542 & n1543 ;
  assign n1545 = ( ~n192 & n813 ) | ( ~n192 & n863 ) | ( n813 & n863 ) ;
  assign n1546 = ( n192 & n813 ) | ( n192 & ~n863 ) | ( n813 & ~n863 ) ;
  assign n1547 = n1545 & n1546 ;
  assign n1548 = ( n483 & n967 ) | ( n483 & ~n1547 ) | ( n967 & ~n1547 ) ;
  assign n1549 = ( n483 & ~n969 ) | ( n483 & n1547 ) | ( ~n969 & n1547 ) ;
  assign n1550 = n1548 & ~n1549 ;
  assign n1551 = ( n1459 & n1544 ) | ( n1459 & n1550 ) | ( n1544 & n1550 ) ;
  assign n1552 = ( ~n1459 & n1544 ) | ( ~n1459 & n1550 ) | ( n1544 & n1550 ) ;
  assign n1553 = ( n1459 & ~n1551 ) | ( n1459 & n1552 ) | ( ~n1551 & n1552 ) ;
  assign n1554 = ( n631 & ~n687 ) | ( n631 & n939 ) | ( ~n687 & n939 ) ;
  assign n1555 = ( n631 & n687 ) | ( n631 & ~n939 ) | ( n687 & ~n939 ) ;
  assign n1556 = n1554 & n1555 ;
  assign n1557 = ( n696 & n819 ) | ( n696 & ~n1556 ) | ( n819 & ~n1556 ) ;
  assign n1558 = ( ~n698 & n819 ) | ( ~n698 & n1556 ) | ( n819 & n1556 ) ;
  assign n1559 = n1557 & ~n1558 ;
  assign n1560 = ( n751 & n758 ) | ( n751 & ~n1466 ) | ( n758 & ~n1466 ) ;
  assign n1561 = ( n758 & ~n1370 ) | ( n758 & n1560 ) | ( ~n1370 & n1560 ) ;
  assign n1562 = ( ~n1379 & n1559 ) | ( ~n1379 & n1561 ) | ( n1559 & n1561 ) ;
  assign n1563 = ( n1559 & n1561 ) | ( n1559 & ~n1562 ) | ( n1561 & ~n1562 ) ;
  assign n1564 = ( n1379 & n1562 ) | ( n1379 & ~n1563 ) | ( n1562 & ~n1563 ) ;
  assign n1565 = ( n1482 & n1553 ) | ( n1482 & ~n1564 ) | ( n1553 & ~n1564 ) ;
  assign n1566 = ( ~n1482 & n1553 ) | ( ~n1482 & n1564 ) | ( n1553 & n1564 ) ;
  assign n1567 = ( ~n1553 & n1565 ) | ( ~n1553 & n1566 ) | ( n1565 & n1566 ) ;
  assign n1568 = ( n1462 & n1485 ) | ( n1462 & ~n1567 ) | ( n1485 & ~n1567 ) ;
  assign n1569 = ( n1462 & n1485 ) | ( n1462 & n1567 ) | ( n1485 & n1567 ) ;
  assign n1570 = ( n1567 & n1568 ) | ( n1567 & ~n1569 ) | ( n1568 & ~n1569 ) ;
  assign n1571 = ( ~n1488 & n1491 ) | ( ~n1488 & n1570 ) | ( n1491 & n1570 ) ;
  assign n1572 = ( n1491 & n1570 ) | ( n1491 & ~n1571 ) | ( n1570 & ~n1571 ) ;
  assign n1573 = ( n1488 & n1571 ) | ( n1488 & ~n1572 ) | ( n1571 & ~n1572 ) ;
  assign n1574 = n104 & n202 ;
  assign n1575 = n533 | n1574 ;
  assign n1576 = n573 | n1575 ;
  assign n1577 = ( n224 & n253 ) | ( n224 & ~n386 ) | ( n253 & ~n386 ) ;
  assign n1578 = ( n265 & n276 ) | ( n265 & ~n1577 ) | ( n276 & ~n1577 ) ;
  assign n1579 = n1577 | n1578 ;
  assign n1580 = n229 | n428 ;
  assign n1581 = n656 | n1580 ;
  assign n1582 = ( n1576 & ~n1579 ) | ( n1576 & n1581 ) | ( ~n1579 & n1581 ) ;
  assign n1583 = ( n438 & n1579 ) | ( n438 & ~n1582 ) | ( n1579 & ~n1582 ) ;
  assign n1584 = n1582 | n1583 ;
  assign n1585 = ( n164 & n283 ) | ( n164 & ~n602 ) | ( n283 & ~n602 ) ;
  assign n1586 = ( n109 & n270 ) | ( n109 & ~n1585 ) | ( n270 & ~n1585 ) ;
  assign n1587 = n1585 | n1586 ;
  assign n1588 = ( n387 & n454 ) | ( n387 & ~n1587 ) | ( n454 & ~n1587 ) ;
  assign n1589 = n1587 | n1588 ;
  assign n1590 = n278 | n363 ;
  assign n1591 = n850 | n1590 ;
  assign n1592 = ( n115 & n201 ) | ( n115 & n539 ) | ( n201 & n539 ) ;
  assign n1593 = ( n132 & n539 ) | ( n132 & ~n1592 ) | ( n539 & ~n1592 ) ;
  assign n1594 = n1592 | n1593 ;
  assign n1595 = ( ~n1589 & n1591 ) | ( ~n1589 & n1594 ) | ( n1591 & n1594 ) ;
  assign n1596 = n1589 | n1595 ;
  assign n1597 = ( n56 & n189 ) | ( n56 & n237 ) | ( n189 & n237 ) ;
  assign n1598 = ( n84 & ~n174 ) | ( n84 & n202 ) | ( ~n174 & n202 ) ;
  assign n1599 = ( n127 & ~n226 ) | ( n127 & n1598 ) | ( ~n226 & n1598 ) ;
  assign n1600 = n226 | n1599 ;
  assign n1601 = ( n385 & n651 ) | ( n385 & ~n1597 ) | ( n651 & ~n1597 ) ;
  assign n1602 = ( n1597 & ~n1600 ) | ( n1597 & n1601 ) | ( ~n1600 & n1601 ) ;
  assign n1603 = n133 | n800 ;
  assign n1604 = ( n342 & ~n1597 ) | ( n342 & n1603 ) | ( ~n1597 & n1603 ) ;
  assign n1605 = n1600 | n1604 ;
  assign n1606 = n1602 | n1605 ;
  assign n1607 = ( ~n442 & n670 ) | ( ~n442 & n1606 ) | ( n670 & n1606 ) ;
  assign n1608 = n442 | n1607 ;
  assign n1609 = ( ~n1584 & n1596 ) | ( ~n1584 & n1608 ) | ( n1596 & n1608 ) ;
  assign n1610 = n1584 | n1609 ;
  assign n1611 = ( n1508 & n1573 ) | ( n1508 & ~n1610 ) | ( n1573 & ~n1610 ) ;
  assign n1612 = ( ~n1508 & n1573 ) | ( ~n1508 & n1610 ) | ( n1573 & n1610 ) ;
  assign n1613 = ( ~n1573 & n1611 ) | ( ~n1573 & n1612 ) | ( n1611 & n1612 ) ;
  assign n1614 = ( n1510 & n1515 ) | ( n1510 & n1613 ) | ( n1515 & n1613 ) ;
  assign n1615 = ( ~n1510 & n1515 ) | ( ~n1510 & n1613 ) | ( n1515 & n1613 ) ;
  assign n1616 = ( n1510 & ~n1614 ) | ( n1510 & n1615 ) | ( ~n1614 & n1615 ) ;
  assign n1617 = n1439 & n1616 ;
  assign n1618 = n1449 & n1613 ;
  assign n1619 = n1450 & n1510 ;
  assign n1620 = n1260 | n1431 ;
  assign n1621 = ( ~n1431 & n1619 ) | ( ~n1431 & n1620 ) | ( n1619 & n1620 ) ;
  assign n1622 = ( ~n1617 & n1618 ) | ( ~n1617 & n1621 ) | ( n1618 & n1621 ) ;
  assign n1623 = ( ~n1262 & n1617 ) | ( ~n1262 & n1622 ) | ( n1617 & n1622 ) ;
  assign n1624 = ( n1617 & n1622 ) | ( n1617 & ~n1623 ) | ( n1622 & ~n1623 ) ;
  assign n1625 = ( n1262 & n1623 ) | ( n1262 & ~n1624 ) | ( n1623 & ~n1624 ) ;
  assign n1626 = ( n1523 & n1538 ) | ( n1523 & n1625 ) | ( n1538 & n1625 ) ;
  assign n1627 = n1266 | n1528 ;
  assign n1628 = n1534 | n1627 ;
  assign n1629 = n1265 & ~n1526 ;
  assign n1630 = ( n199 & n500 ) | ( n199 & ~n1265 ) | ( n500 & ~n1265 ) ;
  assign n1631 = ( ~n1134 & n1524 ) | ( ~n1134 & n1630 ) | ( n1524 & n1630 ) ;
  assign n1632 = ( n1258 & n1259 ) | ( n1258 & n1631 ) | ( n1259 & n1631 ) ;
  assign n1633 = n1440 & n1531 ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = ( ~n1431 & n1629 ) | ( ~n1431 & n1634 ) | ( n1629 & n1634 ) ;
  assign n1636 = n1431 | n1434 ;
  assign n1637 = ( n1513 & n1527 ) | ( n1513 & ~n1636 ) | ( n1527 & ~n1636 ) ;
  assign n1638 = ( n1634 & ~n1635 ) | ( n1634 & n1637 ) | ( ~n1635 & n1637 ) ;
  assign n1639 = n1635 | n1638 ;
  assign n1640 = ( n500 & n1628 ) | ( n500 & ~n1639 ) | ( n1628 & ~n1639 ) ;
  assign n1641 = n500 | n1639 ;
  assign n1642 = n1628 & ~n1639 ;
  assign n1643 = ( ~n1640 & n1641 ) | ( ~n1640 & n1642 ) | ( n1641 & n1642 ) ;
  assign n1644 = ( ~n758 & n1379 ) | ( ~n758 & n1470 ) | ( n1379 & n1470 ) ;
  assign n1645 = ( n1379 & n1470 ) | ( n1379 & ~n1644 ) | ( n1470 & ~n1644 ) ;
  assign n1646 = ( n758 & n1644 ) | ( n758 & ~n1645 ) | ( n1644 & ~n1645 ) ;
  assign n1647 = ( n1551 & n1562 ) | ( n1551 & ~n1646 ) | ( n1562 & ~n1646 ) ;
  assign n1648 = ( ~n1551 & n1562 ) | ( ~n1551 & n1646 ) | ( n1562 & n1646 ) ;
  assign n1649 = ( ~n1562 & n1647 ) | ( ~n1562 & n1648 ) | ( n1647 & n1648 ) ;
  assign n1650 = ( n192 & n813 ) | ( n192 & ~n819 ) | ( n813 & ~n819 ) ;
  assign n1651 = ( ~n192 & n813 ) | ( ~n192 & n819 ) | ( n813 & n819 ) ;
  assign n1652 = n1650 & n1651 ;
  assign n1653 = ( n863 & n967 ) | ( n863 & ~n1652 ) | ( n967 & ~n1652 ) ;
  assign n1654 = ( n863 & ~n969 ) | ( n863 & n1652 ) | ( ~n969 & n1652 ) ;
  assign n1655 = n1653 & ~n1654 ;
  assign n1656 = ( n631 & ~n687 ) | ( n631 & n943 ) | ( ~n687 & n943 ) ;
  assign n1657 = ( n631 & n687 ) | ( n631 & ~n943 ) | ( n687 & ~n943 ) ;
  assign n1658 = n1656 & n1657 ;
  assign n1659 = ( n696 & n939 ) | ( n696 & ~n1658 ) | ( n939 & ~n1658 ) ;
  assign n1660 = ( ~n698 & n939 ) | ( ~n698 & n1658 ) | ( n939 & n1658 ) ;
  assign n1661 = n1659 & ~n1660 ;
  assign n1662 = n483 & n918 ;
  assign n1663 = ( n194 & ~n483 ) | ( n194 & n918 ) | ( ~n483 & n918 ) ;
  assign n1664 = ( ~n918 & n1662 ) | ( ~n918 & n1663 ) | ( n1662 & n1663 ) ;
  assign n1665 = ( n489 & n927 ) | ( n489 & ~n1664 ) | ( n927 & ~n1664 ) ;
  assign n1666 = ( ~n193 & n489 ) | ( ~n193 & n1664 ) | ( n489 & n1664 ) ;
  assign n1667 = n1665 & ~n1666 ;
  assign n1668 = ( n1655 & n1661 ) | ( n1655 & n1667 ) | ( n1661 & n1667 ) ;
  assign n1669 = ( ~n1655 & n1661 ) | ( ~n1655 & n1667 ) | ( n1661 & n1667 ) ;
  assign n1670 = ( n1655 & ~n1668 ) | ( n1655 & n1669 ) | ( ~n1668 & n1669 ) ;
  assign n1671 = ( n1565 & ~n1649 ) | ( n1565 & n1670 ) | ( ~n1649 & n1670 ) ;
  assign n1672 = ( n1565 & n1649 ) | ( n1565 & n1670 ) | ( n1649 & n1670 ) ;
  assign n1673 = ( n1649 & n1671 ) | ( n1649 & ~n1672 ) | ( n1671 & ~n1672 ) ;
  assign n1674 = ( ~n1568 & n1571 ) | ( ~n1568 & n1673 ) | ( n1571 & n1673 ) ;
  assign n1675 = ( n1571 & n1673 ) | ( n1571 & ~n1674 ) | ( n1673 & ~n1674 ) ;
  assign n1676 = ( n1568 & n1674 ) | ( n1568 & ~n1675 ) | ( n1674 & ~n1675 ) ;
  assign n1677 = ( ~n405 & n721 ) | ( ~n405 & n1274 ) | ( n721 & n1274 ) ;
  assign n1678 = n154 | n309 ;
  assign n1679 = n121 | n504 ;
  assign n1680 = n1399 | n1679 ;
  assign n1681 = ( n570 & ~n1678 ) | ( n570 & n1680 ) | ( ~n1678 & n1680 ) ;
  assign n1682 = n1678 | n1681 ;
  assign n1683 = ( n56 & n281 ) | ( n56 & n565 ) | ( n281 & n565 ) ;
  assign n1684 = n133 | n328 ;
  assign n1685 = ( n106 & n422 ) | ( n106 & ~n661 ) | ( n422 & ~n661 ) ;
  assign n1686 = ( ~n215 & n1684 ) | ( ~n215 & n1685 ) | ( n1684 & n1685 ) ;
  assign n1687 = ( n215 & ~n1683 ) | ( n215 & n1686 ) | ( ~n1683 & n1686 ) ;
  assign n1688 = n1683 | n1687 ;
  assign n1689 = ( ~n1274 & n1682 ) | ( ~n1274 & n1688 ) | ( n1682 & n1688 ) ;
  assign n1690 = ( ~n405 & n1677 ) | ( ~n405 & n1689 ) | ( n1677 & n1689 ) ;
  assign n1691 = n405 | n1690 ;
  assign n1692 = ( n1611 & n1676 ) | ( n1611 & ~n1691 ) | ( n1676 & ~n1691 ) ;
  assign n1693 = ( ~n1611 & n1676 ) | ( ~n1611 & n1691 ) | ( n1676 & n1691 ) ;
  assign n1694 = ( ~n1676 & n1692 ) | ( ~n1676 & n1693 ) | ( n1692 & n1693 ) ;
  assign n1695 = ( n1613 & n1614 ) | ( n1613 & n1694 ) | ( n1614 & n1694 ) ;
  assign n1696 = ( ~n1613 & n1614 ) | ( ~n1613 & n1694 ) | ( n1614 & n1694 ) ;
  assign n1697 = ( n1613 & ~n1695 ) | ( n1613 & n1696 ) | ( ~n1695 & n1696 ) ;
  assign n1698 = n1439 & n1697 ;
  assign n1699 = n1449 & n1694 ;
  assign n1700 = n1450 & n1613 ;
  assign n1701 = ~n1260 & n1510 ;
  assign n1702 = ( n1510 & n1700 ) | ( n1510 & ~n1701 ) | ( n1700 & ~n1701 ) ;
  assign n1703 = ( ~n1698 & n1699 ) | ( ~n1698 & n1702 ) | ( n1699 & n1702 ) ;
  assign n1704 = ( ~n1262 & n1698 ) | ( ~n1262 & n1703 ) | ( n1698 & n1703 ) ;
  assign n1705 = ( n1698 & n1703 ) | ( n1698 & ~n1704 ) | ( n1703 & ~n1704 ) ;
  assign n1706 = ( n1262 & n1704 ) | ( n1262 & ~n1705 ) | ( n1704 & ~n1705 ) ;
  assign n1707 = ( n1626 & n1643 ) | ( n1626 & n1706 ) | ( n1643 & n1706 ) ;
  assign n1708 = ( ~n192 & n813 ) | ( ~n192 & n939 ) | ( n813 & n939 ) ;
  assign n1709 = ( n192 & n813 ) | ( n192 & ~n939 ) | ( n813 & ~n939 ) ;
  assign n1710 = n1708 & n1709 ;
  assign n1711 = ( n819 & n967 ) | ( n819 & ~n1710 ) | ( n967 & ~n1710 ) ;
  assign n1712 = ( n819 & ~n969 ) | ( n819 & n1710 ) | ( ~n969 & n1710 ) ;
  assign n1713 = n1711 & ~n1712 ;
  assign n1714 = ( n629 & n695 ) | ( n629 & n1656 ) | ( n695 & n1656 ) ;
  assign n1715 = ( n695 & ~n1465 ) | ( n695 & n1714 ) | ( ~n1465 & n1714 ) ;
  assign n1716 = ( ~n1539 & n1713 ) | ( ~n1539 & n1715 ) | ( n1713 & n1715 ) ;
  assign n1717 = ( n1713 & n1715 ) | ( n1713 & ~n1716 ) | ( n1715 & ~n1716 ) ;
  assign n1718 = ( n1539 & n1716 ) | ( n1539 & ~n1717 ) | ( n1716 & ~n1717 ) ;
  assign n1719 = n194 & ~n863 ;
  assign n1720 = ( ~n193 & n483 ) | ( ~n193 & n1719 ) | ( n483 & n1719 ) ;
  assign n1721 = ( n483 & n927 ) | ( n483 & ~n1719 ) | ( n927 & ~n1719 ) ;
  assign n1722 = ~n1720 & n1721 ;
  assign n1723 = ( n1644 & n1668 ) | ( n1644 & n1722 ) | ( n1668 & n1722 ) ;
  assign n1724 = ( n1644 & ~n1668 ) | ( n1644 & n1722 ) | ( ~n1668 & n1722 ) ;
  assign n1725 = ( n1668 & ~n1723 ) | ( n1668 & n1724 ) | ( ~n1723 & n1724 ) ;
  assign n1726 = ( n1647 & ~n1718 ) | ( n1647 & n1725 ) | ( ~n1718 & n1725 ) ;
  assign n1727 = ( n1647 & n1718 ) | ( n1647 & n1725 ) | ( n1718 & n1725 ) ;
  assign n1728 = ( n1718 & n1726 ) | ( n1718 & ~n1727 ) | ( n1726 & ~n1727 ) ;
  assign n1729 = ( ~n1671 & n1674 ) | ( ~n1671 & n1728 ) | ( n1674 & n1728 ) ;
  assign n1730 = ( n1674 & n1728 ) | ( n1674 & ~n1729 ) | ( n1728 & ~n1729 ) ;
  assign n1731 = ( n1671 & n1729 ) | ( n1671 & ~n1730 ) | ( n1729 & ~n1730 ) ;
  assign n1732 = n133 | n565 ;
  assign n1733 = ( ~n246 & n329 ) | ( ~n246 & n1732 ) | ( n329 & n1732 ) ;
  assign n1734 = ( n84 & n163 ) | ( n84 & n246 ) | ( n163 & n246 ) ;
  assign n1735 = n1733 | n1734 ;
  assign n1736 = n328 | n529 ;
  assign n1737 = n736 | n835 ;
  assign n1738 = ( n56 & n220 ) | ( n56 & n378 ) | ( n220 & n378 ) ;
  assign n1739 = ( ~n1736 & n1737 ) | ( ~n1736 & n1738 ) | ( n1737 & n1738 ) ;
  assign n1740 = n1736 | n1739 ;
  assign n1741 = ( n57 & n135 ) | ( n57 & n252 ) | ( n135 & n252 ) ;
  assign n1742 = ( n98 & n126 ) | ( n98 & n206 ) | ( n126 & n206 ) ;
  assign n1743 = ( n104 & n105 ) | ( n104 & n202 ) | ( n105 & n202 ) ;
  assign n1744 = n1742 | n1743 ;
  assign n1745 = ( n186 & ~n1741 ) | ( n186 & n1744 ) | ( ~n1741 & n1744 ) ;
  assign n1746 = n1741 | n1745 ;
  assign n1747 = ( ~n1735 & n1740 ) | ( ~n1735 & n1746 ) | ( n1740 & n1746 ) ;
  assign n1748 = ( n91 & n111 ) | ( n91 & ~n174 ) | ( n111 & ~n174 ) ;
  assign n1749 = n464 | n1748 ;
  assign n1750 = ( n122 & n387 ) | ( n122 & ~n617 ) | ( n387 & ~n617 ) ;
  assign n1751 = n617 | n1750 ;
  assign n1752 = ( n212 & n772 ) | ( n212 & ~n1751 ) | ( n772 & ~n1751 ) ;
  assign n1753 = n1751 | n1752 ;
  assign n1754 = ( n425 & n1598 ) | ( n425 & ~n1751 ) | ( n1598 & ~n1751 ) ;
  assign n1755 = n468 | n509 ;
  assign n1756 = n1754 | n1755 ;
  assign n1757 = n1753 | n1756 ;
  assign n1758 = ( n1735 & ~n1749 ) | ( n1735 & n1757 ) | ( ~n1749 & n1757 ) ;
  assign n1759 = ( ~n1747 & n1749 ) | ( ~n1747 & n1758 ) | ( n1749 & n1758 ) ;
  assign n1760 = n1747 | n1759 ;
  assign n1761 = ( n1692 & n1731 ) | ( n1692 & ~n1760 ) | ( n1731 & ~n1760 ) ;
  assign n1762 = ( ~n1692 & n1731 ) | ( ~n1692 & n1760 ) | ( n1731 & n1760 ) ;
  assign n1763 = ( ~n1731 & n1761 ) | ( ~n1731 & n1762 ) | ( n1761 & n1762 ) ;
  assign n1764 = ( n1694 & n1695 ) | ( n1694 & n1763 ) | ( n1695 & n1763 ) ;
  assign n1765 = ( ~n1694 & n1695 ) | ( ~n1694 & n1763 ) | ( n1695 & n1763 ) ;
  assign n1766 = ( n1694 & ~n1764 ) | ( n1694 & n1765 ) | ( ~n1764 & n1765 ) ;
  assign n1767 = n1439 & n1766 ;
  assign n1768 = n1449 & n1763 ;
  assign n1769 = n1450 & n1694 ;
  assign n1770 = ~n1260 & n1613 ;
  assign n1771 = ( n1613 & n1769 ) | ( n1613 & ~n1770 ) | ( n1769 & ~n1770 ) ;
  assign n1772 = ( ~n1767 & n1768 ) | ( ~n1767 & n1771 ) | ( n1768 & n1771 ) ;
  assign n1773 = ( ~n1262 & n1767 ) | ( ~n1262 & n1772 ) | ( n1767 & n1772 ) ;
  assign n1774 = ( n1767 & n1772 ) | ( n1767 & ~n1773 ) | ( n1772 & ~n1773 ) ;
  assign n1775 = ( n1262 & n1773 ) | ( n1262 & ~n1774 ) | ( n1773 & ~n1774 ) ;
  assign n1776 = ~n1628 & n1640 ;
  assign n1777 = n500 | n691 ;
  assign n1778 = n500 & n691 ;
  assign n1779 = n1777 & ~n1778 ;
  assign n1780 = ( n1258 & n1259 ) | ( n1258 & n1779 ) | ( n1259 & n1779 ) ;
  assign n1781 = ~n1517 & n1527 ;
  assign n1782 = n1510 & n1629 ;
  assign n1783 = n1440 & n1631 ;
  assign n1784 = ~n1431 & n1531 ;
  assign n1785 = n1783 | n1784 ;
  assign n1786 = ( ~n1781 & n1782 ) | ( ~n1781 & n1785 ) | ( n1782 & n1785 ) ;
  assign n1787 = ( ~n500 & n1781 ) | ( ~n500 & n1786 ) | ( n1781 & n1786 ) ;
  assign n1788 = ( n1781 & n1786 ) | ( n1781 & ~n1787 ) | ( n1786 & ~n1787 ) ;
  assign n1789 = ( n500 & n1787 ) | ( n500 & ~n1788 ) | ( n1787 & ~n1788 ) ;
  assign n1790 = ( n1776 & n1780 ) | ( n1776 & n1789 ) | ( n1780 & n1789 ) ;
  assign n1791 = ( ~n1776 & n1780 ) | ( ~n1776 & n1789 ) | ( n1780 & n1789 ) ;
  assign n1792 = ( n1776 & ~n1790 ) | ( n1776 & n1791 ) | ( ~n1790 & n1791 ) ;
  assign n1793 = ( n1707 & n1775 ) | ( n1707 & n1792 ) | ( n1775 & n1792 ) ;
  assign n1794 = n1527 & n1616 ;
  assign n1795 = n1613 & n1629 ;
  assign n1796 = ~n1431 & n1631 ;
  assign n1797 = n1510 & n1531 ;
  assign n1798 = n1796 | n1797 ;
  assign n1799 = ( ~n1794 & n1795 ) | ( ~n1794 & n1798 ) | ( n1795 & n1798 ) ;
  assign n1800 = ( ~n500 & n1794 ) | ( ~n500 & n1799 ) | ( n1794 & n1799 ) ;
  assign n1801 = ( n1794 & n1799 ) | ( n1794 & ~n1800 ) | ( n1799 & ~n1800 ) ;
  assign n1802 = ( n500 & n1800 ) | ( n500 & ~n1801 ) | ( n1800 & ~n1801 ) ;
  assign n1803 = n705 & ~n1780 ;
  assign n1804 = n705 & ~n756 ;
  assign n1805 = ~n705 & n756 ;
  assign n1806 = ( n1779 & n1804 ) | ( n1779 & n1805 ) | ( n1804 & n1805 ) ;
  assign n1807 = ( n1434 & n1441 ) | ( n1434 & n1806 ) | ( n1441 & n1806 ) ;
  assign n1808 = n1779 & ~n1806 ;
  assign n1809 = ( n1440 & n1807 ) | ( n1440 & n1808 ) | ( n1807 & n1808 ) ;
  assign n1810 = n691 | n756 ;
  assign n1811 = n500 & ~n756 ;
  assign n1812 = ( ~n1777 & n1810 ) | ( ~n1777 & n1811 ) | ( n1810 & n1811 ) ;
  assign n1813 = ( n1258 & n1259 ) | ( n1258 & n1812 ) | ( n1259 & n1812 ) ;
  assign n1814 = ( n1807 & ~n1809 ) | ( n1807 & n1813 ) | ( ~n1809 & n1813 ) ;
  assign n1815 = n1809 | n1814 ;
  assign n1816 = ( n705 & n1803 ) | ( n705 & n1815 ) | ( n1803 & n1815 ) ;
  assign n1817 = ( n705 & ~n1803 ) | ( n705 & n1815 ) | ( ~n1803 & n1815 ) ;
  assign n1818 = ( n1803 & ~n1816 ) | ( n1803 & n1817 ) | ( ~n1816 & n1817 ) ;
  assign n1819 = ( n1790 & n1802 ) | ( n1790 & n1818 ) | ( n1802 & n1818 ) ;
  assign n1820 = ( ~n1790 & n1802 ) | ( ~n1790 & n1818 ) | ( n1802 & n1818 ) ;
  assign n1821 = ( n1790 & ~n1819 ) | ( n1790 & n1820 ) | ( ~n1819 & n1820 ) ;
  assign n1822 = ( ~n695 & n1539 ) | ( ~n695 & n1662 ) | ( n1539 & n1662 ) ;
  assign n1823 = ( n1539 & n1662 ) | ( n1539 & ~n1822 ) | ( n1662 & ~n1822 ) ;
  assign n1824 = ( n695 & n1822 ) | ( n695 & ~n1823 ) | ( n1822 & ~n1823 ) ;
  assign n1825 = n819 & n918 ;
  assign n1826 = ( n194 & ~n819 ) | ( n194 & n918 ) | ( ~n819 & n918 ) ;
  assign n1827 = ( ~n918 & n1825 ) | ( ~n918 & n1826 ) | ( n1825 & n1826 ) ;
  assign n1828 = ( n863 & n927 ) | ( n863 & ~n1827 ) | ( n927 & ~n1827 ) ;
  assign n1829 = ( ~n193 & n863 ) | ( ~n193 & n1827 ) | ( n863 & n1827 ) ;
  assign n1830 = n1828 & ~n1829 ;
  assign n1831 = ( ~n192 & n813 ) | ( ~n192 & n943 ) | ( n813 & n943 ) ;
  assign n1832 = ( n192 & n813 ) | ( n192 & ~n943 ) | ( n813 & ~n943 ) ;
  assign n1833 = n1831 & n1832 ;
  assign n1834 = ( n939 & n967 ) | ( n939 & ~n1833 ) | ( n967 & ~n1833 ) ;
  assign n1835 = ( n939 & ~n969 ) | ( n939 & n1833 ) | ( ~n969 & n1833 ) ;
  assign n1836 = n1834 & ~n1835 ;
  assign n1837 = ( n1716 & n1830 ) | ( n1716 & n1836 ) | ( n1830 & n1836 ) ;
  assign n1838 = ( n1716 & ~n1830 ) | ( n1716 & n1836 ) | ( ~n1830 & n1836 ) ;
  assign n1839 = ( n1830 & ~n1837 ) | ( n1830 & n1838 ) | ( ~n1837 & n1838 ) ;
  assign n1840 = ( n1723 & ~n1824 ) | ( n1723 & n1839 ) | ( ~n1824 & n1839 ) ;
  assign n1841 = ( n1723 & n1824 ) | ( n1723 & n1839 ) | ( n1824 & n1839 ) ;
  assign n1842 = ( n1824 & n1840 ) | ( n1824 & ~n1841 ) | ( n1840 & ~n1841 ) ;
  assign n1843 = ( ~n1726 & n1729 ) | ( ~n1726 & n1842 ) | ( n1729 & n1842 ) ;
  assign n1844 = ( n1729 & n1842 ) | ( n1729 & ~n1843 ) | ( n1842 & ~n1843 ) ;
  assign n1845 = ( n1726 & n1843 ) | ( n1726 & ~n1844 ) | ( n1843 & ~n1844 ) ;
  assign n1846 = n207 | n270 ;
  assign n1847 = ( n380 & n617 ) | ( n380 & ~n1846 ) | ( n617 & ~n1846 ) ;
  assign n1848 = n1846 | n1847 ;
  assign n1849 = ( n406 & n598 ) | ( n406 & ~n1848 ) | ( n598 & ~n1848 ) ;
  assign n1850 = n1848 | n1849 ;
  assign n1851 = n106 | n363 ;
  assign n1852 = ( n308 & n410 ) | ( n308 & ~n1851 ) | ( n410 & ~n1851 ) ;
  assign n1853 = n1851 | n1852 ;
  assign n1854 = ( n222 & ~n286 ) | ( n222 & n1853 ) | ( ~n286 & n1853 ) ;
  assign n1855 = ~n1853 & n1854 ;
  assign n1856 = ( n842 & n1406 ) | ( n842 & n1855 ) | ( n1406 & n1855 ) ;
  assign n1857 = ( n1850 & n1855 ) | ( n1850 & ~n1856 ) | ( n1855 & ~n1856 ) ;
  assign n1858 = n255 | n364 ;
  assign n1859 = ( n56 & n227 ) | ( n56 & n283 ) | ( n227 & n283 ) ;
  assign n1860 = ( n111 & n395 ) | ( n111 & n396 ) | ( n395 & n396 ) ;
  assign n1861 = ( n340 & ~n1859 ) | ( n340 & n1860 ) | ( ~n1859 & n1860 ) ;
  assign n1862 = ( n651 & ~n1859 ) | ( n651 & n1861 ) | ( ~n1859 & n1861 ) ;
  assign n1863 = ( n73 & n105 ) | ( n73 & n202 ) | ( n105 & n202 ) ;
  assign n1864 = n187 | n1863 ;
  assign n1865 = n236 | n248 ;
  assign n1866 = ( n467 & n1231 ) | ( n467 & ~n1865 ) | ( n1231 & ~n1865 ) ;
  assign n1867 = n1865 | n1866 ;
  assign n1868 = ( n50 & ~n56 ) | ( n50 & n91 ) | ( ~n56 & n91 ) ;
  assign n1869 = ( n101 & n609 ) | ( n101 & n1868 ) | ( n609 & n1868 ) ;
  assign n1870 = ( n100 & n428 ) | ( n100 & n1869 ) | ( n428 & n1869 ) ;
  assign n1871 = ( ~n1864 & n1867 ) | ( ~n1864 & n1870 ) | ( n1867 & n1870 ) ;
  assign n1872 = ( ~n651 & n1864 ) | ( ~n651 & n1871 ) | ( n1864 & n1871 ) ;
  assign n1873 = ( n1859 & ~n1862 ) | ( n1859 & n1872 ) | ( ~n1862 & n1872 ) ;
  assign n1874 = n1862 | n1873 ;
  assign n1875 = ( n379 & ~n1858 ) | ( n379 & n1874 ) | ( ~n1858 & n1874 ) ;
  assign n1876 = n1858 | n1875 ;
  assign n1877 = n211 | n895 ;
  assign n1878 = ( ~n56 & n226 ) | ( ~n56 & n281 ) | ( n226 & n281 ) ;
  assign n1879 = ( ~n138 & n1877 ) | ( ~n138 & n1878 ) | ( n1877 & n1878 ) ;
  assign n1880 = ( ~n56 & n151 ) | ( ~n56 & n408 ) | ( n151 & n408 ) ;
  assign n1881 = n564 | n1880 ;
  assign n1882 = ( ~n56 & n243 ) | ( ~n56 & n796 ) | ( n243 & n796 ) ;
  assign n1883 = n526 | n1882 ;
  assign n1884 = ( ~n895 & n1881 ) | ( ~n895 & n1883 ) | ( n1881 & n1883 ) ;
  assign n1885 = ( n138 & ~n1879 ) | ( n138 & n1884 ) | ( ~n1879 & n1884 ) ;
  assign n1886 = n1879 | n1885 ;
  assign n1887 = ( n1850 & ~n1876 ) | ( n1850 & n1886 ) | ( ~n1876 & n1886 ) ;
  assign n1888 = ( n1857 & n1876 ) | ( n1857 & n1887 ) | ( n1876 & n1887 ) ;
  assign n1889 = n1857 & ~n1888 ;
  assign n1890 = ( n1761 & n1845 ) | ( n1761 & n1889 ) | ( n1845 & n1889 ) ;
  assign n1891 = ( ~n1761 & n1845 ) | ( ~n1761 & n1889 ) | ( n1845 & n1889 ) ;
  assign n1892 = ( n1761 & ~n1890 ) | ( n1761 & n1891 ) | ( ~n1890 & n1891 ) ;
  assign n1893 = ( n1763 & n1764 ) | ( n1763 & ~n1892 ) | ( n1764 & ~n1892 ) ;
  assign n1894 = ( ~n1763 & n1764 ) | ( ~n1763 & n1892 ) | ( n1764 & n1892 ) ;
  assign n1895 = ( ~n1764 & n1893 ) | ( ~n1764 & n1894 ) | ( n1893 & n1894 ) ;
  assign n1896 = n1439 & ~n1895 ;
  assign n1897 = n1449 & ~n1892 ;
  assign n1898 = n1450 & n1763 ;
  assign n1899 = ~n1260 & n1694 ;
  assign n1900 = ( n1694 & n1898 ) | ( n1694 & ~n1899 ) | ( n1898 & ~n1899 ) ;
  assign n1901 = ( ~n1896 & n1897 ) | ( ~n1896 & n1900 ) | ( n1897 & n1900 ) ;
  assign n1902 = ( ~n1262 & n1896 ) | ( ~n1262 & n1901 ) | ( n1896 & n1901 ) ;
  assign n1903 = ( n1896 & n1901 ) | ( n1896 & ~n1902 ) | ( n1901 & ~n1902 ) ;
  assign n1904 = ( n1262 & n1902 ) | ( n1262 & ~n1903 ) | ( n1902 & ~n1903 ) ;
  assign n1905 = ( n1793 & n1821 ) | ( n1793 & n1904 ) | ( n1821 & n1904 ) ;
  assign n1906 = n1527 & n1697 ;
  assign n1907 = n1629 & n1694 ;
  assign n1908 = n1510 & n1631 ;
  assign n1909 = n1531 & n1613 ;
  assign n1910 = n1908 | n1909 ;
  assign n1911 = ( ~n1906 & n1907 ) | ( ~n1906 & n1910 ) | ( n1907 & n1910 ) ;
  assign n1912 = ( ~n500 & n1906 ) | ( ~n500 & n1911 ) | ( n1906 & n1911 ) ;
  assign n1913 = ( n1906 & n1911 ) | ( n1906 & ~n1912 ) | ( n1911 & ~n1912 ) ;
  assign n1914 = ( n500 & n1912 ) | ( n500 & ~n1913 ) | ( n1912 & ~n1913 ) ;
  assign n1915 = n500 & n705 ;
  assign n1916 = ( n705 & n1805 ) | ( n705 & ~n1915 ) | ( n1805 & ~n1915 ) ;
  assign n1917 = ( n1778 & ~n1810 ) | ( n1778 & n1916 ) | ( ~n1810 & n1916 ) ;
  assign n1918 = ( n1258 & n1259 ) | ( n1258 & n1917 ) | ( n1259 & n1917 ) ;
  assign n1919 = n1440 & n1812 ;
  assign n1920 = n1918 | n1919 ;
  assign n1921 = ( ~n1431 & n1808 ) | ( ~n1431 & n1920 ) | ( n1808 & n1920 ) ;
  assign n1922 = ( n1513 & ~n1636 ) | ( n1513 & n1806 ) | ( ~n1636 & n1806 ) ;
  assign n1923 = ( n1920 & ~n1921 ) | ( n1920 & n1922 ) | ( ~n1921 & n1922 ) ;
  assign n1924 = n1921 | n1923 ;
  assign n1925 = n705 & n1817 ;
  assign n1926 = n1924 | n1925 ;
  assign n1927 = ( n1924 & n1925 ) | ( n1924 & ~n1926 ) | ( n1925 & ~n1926 ) ;
  assign n1928 = n1926 & ~n1927 ;
  assign n1929 = ( n1819 & n1914 ) | ( n1819 & n1928 ) | ( n1914 & n1928 ) ;
  assign n1930 = ( ~n1819 & n1914 ) | ( ~n1819 & n1928 ) | ( n1914 & n1928 ) ;
  assign n1931 = ( n1819 & ~n1929 ) | ( n1819 & n1930 ) | ( ~n1929 & n1930 ) ;
  assign n1932 = n863 & n918 ;
  assign n1933 = ~n810 & n943 ;
  assign n1934 = n943 & n969 ;
  assign n1935 = ( n811 & ~n1933 ) | ( n811 & n1934 ) | ( ~n1933 & n1934 ) ;
  assign n1936 = n194 & ~n939 ;
  assign n1937 = ( ~n193 & n819 ) | ( ~n193 & n1936 ) | ( n819 & n1936 ) ;
  assign n1938 = ( n819 & n927 ) | ( n819 & ~n1936 ) | ( n927 & ~n1936 ) ;
  assign n1939 = ~n1937 & n1938 ;
  assign n1940 = ( ~n1932 & n1935 ) | ( ~n1932 & n1939 ) | ( n1935 & n1939 ) ;
  assign n1941 = ( n1935 & n1939 ) | ( n1935 & ~n1940 ) | ( n1939 & ~n1940 ) ;
  assign n1942 = ( n1932 & n1940 ) | ( n1932 & ~n1941 ) | ( n1940 & ~n1941 ) ;
  assign n1943 = ( n1822 & n1837 ) | ( n1822 & ~n1942 ) | ( n1837 & ~n1942 ) ;
  assign n1944 = ( ~n1822 & n1837 ) | ( ~n1822 & n1942 ) | ( n1837 & n1942 ) ;
  assign n1945 = ( ~n1837 & n1943 ) | ( ~n1837 & n1944 ) | ( n1943 & n1944 ) ;
  assign n1946 = ( ~n1840 & n1843 ) | ( ~n1840 & n1945 ) | ( n1843 & n1945 ) ;
  assign n1947 = ( n1843 & n1945 ) | ( n1843 & ~n1946 ) | ( n1945 & ~n1946 ) ;
  assign n1948 = ( n1840 & n1946 ) | ( n1840 & ~n1947 ) | ( n1946 & ~n1947 ) ;
  assign n1949 = n229 | n670 ;
  assign n1950 = ( n1244 & ~n1883 ) | ( n1244 & n1949 ) | ( ~n1883 & n1949 ) ;
  assign n1951 = n1883 | n1950 ;
  assign n1952 = n169 | n205 ;
  assign n1953 = ( n665 & n772 ) | ( n665 & ~n1952 ) | ( n772 & ~n1952 ) ;
  assign n1954 = n1952 | n1953 ;
  assign n1955 = ( ~n1874 & n1951 ) | ( ~n1874 & n1954 ) | ( n1951 & n1954 ) ;
  assign n1956 = n228 | n234 ;
  assign n1957 = n144 | n150 ;
  assign n1958 = n520 | n1957 ;
  assign n1959 = ( n468 & ~n1956 ) | ( n468 & n1958 ) | ( ~n1956 & n1958 ) ;
  assign n1960 = n1956 | n1959 ;
  assign n1961 = ( n283 & n347 ) | ( n283 & ~n602 ) | ( n347 & ~n602 ) ;
  assign n1962 = ( n789 & n1738 ) | ( n789 & ~n1961 ) | ( n1738 & ~n1961 ) ;
  assign n1963 = n1961 | n1962 ;
  assign n1964 = ( n683 & ~n1960 ) | ( n683 & n1963 ) | ( ~n1960 & n1963 ) ;
  assign n1965 = n1960 | n1964 ;
  assign n1966 = ( n1874 & ~n1955 ) | ( n1874 & n1965 ) | ( ~n1955 & n1965 ) ;
  assign n1967 = n1955 | n1966 ;
  assign n1968 = ( n1890 & n1948 ) | ( n1890 & ~n1967 ) | ( n1948 & ~n1967 ) ;
  assign n1969 = ( ~n1890 & n1948 ) | ( ~n1890 & n1967 ) | ( n1948 & n1967 ) ;
  assign n1970 = ( ~n1948 & n1968 ) | ( ~n1948 & n1969 ) | ( n1968 & n1969 ) ;
  assign n1971 = ( ~n1892 & n1893 ) | ( ~n1892 & n1970 ) | ( n1893 & n1970 ) ;
  assign n1972 = ( n1892 & n1893 ) | ( n1892 & ~n1970 ) | ( n1893 & ~n1970 ) ;
  assign n1973 = ( ~n1893 & n1971 ) | ( ~n1893 & n1972 ) | ( n1971 & n1972 ) ;
  assign n1974 = n1439 & ~n1973 ;
  assign n1975 = ~n25 & n1763 ;
  assign n1976 = ( n1262 & n1974 ) | ( n1262 & ~n1975 ) | ( n1974 & ~n1975 ) ;
  assign n1977 = n1450 & ~n1892 ;
  assign n1978 = n1449 & n1970 ;
  assign n1979 = n1977 | n1978 ;
  assign n1980 = ( ~n1974 & n1976 ) | ( ~n1974 & n1979 ) | ( n1976 & n1979 ) ;
  assign n1981 = n1976 & ~n1979 ;
  assign n1982 = ( ~n1262 & n1980 ) | ( ~n1262 & n1981 ) | ( n1980 & n1981 ) ;
  assign n1983 = ( n1905 & n1931 ) | ( n1905 & n1982 ) | ( n1931 & n1982 ) ;
  assign n1984 = n1527 & n1766 ;
  assign n1985 = n1629 & n1763 ;
  assign n1986 = n1613 & n1631 ;
  assign n1987 = n1531 & n1694 ;
  assign n1988 = n1986 | n1987 ;
  assign n1989 = ( ~n1984 & n1985 ) | ( ~n1984 & n1988 ) | ( n1985 & n1988 ) ;
  assign n1990 = ( ~n500 & n1984 ) | ( ~n500 & n1989 ) | ( n1984 & n1989 ) ;
  assign n1991 = ( n1984 & n1989 ) | ( n1984 & ~n1990 ) | ( n1989 & ~n1990 ) ;
  assign n1992 = ( n500 & n1990 ) | ( n500 & ~n1991 ) | ( n1990 & ~n1991 ) ;
  assign n1993 = n1803 & ~n1815 ;
  assign n1994 = ~n1924 & n1993 ;
  assign n1995 = ( ~n481 & n487 ) | ( ~n481 & n705 ) | ( n487 & n705 ) ;
  assign n1996 = n489 & n705 ;
  assign n1997 = ( n489 & n1995 ) | ( n489 & ~n1996 ) | ( n1995 & ~n1996 ) ;
  assign n1998 = ( n1258 & n1259 ) | ( n1258 & n1997 ) | ( n1259 & n1997 ) ;
  assign n1999 = ~n1517 & n1806 ;
  assign n2000 = n1510 & n1808 ;
  assign n2001 = n1431 | n1812 ;
  assign n2002 = n1440 & n1917 ;
  assign n2003 = ( ~n1431 & n2001 ) | ( ~n1431 & n2002 ) | ( n2001 & n2002 ) ;
  assign n2004 = ( ~n1999 & n2000 ) | ( ~n1999 & n2003 ) | ( n2000 & n2003 ) ;
  assign n2005 = ( n705 & ~n1999 ) | ( n705 & n2004 ) | ( ~n1999 & n2004 ) ;
  assign n2006 = ( n705 & n2004 ) | ( n705 & ~n2005 ) | ( n2004 & ~n2005 ) ;
  assign n2007 = ( n1999 & n2005 ) | ( n1999 & ~n2006 ) | ( n2005 & ~n2006 ) ;
  assign n2008 = ( n1994 & n1998 ) | ( n1994 & n2007 ) | ( n1998 & n2007 ) ;
  assign n2009 = ( ~n1994 & n1998 ) | ( ~n1994 & n2007 ) | ( n1998 & n2007 ) ;
  assign n2010 = ( n1994 & ~n2008 ) | ( n1994 & n2009 ) | ( ~n2008 & n2009 ) ;
  assign n2011 = ( n1929 & n1992 ) | ( n1929 & n2010 ) | ( n1992 & n2010 ) ;
  assign n2012 = ( ~n1929 & n1992 ) | ( ~n1929 & n2010 ) | ( n1992 & n2010 ) ;
  assign n2013 = ( n1929 & ~n2011 ) | ( n1929 & n2012 ) | ( ~n2011 & n2012 ) ;
  assign n2014 = ( ~n811 & n1825 ) | ( ~n811 & n1932 ) | ( n1825 & n1932 ) ;
  assign n2015 = ( n1825 & n1932 ) | ( n1825 & ~n2014 ) | ( n1932 & ~n2014 ) ;
  assign n2016 = ( n811 & n2014 ) | ( n811 & ~n2015 ) | ( n2014 & ~n2015 ) ;
  assign n2017 = n918 & n943 ;
  assign n2018 = ( n194 & n918 ) | ( n194 & ~n943 ) | ( n918 & ~n943 ) ;
  assign n2019 = ( ~n918 & n2017 ) | ( ~n918 & n2018 ) | ( n2017 & n2018 ) ;
  assign n2020 = ( n927 & n939 ) | ( n927 & ~n2019 ) | ( n939 & ~n2019 ) ;
  assign n2021 = ( ~n193 & n939 ) | ( ~n193 & n2019 ) | ( n939 & n2019 ) ;
  assign n2022 = n2020 & ~n2021 ;
  assign n2023 = ( n1940 & ~n2016 ) | ( n1940 & n2022 ) | ( ~n2016 & n2022 ) ;
  assign n2024 = ( n1940 & n2016 ) | ( n1940 & n2022 ) | ( n2016 & n2022 ) ;
  assign n2025 = ( n2016 & n2023 ) | ( n2016 & ~n2024 ) | ( n2023 & ~n2024 ) ;
  assign n2026 = ( ~n1943 & n1946 ) | ( ~n1943 & n2025 ) | ( n1946 & n2025 ) ;
  assign n2027 = ( n1946 & n2025 ) | ( n1946 & ~n2026 ) | ( n2025 & ~n2026 ) ;
  assign n2028 = ( n1943 & n2026 ) | ( n1943 & ~n2027 ) | ( n2026 & ~n2027 ) ;
  assign n2029 = n297 | n533 ;
  assign n2030 = ( n517 & n617 ) | ( n517 & ~n2029 ) | ( n617 & ~n2029 ) ;
  assign n2031 = n2029 | n2030 ;
  assign n2032 = n340 | n608 ;
  assign n2033 = n741 | n2032 ;
  assign n2034 = ( n433 & n460 ) | ( n433 & ~n608 ) | ( n460 & ~n608 ) ;
  assign n2035 = n137 | n166 ;
  assign n2036 = n529 | n2035 ;
  assign n2037 = ( ~n2032 & n2034 ) | ( ~n2032 & n2036 ) | ( n2034 & n2036 ) ;
  assign n2038 = ( ~n2031 & n2033 ) | ( ~n2031 & n2037 ) | ( n2033 & n2037 ) ;
  assign n2039 = n2031 | n2038 ;
  assign n2040 = ( n292 & n804 ) | ( n292 & ~n2039 ) | ( n804 & ~n2039 ) ;
  assign n2041 = n2039 | n2040 ;
  assign n2042 = ( n1968 & n2028 ) | ( n1968 & ~n2041 ) | ( n2028 & ~n2041 ) ;
  assign n2043 = ( ~n1968 & n2028 ) | ( ~n1968 & n2041 ) | ( n2028 & n2041 ) ;
  assign n2044 = ( ~n2028 & n2042 ) | ( ~n2028 & n2043 ) | ( n2042 & n2043 ) ;
  assign n2045 = ( n1970 & n1971 ) | ( n1970 & n2044 ) | ( n1971 & n2044 ) ;
  assign n2046 = ( ~n1970 & n1971 ) | ( ~n1970 & n2044 ) | ( n1971 & n2044 ) ;
  assign n2047 = ( n1970 & ~n2045 ) | ( n1970 & n2046 ) | ( ~n2045 & n2046 ) ;
  assign n2048 = n1439 & n2047 ;
  assign n2049 = n1449 & n2044 ;
  assign n2050 = n1450 & n1970 ;
  assign n2051 = n1260 | n1892 ;
  assign n2052 = ( ~n1892 & n2050 ) | ( ~n1892 & n2051 ) | ( n2050 & n2051 ) ;
  assign n2053 = ( ~n2048 & n2049 ) | ( ~n2048 & n2052 ) | ( n2049 & n2052 ) ;
  assign n2054 = ( ~n1262 & n2048 ) | ( ~n1262 & n2053 ) | ( n2048 & n2053 ) ;
  assign n2055 = ( n2048 & n2053 ) | ( n2048 & ~n2054 ) | ( n2053 & ~n2054 ) ;
  assign n2056 = ( n1262 & n2054 ) | ( n1262 & ~n2055 ) | ( n2054 & ~n2055 ) ;
  assign n2057 = ( n1983 & n2013 ) | ( n1983 & n2056 ) | ( n2013 & n2056 ) ;
  assign n2058 = n1527 & ~n1895 ;
  assign n2059 = n1629 & ~n1892 ;
  assign n2060 = n1631 & n1694 ;
  assign n2061 = n1531 & n1763 ;
  assign n2062 = n2060 | n2061 ;
  assign n2063 = ( ~n2058 & n2059 ) | ( ~n2058 & n2062 ) | ( n2059 & n2062 ) ;
  assign n2064 = ( ~n500 & n2058 ) | ( ~n500 & n2063 ) | ( n2058 & n2063 ) ;
  assign n2065 = ( n2058 & n2063 ) | ( n2058 & ~n2064 ) | ( n2063 & ~n2064 ) ;
  assign n2066 = ( n500 & n2064 ) | ( n500 & ~n2065 ) | ( n2064 & ~n2065 ) ;
  assign n2067 = n1616 & n1806 ;
  assign n2068 = n1613 & n1808 ;
  assign n2069 = n1510 & ~n1812 ;
  assign n2070 = ~n1431 & n1917 ;
  assign n2071 = ( n1510 & ~n2069 ) | ( n1510 & n2070 ) | ( ~n2069 & n2070 ) ;
  assign n2072 = ( ~n2067 & n2068 ) | ( ~n2067 & n2071 ) | ( n2068 & n2071 ) ;
  assign n2073 = ( n705 & ~n2067 ) | ( n705 & n2072 ) | ( ~n2067 & n2072 ) ;
  assign n2074 = ( n705 & n2072 ) | ( n705 & ~n2073 ) | ( n2072 & ~n2073 ) ;
  assign n2075 = ( n2067 & n2073 ) | ( n2067 & ~n2074 ) | ( n2073 & ~n2074 ) ;
  assign n2076 = ( n483 & ~n860 ) | ( n483 & n862 ) | ( ~n860 & n862 ) ;
  assign n2077 = ( n483 & ~n863 ) | ( n483 & n1997 ) | ( ~n863 & n1997 ) ;
  assign n2078 = ~n2076 & n2077 ;
  assign n2079 = n1997 & ~n2078 ;
  assign n2080 = ( n1434 & n1441 ) | ( n1434 & n2079 ) | ( n1441 & n2079 ) ;
  assign n2081 = n863 & n1998 ;
  assign n2082 = n483 | n489 ;
  assign n2083 = ( n483 & n489 ) | ( n483 & n1997 ) | ( n489 & n1997 ) ;
  assign n2084 = n2082 & ~n2083 ;
  assign n2085 = ( n1258 & n1259 ) | ( n1258 & n2084 ) | ( n1259 & n2084 ) ;
  assign n2086 = n1440 & ~n2078 ;
  assign n2087 = ( n1440 & n2085 ) | ( n1440 & ~n2086 ) | ( n2085 & ~n2086 ) ;
  assign n2088 = ( ~n2080 & n2081 ) | ( ~n2080 & n2087 ) | ( n2081 & n2087 ) ;
  assign n2089 = ( n2080 & n2081 ) | ( n2080 & n2087 ) | ( n2081 & n2087 ) ;
  assign n2090 = n2080 & ~n2081 ;
  assign n2091 = ( n2088 & ~n2089 ) | ( n2088 & n2090 ) | ( ~n2089 & n2090 ) ;
  assign n2092 = ( n2008 & n2075 ) | ( n2008 & n2091 ) | ( n2075 & n2091 ) ;
  assign n2093 = ( ~n2008 & n2075 ) | ( ~n2008 & n2091 ) | ( n2075 & n2091 ) ;
  assign n2094 = ( n2008 & ~n2092 ) | ( n2008 & n2093 ) | ( ~n2092 & n2093 ) ;
  assign n2095 = ( n2011 & n2066 ) | ( n2011 & n2094 ) | ( n2066 & n2094 ) ;
  assign n2096 = ( ~n2011 & n2066 ) | ( ~n2011 & n2094 ) | ( n2066 & n2094 ) ;
  assign n2097 = ( n2011 & ~n2095 ) | ( n2011 & n2096 ) | ( ~n2095 & n2096 ) ;
  assign n2098 = n546 | n668 ;
  assign n2099 = n890 | n2098 ;
  assign n2100 = n88 | n329 ;
  assign n2101 = ( ~n163 & n173 ) | ( ~n163 & n609 ) | ( n173 & n609 ) ;
  assign n2102 = ( n1864 & ~n2100 ) | ( n1864 & n2101 ) | ( ~n2100 & n2101 ) ;
  assign n2103 = n2100 | n2102 ;
  assign n2104 = ( n586 & ~n2099 ) | ( n586 & n2103 ) | ( ~n2099 & n2103 ) ;
  assign n2105 = n2099 | n2104 ;
  assign n2106 = ( n532 & n1236 ) | ( n532 & ~n1850 ) | ( n1236 & ~n1850 ) ;
  assign n2107 = n1850 | n2106 ;
  assign n2108 = ( n57 & n294 ) | ( n57 & n885 ) | ( n294 & n885 ) ;
  assign n2109 = ( n294 & n347 ) | ( n294 & ~n2108 ) | ( n347 & ~n2108 ) ;
  assign n2110 = n2108 | n2109 ;
  assign n2111 = ( ~n50 & n422 ) | ( ~n50 & n1868 ) | ( n422 & n1868 ) ;
  assign n2112 = ( n297 & n520 ) | ( n297 & ~n2111 ) | ( n520 & ~n2111 ) ;
  assign n2113 = n2111 | n2112 ;
  assign n2114 = n1590 | n2113 ;
  assign n2115 = ( ~n56 & n132 ) | ( ~n56 & n237 ) | ( n132 & n237 ) ;
  assign n2116 = ( n618 & ~n1590 ) | ( n618 & n2115 ) | ( ~n1590 & n2115 ) ;
  assign n2117 = ( ~n2110 & n2114 ) | ( ~n2110 & n2116 ) | ( n2114 & n2116 ) ;
  assign n2118 = n2110 | n2117 ;
  assign n2119 = ( ~n2105 & n2107 ) | ( ~n2105 & n2118 ) | ( n2107 & n2118 ) ;
  assign n2120 = n2105 | n2119 ;
  assign n2121 = n918 & n939 ;
  assign n2122 = ( n149 & n943 ) | ( n149 & n2019 ) | ( n943 & n2019 ) ;
  assign n2123 = ( n918 & ~n2017 ) | ( n918 & n2122 ) | ( ~n2017 & n2122 ) ;
  assign n2124 = ( n2014 & ~n2121 ) | ( n2014 & n2123 ) | ( ~n2121 & n2123 ) ;
  assign n2125 = ( n2014 & n2123 ) | ( n2014 & ~n2124 ) | ( n2123 & ~n2124 ) ;
  assign n2126 = ( n2121 & n2124 ) | ( n2121 & ~n2125 ) | ( n2124 & ~n2125 ) ;
  assign n2127 = ( ~n2023 & n2026 ) | ( ~n2023 & n2126 ) | ( n2026 & n2126 ) ;
  assign n2128 = ( n2026 & n2126 ) | ( n2026 & ~n2127 ) | ( n2126 & ~n2127 ) ;
  assign n2129 = ( n2023 & n2127 ) | ( n2023 & ~n2128 ) | ( n2127 & ~n2128 ) ;
  assign n2130 = ( n2042 & ~n2120 ) | ( n2042 & n2129 ) | ( ~n2120 & n2129 ) ;
  assign n2131 = ( n2042 & n2120 ) | ( n2042 & n2129 ) | ( n2120 & n2129 ) ;
  assign n2132 = ( n2120 & n2130 ) | ( n2120 & ~n2131 ) | ( n2130 & ~n2131 ) ;
  assign n2133 = ( n2044 & n2045 ) | ( n2044 & n2132 ) | ( n2045 & n2132 ) ;
  assign n2134 = ( ~n2044 & n2045 ) | ( ~n2044 & n2132 ) | ( n2045 & n2132 ) ;
  assign n2135 = ( n2044 & ~n2133 ) | ( n2044 & n2134 ) | ( ~n2133 & n2134 ) ;
  assign n2136 = n1439 & n2135 ;
  assign n2137 = ~n25 & n1970 ;
  assign n2138 = ( n1262 & n2136 ) | ( n1262 & ~n2137 ) | ( n2136 & ~n2137 ) ;
  assign n2139 = n1450 & n2044 ;
  assign n2140 = n1449 & n2132 ;
  assign n2141 = n2139 | n2140 ;
  assign n2142 = ( ~n2136 & n2138 ) | ( ~n2136 & n2141 ) | ( n2138 & n2141 ) ;
  assign n2143 = n2138 & ~n2141 ;
  assign n2144 = ( ~n1262 & n2142 ) | ( ~n1262 & n2143 ) | ( n2142 & n2143 ) ;
  assign n2145 = ( n2057 & n2097 ) | ( n2057 & n2144 ) | ( n2097 & n2144 ) ;
  assign n2146 = ( n863 & ~n1995 ) | ( n863 & n1996 ) | ( ~n1995 & n1996 ) ;
  assign n2147 = ( n2076 & ~n2082 ) | ( n2076 & n2146 ) | ( ~n2082 & n2146 ) ;
  assign n2148 = ( n1258 & n1259 ) | ( n1258 & n2147 ) | ( n1259 & n2147 ) ;
  assign n2149 = ( ~n1440 & n2082 ) | ( ~n1440 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2150 = ( n2082 & n2148 ) | ( n2082 & ~n2149 ) | ( n2148 & ~n2149 ) ;
  assign n2151 = ( ~n1431 & n2078 ) | ( ~n1431 & n2150 ) | ( n2078 & n2150 ) ;
  assign n2152 = ( n1513 & ~n1636 ) | ( n1513 & n2079 ) | ( ~n1636 & n2079 ) ;
  assign n2153 = ( n2150 & ~n2151 ) | ( n2150 & n2152 ) | ( ~n2151 & n2152 ) ;
  assign n2154 = n2151 | n2153 ;
  assign n2155 = n1998 | n2080 ;
  assign n2156 = n2087 | n2155 ;
  assign n2157 = ( n863 & ~n2154 ) | ( n863 & n2156 ) | ( ~n2154 & n2156 ) ;
  assign n2158 = n863 | n2154 ;
  assign n2159 = ~n2154 & n2156 ;
  assign n2160 = ( ~n2157 & n2158 ) | ( ~n2157 & n2159 ) | ( n2158 & n2159 ) ;
  assign n2161 = n1697 & n1806 ;
  assign n2162 = n1694 & n1808 ;
  assign n2163 = n1613 & ~n1812 ;
  assign n2164 = n1510 & n1917 ;
  assign n2165 = ( n1613 & ~n2163 ) | ( n1613 & n2164 ) | ( ~n2163 & n2164 ) ;
  assign n2166 = ( ~n2161 & n2162 ) | ( ~n2161 & n2165 ) | ( n2162 & n2165 ) ;
  assign n2167 = ( n705 & ~n2161 ) | ( n705 & n2166 ) | ( ~n2161 & n2166 ) ;
  assign n2168 = ( n705 & n2166 ) | ( n705 & ~n2167 ) | ( n2166 & ~n2167 ) ;
  assign n2169 = ( n2161 & n2167 ) | ( n2161 & ~n2168 ) | ( n2167 & ~n2168 ) ;
  assign n2170 = ( n2092 & n2160 ) | ( n2092 & n2169 ) | ( n2160 & n2169 ) ;
  assign n2171 = ( ~n2092 & n2160 ) | ( ~n2092 & n2169 ) | ( n2160 & n2169 ) ;
  assign n2172 = ( n2092 & ~n2170 ) | ( n2092 & n2171 ) | ( ~n2170 & n2171 ) ;
  assign n2173 = n1527 & ~n1973 ;
  assign n2174 = n1629 & n1970 ;
  assign n2175 = n1631 & n1763 ;
  assign n2176 = n1531 & ~n1892 ;
  assign n2177 = n2175 | n2176 ;
  assign n2178 = ( ~n2173 & n2174 ) | ( ~n2173 & n2177 ) | ( n2174 & n2177 ) ;
  assign n2179 = ( ~n500 & n2173 ) | ( ~n500 & n2178 ) | ( n2173 & n2178 ) ;
  assign n2180 = ( n2173 & n2178 ) | ( n2173 & ~n2179 ) | ( n2178 & ~n2179 ) ;
  assign n2181 = ( n500 & n2179 ) | ( n500 & ~n2180 ) | ( n2179 & ~n2180 ) ;
  assign n2182 = ( n2095 & n2172 ) | ( n2095 & n2181 ) | ( n2172 & n2181 ) ;
  assign n2183 = ( ~n2095 & n2172 ) | ( ~n2095 & n2181 ) | ( n2172 & n2181 ) ;
  assign n2184 = ( n2095 & ~n2182 ) | ( n2095 & n2183 ) | ( ~n2182 & n2183 ) ;
  assign n2185 = ( n224 & n356 ) | ( n224 & ~n386 ) | ( n356 & ~n386 ) ;
  assign n2186 = n337 | n707 ;
  assign n2187 = n2185 | n2186 ;
  assign n2188 = n326 | n440 ;
  assign n2189 = n1289 | n2188 ;
  assign n2190 = ( ~n56 & n204 ) | ( ~n56 & n427 ) | ( n204 & n427 ) ;
  assign n2191 = ( ~n1685 & n2189 ) | ( ~n1685 & n2190 ) | ( n2189 & n2190 ) ;
  assign n2192 = n1685 | n2191 ;
  assign n2193 = ( ~n123 & n222 ) | ( ~n123 & n2192 ) | ( n222 & n2192 ) ;
  assign n2194 = ~n2192 & n2193 ;
  assign n2195 = n265 | n325 ;
  assign n2196 = ( n529 & n1870 ) | ( n529 & ~n2195 ) | ( n1870 & ~n2195 ) ;
  assign n2197 = n2195 | n2196 ;
  assign n2198 = ( n2187 & n2194 ) | ( n2187 & ~n2197 ) | ( n2194 & ~n2197 ) ;
  assign n2199 = ~n2187 & n2198 ;
  assign n2200 = n263 | n462 ;
  assign n2201 = ( n1608 & n2199 ) | ( n1608 & n2200 ) | ( n2199 & n2200 ) ;
  assign n2202 = n2199 & ~n2201 ;
  assign n2203 = ~n939 & n943 ;
  assign n2204 = ( ~n54 & n939 ) | ( ~n54 & n941 ) | ( n939 & n941 ) ;
  assign n2205 = n2203 | n2204 ;
  assign n2206 = ( n900 & n917 ) | ( n900 & ~n2205 ) | ( n917 & ~n2205 ) ;
  assign n2207 = ( ~n2124 & n2127 ) | ( ~n2124 & n2206 ) | ( n2127 & n2206 ) ;
  assign n2208 = ( n2127 & n2206 ) | ( n2127 & ~n2207 ) | ( n2206 & ~n2207 ) ;
  assign n2209 = ( n2124 & n2207 ) | ( n2124 & ~n2208 ) | ( n2207 & ~n2208 ) ;
  assign n2210 = ( n2130 & n2202 ) | ( n2130 & n2209 ) | ( n2202 & n2209 ) ;
  assign n2211 = ( n2130 & ~n2202 ) | ( n2130 & n2209 ) | ( ~n2202 & n2209 ) ;
  assign n2212 = ( n2202 & ~n2210 ) | ( n2202 & n2211 ) | ( ~n2210 & n2211 ) ;
  assign n2213 = ( n2132 & n2133 ) | ( n2132 & ~n2212 ) | ( n2133 & ~n2212 ) ;
  assign n2214 = ( n2045 & ~n2134 ) | ( n2045 & n2212 ) | ( ~n2134 & n2212 ) ;
  assign n2215 = ( ~n2133 & n2213 ) | ( ~n2133 & n2214 ) | ( n2213 & n2214 ) ;
  assign n2216 = n1439 & ~n2215 ;
  assign n2217 = n1449 & ~n2212 ;
  assign n2218 = n1450 & n2132 ;
  assign n2219 = ~n1260 & n2044 ;
  assign n2220 = ( n2044 & n2218 ) | ( n2044 & ~n2219 ) | ( n2218 & ~n2219 ) ;
  assign n2221 = ( ~n2216 & n2217 ) | ( ~n2216 & n2220 ) | ( n2217 & n2220 ) ;
  assign n2222 = ( ~n1262 & n2216 ) | ( ~n1262 & n2221 ) | ( n2216 & n2221 ) ;
  assign n2223 = ( n2216 & n2221 ) | ( n2216 & ~n2222 ) | ( n2221 & ~n2222 ) ;
  assign n2224 = ( n1262 & n2222 ) | ( n1262 & ~n2223 ) | ( n2222 & ~n2223 ) ;
  assign n2225 = ( n2145 & n2184 ) | ( n2145 & n2224 ) | ( n2184 & n2224 ) ;
  assign n2226 = n1527 & n2047 ;
  assign n2227 = n1629 & n2044 ;
  assign n2228 = n1631 & ~n1892 ;
  assign n2229 = n1531 & n1970 ;
  assign n2230 = n2228 | n2229 ;
  assign n2231 = ( ~n2226 & n2227 ) | ( ~n2226 & n2230 ) | ( n2227 & n2230 ) ;
  assign n2232 = ( ~n500 & n2226 ) | ( ~n500 & n2231 ) | ( n2226 & n2231 ) ;
  assign n2233 = ( n2226 & n2231 ) | ( n2226 & ~n2232 ) | ( n2231 & ~n2232 ) ;
  assign n2234 = ( n500 & n2232 ) | ( n500 & ~n2233 ) | ( n2232 & ~n2233 ) ;
  assign n2235 = n1766 & n1806 ;
  assign n2236 = n1763 & n1808 ;
  assign n2237 = ~n1694 & n1812 ;
  assign n2238 = n1613 & n1917 ;
  assign n2239 = ( n1812 & ~n2237 ) | ( n1812 & n2238 ) | ( ~n2237 & n2238 ) ;
  assign n2240 = ( ~n2235 & n2236 ) | ( ~n2235 & n2239 ) | ( n2236 & n2239 ) ;
  assign n2241 = ( n705 & ~n2235 ) | ( n705 & n2240 ) | ( ~n2235 & n2240 ) ;
  assign n2242 = ( n705 & n2240 ) | ( n705 & ~n2241 ) | ( n2240 & ~n2241 ) ;
  assign n2243 = ( n2235 & n2241 ) | ( n2235 & ~n2242 ) | ( n2241 & ~n2242 ) ;
  assign n2244 = ~n2156 & n2157 ;
  assign n2245 = n819 | n863 ;
  assign n2246 = ( n819 & n863 ) | ( n819 & ~n2245 ) | ( n863 & ~n2245 ) ;
  assign n2247 = n2245 & ~n2246 ;
  assign n2248 = ( n1258 & n1259 ) | ( n1258 & n2247 ) | ( n1259 & n2247 ) ;
  assign n2249 = ~n1517 & n2079 ;
  assign n2250 = n1510 & n2078 ;
  assign n2251 = n1440 & n2147 ;
  assign n2252 = ( ~n1431 & n2082 ) | ( ~n1431 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2253 = ( ~n2083 & n2251 ) | ( ~n2083 & n2252 ) | ( n2251 & n2252 ) ;
  assign n2254 = ( ~n2249 & n2250 ) | ( ~n2249 & n2253 ) | ( n2250 & n2253 ) ;
  assign n2255 = ( ~n863 & n2249 ) | ( ~n863 & n2254 ) | ( n2249 & n2254 ) ;
  assign n2256 = ( n2249 & n2254 ) | ( n2249 & ~n2255 ) | ( n2254 & ~n2255 ) ;
  assign n2257 = ( n863 & n2255 ) | ( n863 & ~n2256 ) | ( n2255 & ~n2256 ) ;
  assign n2258 = ( n2244 & n2248 ) | ( n2244 & n2257 ) | ( n2248 & n2257 ) ;
  assign n2259 = ( ~n2244 & n2248 ) | ( ~n2244 & n2257 ) | ( n2248 & n2257 ) ;
  assign n2260 = ( n2244 & ~n2258 ) | ( n2244 & n2259 ) | ( ~n2258 & n2259 ) ;
  assign n2261 = ( n2170 & n2243 ) | ( n2170 & n2260 ) | ( n2243 & n2260 ) ;
  assign n2262 = ( ~n2170 & n2243 ) | ( ~n2170 & n2260 ) | ( n2243 & n2260 ) ;
  assign n2263 = ( n2170 & ~n2261 ) | ( n2170 & n2262 ) | ( ~n2261 & n2262 ) ;
  assign n2264 = ( n2182 & n2234 ) | ( n2182 & n2263 ) | ( n2234 & n2263 ) ;
  assign n2265 = ( ~n2182 & n2234 ) | ( ~n2182 & n2263 ) | ( n2234 & n2263 ) ;
  assign n2266 = ( n2182 & ~n2264 ) | ( n2182 & n2265 ) | ( ~n2264 & n2265 ) ;
  assign n2267 = ( ~n56 & n342 ) | ( ~n56 & n371 ) | ( n342 & n371 ) ;
  assign n2268 = n569 | n2267 ;
  assign n2269 = ( ~n56 & n184 ) | ( ~n56 & n224 ) | ( n184 & n224 ) ;
  assign n2270 = ( n605 & ~n2268 ) | ( n605 & n2269 ) | ( ~n2268 & n2269 ) ;
  assign n2271 = n2268 | n2270 ;
  assign n2272 = ( n769 & n849 ) | ( n769 & ~n1274 ) | ( n849 & ~n1274 ) ;
  assign n2273 = n1274 | n2272 ;
  assign n2274 = n169 | n269 ;
  assign n2275 = n189 | n229 ;
  assign n2276 = ( n345 & ~n469 ) | ( n345 & n2275 ) | ( ~n469 & n2275 ) ;
  assign n2277 = n469 | n2276 ;
  assign n2278 = ( n282 & ~n2274 ) | ( n282 & n2277 ) | ( ~n2274 & n2277 ) ;
  assign n2279 = n2274 | n2278 ;
  assign n2280 = ( ~n2271 & n2273 ) | ( ~n2271 & n2279 ) | ( n2273 & n2279 ) ;
  assign n2281 = n2271 | n2280 ;
  assign n2282 = n2210 & ~n2281 ;
  assign n2283 = ~n2210 & n2281 ;
  assign n2284 = n2282 | n2283 ;
  assign n2285 = ( ~n2212 & n2213 ) | ( ~n2212 & n2284 ) | ( n2213 & n2284 ) ;
  assign n2286 = ( n2132 & n2214 ) | ( n2132 & ~n2284 ) | ( n2214 & ~n2284 ) ;
  assign n2287 = ( ~n2213 & n2285 ) | ( ~n2213 & n2286 ) | ( n2285 & n2286 ) ;
  assign n2288 = n1439 & ~n2287 ;
  assign n2289 = ~n25 & n2132 ;
  assign n2290 = ( n1262 & n2288 ) | ( n1262 & ~n2289 ) | ( n2288 & ~n2289 ) ;
  assign n2291 = ( n1449 & n2282 ) | ( n1449 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2292 = n1450 & n2212 ;
  assign n2293 = ( n1450 & n2291 ) | ( n1450 & ~n2292 ) | ( n2291 & ~n2292 ) ;
  assign n2294 = ( ~n2288 & n2290 ) | ( ~n2288 & n2293 ) | ( n2290 & n2293 ) ;
  assign n2295 = n2290 & ~n2293 ;
  assign n2296 = ( ~n1262 & n2294 ) | ( ~n1262 & n2295 ) | ( n2294 & n2295 ) ;
  assign n2297 = ( n2225 & n2266 ) | ( n2225 & n2296 ) | ( n2266 & n2296 ) ;
  assign n2298 = n1806 & ~n1895 ;
  assign n2299 = n1808 & ~n1892 ;
  assign n2300 = n1763 & n1812 ;
  assign n2301 = n1694 & ~n1917 ;
  assign n2302 = ( n1694 & n2300 ) | ( n1694 & ~n2301 ) | ( n2300 & ~n2301 ) ;
  assign n2303 = ( ~n2298 & n2299 ) | ( ~n2298 & n2302 ) | ( n2299 & n2302 ) ;
  assign n2304 = ( n705 & ~n2298 ) | ( n705 & n2303 ) | ( ~n2298 & n2303 ) ;
  assign n2305 = ( n705 & n2303 ) | ( n705 & ~n2304 ) | ( n2303 & ~n2304 ) ;
  assign n2306 = ( n2298 & n2304 ) | ( n2298 & ~n2305 ) | ( n2304 & ~n2305 ) ;
  assign n2307 = n1616 & n2079 ;
  assign n2308 = n1613 & n2078 ;
  assign n2309 = ~n1431 & n2147 ;
  assign n2310 = ( n1510 & n2082 ) | ( n1510 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2311 = ( ~n2083 & n2309 ) | ( ~n2083 & n2310 ) | ( n2309 & n2310 ) ;
  assign n2312 = ( ~n2307 & n2308 ) | ( ~n2307 & n2311 ) | ( n2308 & n2311 ) ;
  assign n2313 = ( ~n863 & n2307 ) | ( ~n863 & n2312 ) | ( n2307 & n2312 ) ;
  assign n2314 = ( n2307 & n2312 ) | ( n2307 & ~n2313 ) | ( n2312 & ~n2313 ) ;
  assign n2315 = ( n863 & n2313 ) | ( n863 & ~n2314 ) | ( n2313 & ~n2314 ) ;
  assign n2316 = ( n2203 & n2204 ) | ( n2203 & n2247 ) | ( n2204 & n2247 ) ;
  assign n2317 = ( n1434 & n1441 ) | ( n1434 & n2316 ) | ( n1441 & n2316 ) ;
  assign n2318 = ( n943 & n1258 ) | ( n943 & n1259 ) | ( n1258 & n1259 ) ;
  assign n2319 = n2247 & n2318 ;
  assign n2320 = n863 & n939 ;
  assign n2321 = ( n938 & n939 ) | ( n938 & ~n2245 ) | ( n939 & ~n2245 ) ;
  assign n2322 = ( n2246 & ~n2320 ) | ( n2246 & n2321 ) | ( ~n2320 & n2321 ) ;
  assign n2323 = ( n1258 & n1259 ) | ( n1258 & n2322 ) | ( n1259 & n2322 ) ;
  assign n2324 = n2247 & ~n2316 ;
  assign n2325 = n1440 & n2324 ;
  assign n2326 = n2323 | n2325 ;
  assign n2327 = ( ~n2317 & n2319 ) | ( ~n2317 & n2326 ) | ( n2319 & n2326 ) ;
  assign n2328 = ( n2319 & n2326 ) | ( n2319 & ~n2327 ) | ( n2326 & ~n2327 ) ;
  assign n2329 = ( n2317 & n2327 ) | ( n2317 & ~n2328 ) | ( n2327 & ~n2328 ) ;
  assign n2330 = ( n2258 & n2315 ) | ( n2258 & n2329 ) | ( n2315 & n2329 ) ;
  assign n2331 = ( ~n2258 & n2315 ) | ( ~n2258 & n2329 ) | ( n2315 & n2329 ) ;
  assign n2332 = ( n2258 & ~n2330 ) | ( n2258 & n2331 ) | ( ~n2330 & n2331 ) ;
  assign n2333 = ( n2261 & n2306 ) | ( n2261 & n2332 ) | ( n2306 & n2332 ) ;
  assign n2334 = ( ~n2261 & n2306 ) | ( ~n2261 & n2332 ) | ( n2306 & n2332 ) ;
  assign n2335 = ( n2261 & ~n2333 ) | ( n2261 & n2334 ) | ( ~n2333 & n2334 ) ;
  assign n2336 = n1527 & n2135 ;
  assign n2337 = n1629 & n2132 ;
  assign n2338 = n1631 & n1970 ;
  assign n2339 = n1531 & n2044 ;
  assign n2340 = n2338 | n2339 ;
  assign n2341 = ( ~n2336 & n2337 ) | ( ~n2336 & n2340 ) | ( n2337 & n2340 ) ;
  assign n2342 = ( ~n500 & n2336 ) | ( ~n500 & n2341 ) | ( n2336 & n2341 ) ;
  assign n2343 = ( n2336 & n2341 ) | ( n2336 & ~n2342 ) | ( n2341 & ~n2342 ) ;
  assign n2344 = ( n500 & n2342 ) | ( n500 & ~n2343 ) | ( n2342 & ~n2343 ) ;
  assign n2345 = ( n2264 & n2335 ) | ( n2264 & n2344 ) | ( n2335 & n2344 ) ;
  assign n2346 = ( ~n2264 & n2335 ) | ( ~n2264 & n2344 ) | ( n2335 & n2344 ) ;
  assign n2347 = ( n2264 & ~n2345 ) | ( n2264 & n2346 ) | ( ~n2345 & n2346 ) ;
  assign n2348 = n503 | n1239 ;
  assign n2349 = ( ~n56 & n120 ) | ( ~n56 & n237 ) | ( n120 & n237 ) ;
  assign n2350 = n2348 | n2349 ;
  assign n2351 = n338 | n468 ;
  assign n2352 = ( n281 & n422 ) | ( n281 & ~n426 ) | ( n422 & ~n426 ) ;
  assign n2353 = ( ~n2348 & n2351 ) | ( ~n2348 & n2352 ) | ( n2351 & n2352 ) ;
  assign n2354 = ( n83 & n107 ) | ( n83 & n126 ) | ( n107 & n126 ) ;
  assign n2355 = n1864 | n2354 ;
  assign n2356 = ( n247 & n325 ) | ( n247 & ~n586 ) | ( n325 & ~n586 ) ;
  assign n2357 = n586 | n2356 ;
  assign n2358 = ( ~n2349 & n2355 ) | ( ~n2349 & n2357 ) | ( n2355 & n2357 ) ;
  assign n2359 = n2353 | n2358 ;
  assign n2360 = n253 | n310 ;
  assign n2361 = ( n1253 & n1574 ) | ( n1253 & ~n2360 ) | ( n1574 & ~n2360 ) ;
  assign n2362 = n2360 | n2361 ;
  assign n2363 = ( ~n2350 & n2359 ) | ( ~n2350 & n2362 ) | ( n2359 & n2362 ) ;
  assign n2364 = n2350 | n2363 ;
  assign n2365 = ( n236 & n458 ) | ( n236 & ~n765 ) | ( n458 & ~n765 ) ;
  assign n2366 = n765 | n2365 ;
  assign n2367 = ( n78 & n202 ) | ( n78 & n378 ) | ( n202 & n378 ) ;
  assign n2368 = ( n92 & n142 ) | ( n92 & ~n2367 ) | ( n142 & ~n2367 ) ;
  assign n2369 = n2367 | n2368 ;
  assign n2370 = n326 | n449 ;
  assign n2371 = n670 | n2370 ;
  assign n2372 = ( n134 & n163 ) | ( n134 & n202 ) | ( n163 & n202 ) ;
  assign n2373 = ( n514 & ~n2371 ) | ( n514 & n2372 ) | ( ~n2371 & n2372 ) ;
  assign n2374 = n2371 | n2373 ;
  assign n2375 = ( ~n2366 & n2369 ) | ( ~n2366 & n2374 ) | ( n2369 & n2374 ) ;
  assign n2376 = ( n552 & n1581 ) | ( n552 & ~n2366 ) | ( n1581 & ~n2366 ) ;
  assign n2377 = n2366 | n2376 ;
  assign n2378 = ( ~n2364 & n2375 ) | ( ~n2364 & n2377 ) | ( n2375 & n2377 ) ;
  assign n2379 = n2364 | n2378 ;
  assign n2380 = n2282 & ~n2379 ;
  assign n2381 = ~n2282 & n2379 ;
  assign n2382 = n2380 | n2381 ;
  assign n2383 = ( n2284 & n2285 ) | ( n2284 & n2382 ) | ( n2285 & n2382 ) ;
  assign n2384 = ( ~n2212 & n2286 ) | ( ~n2212 & n2382 ) | ( n2286 & n2382 ) ;
  assign n2385 = ( n2284 & ~n2383 ) | ( n2284 & n2384 ) | ( ~n2383 & n2384 ) ;
  assign n2386 = n1439 & n2385 ;
  assign n2387 = ( n1449 & n2380 ) | ( n1449 & n2381 ) | ( n2380 & n2381 ) ;
  assign n2388 = ( n1450 & n2282 ) | ( n1450 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2389 = n1260 & n2212 ;
  assign n2390 = ( n1260 & n2388 ) | ( n1260 & ~n2389 ) | ( n2388 & ~n2389 ) ;
  assign n2391 = ( ~n2386 & n2387 ) | ( ~n2386 & n2390 ) | ( n2387 & n2390 ) ;
  assign n2392 = ( ~n1262 & n2386 ) | ( ~n1262 & n2391 ) | ( n2386 & n2391 ) ;
  assign n2393 = ( n2386 & n2391 ) | ( n2386 & ~n2392 ) | ( n2391 & ~n2392 ) ;
  assign n2394 = ( n1262 & n2392 ) | ( n1262 & ~n2393 ) | ( n2392 & ~n2393 ) ;
  assign n2395 = ( n2297 & n2347 ) | ( n2297 & n2394 ) | ( n2347 & n2394 ) ;
  assign n2396 = n1527 & ~n2215 ;
  assign n2397 = n1629 & ~n2212 ;
  assign n2398 = n1631 & n2044 ;
  assign n2399 = n1531 & n2132 ;
  assign n2400 = n2398 | n2399 ;
  assign n2401 = ( ~n2396 & n2397 ) | ( ~n2396 & n2400 ) | ( n2397 & n2400 ) ;
  assign n2402 = ( ~n500 & n2396 ) | ( ~n500 & n2401 ) | ( n2396 & n2401 ) ;
  assign n2403 = ( n2396 & n2401 ) | ( n2396 & ~n2402 ) | ( n2401 & ~n2402 ) ;
  assign n2404 = ( n500 & n2402 ) | ( n500 & ~n2403 ) | ( n2402 & ~n2403 ) ;
  assign n2405 = n1697 & n2079 ;
  assign n2406 = n1694 & n2078 ;
  assign n2407 = n1510 & n2147 ;
  assign n2408 = ( n1613 & n2082 ) | ( n1613 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2409 = ( ~n2083 & n2407 ) | ( ~n2083 & n2408 ) | ( n2407 & n2408 ) ;
  assign n2410 = ( ~n2405 & n2406 ) | ( ~n2405 & n2409 ) | ( n2406 & n2409 ) ;
  assign n2411 = ( ~n863 & n2405 ) | ( ~n863 & n2410 ) | ( n2405 & n2410 ) ;
  assign n2412 = ( n2405 & n2410 ) | ( n2405 & ~n2411 ) | ( n2410 & ~n2411 ) ;
  assign n2413 = ( n863 & n2411 ) | ( n863 & ~n2412 ) | ( n2411 & ~n2412 ) ;
  assign n2414 = n943 & ~n2248 ;
  assign n2415 = ( ~n2317 & n2326 ) | ( ~n2317 & n2414 ) | ( n2326 & n2414 ) ;
  assign n2416 = ~n2326 & n2415 ;
  assign n2417 = ( n819 & ~n939 ) | ( n819 & n2205 ) | ( ~n939 & n2205 ) ;
  assign n2418 = ( ~n2245 & n2320 ) | ( ~n2245 & n2417 ) | ( n2320 & n2417 ) ;
  assign n2419 = ( n1258 & n1259 ) | ( n1258 & n2418 ) | ( n1259 & n2418 ) ;
  assign n2420 = n1440 & n2322 ;
  assign n2421 = n2419 | n2420 ;
  assign n2422 = ( ~n1431 & n2324 ) | ( ~n1431 & n2421 ) | ( n2324 & n2421 ) ;
  assign n2423 = ( n1513 & ~n1636 ) | ( n1513 & n2316 ) | ( ~n1636 & n2316 ) ;
  assign n2424 = ( n2421 & ~n2422 ) | ( n2421 & n2423 ) | ( ~n2422 & n2423 ) ;
  assign n2425 = n2422 | n2424 ;
  assign n2426 = ( ~n943 & n2416 ) | ( ~n943 & n2425 ) | ( n2416 & n2425 ) ;
  assign n2427 = ( n2416 & n2425 ) | ( n2416 & ~n2426 ) | ( n2425 & ~n2426 ) ;
  assign n2428 = ( n943 & n2426 ) | ( n943 & ~n2427 ) | ( n2426 & ~n2427 ) ;
  assign n2429 = ( n2330 & n2413 ) | ( n2330 & n2428 ) | ( n2413 & n2428 ) ;
  assign n2430 = ( n2330 & ~n2413 ) | ( n2330 & n2428 ) | ( ~n2413 & n2428 ) ;
  assign n2431 = ( n2413 & ~n2429 ) | ( n2413 & n2430 ) | ( ~n2429 & n2430 ) ;
  assign n2432 = n1806 & ~n1973 ;
  assign n2433 = n1808 & n1970 ;
  assign n2434 = n1763 & n1917 ;
  assign n2435 = n1812 & ~n1892 ;
  assign n2436 = n2434 | n2435 ;
  assign n2437 = ( ~n2432 & n2433 ) | ( ~n2432 & n2436 ) | ( n2433 & n2436 ) ;
  assign n2438 = ( n705 & ~n2432 ) | ( n705 & n2437 ) | ( ~n2432 & n2437 ) ;
  assign n2439 = ( n705 & n2437 ) | ( n705 & ~n2438 ) | ( n2437 & ~n2438 ) ;
  assign n2440 = ( n2432 & n2438 ) | ( n2432 & ~n2439 ) | ( n2438 & ~n2439 ) ;
  assign n2441 = ( n2333 & n2431 ) | ( n2333 & n2440 ) | ( n2431 & n2440 ) ;
  assign n2442 = ( ~n2333 & n2431 ) | ( ~n2333 & n2440 ) | ( n2431 & n2440 ) ;
  assign n2443 = ( n2333 & ~n2441 ) | ( n2333 & n2442 ) | ( ~n2441 & n2442 ) ;
  assign n2444 = ( n2345 & n2404 ) | ( n2345 & n2443 ) | ( n2404 & n2443 ) ;
  assign n2445 = ( ~n2345 & n2404 ) | ( ~n2345 & n2443 ) | ( n2404 & n2443 ) ;
  assign n2446 = ( n2345 & ~n2444 ) | ( n2345 & n2445 ) | ( ~n2444 & n2445 ) ;
  assign n2447 = ( n360 & ~n619 ) | ( n360 & n1395 ) | ( ~n619 & n1395 ) ;
  assign n2448 = ~n1395 & n2447 ;
  assign n2449 = ( n57 & n114 ) | ( n57 & n137 ) | ( n114 & n137 ) ;
  assign n2450 = n533 | n2449 ;
  assign n2451 = n742 | n2450 ;
  assign n2452 = n2448 & ~n2451 ;
  assign n2453 = ( ~n179 & n1960 ) | ( ~n179 & n2452 ) | ( n1960 & n2452 ) ;
  assign n2454 = ( ~n916 & n1960 ) | ( ~n916 & n2453 ) | ( n1960 & n2453 ) ;
  assign n2455 = ( n1399 & n1960 ) | ( n1399 & n2454 ) | ( n1960 & n2454 ) ;
  assign n2456 = n2454 & ~n2455 ;
  assign n2457 = n2380 & n2456 ;
  assign n2458 = n2380 | n2456 ;
  assign n2459 = ( n1449 & n2457 ) | ( n1449 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n2460 = n2381 | n2456 ;
  assign n2461 = n2381 & n2456 ;
  assign n2462 = ( n2383 & n2460 ) | ( n2383 & ~n2461 ) | ( n2460 & ~n2461 ) ;
  assign n2463 = ( n2381 & ~n2383 ) | ( n2381 & n2456 ) | ( ~n2383 & n2456 ) ;
  assign n2464 = n2460 & ~n2463 ;
  assign n2465 = ( n1439 & ~n2462 ) | ( n1439 & n2464 ) | ( ~n2462 & n2464 ) ;
  assign n2466 = ( n1260 & n2282 ) | ( n1260 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2467 = ( x0 & x1 ) | ( x0 & ~n2382 ) | ( x1 & ~n2382 ) ;
  assign n2468 = ( x1 & n2466 ) | ( x1 & ~n2467 ) | ( n2466 & ~n2467 ) ;
  assign n2469 = ( ~n2459 & n2465 ) | ( ~n2459 & n2468 ) | ( n2465 & n2468 ) ;
  assign n2470 = ( ~n1262 & n2459 ) | ( ~n1262 & n2469 ) | ( n2459 & n2469 ) ;
  assign n2471 = ( n2459 & n2469 ) | ( n2459 & ~n2470 ) | ( n2469 & ~n2470 ) ;
  assign n2472 = ( n1262 & n2470 ) | ( n1262 & ~n2471 ) | ( n2470 & ~n2471 ) ;
  assign n2473 = ( n2395 & n2446 ) | ( n2395 & n2472 ) | ( n2446 & n2472 ) ;
  assign n2474 = n1527 & ~n2287 ;
  assign n2475 = ( n1629 & n2282 ) | ( n1629 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2476 = n1631 & n2132 ;
  assign n2477 = n1531 & ~n2212 ;
  assign n2478 = n2476 | n2477 ;
  assign n2479 = ( ~n2474 & n2475 ) | ( ~n2474 & n2478 ) | ( n2475 & n2478 ) ;
  assign n2480 = ( ~n500 & n2474 ) | ( ~n500 & n2479 ) | ( n2474 & n2479 ) ;
  assign n2481 = ( n2474 & n2479 ) | ( n2474 & ~n2480 ) | ( n2479 & ~n2480 ) ;
  assign n2482 = ( n500 & n2480 ) | ( n500 & ~n2481 ) | ( n2480 & ~n2481 ) ;
  assign n2483 = n1766 & n2079 ;
  assign n2484 = n1763 & n2078 ;
  assign n2485 = n1613 & n2147 ;
  assign n2486 = ( n1694 & n2082 ) | ( n1694 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2487 = ( ~n2083 & n2485 ) | ( ~n2083 & n2486 ) | ( n2485 & n2486 ) ;
  assign n2488 = ( ~n2483 & n2484 ) | ( ~n2483 & n2487 ) | ( n2484 & n2487 ) ;
  assign n2489 = ( ~n863 & n2483 ) | ( ~n863 & n2488 ) | ( n2483 & n2488 ) ;
  assign n2490 = ( n2483 & n2488 ) | ( n2483 & ~n2489 ) | ( n2488 & ~n2489 ) ;
  assign n2491 = ( n863 & n2489 ) | ( n863 & ~n2490 ) | ( n2489 & ~n2490 ) ;
  assign n2492 = n2416 & ~n2425 ;
  assign n2493 = ~n1517 & n2316 ;
  assign n2494 = n1510 & n2324 ;
  assign n2495 = n1440 & n2418 ;
  assign n2496 = ~n1431 & n2322 ;
  assign n2497 = n2495 | n2496 ;
  assign n2498 = ( ~n2493 & n2494 ) | ( ~n2493 & n2497 ) | ( n2494 & n2497 ) ;
  assign n2499 = ( ~n943 & n2493 ) | ( ~n943 & n2498 ) | ( n2493 & n2498 ) ;
  assign n2500 = ( n2493 & n2498 ) | ( n2493 & ~n2499 ) | ( n2498 & ~n2499 ) ;
  assign n2501 = ( n943 & n2499 ) | ( n943 & ~n2500 ) | ( n2499 & ~n2500 ) ;
  assign n2502 = ( n2318 & n2492 ) | ( n2318 & n2501 ) | ( n2492 & n2501 ) ;
  assign n2503 = ( n2318 & ~n2492 ) | ( n2318 & n2501 ) | ( ~n2492 & n2501 ) ;
  assign n2504 = ( n2492 & ~n2502 ) | ( n2492 & n2503 ) | ( ~n2502 & n2503 ) ;
  assign n2505 = ( n2429 & n2491 ) | ( n2429 & n2504 ) | ( n2491 & n2504 ) ;
  assign n2506 = ( n2429 & ~n2491 ) | ( n2429 & n2504 ) | ( ~n2491 & n2504 ) ;
  assign n2507 = ( n2491 & ~n2505 ) | ( n2491 & n2506 ) | ( ~n2505 & n2506 ) ;
  assign n2508 = n1806 & n2047 ;
  assign n2509 = n1808 & n2044 ;
  assign n2510 = ~n1892 & n1917 ;
  assign n2511 = n1812 & n1970 ;
  assign n2512 = n2510 | n2511 ;
  assign n2513 = ( ~n2508 & n2509 ) | ( ~n2508 & n2512 ) | ( n2509 & n2512 ) ;
  assign n2514 = ( n705 & ~n2508 ) | ( n705 & n2513 ) | ( ~n2508 & n2513 ) ;
  assign n2515 = ( n705 & n2513 ) | ( n705 & ~n2514 ) | ( n2513 & ~n2514 ) ;
  assign n2516 = ( n2508 & n2514 ) | ( n2508 & ~n2515 ) | ( n2514 & ~n2515 ) ;
  assign n2517 = ( n2441 & n2507 ) | ( n2441 & n2516 ) | ( n2507 & n2516 ) ;
  assign n2518 = ( n2441 & ~n2507 ) | ( n2441 & n2516 ) | ( ~n2507 & n2516 ) ;
  assign n2519 = ( n2507 & ~n2517 ) | ( n2507 & n2518 ) | ( ~n2517 & n2518 ) ;
  assign n2520 = ( n2444 & n2482 ) | ( n2444 & n2519 ) | ( n2482 & n2519 ) ;
  assign n2521 = ( n2444 & ~n2482 ) | ( n2444 & n2519 ) | ( ~n2482 & n2519 ) ;
  assign n2522 = ( n2482 & ~n2520 ) | ( n2482 & n2521 ) | ( ~n2520 & n2521 ) ;
  assign n2523 = ~n2457 & n2458 ;
  assign n2524 = ( n2382 & n2383 ) | ( n2382 & ~n2523 ) | ( n2383 & ~n2523 ) ;
  assign n2525 = n373 | n891 ;
  assign n2526 = ( n73 & n98 ) | ( n73 & n202 ) | ( n98 & n202 ) ;
  assign n2527 = n123 | n2526 ;
  assign n2528 = ( ~n140 & n309 ) | ( ~n140 & n2527 ) | ( n309 & n2527 ) ;
  assign n2529 = n140 | n2528 ;
  assign n2530 = ( n889 & ~n2525 ) | ( n889 & n2529 ) | ( ~n2525 & n2529 ) ;
  assign n2531 = n2525 | n2530 ;
  assign n2532 = ( n158 & ~n179 ) | ( n158 & n2531 ) | ( ~n179 & n2531 ) ;
  assign n2533 = ( n179 & n914 ) | ( n179 & ~n2532 ) | ( n914 & ~n2532 ) ;
  assign n2534 = n2532 | n2533 ;
  assign n2535 = ( ~n2458 & n2524 ) | ( ~n2458 & n2534 ) | ( n2524 & n2534 ) ;
  assign n2536 = ( n2524 & n2534 ) | ( n2524 & ~n2535 ) | ( n2534 & ~n2535 ) ;
  assign n2537 = ( n2458 & n2535 ) | ( n2458 & ~n2536 ) | ( n2535 & ~n2536 ) ;
  assign n2538 = n1439 & ~n2537 ;
  assign n2539 = n2457 & ~n2534 ;
  assign n2540 = ~n2457 & n2534 ;
  assign n2541 = ( n1449 & n2539 ) | ( n1449 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2542 = ( n1260 & n2380 ) | ( n1260 & n2381 ) | ( n2380 & n2381 ) ;
  assign n2543 = ( x0 & x1 ) | ( x0 & n2523 ) | ( x1 & n2523 ) ;
  assign n2544 = ( x1 & n2542 ) | ( x1 & ~n2543 ) | ( n2542 & ~n2543 ) ;
  assign n2545 = ( ~n2538 & n2541 ) | ( ~n2538 & n2544 ) | ( n2541 & n2544 ) ;
  assign n2546 = ( ~n1262 & n2538 ) | ( ~n1262 & n2545 ) | ( n2538 & n2545 ) ;
  assign n2547 = ( n2538 & n2545 ) | ( n2538 & ~n2546 ) | ( n2545 & ~n2546 ) ;
  assign n2548 = ( n1262 & n2546 ) | ( n1262 & ~n2547 ) | ( n2546 & ~n2547 ) ;
  assign n2549 = ( n2473 & n2522 ) | ( n2473 & n2548 ) | ( n2522 & n2548 ) ;
  assign n2550 = ( ~n2473 & n2522 ) | ( ~n2473 & n2548 ) | ( n2522 & n2548 ) ;
  assign n2551 = ( n2473 & ~n2549 ) | ( n2473 & n2550 ) | ( ~n2549 & n2550 ) ;
  assign n2552 = n133 | n1284 ;
  assign n2553 = n256 | n341 ;
  assign n2554 = ( n137 & n286 ) | ( n137 & ~n520 ) | ( n286 & ~n520 ) ;
  assign n2555 = n520 | n2554 ;
  assign n2556 = ( n725 & n2352 ) | ( n725 & ~n2555 ) | ( n2352 & ~n2555 ) ;
  assign n2557 = n2555 | n2556 ;
  assign n2558 = ( ~n1284 & n2553 ) | ( ~n1284 & n2557 ) | ( n2553 & n2557 ) ;
  assign n2559 = n599 | n2370 ;
  assign n2560 = n112 | n308 ;
  assign n2561 = ( n87 & n131 ) | ( n87 & n163 ) | ( n131 & n163 ) ;
  assign n2562 = n347 | n796 ;
  assign n2563 = ( n1239 & ~n2561 ) | ( n1239 & n2562 ) | ( ~n2561 & n2562 ) ;
  assign n2564 = n2561 | n2563 ;
  assign n2565 = ( n1880 & ~n2560 ) | ( n1880 & n2564 ) | ( ~n2560 & n2564 ) ;
  assign n2566 = n2560 | n2565 ;
  assign n2567 = ( n588 & ~n2559 ) | ( n588 & n2566 ) | ( ~n2559 & n2566 ) ;
  assign n2568 = n2559 | n2567 ;
  assign n2569 = ( n2552 & n2558 ) | ( n2552 & ~n2568 ) | ( n2558 & ~n2568 ) ;
  assign n2570 = n252 | n284 ;
  assign n2571 = n186 | n364 ;
  assign n2572 = ( ~n324 & n1683 ) | ( ~n324 & n2571 ) | ( n1683 & n2571 ) ;
  assign n2573 = n89 | n2572 ;
  assign n2574 = n270 | n428 ;
  assign n2575 = ( n526 & n1600 ) | ( n526 & ~n2574 ) | ( n1600 & ~n2574 ) ;
  assign n2576 = n2574 | n2575 ;
  assign n2577 = ( n324 & ~n2573 ) | ( n324 & n2576 ) | ( ~n2573 & n2576 ) ;
  assign n2578 = n2573 | n2577 ;
  assign n2579 = ( n585 & ~n2570 ) | ( n585 & n2578 ) | ( ~n2570 & n2578 ) ;
  assign n2580 = n2570 | n2579 ;
  assign n2581 = ( n2568 & ~n2569 ) | ( n2568 & n2580 ) | ( ~n2569 & n2580 ) ;
  assign n2582 = n2569 | n2581 ;
  assign n2583 = ( ~n2395 & n2446 ) | ( ~n2395 & n2472 ) | ( n2446 & n2472 ) ;
  assign n2584 = ( n2395 & ~n2473 ) | ( n2395 & n2583 ) | ( ~n2473 & n2583 ) ;
  assign n2585 = ( n87 & n202 ) | ( n87 & n669 ) | ( n202 & n669 ) ;
  assign n2586 = n623 | n2187 ;
  assign n2587 = n2585 | n2586 ;
  assign n2588 = ( ~n331 & n836 ) | ( ~n331 & n890 ) | ( n836 & n890 ) ;
  assign n2589 = ( n134 & n163 ) | ( n134 & n432 ) | ( n163 & n432 ) ;
  assign n2590 = n2588 | n2589 ;
  assign n2591 = ( n1406 & ~n1740 ) | ( n1406 & n2590 ) | ( ~n1740 & n2590 ) ;
  assign n2592 = n1740 | n2591 ;
  assign n2593 = n2587 | n2592 ;
  assign n2594 = ( n129 & ~n1291 ) | ( n129 & n1417 ) | ( ~n1291 & n1417 ) ;
  assign n2595 = ( n1291 & ~n1685 ) | ( n1291 & n2594 ) | ( ~n1685 & n2594 ) ;
  assign n2596 = n1685 | n2595 ;
  assign n2597 = ( n56 & n224 ) | ( n56 & n250 ) | ( n224 & n250 ) ;
  assign n2598 = ( n294 & n338 ) | ( n294 & ~n2597 ) | ( n338 & ~n2597 ) ;
  assign n2599 = n2597 | n2598 ;
  assign n2600 = ( n1589 & ~n2596 ) | ( n1589 & n2599 ) | ( ~n2596 & n2599 ) ;
  assign n2601 = ( ~n107 & n203 ) | ( ~n107 & n326 ) | ( n203 & n326 ) ;
  assign n2602 = n342 | n2601 ;
  assign n2603 = ( n2596 & ~n2600 ) | ( n2596 & n2602 ) | ( ~n2600 & n2602 ) ;
  assign n2604 = ( ~n2593 & n2600 ) | ( ~n2593 & n2603 ) | ( n2600 & n2603 ) ;
  assign n2605 = ( n2584 & n2593 ) | ( n2584 & n2604 ) | ( n2593 & n2604 ) ;
  assign n2606 = ( n2551 & n2582 ) | ( n2551 & n2605 ) | ( n2582 & n2605 ) ;
  assign n2607 = n1527 & n2385 ;
  assign n2608 = ( n1629 & n2380 ) | ( n1629 & n2381 ) | ( n2380 & n2381 ) ;
  assign n2609 = ( n1531 & n2282 ) | ( n1531 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2610 = n1631 & n2212 ;
  assign n2611 = ( n1631 & n2609 ) | ( n1631 & ~n2610 ) | ( n2609 & ~n2610 ) ;
  assign n2612 = ( ~n2607 & n2608 ) | ( ~n2607 & n2611 ) | ( n2608 & n2611 ) ;
  assign n2613 = ( ~n500 & n2607 ) | ( ~n500 & n2612 ) | ( n2607 & n2612 ) ;
  assign n2614 = ( n2607 & n2612 ) | ( n2607 & ~n2613 ) | ( n2612 & ~n2613 ) ;
  assign n2615 = ( n500 & n2613 ) | ( n500 & ~n2614 ) | ( n2613 & ~n2614 ) ;
  assign n2616 = n1806 & n2135 ;
  assign n2617 = n1808 & n2132 ;
  assign n2618 = n1917 & n1970 ;
  assign n2619 = n1812 & n2044 ;
  assign n2620 = n2618 | n2619 ;
  assign n2621 = ( ~n2616 & n2617 ) | ( ~n2616 & n2620 ) | ( n2617 & n2620 ) ;
  assign n2622 = ( n705 & ~n2616 ) | ( n705 & n2621 ) | ( ~n2616 & n2621 ) ;
  assign n2623 = ( n705 & n2621 ) | ( n705 & ~n2622 ) | ( n2621 & ~n2622 ) ;
  assign n2624 = ( n2616 & n2622 ) | ( n2616 & ~n2623 ) | ( n2622 & ~n2623 ) ;
  assign n2625 = ~n1895 & n2079 ;
  assign n2626 = ~n1892 & n2078 ;
  assign n2627 = n1694 & n2147 ;
  assign n2628 = ( n1763 & n2082 ) | ( n1763 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2629 = ( ~n2083 & n2627 ) | ( ~n2083 & n2628 ) | ( n2627 & n2628 ) ;
  assign n2630 = ( ~n2625 & n2626 ) | ( ~n2625 & n2629 ) | ( n2626 & n2629 ) ;
  assign n2631 = ( ~n863 & n2625 ) | ( ~n863 & n2630 ) | ( n2625 & n2630 ) ;
  assign n2632 = ( n2625 & n2630 ) | ( n2625 & ~n2631 ) | ( n2630 & ~n2631 ) ;
  assign n2633 = ( n863 & n2631 ) | ( n863 & ~n2632 ) | ( n2631 & ~n2632 ) ;
  assign n2634 = n943 & ~n1440 ;
  assign n2635 = ~n1431 & n2418 ;
  assign n2636 = n1510 & n2322 ;
  assign n2637 = n2635 | n2636 ;
  assign n2638 = n1613 & ~n2324 ;
  assign n2639 = ( n1613 & n2637 ) | ( n1613 & ~n2638 ) | ( n2637 & ~n2638 ) ;
  assign n2640 = n1616 & n2316 ;
  assign n2641 = n2639 | n2640 ;
  assign n2642 = ( ~n2502 & n2634 ) | ( ~n2502 & n2641 ) | ( n2634 & n2641 ) ;
  assign n2643 = ( n2634 & n2641 ) | ( n2634 & ~n2642 ) | ( n2641 & ~n2642 ) ;
  assign n2644 = ( n2502 & n2642 ) | ( n2502 & ~n2643 ) | ( n2642 & ~n2643 ) ;
  assign n2645 = ( n2505 & n2633 ) | ( n2505 & n2644 ) | ( n2633 & n2644 ) ;
  assign n2646 = ( n2505 & ~n2633 ) | ( n2505 & n2644 ) | ( ~n2633 & n2644 ) ;
  assign n2647 = ( n2633 & ~n2645 ) | ( n2633 & n2646 ) | ( ~n2645 & n2646 ) ;
  assign n2648 = ( n2517 & n2624 ) | ( n2517 & n2647 ) | ( n2624 & n2647 ) ;
  assign n2649 = ( n2517 & ~n2624 ) | ( n2517 & n2647 ) | ( ~n2624 & n2647 ) ;
  assign n2650 = ( n2624 & ~n2648 ) | ( n2624 & n2649 ) | ( ~n2648 & n2649 ) ;
  assign n2651 = ( n2520 & n2615 ) | ( n2520 & n2650 ) | ( n2615 & n2650 ) ;
  assign n2652 = ( n2520 & ~n2615 ) | ( n2520 & n2650 ) | ( ~n2615 & n2650 ) ;
  assign n2653 = ( n2615 & ~n2651 ) | ( n2615 & n2652 ) | ( ~n2651 & n2652 ) ;
  assign n2654 = ( ~n2523 & n2524 ) | ( ~n2523 & n2534 ) | ( n2524 & n2534 ) ;
  assign n2655 = n109 | n224 ;
  assign n2656 = n121 | n159 ;
  assign n2657 = n2655 | n2656 ;
  assign n2658 = n97 | n179 ;
  assign n2659 = n907 | n2658 ;
  assign n2660 = ( n899 & ~n2657 ) | ( n899 & n2659 ) | ( ~n2657 & n2659 ) ;
  assign n2661 = n2657 | n2660 ;
  assign n2662 = ( ~n2540 & n2654 ) | ( ~n2540 & n2661 ) | ( n2654 & n2661 ) ;
  assign n2663 = n2539 | n2540 ;
  assign n2664 = ( n2654 & n2661 ) | ( n2654 & n2663 ) | ( n2661 & n2663 ) ;
  assign n2665 = ( n2540 & n2662 ) | ( n2540 & ~n2664 ) | ( n2662 & ~n2664 ) ;
  assign n2666 = n1439 & n2665 ;
  assign n2667 = ~n2539 & n2661 ;
  assign n2668 = n1449 & n2667 ;
  assign n2669 = ( n1260 & n2457 ) | ( n1260 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n2670 = ( x0 & x1 ) | ( x0 & ~n2663 ) | ( x1 & ~n2663 ) ;
  assign n2671 = ( x1 & n2669 ) | ( x1 & ~n2670 ) | ( n2669 & ~n2670 ) ;
  assign n2672 = ( ~n2666 & n2668 ) | ( ~n2666 & n2671 ) | ( n2668 & n2671 ) ;
  assign n2673 = ( ~n1262 & n2666 ) | ( ~n1262 & n2672 ) | ( n2666 & n2672 ) ;
  assign n2674 = ( n2666 & n2672 ) | ( n2666 & ~n2673 ) | ( n2672 & ~n2673 ) ;
  assign n2675 = ( n1262 & n2673 ) | ( n1262 & ~n2674 ) | ( n2673 & ~n2674 ) ;
  assign n2676 = ( n2549 & n2653 ) | ( n2549 & n2675 ) | ( n2653 & n2675 ) ;
  assign n2677 = ( n2549 & ~n2653 ) | ( n2549 & n2675 ) | ( ~n2653 & n2675 ) ;
  assign n2678 = ( n2653 & ~n2676 ) | ( n2653 & n2677 ) | ( ~n2676 & n2677 ) ;
  assign n2679 = ( n234 & n363 ) | ( n234 & ~n820 ) | ( n363 & ~n820 ) ;
  assign n2680 = n820 | n2679 ;
  assign n2681 = n644 | n2362 ;
  assign n2682 = n2680 | n2681 ;
  assign n2683 = n709 | n2348 ;
  assign n2684 = n220 | n610 ;
  assign n2685 = ( n2190 & ~n2683 ) | ( n2190 & n2684 ) | ( ~n2683 & n2684 ) ;
  assign n2686 = n143 | n154 ;
  assign n2687 = ( n314 & n2366 ) | ( n314 & ~n2686 ) | ( n2366 & ~n2686 ) ;
  assign n2688 = n2686 | n2687 ;
  assign n2689 = ( n2683 & n2685 ) | ( n2683 & ~n2688 ) | ( n2685 & ~n2688 ) ;
  assign n2690 = ( n679 & n2688 ) | ( n679 & ~n2689 ) | ( n2688 & ~n2689 ) ;
  assign n2691 = n2689 | n2690 ;
  assign n2692 = n246 | n786 ;
  assign n2693 = n116 | n120 ;
  assign n2694 = ( n56 & n189 ) | ( n56 & n283 ) | ( n189 & n283 ) ;
  assign n2695 = ( n109 & ~n378 ) | ( n109 & n2694 ) | ( ~n378 & n2694 ) ;
  assign n2696 = ( ~n569 & n1494 ) | ( ~n569 & n2695 ) | ( n1494 & n2695 ) ;
  assign n2697 = n569 | n2696 ;
  assign n2698 = ( n294 & n364 ) | ( n294 & ~n647 ) | ( n364 & ~n647 ) ;
  assign n2699 = n647 | n2698 ;
  assign n2700 = ( n105 & n126 ) | ( n105 & n163 ) | ( n126 & n163 ) ;
  assign n2701 = ( n1860 & ~n2699 ) | ( n1860 & n2700 ) | ( ~n2699 & n2700 ) ;
  assign n2702 = n2699 | n2701 ;
  assign n2703 = ( n78 & n202 ) | ( n78 & n227 ) | ( n202 & n227 ) ;
  assign n2704 = n386 | n439 ;
  assign n2705 = n2703 | n2704 ;
  assign n2706 = ( ~n2697 & n2702 ) | ( ~n2697 & n2705 ) | ( n2702 & n2705 ) ;
  assign n2707 = n2697 | n2706 ;
  assign n2708 = ( ~n2692 & n2693 ) | ( ~n2692 & n2707 ) | ( n2693 & n2707 ) ;
  assign n2709 = n2692 | n2708 ;
  assign n2710 = ( ~n2682 & n2691 ) | ( ~n2682 & n2709 ) | ( n2691 & n2709 ) ;
  assign n2711 = n2682 | n2710 ;
  assign n2712 = ( ~n2606 & n2678 ) | ( ~n2606 & n2711 ) | ( n2678 & n2711 ) ;
  assign n2713 = ( n2606 & n2678 ) | ( n2606 & n2711 ) | ( n2678 & n2711 ) ;
  assign n2714 = ( n2606 & n2712 ) | ( n2606 & ~n2713 ) | ( n2712 & ~n2713 ) ;
  assign n2715 = n273 | n842 ;
  assign n2716 = ( n150 & ~n428 ) | ( n150 & n440 ) | ( ~n428 & n440 ) ;
  assign n2717 = n428 | n2716 ;
  assign n2718 = n588 | n2700 ;
  assign n2719 = ( n781 & ~n2717 ) | ( n781 & n2718 ) | ( ~n2717 & n2718 ) ;
  assign n2720 = n2717 | n2719 ;
  assign n2721 = ( n2366 & ~n2715 ) | ( n2366 & n2720 ) | ( ~n2715 & n2720 ) ;
  assign n2722 = n2715 | n2721 ;
  assign n2723 = ( n580 & n1757 ) | ( n580 & ~n2722 ) | ( n1757 & ~n2722 ) ;
  assign n2724 = n2722 | n2723 ;
  assign n2725 = n1806 & ~n2215 ;
  assign n2726 = n1808 & ~n2212 ;
  assign n2727 = n1917 & n2044 ;
  assign n2728 = n1812 & n2132 ;
  assign n2729 = n2727 | n2728 ;
  assign n2730 = ( ~n2725 & n2726 ) | ( ~n2725 & n2729 ) | ( n2726 & n2729 ) ;
  assign n2731 = ( n705 & ~n2725 ) | ( n705 & n2730 ) | ( ~n2725 & n2730 ) ;
  assign n2732 = ( n705 & n2730 ) | ( n705 & ~n2731 ) | ( n2730 & ~n2731 ) ;
  assign n2733 = ( n2725 & n2731 ) | ( n2725 & ~n2732 ) | ( n2731 & ~n2732 ) ;
  assign n2734 = n1510 & n2418 ;
  assign n2735 = n1613 & n2322 ;
  assign n2736 = n2734 | n2735 ;
  assign n2737 = n1694 & ~n2324 ;
  assign n2738 = ( n1694 & n2736 ) | ( n1694 & ~n2737 ) | ( n2736 & ~n2737 ) ;
  assign n2739 = n1697 & n2316 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n943 & n1431 ;
  assign n2742 = ~n943 & n2641 ;
  assign n2743 = ( n943 & ~n2642 ) | ( n943 & n2742 ) | ( ~n2642 & n2742 ) ;
  assign n2744 = ( n2740 & n2741 ) | ( n2740 & ~n2743 ) | ( n2741 & ~n2743 ) ;
  assign n2745 = ( n2740 & ~n2741 ) | ( n2740 & n2743 ) | ( ~n2741 & n2743 ) ;
  assign n2746 = ( ~n2740 & n2744 ) | ( ~n2740 & n2745 ) | ( n2744 & n2745 ) ;
  assign n2747 = ~n1973 & n2079 ;
  assign n2748 = n1970 & n2078 ;
  assign n2749 = n1763 & n2147 ;
  assign n2750 = ( ~n1892 & n2082 ) | ( ~n1892 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2751 = ( ~n2083 & n2749 ) | ( ~n2083 & n2750 ) | ( n2749 & n2750 ) ;
  assign n2752 = ( ~n2747 & n2748 ) | ( ~n2747 & n2751 ) | ( n2748 & n2751 ) ;
  assign n2753 = ( ~n863 & n2747 ) | ( ~n863 & n2752 ) | ( n2747 & n2752 ) ;
  assign n2754 = ( n2747 & n2752 ) | ( n2747 & ~n2753 ) | ( n2752 & ~n2753 ) ;
  assign n2755 = ( n863 & n2753 ) | ( n863 & ~n2754 ) | ( n2753 & ~n2754 ) ;
  assign n2756 = ( n2645 & n2746 ) | ( n2645 & n2755 ) | ( n2746 & n2755 ) ;
  assign n2757 = ( n2645 & ~n2746 ) | ( n2645 & n2755 ) | ( ~n2746 & n2755 ) ;
  assign n2758 = ( n2746 & ~n2756 ) | ( n2746 & n2757 ) | ( ~n2756 & n2757 ) ;
  assign n2759 = ( n2648 & n2733 ) | ( n2648 & n2758 ) | ( n2733 & n2758 ) ;
  assign n2760 = ( n2648 & ~n2733 ) | ( n2648 & n2758 ) | ( ~n2733 & n2758 ) ;
  assign n2761 = ( n2733 & ~n2759 ) | ( n2733 & n2760 ) | ( ~n2759 & n2760 ) ;
  assign n2762 = ( n1629 & n2457 ) | ( n1629 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n2763 = ( n1631 & n2282 ) | ( n1631 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2764 = ( n1531 & n2380 ) | ( n1531 & n2381 ) | ( n2380 & n2381 ) ;
  assign n2765 = n2763 | n2764 ;
  assign n2766 = ( n1527 & ~n2462 ) | ( n1527 & n2464 ) | ( ~n2462 & n2464 ) ;
  assign n2767 = ( ~n2762 & n2765 ) | ( ~n2762 & n2766 ) | ( n2765 & n2766 ) ;
  assign n2768 = ( ~n500 & n2762 ) | ( ~n500 & n2767 ) | ( n2762 & n2767 ) ;
  assign n2769 = ( n2762 & n2767 ) | ( n2762 & ~n2768 ) | ( n2767 & ~n2768 ) ;
  assign n2770 = ( n500 & n2768 ) | ( n500 & ~n2769 ) | ( n2768 & ~n2769 ) ;
  assign n2771 = ( n2651 & n2761 ) | ( n2651 & n2770 ) | ( n2761 & n2770 ) ;
  assign n2772 = ( n2651 & ~n2761 ) | ( n2651 & n2770 ) | ( ~n2761 & n2770 ) ;
  assign n2773 = ( n2761 & ~n2771 ) | ( n2761 & n2772 ) | ( ~n2771 & n2772 ) ;
  assign n2774 = n654 | n1243 ;
  assign n2775 = n220 | n266 ;
  assign n2776 = n442 | n458 ;
  assign n2777 = n2775 | n2776 ;
  assign n2778 = ( n2700 & ~n2774 ) | ( n2700 & n2777 ) | ( ~n2774 & n2777 ) ;
  assign n2779 = n2774 | n2778 ;
  assign n2780 = n1395 | n2275 ;
  assign n2781 = ( n78 & n91 ) | ( n78 & n163 ) | ( n91 & n163 ) ;
  assign n2782 = n420 | n2781 ;
  assign n2783 = n187 | n203 ;
  assign n2784 = ( n439 & n650 ) | ( n439 & ~n2783 ) | ( n650 & ~n2783 ) ;
  assign n2785 = n2783 | n2784 ;
  assign n2786 = ( ~n2780 & n2782 ) | ( ~n2780 & n2785 ) | ( n2782 & n2785 ) ;
  assign n2787 = n2780 | n2786 ;
  assign n2788 = ( n368 & n2197 ) | ( n368 & n2787 ) | ( n2197 & n2787 ) ;
  assign n2789 = ( n368 & n2779 ) | ( n368 & ~n2788 ) | ( n2779 & ~n2788 ) ;
  assign n2790 = ~n2779 & n2789 ;
  assign n2791 = ( n2664 & ~n2667 ) | ( n2664 & n2790 ) | ( ~n2667 & n2790 ) ;
  assign n2792 = ( n2664 & n2790 ) | ( n2664 & ~n2791 ) | ( n2790 & ~n2791 ) ;
  assign n2793 = ( n2667 & n2791 ) | ( n2667 & ~n2792 ) | ( n2791 & ~n2792 ) ;
  assign n2794 = n1439 & ~n2793 ;
  assign n2795 = n1449 & ~n2790 ;
  assign n2796 = ( n1260 & n2539 ) | ( n1260 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2797 = n1450 & n2667 ;
  assign n2798 = n2796 | n2797 ;
  assign n2799 = ( ~n2794 & n2795 ) | ( ~n2794 & n2798 ) | ( n2795 & n2798 ) ;
  assign n2800 = ( ~n1262 & n2794 ) | ( ~n1262 & n2799 ) | ( n2794 & n2799 ) ;
  assign n2801 = ( n2794 & n2799 ) | ( n2794 & ~n2800 ) | ( n2799 & ~n2800 ) ;
  assign n2802 = ( n1262 & n2800 ) | ( n1262 & ~n2801 ) | ( n2800 & ~n2801 ) ;
  assign n2803 = ( n2676 & n2773 ) | ( n2676 & n2802 ) | ( n2773 & n2802 ) ;
  assign n2804 = ( n2676 & ~n2773 ) | ( n2676 & n2802 ) | ( ~n2773 & n2802 ) ;
  assign n2805 = ( n2773 & ~n2803 ) | ( n2773 & n2804 ) | ( ~n2803 & n2804 ) ;
  assign n2806 = ( n2713 & n2724 ) | ( n2713 & n2805 ) | ( n2724 & n2805 ) ;
  assign n2807 = ( ~n2713 & n2724 ) | ( ~n2713 & n2805 ) | ( n2724 & n2805 ) ;
  assign n2808 = ( n2713 & ~n2806 ) | ( n2713 & n2807 ) | ( ~n2806 & n2807 ) ;
  assign n2809 = n2714 & n2808 ;
  assign n2810 = n2808 & ~n2809 ;
  assign n2811 = ( n2714 & ~n2809 ) | ( n2714 & n2810 ) | ( ~n2809 & n2810 ) ;
  assign n2812 = x22 | x23 ;
  assign n2813 = ( x22 & x23 ) | ( x22 & ~n2812 ) | ( x23 & ~n2812 ) ;
  assign n2814 = n2812 & ~n2813 ;
  assign n2815 = ( n2664 & n2667 ) | ( n2664 & ~n2790 ) | ( n2667 & ~n2790 ) ;
  assign n2816 = n838 & ~n1410 ;
  assign n2817 = n230 | n325 ;
  assign n2818 = ( n281 & ~n337 ) | ( n281 & n341 ) | ( ~n337 & n341 ) ;
  assign n2819 = ( n226 & ~n230 ) | ( n226 & n2818 ) | ( ~n230 & n2818 ) ;
  assign n2820 = n455 | n742 ;
  assign n2821 = ( ~n230 & n624 ) | ( ~n230 & n2820 ) | ( n624 & n2820 ) ;
  assign n2822 = ( ~n2817 & n2819 ) | ( ~n2817 & n2821 ) | ( n2819 & n2821 ) ;
  assign n2823 = n2817 | n2822 ;
  assign n2824 = n639 | n1417 ;
  assign n2825 = n154 | n234 ;
  assign n2826 = ( n118 & n539 ) | ( n118 & ~n2825 ) | ( n539 & ~n2825 ) ;
  assign n2827 = n2825 | n2826 ;
  assign n2828 = ( n1860 & ~n2824 ) | ( n1860 & n2827 ) | ( ~n2824 & n2827 ) ;
  assign n2829 = n2824 | n2828 ;
  assign n2830 = ( n2816 & n2823 ) | ( n2816 & n2829 ) | ( n2823 & n2829 ) ;
  assign n2831 = n2816 & ~n2830 ;
  assign n2832 = ( n2790 & n2815 ) | ( n2790 & n2831 ) | ( n2815 & n2831 ) ;
  assign n2833 = ( ~n2790 & n2815 ) | ( ~n2790 & n2831 ) | ( n2815 & n2831 ) ;
  assign n2834 = ( n2790 & ~n2832 ) | ( n2790 & n2833 ) | ( ~n2832 & n2833 ) ;
  assign n2835 = n1439 & n2834 ;
  assign n2836 = n1449 & ~n2831 ;
  assign n2837 = n1260 & n2667 ;
  assign n2838 = n1450 & ~n2790 ;
  assign n2839 = n2837 | n2838 ;
  assign n2840 = ( ~n2835 & n2836 ) | ( ~n2835 & n2839 ) | ( n2836 & n2839 ) ;
  assign n2841 = ( ~n1262 & n2835 ) | ( ~n1262 & n2840 ) | ( n2835 & n2840 ) ;
  assign n2842 = ( n2835 & n2840 ) | ( n2835 & ~n2841 ) | ( n2840 & ~n2841 ) ;
  assign n2843 = ( n1262 & n2841 ) | ( n1262 & ~n2842 ) | ( n2841 & ~n2842 ) ;
  assign n2844 = n1806 & ~n2287 ;
  assign n2845 = ( n1808 & n2282 ) | ( n1808 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2846 = n1917 & n2132 ;
  assign n2847 = n1812 & ~n2212 ;
  assign n2848 = n2846 | n2847 ;
  assign n2849 = ( ~n2844 & n2845 ) | ( ~n2844 & n2848 ) | ( n2845 & n2848 ) ;
  assign n2850 = ( n705 & ~n2844 ) | ( n705 & n2849 ) | ( ~n2844 & n2849 ) ;
  assign n2851 = ( n705 & n2849 ) | ( n705 & ~n2850 ) | ( n2849 & ~n2850 ) ;
  assign n2852 = ( n2844 & n2850 ) | ( n2844 & ~n2851 ) | ( n2850 & ~n2851 ) ;
  assign n2853 = n2047 & n2079 ;
  assign n2854 = n2044 & n2078 ;
  assign n2855 = ~n1892 & n2147 ;
  assign n2856 = ( n1970 & n2082 ) | ( n1970 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2857 = ( ~n2083 & n2855 ) | ( ~n2083 & n2856 ) | ( n2855 & n2856 ) ;
  assign n2858 = ( ~n2853 & n2854 ) | ( ~n2853 & n2857 ) | ( n2854 & n2857 ) ;
  assign n2859 = ( ~n863 & n2853 ) | ( ~n863 & n2858 ) | ( n2853 & n2858 ) ;
  assign n2860 = ( n2853 & n2858 ) | ( n2853 & ~n2859 ) | ( n2858 & ~n2859 ) ;
  assign n2861 = ( n863 & n2859 ) | ( n863 & ~n2860 ) | ( n2859 & ~n2860 ) ;
  assign n2862 = n1613 & n2418 ;
  assign n2863 = n1694 & n2322 ;
  assign n2864 = n2862 | n2863 ;
  assign n2865 = n1763 & ~n2324 ;
  assign n2866 = ( n1763 & n2864 ) | ( n1763 & ~n2865 ) | ( n2864 & ~n2865 ) ;
  assign n2867 = n1766 & n2316 ;
  assign n2868 = n2866 | n2867 ;
  assign n2869 = n943 & ~n1510 ;
  assign n2870 = n943 | n2740 ;
  assign n2871 = ~n2744 & n2870 ;
  assign n2872 = ( ~n2868 & n2869 ) | ( ~n2868 & n2871 ) | ( n2869 & n2871 ) ;
  assign n2873 = ( n2868 & n2869 ) | ( n2868 & n2871 ) | ( n2869 & n2871 ) ;
  assign n2874 = ( n2868 & n2872 ) | ( n2868 & ~n2873 ) | ( n2872 & ~n2873 ) ;
  assign n2875 = ( n2756 & n2861 ) | ( n2756 & n2874 ) | ( n2861 & n2874 ) ;
  assign n2876 = ( n2756 & ~n2861 ) | ( n2756 & n2874 ) | ( ~n2861 & n2874 ) ;
  assign n2877 = ( n2861 & ~n2875 ) | ( n2861 & n2876 ) | ( ~n2875 & n2876 ) ;
  assign n2878 = ( n2759 & n2852 ) | ( n2759 & n2877 ) | ( n2852 & n2877 ) ;
  assign n2879 = ( n2759 & ~n2852 ) | ( n2759 & n2877 ) | ( ~n2852 & n2877 ) ;
  assign n2880 = ( n2852 & ~n2878 ) | ( n2852 & n2879 ) | ( ~n2878 & n2879 ) ;
  assign n2881 = n1527 & ~n2537 ;
  assign n2882 = ( n1629 & n2539 ) | ( n1629 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2883 = ( n1631 & n2380 ) | ( n1631 & n2381 ) | ( n2380 & n2381 ) ;
  assign n2884 = ( n1531 & n2457 ) | ( n1531 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n2885 = n2883 | n2884 ;
  assign n2886 = ( ~n2881 & n2882 ) | ( ~n2881 & n2885 ) | ( n2882 & n2885 ) ;
  assign n2887 = ( ~n500 & n2881 ) | ( ~n500 & n2886 ) | ( n2881 & n2886 ) ;
  assign n2888 = ( n2881 & n2886 ) | ( n2881 & ~n2887 ) | ( n2886 & ~n2887 ) ;
  assign n2889 = ( n500 & n2887 ) | ( n500 & ~n2888 ) | ( n2887 & ~n2888 ) ;
  assign n2890 = ( n2771 & n2880 ) | ( n2771 & n2889 ) | ( n2880 & n2889 ) ;
  assign n2891 = ( n2771 & ~n2880 ) | ( n2771 & n2889 ) | ( ~n2880 & n2889 ) ;
  assign n2892 = ( n2880 & ~n2890 ) | ( n2880 & n2891 ) | ( ~n2890 & n2891 ) ;
  assign n2893 = ( n2803 & n2843 ) | ( n2803 & n2892 ) | ( n2843 & n2892 ) ;
  assign n2894 = ( n2803 & ~n2843 ) | ( n2803 & n2892 ) | ( ~n2843 & n2892 ) ;
  assign n2895 = ( n2843 & ~n2893 ) | ( n2843 & n2894 ) | ( ~n2893 & n2894 ) ;
  assign n2896 = n340 | n1684 ;
  assign n2897 = n186 | n253 ;
  assign n2898 = ( n539 & ~n1684 ) | ( n539 & n2897 ) | ( ~n1684 & n2897 ) ;
  assign n2899 = ( ~n2357 & n2896 ) | ( ~n2357 & n2898 ) | ( n2896 & n2898 ) ;
  assign n2900 = ( n111 & n136 ) | ( n111 & n202 ) | ( n136 & n202 ) ;
  assign n2901 = ( n154 & n265 ) | ( n154 & ~n2900 ) | ( n265 & ~n2900 ) ;
  assign n2902 = n2900 | n2901 ;
  assign n2903 = n209 | n825 ;
  assign n2904 = ( n2366 & ~n2902 ) | ( n2366 & n2903 ) | ( ~n2902 & n2903 ) ;
  assign n2905 = ( ~n2357 & n2902 ) | ( ~n2357 & n2904 ) | ( n2902 & n2904 ) ;
  assign n2906 = ( n2357 & ~n2899 ) | ( n2357 & n2905 ) | ( ~n2899 & n2905 ) ;
  assign n2907 = n2899 | n2906 ;
  assign n2908 = ( n1886 & n2707 ) | ( n1886 & ~n2907 ) | ( n2707 & ~n2907 ) ;
  assign n2909 = n2907 | n2908 ;
  assign n2910 = ( n2806 & n2895 ) | ( n2806 & n2909 ) | ( n2895 & n2909 ) ;
  assign n2911 = ( n2806 & ~n2895 ) | ( n2806 & n2909 ) | ( ~n2895 & n2909 ) ;
  assign n2912 = ( n2895 & ~n2910 ) | ( n2895 & n2911 ) | ( ~n2910 & n2911 ) ;
  assign n2913 = ( n2809 & n2811 ) | ( n2809 & ~n2912 ) | ( n2811 & ~n2912 ) ;
  assign n2914 = n2809 & n2912 ;
  assign n2915 = ( n2912 & n2913 ) | ( n2912 & ~n2914 ) | ( n2913 & ~n2914 ) ;
  assign n2916 = ( ~n2814 & n2913 ) | ( ~n2814 & n2915 ) | ( n2913 & n2915 ) ;
  assign n2917 = n2814 & n2915 ;
  assign n2918 = ( n2912 & n2915 ) | ( n2912 & n2917 ) | ( n2915 & n2917 ) ;
  assign n2919 = ( ~n2811 & n2916 ) | ( ~n2811 & n2918 ) | ( n2916 & n2918 ) ;
  assign n2920 = n1806 & n2385 ;
  assign n2921 = ( n1808 & n2380 ) | ( n1808 & n2381 ) | ( n2380 & n2381 ) ;
  assign n2922 = ( n1812 & n2282 ) | ( n1812 & n2283 ) | ( n2282 & n2283 ) ;
  assign n2923 = n1917 & n2212 ;
  assign n2924 = ( n1917 & n2922 ) | ( n1917 & ~n2923 ) | ( n2922 & ~n2923 ) ;
  assign n2925 = ( ~n2920 & n2921 ) | ( ~n2920 & n2924 ) | ( n2921 & n2924 ) ;
  assign n2926 = ( n705 & ~n2920 ) | ( n705 & n2925 ) | ( ~n2920 & n2925 ) ;
  assign n2927 = ( n705 & n2925 ) | ( n705 & ~n2926 ) | ( n2925 & ~n2926 ) ;
  assign n2928 = ( n2920 & n2926 ) | ( n2920 & ~n2927 ) | ( n2926 & ~n2927 ) ;
  assign n2929 = n2079 & n2135 ;
  assign n2930 = n2078 & n2132 ;
  assign n2931 = n1970 & n2147 ;
  assign n2932 = ( n2044 & n2082 ) | ( n2044 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2933 = ( ~n2083 & n2931 ) | ( ~n2083 & n2932 ) | ( n2931 & n2932 ) ;
  assign n2934 = ( ~n2929 & n2930 ) | ( ~n2929 & n2933 ) | ( n2930 & n2933 ) ;
  assign n2935 = ( ~n863 & n2929 ) | ( ~n863 & n2934 ) | ( n2929 & n2934 ) ;
  assign n2936 = ( n2929 & n2934 ) | ( n2929 & ~n2935 ) | ( n2934 & ~n2935 ) ;
  assign n2937 = ( n863 & n2935 ) | ( n863 & ~n2936 ) | ( n2935 & ~n2936 ) ;
  assign n2938 = n1694 & n2418 ;
  assign n2939 = n1763 & n2322 ;
  assign n2940 = n2938 | n2939 ;
  assign n2941 = n1892 | n2324 ;
  assign n2942 = ( ~n1892 & n2940 ) | ( ~n1892 & n2941 ) | ( n2940 & n2941 ) ;
  assign n2943 = ~n1895 & n2316 ;
  assign n2944 = n2942 | n2943 ;
  assign n2945 = n943 & ~n1613 ;
  assign n2946 = n943 & ~n2868 ;
  assign n2947 = ( ~n2869 & n2873 ) | ( ~n2869 & n2946 ) | ( n2873 & n2946 ) ;
  assign n2948 = ( n2944 & n2945 ) | ( n2944 & ~n2947 ) | ( n2945 & ~n2947 ) ;
  assign n2949 = ( n2944 & ~n2945 ) | ( n2944 & n2947 ) | ( ~n2945 & n2947 ) ;
  assign n2950 = ( ~n2944 & n2948 ) | ( ~n2944 & n2949 ) | ( n2948 & n2949 ) ;
  assign n2951 = ( n2875 & n2937 ) | ( n2875 & n2950 ) | ( n2937 & n2950 ) ;
  assign n2952 = ( n2875 & ~n2937 ) | ( n2875 & n2950 ) | ( ~n2937 & n2950 ) ;
  assign n2953 = ( n2937 & ~n2951 ) | ( n2937 & n2952 ) | ( ~n2951 & n2952 ) ;
  assign n2954 = ( n2878 & n2928 ) | ( n2878 & n2953 ) | ( n2928 & n2953 ) ;
  assign n2955 = ( n2878 & ~n2928 ) | ( n2878 & n2953 ) | ( ~n2928 & n2953 ) ;
  assign n2956 = ( n2928 & ~n2954 ) | ( n2928 & n2955 ) | ( ~n2954 & n2955 ) ;
  assign n2957 = n1527 & n2665 ;
  assign n2958 = n1629 & n2667 ;
  assign n2959 = ( n1631 & n2457 ) | ( n1631 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n2960 = ( n1531 & n2539 ) | ( n1531 & n2540 ) | ( n2539 & n2540 ) ;
  assign n2961 = n2959 | n2960 ;
  assign n2962 = ( ~n2957 & n2958 ) | ( ~n2957 & n2961 ) | ( n2958 & n2961 ) ;
  assign n2963 = ( ~n500 & n2957 ) | ( ~n500 & n2962 ) | ( n2957 & n2962 ) ;
  assign n2964 = ( n2957 & n2962 ) | ( n2957 & ~n2963 ) | ( n2962 & ~n2963 ) ;
  assign n2965 = ( n500 & n2963 ) | ( n500 & ~n2964 ) | ( n2963 & ~n2964 ) ;
  assign n2966 = ( n2890 & n2956 ) | ( n2890 & n2965 ) | ( n2956 & n2965 ) ;
  assign n2967 = ( n2890 & ~n2956 ) | ( n2890 & n2965 ) | ( ~n2956 & n2965 ) ;
  assign n2968 = ( n2956 & ~n2966 ) | ( n2956 & n2967 ) | ( ~n2966 & n2967 ) ;
  assign n2969 = n1260 & ~n2790 ;
  assign n2970 = n1450 & ~n2831 ;
  assign n2971 = n2790 & ~n2815 ;
  assign n2972 = ~n2815 & n2831 ;
  assign n2973 = ~n2790 & n2831 ;
  assign n2974 = ( n2971 & ~n2972 ) | ( n2971 & n2973 ) | ( ~n2972 & n2973 ) ;
  assign n2975 = n2970 | n2974 ;
  assign n2976 = ( n1439 & n2970 ) | ( n1439 & n2975 ) | ( n2970 & n2975 ) ;
  assign n2977 = ( n1262 & ~n2969 ) | ( n1262 & n2976 ) | ( ~n2969 & n2976 ) ;
  assign n2978 = n1262 & ~n2976 ;
  assign n2979 = ( ~n1262 & n2977 ) | ( ~n1262 & n2978 ) | ( n2977 & n2978 ) ;
  assign n2980 = ( n2893 & n2968 ) | ( n2893 & n2979 ) | ( n2968 & n2979 ) ;
  assign n2981 = ( n2893 & ~n2968 ) | ( n2893 & n2979 ) | ( ~n2968 & n2979 ) ;
  assign n2982 = ( n2968 & ~n2980 ) | ( n2968 & n2981 ) | ( ~n2980 & n2981 ) ;
  assign n2983 = n112 | n538 ;
  assign n2984 = ( n98 & n111 ) | ( n98 & n206 ) | ( n111 & n206 ) ;
  assign n2985 = n329 | n2984 ;
  assign n2986 = ( n2188 & ~n2983 ) | ( n2188 & n2985 ) | ( ~n2983 & n2985 ) ;
  assign n2987 = n2983 | n2986 ;
  assign n2988 = n133 | n325 ;
  assign n2989 = ( n617 & n785 ) | ( n617 & ~n2988 ) | ( n785 & ~n2988 ) ;
  assign n2990 = n2988 | n2989 ;
  assign n2991 = n88 | n308 ;
  assign n2992 = ( n797 & n901 ) | ( n797 & ~n2991 ) | ( n901 & ~n2991 ) ;
  assign n2993 = n2991 | n2992 ;
  assign n2994 = ( ~n2987 & n2990 ) | ( ~n2987 & n2993 ) | ( n2990 & n2993 ) ;
  assign n2995 = ( ~n616 & n2987 ) | ( ~n616 & n2994 ) | ( n2987 & n2994 ) ;
  assign n2996 = ( n616 & n2592 ) | ( n616 & ~n2995 ) | ( n2592 & ~n2995 ) ;
  assign n2997 = n2995 | n2996 ;
  assign n2998 = ( n2910 & n2982 ) | ( n2910 & n2997 ) | ( n2982 & n2997 ) ;
  assign n2999 = ( n2910 & ~n2982 ) | ( n2910 & n2997 ) | ( ~n2982 & n2997 ) ;
  assign n3000 = ( n2982 & ~n2998 ) | ( n2982 & n2999 ) | ( ~n2998 & n2999 ) ;
  assign n3001 = ( ~n2914 & n2917 ) | ( ~n2914 & n3000 ) | ( n2917 & n3000 ) ;
  assign n3002 = ( n2917 & n3000 ) | ( n2917 & ~n3001 ) | ( n3000 & ~n3001 ) ;
  assign n3003 = ( n2914 & n3001 ) | ( n2914 & ~n3002 ) | ( n3001 & ~n3002 ) ;
  assign n3004 = n2914 & n3000 ;
  assign n3005 = ( n2915 & n3000 ) | ( n2915 & ~n3004 ) | ( n3000 & ~n3004 ) ;
  assign n3006 = ( n2914 & ~n3004 ) | ( n2914 & n3005 ) | ( ~n3004 & n3005 ) ;
  assign n3007 = n2814 & n3006 ;
  assign n3008 = ( n1808 & n2457 ) | ( n1808 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3009 = ( n1917 & n2282 ) | ( n1917 & n2283 ) | ( n2282 & n2283 ) ;
  assign n3010 = ( n1812 & n2380 ) | ( n1812 & n2381 ) | ( n2380 & n2381 ) ;
  assign n3011 = n3009 | n3010 ;
  assign n3012 = ( n1806 & ~n2462 ) | ( n1806 & n2464 ) | ( ~n2462 & n2464 ) ;
  assign n3013 = ( ~n3008 & n3011 ) | ( ~n3008 & n3012 ) | ( n3011 & n3012 ) ;
  assign n3014 = ( n705 & ~n3008 ) | ( n705 & n3013 ) | ( ~n3008 & n3013 ) ;
  assign n3015 = ( n705 & n3013 ) | ( n705 & ~n3014 ) | ( n3013 & ~n3014 ) ;
  assign n3016 = ( n3008 & n3014 ) | ( n3008 & ~n3015 ) | ( n3014 & ~n3015 ) ;
  assign n3017 = n2079 & ~n2215 ;
  assign n3018 = n2078 & ~n2212 ;
  assign n3019 = n2044 & n2147 ;
  assign n3020 = ( n2082 & n2083 ) | ( n2082 & n2132 ) | ( n2083 & n2132 ) ;
  assign n3021 = ( ~n2083 & n3019 ) | ( ~n2083 & n3020 ) | ( n3019 & n3020 ) ;
  assign n3022 = ( ~n3017 & n3018 ) | ( ~n3017 & n3021 ) | ( n3018 & n3021 ) ;
  assign n3023 = ( ~n863 & n3017 ) | ( ~n863 & n3022 ) | ( n3017 & n3022 ) ;
  assign n3024 = ( n3017 & n3022 ) | ( n3017 & ~n3023 ) | ( n3022 & ~n3023 ) ;
  assign n3025 = ( n863 & n3023 ) | ( n863 & ~n3024 ) | ( n3023 & ~n3024 ) ;
  assign n3026 = n1763 & n2418 ;
  assign n3027 = ~n1892 & n2322 ;
  assign n3028 = n3026 | n3027 ;
  assign n3029 = n1970 & ~n2324 ;
  assign n3030 = ( n1970 & n3028 ) | ( n1970 & ~n3029 ) | ( n3028 & ~n3029 ) ;
  assign n3031 = ~n1973 & n2316 ;
  assign n3032 = n3030 | n3031 ;
  assign n3033 = n943 & ~n1694 ;
  assign n3034 = n943 | n2944 ;
  assign n3035 = ~n2948 & n3034 ;
  assign n3036 = ( ~n3032 & n3033 ) | ( ~n3032 & n3035 ) | ( n3033 & n3035 ) ;
  assign n3037 = ( n3032 & n3033 ) | ( n3032 & n3035 ) | ( n3033 & n3035 ) ;
  assign n3038 = ( n3032 & n3036 ) | ( n3032 & ~n3037 ) | ( n3036 & ~n3037 ) ;
  assign n3039 = ( n2951 & n3025 ) | ( n2951 & n3038 ) | ( n3025 & n3038 ) ;
  assign n3040 = ( n2951 & ~n3025 ) | ( n2951 & n3038 ) | ( ~n3025 & n3038 ) ;
  assign n3041 = ( n3025 & ~n3039 ) | ( n3025 & n3040 ) | ( ~n3039 & n3040 ) ;
  assign n3042 = ( n2954 & n3016 ) | ( n2954 & n3041 ) | ( n3016 & n3041 ) ;
  assign n3043 = ( n2954 & ~n3016 ) | ( n2954 & n3041 ) | ( ~n3016 & n3041 ) ;
  assign n3044 = ( n3016 & ~n3042 ) | ( n3016 & n3043 ) | ( ~n3042 & n3043 ) ;
  assign n3045 = ( n2790 & n2831 ) | ( n2790 & n2971 ) | ( n2831 & n2971 ) ;
  assign n3046 = n1439 & ~n3045 ;
  assign n3047 = ( n1260 & ~n2831 ) | ( n1260 & n3046 ) | ( ~n2831 & n3046 ) ;
  assign n3048 = n1262 | n3047 ;
  assign n3049 = ( n1262 & n3047 ) | ( n1262 & ~n3048 ) | ( n3047 & ~n3048 ) ;
  assign n3050 = n3048 & ~n3049 ;
  assign n3051 = n1527 & ~n2793 ;
  assign n3052 = n1629 & ~n2790 ;
  assign n3053 = ( n1631 & n2539 ) | ( n1631 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3054 = n1531 & n2667 ;
  assign n3055 = n3053 | n3054 ;
  assign n3056 = ( ~n3051 & n3052 ) | ( ~n3051 & n3055 ) | ( n3052 & n3055 ) ;
  assign n3057 = ( ~n500 & n3051 ) | ( ~n500 & n3056 ) | ( n3051 & n3056 ) ;
  assign n3058 = ( n3051 & n3056 ) | ( n3051 & ~n3057 ) | ( n3056 & ~n3057 ) ;
  assign n3059 = ( n500 & n3057 ) | ( n500 & ~n3058 ) | ( n3057 & ~n3058 ) ;
  assign n3060 = ( n3044 & n3050 ) | ( n3044 & n3059 ) | ( n3050 & n3059 ) ;
  assign n3061 = ( ~n3044 & n3050 ) | ( ~n3044 & n3059 ) | ( n3050 & n3059 ) ;
  assign n3062 = ( n3044 & ~n3060 ) | ( n3044 & n3061 ) | ( ~n3060 & n3061 ) ;
  assign n3063 = ( n2966 & n2980 ) | ( n2966 & n3062 ) | ( n2980 & n3062 ) ;
  assign n3064 = ( n2966 & ~n2980 ) | ( n2966 & n3062 ) | ( ~n2980 & n3062 ) ;
  assign n3065 = ( n2980 & ~n3063 ) | ( n2980 & n3064 ) | ( ~n3063 & n3064 ) ;
  assign n3066 = n651 | n849 ;
  assign n3067 = n2564 | n3066 ;
  assign n3068 = ( n107 & n126 ) | ( n107 & n163 ) | ( n126 & n163 ) ;
  assign n3069 = n890 | n1684 ;
  assign n3070 = n3068 | n3069 ;
  assign n3071 = n470 | n1850 ;
  assign n3072 = ( ~n206 & n243 ) | ( ~n206 & n427 ) | ( n243 & n427 ) ;
  assign n3073 = ( n143 & n203 ) | ( n143 & ~n3072 ) | ( n203 & ~n3072 ) ;
  assign n3074 = n3072 | n3073 ;
  assign n3075 = ( ~n3070 & n3071 ) | ( ~n3070 & n3074 ) | ( n3071 & n3074 ) ;
  assign n3076 = n3070 | n3075 ;
  assign n3077 = ( n558 & ~n3067 ) | ( n558 & n3076 ) | ( ~n3067 & n3076 ) ;
  assign n3078 = n3067 | n3077 ;
  assign n3079 = ( n2998 & n3065 ) | ( n2998 & n3078 ) | ( n3065 & n3078 ) ;
  assign n3080 = ( n2998 & ~n3065 ) | ( n2998 & n3078 ) | ( ~n3065 & n3078 ) ;
  assign n3081 = ( n3065 & ~n3079 ) | ( n3065 & n3080 ) | ( ~n3079 & n3080 ) ;
  assign n3082 = ( n3004 & n3007 ) | ( n3004 & n3081 ) | ( n3007 & n3081 ) ;
  assign n3083 = n3004 | n3081 ;
  assign n3084 = ~n3007 & n3083 ;
  assign n3085 = ( n3007 & ~n3082 ) | ( n3007 & n3084 ) | ( ~n3082 & n3084 ) ;
  assign n3086 = n3004 & n3081 ;
  assign n3087 = ( n3006 & n3083 ) | ( n3006 & ~n3086 ) | ( n3083 & ~n3086 ) ;
  assign n3088 = n2814 & n3087 ;
  assign n3089 = n1806 & ~n2537 ;
  assign n3090 = ( n1808 & n2539 ) | ( n1808 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3091 = ( n1917 & n2380 ) | ( n1917 & n2381 ) | ( n2380 & n2381 ) ;
  assign n3092 = ( n1812 & n2457 ) | ( n1812 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3093 = n3091 | n3092 ;
  assign n3094 = ( ~n3089 & n3090 ) | ( ~n3089 & n3093 ) | ( n3090 & n3093 ) ;
  assign n3095 = ( n705 & ~n3089 ) | ( n705 & n3094 ) | ( ~n3089 & n3094 ) ;
  assign n3096 = ( n705 & n3094 ) | ( n705 & ~n3095 ) | ( n3094 & ~n3095 ) ;
  assign n3097 = ( n3089 & n3095 ) | ( n3089 & ~n3096 ) | ( n3095 & ~n3096 ) ;
  assign n3098 = n943 & n1763 ;
  assign n3099 = n2047 & n2316 ;
  assign n3100 = n2044 & n2324 ;
  assign n3101 = ~n1892 & n2418 ;
  assign n3102 = n1970 & n2322 ;
  assign n3103 = n3101 | n3102 ;
  assign n3104 = ( ~n3099 & n3100 ) | ( ~n3099 & n3103 ) | ( n3100 & n3103 ) ;
  assign n3105 = ( ~n943 & n3099 ) | ( ~n943 & n3104 ) | ( n3099 & n3104 ) ;
  assign n3106 = ( n3099 & n3104 ) | ( n3099 & ~n3105 ) | ( n3104 & ~n3105 ) ;
  assign n3107 = ( n943 & n3105 ) | ( n943 & ~n3106 ) | ( n3105 & ~n3106 ) ;
  assign n3108 = ( n1262 & n3098 ) | ( n1262 & n3107 ) | ( n3098 & n3107 ) ;
  assign n3109 = ( n1262 & ~n3098 ) | ( n1262 & n3107 ) | ( ~n3098 & n3107 ) ;
  assign n3110 = ( n3098 & ~n3108 ) | ( n3098 & n3109 ) | ( ~n3108 & n3109 ) ;
  assign n3111 = n943 & ~n3032 ;
  assign n3112 = ( ~n3033 & n3037 ) | ( ~n3033 & n3111 ) | ( n3037 & n3111 ) ;
  assign n3113 = n2079 & ~n2287 ;
  assign n3114 = ( n2078 & n2282 ) | ( n2078 & n2283 ) | ( n2282 & n2283 ) ;
  assign n3115 = n2132 & n2147 ;
  assign n3116 = ( n2082 & n2083 ) | ( n2082 & ~n2212 ) | ( n2083 & ~n2212 ) ;
  assign n3117 = ( ~n2083 & n3115 ) | ( ~n2083 & n3116 ) | ( n3115 & n3116 ) ;
  assign n3118 = ( ~n3113 & n3114 ) | ( ~n3113 & n3117 ) | ( n3114 & n3117 ) ;
  assign n3119 = ( ~n863 & n3113 ) | ( ~n863 & n3118 ) | ( n3113 & n3118 ) ;
  assign n3120 = ( n3113 & n3118 ) | ( n3113 & ~n3119 ) | ( n3118 & ~n3119 ) ;
  assign n3121 = ( n863 & n3119 ) | ( n863 & ~n3120 ) | ( n3119 & ~n3120 ) ;
  assign n3122 = ( n3110 & n3112 ) | ( n3110 & n3121 ) | ( n3112 & n3121 ) ;
  assign n3123 = ( ~n3110 & n3112 ) | ( ~n3110 & n3121 ) | ( n3112 & n3121 ) ;
  assign n3124 = ( n3110 & ~n3122 ) | ( n3110 & n3123 ) | ( ~n3122 & n3123 ) ;
  assign n3125 = ( n3039 & n3097 ) | ( n3039 & n3124 ) | ( n3097 & n3124 ) ;
  assign n3126 = ( n3039 & ~n3097 ) | ( n3039 & n3124 ) | ( ~n3097 & n3124 ) ;
  assign n3127 = ( n3097 & ~n3125 ) | ( n3097 & n3126 ) | ( ~n3125 & n3126 ) ;
  assign n3128 = n1527 & n2834 ;
  assign n3129 = n1631 & n2667 ;
  assign n3130 = n1531 & ~n2790 ;
  assign n3131 = n3129 | n3130 ;
  assign n3132 = n1629 & ~n2831 ;
  assign n3133 = ( ~n3128 & n3131 ) | ( ~n3128 & n3132 ) | ( n3131 & n3132 ) ;
  assign n3134 = ( ~n500 & n3128 ) | ( ~n500 & n3133 ) | ( n3128 & n3133 ) ;
  assign n3135 = ( n3128 & n3133 ) | ( n3128 & ~n3134 ) | ( n3133 & ~n3134 ) ;
  assign n3136 = ( n500 & n3134 ) | ( n500 & ~n3135 ) | ( n3134 & ~n3135 ) ;
  assign n3137 = ( n3042 & n3127 ) | ( n3042 & n3136 ) | ( n3127 & n3136 ) ;
  assign n3138 = ( n3042 & ~n3127 ) | ( n3042 & n3136 ) | ( ~n3127 & n3136 ) ;
  assign n3139 = ( n3127 & ~n3137 ) | ( n3127 & n3138 ) | ( ~n3137 & n3138 ) ;
  assign n3140 = ( n3060 & n3063 ) | ( n3060 & n3139 ) | ( n3063 & n3139 ) ;
  assign n3141 = ( n3060 & ~n3063 ) | ( n3060 & n3139 ) | ( ~n3063 & n3139 ) ;
  assign n3142 = ( n3063 & ~n3140 ) | ( n3063 & n3141 ) | ( ~n3140 & n3141 ) ;
  assign n3143 = n772 | n1395 ;
  assign n3144 = n154 | n248 ;
  assign n3145 = ( n618 & ~n715 ) | ( n618 & n1574 ) | ( ~n715 & n1574 ) ;
  assign n3146 = n715 | n3145 ;
  assign n3147 = ( n337 & ~n3144 ) | ( n337 & n3146 ) | ( ~n3144 & n3146 ) ;
  assign n3148 = n3144 | n3147 ;
  assign n3149 = ( n2188 & ~n3143 ) | ( n2188 & n3148 ) | ( ~n3143 & n3148 ) ;
  assign n3150 = n3143 | n3149 ;
  assign n3151 = n519 | n729 ;
  assign n3152 = ( n1288 & ~n3150 ) | ( n1288 & n3151 ) | ( ~n3150 & n3151 ) ;
  assign n3153 = n3150 | n3152 ;
  assign n3154 = ( n3079 & n3142 ) | ( n3079 & n3153 ) | ( n3142 & n3153 ) ;
  assign n3155 = ( n3079 & ~n3142 ) | ( n3079 & n3153 ) | ( ~n3142 & n3153 ) ;
  assign n3156 = ( n3142 & ~n3154 ) | ( n3142 & n3155 ) | ( ~n3154 & n3155 ) ;
  assign n3157 = ( ~n3086 & n3088 ) | ( ~n3086 & n3156 ) | ( n3088 & n3156 ) ;
  assign n3158 = ( n3088 & n3156 ) | ( n3088 & ~n3157 ) | ( n3156 & ~n3157 ) ;
  assign n3159 = ( n3086 & n3157 ) | ( n3086 & ~n3158 ) | ( n3157 & ~n3158 ) ;
  assign n3160 = n3086 & n3156 ;
  assign n3161 = n1527 & n2974 ;
  assign n3162 = n1631 & ~n2790 ;
  assign n3163 = n1531 & ~n2831 ;
  assign n3164 = n3162 | n3163 ;
  assign n3165 = ( ~n500 & n3161 ) | ( ~n500 & n3164 ) | ( n3161 & n3164 ) ;
  assign n3166 = ( n3161 & n3164 ) | ( n3161 & ~n3165 ) | ( n3164 & ~n3165 ) ;
  assign n3167 = ( n500 & n3165 ) | ( n500 & ~n3166 ) | ( n3165 & ~n3166 ) ;
  assign n3168 = n1806 & n2665 ;
  assign n3169 = n1808 & n2667 ;
  assign n3170 = ( n1917 & n2457 ) | ( n1917 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3171 = ( n1812 & n2539 ) | ( n1812 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3172 = n3170 | n3171 ;
  assign n3173 = ( ~n3168 & n3169 ) | ( ~n3168 & n3172 ) | ( n3169 & n3172 ) ;
  assign n3174 = ( n705 & ~n3168 ) | ( n705 & n3173 ) | ( ~n3168 & n3173 ) ;
  assign n3175 = ( n705 & n3173 ) | ( n705 & ~n3174 ) | ( n3173 & ~n3174 ) ;
  assign n3176 = ( n3168 & n3174 ) | ( n3168 & ~n3175 ) | ( n3174 & ~n3175 ) ;
  assign n3177 = n2135 & n2316 ;
  assign n3178 = n2132 & n2324 ;
  assign n3179 = n1970 & n2418 ;
  assign n3180 = n2044 & n2322 ;
  assign n3181 = n3179 | n3180 ;
  assign n3182 = ( ~n3177 & n3178 ) | ( ~n3177 & n3181 ) | ( n3178 & n3181 ) ;
  assign n3183 = ( ~n943 & n3177 ) | ( ~n943 & n3182 ) | ( n3177 & n3182 ) ;
  assign n3184 = ( n3177 & n3182 ) | ( n3177 & ~n3183 ) | ( n3182 & ~n3183 ) ;
  assign n3185 = ( n943 & n3183 ) | ( n943 & ~n3184 ) | ( n3183 & ~n3184 ) ;
  assign n3186 = n2079 & n2385 ;
  assign n3187 = ( n2078 & n2380 ) | ( n2078 & n2381 ) | ( n2380 & n2381 ) ;
  assign n3188 = ( n2084 & n2282 ) | ( n2084 & n2283 ) | ( n2282 & n2283 ) ;
  assign n3189 = n2147 & n2212 ;
  assign n3190 = ( n2147 & n3188 ) | ( n2147 & ~n3189 ) | ( n3188 & ~n3189 ) ;
  assign n3191 = ( ~n3186 & n3187 ) | ( ~n3186 & n3190 ) | ( n3187 & n3190 ) ;
  assign n3192 = ( ~n863 & n3186 ) | ( ~n863 & n3191 ) | ( n3186 & n3191 ) ;
  assign n3193 = ( n3186 & n3191 ) | ( n3186 & ~n3192 ) | ( n3191 & ~n3192 ) ;
  assign n3194 = ( n863 & n3192 ) | ( n863 & ~n3193 ) | ( n3192 & ~n3193 ) ;
  assign n3195 = n943 & ~n1892 ;
  assign n3196 = ( n1262 & n3108 ) | ( n1262 & n3195 ) | ( n3108 & n3195 ) ;
  assign n3197 = ( ~n1262 & n3108 ) | ( ~n1262 & n3195 ) | ( n3108 & n3195 ) ;
  assign n3198 = ( n1262 & ~n3196 ) | ( n1262 & n3197 ) | ( ~n3196 & n3197 ) ;
  assign n3199 = ( n3185 & n3194 ) | ( n3185 & n3198 ) | ( n3194 & n3198 ) ;
  assign n3200 = ( ~n3185 & n3194 ) | ( ~n3185 & n3198 ) | ( n3194 & n3198 ) ;
  assign n3201 = ( n3185 & ~n3199 ) | ( n3185 & n3200 ) | ( ~n3199 & n3200 ) ;
  assign n3202 = ( n3122 & n3176 ) | ( n3122 & n3201 ) | ( n3176 & n3201 ) ;
  assign n3203 = ( n3122 & ~n3176 ) | ( n3122 & n3201 ) | ( ~n3176 & n3201 ) ;
  assign n3204 = ( n3176 & ~n3202 ) | ( n3176 & n3203 ) | ( ~n3202 & n3203 ) ;
  assign n3205 = ( n3125 & n3167 ) | ( n3125 & n3204 ) | ( n3167 & n3204 ) ;
  assign n3206 = ( n3125 & ~n3167 ) | ( n3125 & n3204 ) | ( ~n3167 & n3204 ) ;
  assign n3207 = ( n3167 & ~n3205 ) | ( n3167 & n3206 ) | ( ~n3205 & n3206 ) ;
  assign n3208 = ( n3137 & n3140 ) | ( n3137 & n3207 ) | ( n3140 & n3207 ) ;
  assign n3209 = ( n3137 & ~n3140 ) | ( n3137 & n3207 ) | ( ~n3140 & n3207 ) ;
  assign n3210 = ( n3140 & ~n3208 ) | ( n3140 & n3209 ) | ( ~n3208 & n3209 ) ;
  assign n3211 = n820 | n1598 ;
  assign n3212 = n309 | n321 ;
  assign n3213 = n203 | n1401 ;
  assign n3214 = ( n257 & n283 ) | ( n257 & ~n602 ) | ( n283 & ~n602 ) ;
  assign n3215 = n533 | n715 ;
  assign n3216 = n3214 | n3215 ;
  assign n3217 = ( n3212 & ~n3213 ) | ( n3212 & n3216 ) | ( ~n3213 & n3216 ) ;
  assign n3218 = ( n2903 & n3213 ) | ( n2903 & ~n3217 ) | ( n3213 & ~n3217 ) ;
  assign n3219 = n3217 | n3218 ;
  assign n3220 = ( ~n2364 & n3211 ) | ( ~n2364 & n3219 ) | ( n3211 & n3219 ) ;
  assign n3221 = ( ~n1735 & n2364 ) | ( ~n1735 & n3220 ) | ( n2364 & n3220 ) ;
  assign n3222 = ( n1735 & n2829 ) | ( n1735 & ~n3221 ) | ( n2829 & ~n3221 ) ;
  assign n3223 = n3221 | n3222 ;
  assign n3224 = ( n3154 & n3210 ) | ( n3154 & n3223 ) | ( n3210 & n3223 ) ;
  assign n3225 = ( n3154 & ~n3210 ) | ( n3154 & n3223 ) | ( ~n3210 & n3223 ) ;
  assign n3226 = ( n3210 & ~n3224 ) | ( n3210 & n3225 ) | ( ~n3224 & n3225 ) ;
  assign n3227 = ( n2814 & n3088 ) | ( n2814 & n3159 ) | ( n3088 & n3159 ) ;
  assign n3228 = ( ~n3160 & n3226 ) | ( ~n3160 & n3227 ) | ( n3226 & n3227 ) ;
  assign n3229 = ( n3226 & n3227 ) | ( n3226 & ~n3228 ) | ( n3227 & ~n3228 ) ;
  assign n3230 = ( n3160 & n3228 ) | ( n3160 & ~n3229 ) | ( n3228 & ~n3229 ) ;
  assign n3231 = n1527 & ~n3045 ;
  assign n3232 = ( n1631 & ~n2831 ) | ( n1631 & n3231 ) | ( ~n2831 & n3231 ) ;
  assign n3233 = n500 | n3232 ;
  assign n3234 = ( n500 & n3232 ) | ( n500 & ~n3233 ) | ( n3232 & ~n3233 ) ;
  assign n3235 = n3233 & ~n3234 ;
  assign n3236 = n1806 & ~n2793 ;
  assign n3237 = n1808 & ~n2790 ;
  assign n3238 = ( n1917 & n2539 ) | ( n1917 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3239 = n1812 & n2667 ;
  assign n3240 = n3238 | n3239 ;
  assign n3241 = ( ~n3236 & n3237 ) | ( ~n3236 & n3240 ) | ( n3237 & n3240 ) ;
  assign n3242 = ( n705 & ~n3236 ) | ( n705 & n3241 ) | ( ~n3236 & n3241 ) ;
  assign n3243 = ( n705 & n3241 ) | ( n705 & ~n3242 ) | ( n3241 & ~n3242 ) ;
  assign n3244 = ( n3236 & n3242 ) | ( n3236 & ~n3243 ) | ( n3242 & ~n3243 ) ;
  assign n3245 = ~n2215 & n2316 ;
  assign n3246 = ~n2212 & n2324 ;
  assign n3247 = n2044 & n2418 ;
  assign n3248 = n2132 & n2322 ;
  assign n3249 = n3247 | n3248 ;
  assign n3250 = ( ~n3245 & n3246 ) | ( ~n3245 & n3249 ) | ( n3246 & n3249 ) ;
  assign n3251 = ( ~n943 & n3245 ) | ( ~n943 & n3250 ) | ( n3245 & n3250 ) ;
  assign n3252 = ( n3245 & n3250 ) | ( n3245 & ~n3251 ) | ( n3250 & ~n3251 ) ;
  assign n3253 = ( n943 & n3251 ) | ( n943 & ~n3252 ) | ( n3251 & ~n3252 ) ;
  assign n3254 = ( n2078 & n2457 ) | ( n2078 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3255 = ( n2079 & ~n2462 ) | ( n2079 & n2464 ) | ( ~n2462 & n2464 ) ;
  assign n3256 = ( n2147 & n2282 ) | ( n2147 & n2283 ) | ( n2282 & n2283 ) ;
  assign n3257 = ( n2082 & n2083 ) | ( n2082 & n2382 ) | ( n2083 & n2382 ) ;
  assign n3258 = ( ~n2083 & n3256 ) | ( ~n2083 & n3257 ) | ( n3256 & n3257 ) ;
  assign n3259 = ( ~n3254 & n3255 ) | ( ~n3254 & n3258 ) | ( n3255 & n3258 ) ;
  assign n3260 = ( ~n863 & n3254 ) | ( ~n863 & n3259 ) | ( n3254 & n3259 ) ;
  assign n3261 = ( n3254 & n3259 ) | ( n3254 & ~n3260 ) | ( n3259 & ~n3260 ) ;
  assign n3262 = ( n863 & n3260 ) | ( n863 & ~n3261 ) | ( n3260 & ~n3261 ) ;
  assign n3263 = n943 & n1970 ;
  assign n3264 = ( n1262 & n3196 ) | ( n1262 & n3263 ) | ( n3196 & n3263 ) ;
  assign n3265 = ( n1262 & ~n3196 ) | ( n1262 & n3263 ) | ( ~n3196 & n3263 ) ;
  assign n3266 = ( n3196 & ~n3264 ) | ( n3196 & n3265 ) | ( ~n3264 & n3265 ) ;
  assign n3267 = ( n3253 & n3262 ) | ( n3253 & n3266 ) | ( n3262 & n3266 ) ;
  assign n3268 = ( ~n3253 & n3262 ) | ( ~n3253 & n3266 ) | ( n3262 & n3266 ) ;
  assign n3269 = ( n3253 & ~n3267 ) | ( n3253 & n3268 ) | ( ~n3267 & n3268 ) ;
  assign n3270 = ( n3199 & n3244 ) | ( n3199 & n3269 ) | ( n3244 & n3269 ) ;
  assign n3271 = ( n3199 & ~n3244 ) | ( n3199 & n3269 ) | ( ~n3244 & n3269 ) ;
  assign n3272 = ( n3244 & ~n3270 ) | ( n3244 & n3271 ) | ( ~n3270 & n3271 ) ;
  assign n3273 = ( n3202 & n3235 ) | ( n3202 & n3272 ) | ( n3235 & n3272 ) ;
  assign n3274 = ( n3202 & ~n3235 ) | ( n3202 & n3272 ) | ( ~n3235 & n3272 ) ;
  assign n3275 = ( n3235 & ~n3273 ) | ( n3235 & n3274 ) | ( ~n3273 & n3274 ) ;
  assign n3276 = ( n3205 & n3208 ) | ( n3205 & n3275 ) | ( n3208 & n3275 ) ;
  assign n3277 = ( n3205 & ~n3208 ) | ( n3205 & n3275 ) | ( ~n3208 & n3275 ) ;
  assign n3278 = ( n3208 & ~n3276 ) | ( n3208 & n3277 ) | ( ~n3276 & n3277 ) ;
  assign n3279 = ( n726 & n1755 ) | ( n726 & ~n2526 ) | ( n1755 & ~n2526 ) ;
  assign n3280 = n2526 | n3279 ;
  assign n3281 = n311 | n326 ;
  assign n3282 = n150 | n170 ;
  assign n3283 = ( n1278 & ~n3281 ) | ( n1278 & n3282 ) | ( ~n3281 & n3282 ) ;
  assign n3284 = n3281 | n3283 ;
  assign n3285 = ( ~n2709 & n3280 ) | ( ~n2709 & n3284 ) | ( n3280 & n3284 ) ;
  assign n3286 = n670 | n2820 ;
  assign n3287 = n1598 | n1684 ;
  assign n3288 = ( n1282 & n1397 ) | ( n1282 & ~n3287 ) | ( n1397 & ~n3287 ) ;
  assign n3289 = n3287 | n3288 ;
  assign n3290 = n380 | n653 ;
  assign n3291 = ( ~n3286 & n3289 ) | ( ~n3286 & n3290 ) | ( n3289 & n3290 ) ;
  assign n3292 = n3286 | n3291 ;
  assign n3293 = ( n2709 & ~n3285 ) | ( n2709 & n3292 ) | ( ~n3285 & n3292 ) ;
  assign n3294 = n3285 | n3293 ;
  assign n3295 = ( n3224 & n3278 ) | ( n3224 & n3294 ) | ( n3278 & n3294 ) ;
  assign n3296 = ( n3224 & ~n3278 ) | ( n3224 & n3294 ) | ( ~n3278 & n3294 ) ;
  assign n3297 = ( n3278 & ~n3295 ) | ( n3278 & n3296 ) | ( ~n3295 & n3296 ) ;
  assign n3298 = n3160 & n3226 ;
  assign n3299 = n3297 & n3298 ;
  assign n3300 = ~n3160 & n3226 ;
  assign n3301 = ( n3086 & ~n3087 ) | ( n3086 & n3156 ) | ( ~n3087 & n3156 ) ;
  assign n3302 = ( n3087 & ~n3226 ) | ( n3087 & n3301 ) | ( ~n3226 & n3301 ) ;
  assign n3303 = ( n2814 & n3300 ) | ( n2814 & n3302 ) | ( n3300 & n3302 ) ;
  assign n3304 = ( n3297 & n3298 ) | ( n3297 & ~n3303 ) | ( n3298 & ~n3303 ) ;
  assign n3305 = ( n3226 & n3297 ) | ( n3226 & ~n3300 ) | ( n3297 & ~n3300 ) ;
  assign n3306 = ( n3299 & n3303 ) | ( n3299 & ~n3305 ) | ( n3303 & ~n3305 ) ;
  assign n3307 = ( ~n3299 & n3304 ) | ( ~n3299 & n3306 ) | ( n3304 & n3306 ) ;
  assign n3308 = ~n3299 & n3305 ;
  assign n3309 = ( n2814 & n3303 ) | ( n2814 & n3308 ) | ( n3303 & n3308 ) ;
  assign n3310 = n1806 & n2834 ;
  assign n3311 = n1917 & n2667 ;
  assign n3312 = n1812 & ~n2790 ;
  assign n3313 = n3311 | n3312 ;
  assign n3314 = n1808 & ~n2831 ;
  assign n3315 = ( ~n3310 & n3313 ) | ( ~n3310 & n3314 ) | ( n3313 & n3314 ) ;
  assign n3316 = ( n705 & ~n3310 ) | ( n705 & n3315 ) | ( ~n3310 & n3315 ) ;
  assign n3317 = ( n705 & n3315 ) | ( n705 & ~n3316 ) | ( n3315 & ~n3316 ) ;
  assign n3318 = ( n3310 & n3316 ) | ( n3310 & ~n3317 ) | ( n3316 & ~n3317 ) ;
  assign n3319 = n2079 & ~n2537 ;
  assign n3320 = ( n2078 & n2539 ) | ( n2078 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3321 = ( n2147 & n2380 ) | ( n2147 & n2381 ) | ( n2380 & n2381 ) ;
  assign n3322 = ( n2082 & n2083 ) | ( n2082 & ~n2523 ) | ( n2083 & ~n2523 ) ;
  assign n3323 = ( ~n2083 & n3321 ) | ( ~n2083 & n3322 ) | ( n3321 & n3322 ) ;
  assign n3324 = ( ~n3319 & n3320 ) | ( ~n3319 & n3323 ) | ( n3320 & n3323 ) ;
  assign n3325 = ( ~n863 & n3319 ) | ( ~n863 & n3324 ) | ( n3319 & n3324 ) ;
  assign n3326 = ( n3319 & n3324 ) | ( n3319 & ~n3325 ) | ( n3324 & ~n3325 ) ;
  assign n3327 = ( n863 & n3325 ) | ( n863 & ~n3326 ) | ( n3325 & ~n3326 ) ;
  assign n3328 = ~n2287 & n2316 ;
  assign n3329 = ( n2282 & n2283 ) | ( n2282 & n2324 ) | ( n2283 & n2324 ) ;
  assign n3330 = n2132 & n2418 ;
  assign n3331 = ~n2212 & n2322 ;
  assign n3332 = n3330 | n3331 ;
  assign n3333 = ( ~n3328 & n3329 ) | ( ~n3328 & n3332 ) | ( n3329 & n3332 ) ;
  assign n3334 = ( ~n943 & n3328 ) | ( ~n943 & n3333 ) | ( n3328 & n3333 ) ;
  assign n3335 = ( n3328 & n3333 ) | ( n3328 & ~n3334 ) | ( n3333 & ~n3334 ) ;
  assign n3336 = ( n943 & n3334 ) | ( n943 & ~n3335 ) | ( n3334 & ~n3335 ) ;
  assign n3337 = n943 & n2044 ;
  assign n3338 = ( n500 & n1262 ) | ( n500 & ~n3337 ) | ( n1262 & ~n3337 ) ;
  assign n3339 = ( n500 & ~n1262 ) | ( n500 & n3337 ) | ( ~n1262 & n3337 ) ;
  assign n3340 = ( ~n500 & n3338 ) | ( ~n500 & n3339 ) | ( n3338 & n3339 ) ;
  assign n3341 = ( n3264 & n3336 ) | ( n3264 & n3340 ) | ( n3336 & n3340 ) ;
  assign n3342 = ( n3264 & ~n3336 ) | ( n3264 & n3340 ) | ( ~n3336 & n3340 ) ;
  assign n3343 = ( n3336 & ~n3341 ) | ( n3336 & n3342 ) | ( ~n3341 & n3342 ) ;
  assign n3344 = ( n3267 & n3327 ) | ( n3267 & n3343 ) | ( n3327 & n3343 ) ;
  assign n3345 = ( n3267 & ~n3327 ) | ( n3267 & n3343 ) | ( ~n3327 & n3343 ) ;
  assign n3346 = ( n3327 & ~n3344 ) | ( n3327 & n3345 ) | ( ~n3344 & n3345 ) ;
  assign n3347 = ( n3270 & n3318 ) | ( n3270 & n3346 ) | ( n3318 & n3346 ) ;
  assign n3348 = ( n3270 & ~n3318 ) | ( n3270 & n3346 ) | ( ~n3318 & n3346 ) ;
  assign n3349 = ( n3318 & ~n3347 ) | ( n3318 & n3348 ) | ( ~n3347 & n3348 ) ;
  assign n3350 = ( n3273 & n3276 ) | ( n3273 & n3349 ) | ( n3276 & n3349 ) ;
  assign n3351 = ( n3273 & ~n3276 ) | ( n3273 & n3349 ) | ( ~n3276 & n3349 ) ;
  assign n3352 = ( n3276 & ~n3350 ) | ( n3276 & n3351 ) | ( ~n3350 & n3351 ) ;
  assign n3353 = n186 | n314 ;
  assign n3354 = ( n530 & n3213 ) | ( n530 & ~n3353 ) | ( n3213 & ~n3353 ) ;
  assign n3355 = n3353 | n3354 ;
  assign n3356 = n409 | n619 ;
  assign n3357 = n294 | n1574 ;
  assign n3358 = ( ~n83 & n282 ) | ( ~n83 & n3357 ) | ( n282 & n3357 ) ;
  assign n3359 = ( ~n3355 & n3356 ) | ( ~n3355 & n3358 ) | ( n3356 & n3358 ) ;
  assign n3360 = n3355 | n3359 ;
  assign n3361 = n1876 | n3292 ;
  assign n3362 = n3360 | n3361 ;
  assign n3363 = ( n3295 & n3352 ) | ( n3295 & n3362 ) | ( n3352 & n3362 ) ;
  assign n3364 = ( n3295 & ~n3352 ) | ( n3295 & n3362 ) | ( ~n3352 & n3362 ) ;
  assign n3365 = ( n3352 & ~n3363 ) | ( n3352 & n3364 ) | ( ~n3363 & n3364 ) ;
  assign n3366 = ( n3299 & ~n3309 ) | ( n3299 & n3365 ) | ( ~n3309 & n3365 ) ;
  assign n3367 = ( n3299 & n3365 ) | ( n3299 & ~n3366 ) | ( n3365 & ~n3366 ) ;
  assign n3368 = ( n3309 & n3366 ) | ( n3309 & ~n3367 ) | ( n3366 & ~n3367 ) ;
  assign n3369 = n1917 & ~n2790 ;
  assign n3370 = n1806 & n2974 ;
  assign n3371 = n1812 & ~n2831 ;
  assign n3372 = ( ~n3369 & n3370 ) | ( ~n3369 & n3371 ) | ( n3370 & n3371 ) ;
  assign n3373 = ( n705 & ~n3369 ) | ( n705 & n3372 ) | ( ~n3369 & n3372 ) ;
  assign n3374 = ( n705 & n3372 ) | ( n705 & ~n3373 ) | ( n3372 & ~n3373 ) ;
  assign n3375 = ( n3369 & n3373 ) | ( n3369 & ~n3374 ) | ( n3373 & ~n3374 ) ;
  assign n3376 = n2079 & n2665 ;
  assign n3377 = n2078 & n2667 ;
  assign n3378 = ( n2147 & n2457 ) | ( n2147 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3379 = ( n2082 & n2083 ) | ( n2082 & n2663 ) | ( n2083 & n2663 ) ;
  assign n3380 = ( ~n2083 & n3378 ) | ( ~n2083 & n3379 ) | ( n3378 & n3379 ) ;
  assign n3381 = ( ~n3376 & n3377 ) | ( ~n3376 & n3380 ) | ( n3377 & n3380 ) ;
  assign n3382 = ( ~n863 & n3376 ) | ( ~n863 & n3381 ) | ( n3376 & n3381 ) ;
  assign n3383 = ( n3376 & n3381 ) | ( n3376 & ~n3382 ) | ( n3381 & ~n3382 ) ;
  assign n3384 = ( n863 & n3382 ) | ( n863 & ~n3383 ) | ( n3382 & ~n3383 ) ;
  assign n3385 = n943 & n2132 ;
  assign n3386 = n2316 & n2385 ;
  assign n3387 = ( n2324 & n2380 ) | ( n2324 & n2381 ) | ( n2380 & n2381 ) ;
  assign n3388 = ( n2282 & n2283 ) | ( n2282 & n2322 ) | ( n2283 & n2322 ) ;
  assign n3389 = n2212 & n2418 ;
  assign n3390 = ( n2418 & n3388 ) | ( n2418 & ~n3389 ) | ( n3388 & ~n3389 ) ;
  assign n3391 = ( ~n3386 & n3387 ) | ( ~n3386 & n3390 ) | ( n3387 & n3390 ) ;
  assign n3392 = ( ~n943 & n3386 ) | ( ~n943 & n3391 ) | ( n3386 & n3391 ) ;
  assign n3393 = ( n3386 & n3391 ) | ( n3386 & ~n3392 ) | ( n3391 & ~n3392 ) ;
  assign n3394 = ( n943 & n3392 ) | ( n943 & ~n3393 ) | ( n3392 & ~n3393 ) ;
  assign n3395 = ( n3338 & n3385 ) | ( n3338 & ~n3394 ) | ( n3385 & ~n3394 ) ;
  assign n3396 = ( n3338 & ~n3385 ) | ( n3338 & n3394 ) | ( ~n3385 & n3394 ) ;
  assign n3397 = ( ~n3338 & n3395 ) | ( ~n3338 & n3396 ) | ( n3395 & n3396 ) ;
  assign n3398 = ( n3341 & n3384 ) | ( n3341 & n3397 ) | ( n3384 & n3397 ) ;
  assign n3399 = ( n3341 & ~n3384 ) | ( n3341 & n3397 ) | ( ~n3384 & n3397 ) ;
  assign n3400 = ( n3384 & ~n3398 ) | ( n3384 & n3399 ) | ( ~n3398 & n3399 ) ;
  assign n3401 = ( n3344 & n3375 ) | ( n3344 & n3400 ) | ( n3375 & n3400 ) ;
  assign n3402 = ( n3344 & ~n3375 ) | ( n3344 & n3400 ) | ( ~n3375 & n3400 ) ;
  assign n3403 = ( n3375 & ~n3401 ) | ( n3375 & n3402 ) | ( ~n3401 & n3402 ) ;
  assign n3404 = ( n3347 & n3350 ) | ( n3347 & n3403 ) | ( n3350 & n3403 ) ;
  assign n3405 = ( n3347 & ~n3350 ) | ( n3347 & n3403 ) | ( ~n3350 & n3403 ) ;
  assign n3406 = ( n3350 & ~n3404 ) | ( n3350 & n3405 ) | ( ~n3404 & n3405 ) ;
  assign n3407 = ( n56 & n224 ) | ( n56 & n363 ) | ( n224 & n363 ) ;
  assign n3408 = n246 | n3407 ;
  assign n3409 = n144 | n574 ;
  assign n3410 = n1859 | n3409 ;
  assign n3411 = ( n1227 & n3408 ) | ( n1227 & ~n3410 ) | ( n3408 & ~n3410 ) ;
  assign n3412 = ( n679 & n3410 ) | ( n679 & ~n3411 ) | ( n3410 & ~n3411 ) ;
  assign n3413 = n3411 | n3412 ;
  assign n3414 = ( n735 & ~n745 ) | ( n735 & n1679 ) | ( ~n745 & n1679 ) ;
  assign n3415 = n2580 | n3414 ;
  assign n3416 = ( n57 & n84 ) | ( n57 & n91 ) | ( n84 & n91 ) ;
  assign n3417 = n458 | n3416 ;
  assign n3418 = n745 | n3417 ;
  assign n3419 = ( ~n352 & n371 ) | ( ~n352 & n1270 ) | ( n371 & n1270 ) ;
  assign n3420 = n352 | n3419 ;
  assign n3421 = ( ~n3414 & n3418 ) | ( ~n3414 & n3420 ) | ( n3418 & n3420 ) ;
  assign n3422 = ( ~n3413 & n3415 ) | ( ~n3413 & n3421 ) | ( n3415 & n3421 ) ;
  assign n3423 = n3413 | n3422 ;
  assign n3424 = ( n3363 & n3406 ) | ( n3363 & n3423 ) | ( n3406 & n3423 ) ;
  assign n3425 = ( n3363 & ~n3406 ) | ( n3363 & n3423 ) | ( ~n3406 & n3423 ) ;
  assign n3426 = ( n3406 & ~n3424 ) | ( n3406 & n3425 ) | ( ~n3424 & n3425 ) ;
  assign n3427 = n3299 & n3365 ;
  assign n3428 = n3426 & n3427 ;
  assign n3429 = ~n3299 & n3365 ;
  assign n3430 = ( n3226 & ~n3298 ) | ( n3226 & n3302 ) | ( ~n3298 & n3302 ) ;
  assign n3431 = ( n3297 & ~n3298 ) | ( n3297 & n3430 ) | ( ~n3298 & n3430 ) ;
  assign n3432 = ( n3298 & ~n3365 ) | ( n3298 & n3431 ) | ( ~n3365 & n3431 ) ;
  assign n3433 = ( n2814 & n3429 ) | ( n2814 & n3432 ) | ( n3429 & n3432 ) ;
  assign n3434 = ( n3426 & n3427 ) | ( n3426 & ~n3433 ) | ( n3427 & ~n3433 ) ;
  assign n3435 = ( n3365 & n3426 ) | ( n3365 & ~n3429 ) | ( n3426 & ~n3429 ) ;
  assign n3436 = ( n3428 & n3433 ) | ( n3428 & ~n3435 ) | ( n3433 & ~n3435 ) ;
  assign n3437 = ( ~n3428 & n3434 ) | ( ~n3428 & n3436 ) | ( n3434 & n3436 ) ;
  assign n3438 = ~n3428 & n3435 ;
  assign n3439 = ( n2814 & n3433 ) | ( n2814 & n3438 ) | ( n3433 & n3438 ) ;
  assign n3440 = n1806 & ~n3045 ;
  assign n3441 = ( n1917 & ~n2831 ) | ( n1917 & n3440 ) | ( ~n2831 & n3440 ) ;
  assign n3442 = n705 | n3441 ;
  assign n3443 = ( n705 & n3441 ) | ( n705 & ~n3442 ) | ( n3441 & ~n3442 ) ;
  assign n3444 = n3442 & ~n3443 ;
  assign n3445 = ( n943 & n2132 ) | ( n943 & ~n2212 ) | ( n2132 & ~n2212 ) ;
  assign n3446 = n2132 & ~n2212 ;
  assign n3447 = ( n2282 & n2283 ) | ( n2282 & n2418 ) | ( n2283 & n2418 ) ;
  assign n3448 = ( n2322 & n2380 ) | ( n2322 & n2381 ) | ( n2380 & n2381 ) ;
  assign n3449 = n3447 | n3448 ;
  assign n3450 = ( n2324 & n2457 ) | ( n2324 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3451 = ( n2316 & ~n2462 ) | ( n2316 & n2464 ) | ( ~n2462 & n2464 ) ;
  assign n3452 = ( ~n3449 & n3450 ) | ( ~n3449 & n3451 ) | ( n3450 & n3451 ) ;
  assign n3453 = ( ~n943 & n3449 ) | ( ~n943 & n3452 ) | ( n3449 & n3452 ) ;
  assign n3454 = ( n3449 & n3452 ) | ( n3449 & ~n3453 ) | ( n3452 & ~n3453 ) ;
  assign n3455 = ( n943 & n3453 ) | ( n943 & ~n3454 ) | ( n3453 & ~n3454 ) ;
  assign n3456 = ( ~n3445 & n3446 ) | ( ~n3445 & n3455 ) | ( n3446 & n3455 ) ;
  assign n3457 = ( n3446 & n3455 ) | ( n3446 & ~n3456 ) | ( n3455 & ~n3456 ) ;
  assign n3458 = ( n3445 & n3456 ) | ( n3445 & ~n3457 ) | ( n3456 & ~n3457 ) ;
  assign n3459 = n2079 & ~n2793 ;
  assign n3460 = n2078 & ~n2790 ;
  assign n3461 = ( n2147 & n2539 ) | ( n2147 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3462 = ( n2082 & n2083 ) | ( n2082 & n2667 ) | ( n2083 & n2667 ) ;
  assign n3463 = ( ~n2083 & n3461 ) | ( ~n2083 & n3462 ) | ( n3461 & n3462 ) ;
  assign n3464 = ( ~n3459 & n3460 ) | ( ~n3459 & n3463 ) | ( n3460 & n3463 ) ;
  assign n3465 = ( ~n863 & n3459 ) | ( ~n863 & n3464 ) | ( n3459 & n3464 ) ;
  assign n3466 = ( n3459 & n3464 ) | ( n3459 & ~n3465 ) | ( n3464 & ~n3465 ) ;
  assign n3467 = ( n863 & n3465 ) | ( n863 & ~n3466 ) | ( n3465 & ~n3466 ) ;
  assign n3468 = ( n3395 & n3458 ) | ( n3395 & ~n3467 ) | ( n3458 & ~n3467 ) ;
  assign n3469 = ( ~n3395 & n3458 ) | ( ~n3395 & n3467 ) | ( n3458 & n3467 ) ;
  assign n3470 = ( ~n3458 & n3468 ) | ( ~n3458 & n3469 ) | ( n3468 & n3469 ) ;
  assign n3471 = ( n3398 & n3444 ) | ( n3398 & n3470 ) | ( n3444 & n3470 ) ;
  assign n3472 = ( n3398 & ~n3444 ) | ( n3398 & n3470 ) | ( ~n3444 & n3470 ) ;
  assign n3473 = ( n3444 & ~n3471 ) | ( n3444 & n3472 ) | ( ~n3471 & n3472 ) ;
  assign n3474 = ( n3401 & n3404 ) | ( n3401 & n3473 ) | ( n3404 & n3473 ) ;
  assign n3475 = ( n3401 & ~n3404 ) | ( n3401 & n3473 ) | ( ~n3404 & n3473 ) ;
  assign n3476 = ( n3404 & ~n3474 ) | ( n3404 & n3475 ) | ( ~n3474 & n3475 ) ;
  assign n3477 = n165 | n265 ;
  assign n3478 = ( n395 & n2357 ) | ( n395 & ~n3477 ) | ( n2357 & ~n3477 ) ;
  assign n3479 = n3477 | n3478 ;
  assign n3480 = n619 | n2526 ;
  assign n3481 = ( n85 & n237 ) | ( n85 & ~n271 ) | ( n237 & ~n271 ) ;
  assign n3482 = n509 | n602 ;
  assign n3483 = n3481 | n3482 ;
  assign n3484 = ( ~n3479 & n3480 ) | ( ~n3479 & n3483 ) | ( n3480 & n3483 ) ;
  assign n3485 = n3479 | n3484 ;
  assign n3486 = n545 | n1410 ;
  assign n3487 = ( n2682 & ~n3485 ) | ( n2682 & n3486 ) | ( ~n3485 & n3486 ) ;
  assign n3488 = n3485 | n3487 ;
  assign n3489 = ( n3424 & n3476 ) | ( n3424 & n3488 ) | ( n3476 & n3488 ) ;
  assign n3490 = ( n3424 & ~n3476 ) | ( n3424 & n3488 ) | ( ~n3476 & n3488 ) ;
  assign n3491 = ( n3476 & ~n3489 ) | ( n3476 & n3490 ) | ( ~n3489 & n3490 ) ;
  assign n3492 = ( n3428 & ~n3439 ) | ( n3428 & n3491 ) | ( ~n3439 & n3491 ) ;
  assign n3493 = ( n3428 & n3491 ) | ( n3428 & ~n3492 ) | ( n3491 & ~n3492 ) ;
  assign n3494 = ( n3439 & n3492 ) | ( n3439 & ~n3493 ) | ( n3492 & ~n3493 ) ;
  assign n3495 = n2079 & n2834 ;
  assign n3496 = n2078 & ~n2831 ;
  assign n3497 = n2147 & n2667 ;
  assign n3498 = ( n2082 & n2083 ) | ( n2082 & ~n2790 ) | ( n2083 & ~n2790 ) ;
  assign n3499 = ( ~n2083 & n3497 ) | ( ~n2083 & n3498 ) | ( n3497 & n3498 ) ;
  assign n3500 = ( ~n3495 & n3496 ) | ( ~n3495 & n3499 ) | ( n3496 & n3499 ) ;
  assign n3501 = ( ~n863 & n3495 ) | ( ~n863 & n3500 ) | ( n3495 & n3500 ) ;
  assign n3502 = ( n3495 & n3500 ) | ( n3495 & ~n3501 ) | ( n3500 & ~n3501 ) ;
  assign n3503 = ( n863 & n3501 ) | ( n863 & ~n3502 ) | ( n3501 & ~n3502 ) ;
  assign n3504 = ( n943 & n2282 ) | ( n943 & n2283 ) | ( n2282 & n2283 ) ;
  assign n3505 = ( ~n705 & n3385 ) | ( ~n705 & n3504 ) | ( n3385 & n3504 ) ;
  assign n3506 = ( n705 & n3385 ) | ( n705 & ~n3504 ) | ( n3385 & ~n3504 ) ;
  assign n3507 = ( ~n3385 & n3505 ) | ( ~n3385 & n3506 ) | ( n3505 & n3506 ) ;
  assign n3508 = ( n2380 & n2381 ) | ( n2380 & n2418 ) | ( n2381 & n2418 ) ;
  assign n3509 = ( n2322 & n2457 ) | ( n2322 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3510 = n3508 | n3509 ;
  assign n3511 = n2316 & ~n2537 ;
  assign n3512 = ( n2324 & n2539 ) | ( n2324 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3513 = ( ~n3510 & n3511 ) | ( ~n3510 & n3512 ) | ( n3511 & n3512 ) ;
  assign n3514 = ( ~n943 & n3510 ) | ( ~n943 & n3513 ) | ( n3510 & n3513 ) ;
  assign n3515 = ( n3510 & n3513 ) | ( n3510 & ~n3514 ) | ( n3513 & ~n3514 ) ;
  assign n3516 = ( n943 & n3514 ) | ( n943 & ~n3515 ) | ( n3514 & ~n3515 ) ;
  assign n3517 = ( ~n3385 & n3455 ) | ( ~n3385 & n3458 ) | ( n3455 & n3458 ) ;
  assign n3518 = ( ~n3507 & n3516 ) | ( ~n3507 & n3517 ) | ( n3516 & n3517 ) ;
  assign n3519 = ( n3507 & n3516 ) | ( n3507 & n3517 ) | ( n3516 & n3517 ) ;
  assign n3520 = ( n3507 & n3518 ) | ( n3507 & ~n3519 ) | ( n3518 & ~n3519 ) ;
  assign n3521 = ( n3468 & ~n3503 ) | ( n3468 & n3520 ) | ( ~n3503 & n3520 ) ;
  assign n3522 = ( n3468 & n3503 ) | ( n3468 & n3520 ) | ( n3503 & n3520 ) ;
  assign n3523 = ( n3503 & n3521 ) | ( n3503 & ~n3522 ) | ( n3521 & ~n3522 ) ;
  assign n3524 = ( n3471 & n3474 ) | ( n3471 & n3523 ) | ( n3474 & n3523 ) ;
  assign n3525 = ( n3471 & ~n3474 ) | ( n3471 & n3523 ) | ( ~n3474 & n3523 ) ;
  assign n3526 = ( n3474 & ~n3524 ) | ( n3474 & n3525 ) | ( ~n3524 & n3525 ) ;
  assign n3527 = n89 | n2190 ;
  assign n3528 = n172 | n339 ;
  assign n3529 = n315 | n649 ;
  assign n3530 = n3528 | n3529 ;
  assign n3531 = ( n743 & n2366 ) | ( n743 & ~n3530 ) | ( n2366 & ~n3530 ) ;
  assign n3532 = n3530 | n3531 ;
  assign n3533 = ( n2526 & ~n3527 ) | ( n2526 & n3532 ) | ( ~n3527 & n3532 ) ;
  assign n3534 = n3527 | n3533 ;
  assign n3535 = ( n292 & ~n771 ) | ( n292 & n3534 ) | ( ~n771 & n3534 ) ;
  assign n3536 = ( n771 & n2568 ) | ( n771 & ~n3535 ) | ( n2568 & ~n3535 ) ;
  assign n3537 = n3535 | n3536 ;
  assign n3538 = ( n3489 & n3526 ) | ( n3489 & n3537 ) | ( n3526 & n3537 ) ;
  assign n3539 = ( n3489 & ~n3526 ) | ( n3489 & n3537 ) | ( ~n3526 & n3537 ) ;
  assign n3540 = ( n3526 & ~n3538 ) | ( n3526 & n3539 ) | ( ~n3538 & n3539 ) ;
  assign n3541 = n3428 & n3491 ;
  assign n3542 = n3540 & n3541 ;
  assign n3543 = ~n3428 & n3491 ;
  assign n3544 = ( n3426 & n3432 ) | ( n3426 & ~n3491 ) | ( n3432 & ~n3491 ) ;
  assign n3545 = ( n3365 & ~n3491 ) | ( n3365 & n3544 ) | ( ~n3491 & n3544 ) ;
  assign n3546 = ( n2814 & n3543 ) | ( n2814 & n3545 ) | ( n3543 & n3545 ) ;
  assign n3547 = ( n3540 & n3541 ) | ( n3540 & ~n3546 ) | ( n3541 & ~n3546 ) ;
  assign n3548 = ( n3491 & n3540 ) | ( n3491 & ~n3543 ) | ( n3540 & ~n3543 ) ;
  assign n3549 = ( n3542 & n3546 ) | ( n3542 & ~n3548 ) | ( n3546 & ~n3548 ) ;
  assign n3550 = ( ~n3542 & n3547 ) | ( ~n3542 & n3549 ) | ( n3547 & n3549 ) ;
  assign n3551 = ~n3542 & n3548 ;
  assign n3552 = ( n2814 & n3546 ) | ( n2814 & n3551 ) | ( n3546 & n3551 ) ;
  assign n3553 = ( n943 & n2380 ) | ( n943 & n2381 ) | ( n2380 & n2381 ) ;
  assign n3554 = ( n2418 & n2457 ) | ( n2418 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3555 = ( n2322 & n2539 ) | ( n2322 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3556 = n3554 | n3555 ;
  assign n3557 = n2316 & n2665 ;
  assign n3558 = n2324 & n2667 ;
  assign n3559 = ( ~n3556 & n3557 ) | ( ~n3556 & n3558 ) | ( n3557 & n3558 ) ;
  assign n3560 = ( ~n943 & n3556 ) | ( ~n943 & n3559 ) | ( n3556 & n3559 ) ;
  assign n3561 = ( n3556 & n3559 ) | ( n3556 & ~n3560 ) | ( n3559 & ~n3560 ) ;
  assign n3562 = ( n943 & n3560 ) | ( n943 & ~n3561 ) | ( n3560 & ~n3561 ) ;
  assign n3563 = ( n3505 & ~n3553 ) | ( n3505 & n3562 ) | ( ~n3553 & n3562 ) ;
  assign n3564 = ( n3505 & n3553 ) | ( n3505 & n3562 ) | ( n3553 & n3562 ) ;
  assign n3565 = ( n3553 & n3563 ) | ( n3553 & ~n3564 ) | ( n3563 & ~n3564 ) ;
  assign n3566 = n2079 & n2974 ;
  assign n3567 = n2147 & ~n2790 ;
  assign n3568 = ( n2082 & n2083 ) | ( n2082 & ~n2831 ) | ( n2083 & ~n2831 ) ;
  assign n3569 = ( ~n2083 & n3567 ) | ( ~n2083 & n3568 ) | ( n3567 & n3568 ) ;
  assign n3570 = ( ~n863 & n3566 ) | ( ~n863 & n3569 ) | ( n3566 & n3569 ) ;
  assign n3571 = ( n3566 & n3569 ) | ( n3566 & ~n3570 ) | ( n3569 & ~n3570 ) ;
  assign n3572 = ( n863 & n3570 ) | ( n863 & ~n3571 ) | ( n3570 & ~n3571 ) ;
  assign n3573 = ( n3518 & ~n3565 ) | ( n3518 & n3572 ) | ( ~n3565 & n3572 ) ;
  assign n3574 = ( n3518 & n3565 ) | ( n3518 & n3572 ) | ( n3565 & n3572 ) ;
  assign n3575 = ( n3565 & n3573 ) | ( n3565 & ~n3574 ) | ( n3573 & ~n3574 ) ;
  assign n3576 = ( n3521 & ~n3524 ) | ( n3521 & n3575 ) | ( ~n3524 & n3575 ) ;
  assign n3577 = ( n3521 & n3524 ) | ( n3521 & n3575 ) | ( n3524 & n3575 ) ;
  assign n3578 = ( n3524 & n3576 ) | ( n3524 & ~n3577 ) | ( n3576 & ~n3577 ) ;
  assign n3579 = ( n204 & n343 ) | ( n204 & ~n352 ) | ( n343 & ~n352 ) ;
  assign n3580 = n156 | n354 ;
  assign n3581 = ( n140 & ~n3579 ) | ( n140 & n3580 ) | ( ~n3579 & n3580 ) ;
  assign n3582 = n3579 | n3581 ;
  assign n3583 = ( n807 & n2779 ) | ( n807 & ~n3582 ) | ( n2779 & ~n3582 ) ;
  assign n3584 = n3582 | n3583 ;
  assign n3585 = ( n3538 & n3578 ) | ( n3538 & n3584 ) | ( n3578 & n3584 ) ;
  assign n3586 = ( n3538 & ~n3578 ) | ( n3538 & n3584 ) | ( ~n3578 & n3584 ) ;
  assign n3587 = ( n3578 & ~n3585 ) | ( n3578 & n3586 ) | ( ~n3585 & n3586 ) ;
  assign n3588 = ( n3542 & ~n3552 ) | ( n3542 & n3587 ) | ( ~n3552 & n3587 ) ;
  assign n3589 = ( n3542 & n3587 ) | ( n3542 & ~n3588 ) | ( n3587 & ~n3588 ) ;
  assign n3590 = ( n3552 & n3588 ) | ( n3552 & ~n3589 ) | ( n3588 & ~n3589 ) ;
  assign n3591 = ( n943 & ~n2460 ) | ( n943 & n2461 ) | ( ~n2460 & n2461 ) ;
  assign n3592 = n3563 & ~n3591 ;
  assign n3593 = n3563 & n3591 ;
  assign n3594 = ( n3591 & n3592 ) | ( n3591 & ~n3593 ) | ( n3592 & ~n3593 ) ;
  assign n3595 = ( n2418 & n2539 ) | ( n2418 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3596 = n2322 & n2667 ;
  assign n3597 = n3595 | n3596 ;
  assign n3598 = n2316 & ~n2793 ;
  assign n3599 = n2324 & ~n2790 ;
  assign n3600 = ( ~n3597 & n3598 ) | ( ~n3597 & n3599 ) | ( n3598 & n3599 ) ;
  assign n3601 = ( ~n943 & n3597 ) | ( ~n943 & n3600 ) | ( n3597 & n3600 ) ;
  assign n3602 = ( n3597 & n3600 ) | ( n3597 & ~n3601 ) | ( n3600 & ~n3601 ) ;
  assign n3603 = ( n943 & n3601 ) | ( n943 & ~n3602 ) | ( n3601 & ~n3602 ) ;
  assign n3604 = n2079 & ~n3045 ;
  assign n3605 = ( n2147 & ~n2831 ) | ( n2147 & n3604 ) | ( ~n2831 & n3604 ) ;
  assign n3606 = n863 | n3605 ;
  assign n3607 = ( n863 & n3605 ) | ( n863 & ~n3606 ) | ( n3605 & ~n3606 ) ;
  assign n3608 = n3606 & ~n3607 ;
  assign n3609 = ( ~n3594 & n3603 ) | ( ~n3594 & n3608 ) | ( n3603 & n3608 ) ;
  assign n3610 = ( n3603 & n3608 ) | ( n3603 & ~n3609 ) | ( n3608 & ~n3609 ) ;
  assign n3611 = ( n3594 & n3609 ) | ( n3594 & ~n3610 ) | ( n3609 & ~n3610 ) ;
  assign n3612 = ( ~n3573 & n3576 ) | ( ~n3573 & n3611 ) | ( n3576 & n3611 ) ;
  assign n3613 = ( n3576 & n3611 ) | ( n3576 & ~n3612 ) | ( n3611 & ~n3612 ) ;
  assign n3614 = ( n3573 & n3612 ) | ( n3573 & ~n3613 ) | ( n3612 & ~n3613 ) ;
  assign n3615 = ( n246 & n408 ) | ( n246 & ~n1575 ) | ( n408 & ~n1575 ) ;
  assign n3616 = n1575 | n3615 ;
  assign n3617 = n470 | n2987 ;
  assign n3618 = ( n56 & n395 ) | ( n56 & n458 ) | ( n395 & n458 ) ;
  assign n3619 = n337 | n3618 ;
  assign n3620 = ( n244 & n449 ) | ( n244 & ~n3619 ) | ( n449 & ~n3619 ) ;
  assign n3621 = n3619 | n3620 ;
  assign n3622 = ( ~n3616 & n3617 ) | ( ~n3616 & n3621 ) | ( n3617 & n3621 ) ;
  assign n3623 = n3616 | n3622 ;
  assign n3624 = ( n1606 & n1965 ) | ( n1606 & ~n3623 ) | ( n1965 & ~n3623 ) ;
  assign n3625 = n3623 | n3624 ;
  assign n3626 = ( n3585 & n3614 ) | ( n3585 & n3625 ) | ( n3614 & n3625 ) ;
  assign n3627 = ( n3585 & ~n3614 ) | ( n3585 & n3625 ) | ( ~n3614 & n3625 ) ;
  assign n3628 = ( n3614 & ~n3626 ) | ( n3614 & n3627 ) | ( ~n3626 & n3627 ) ;
  assign n3629 = n3542 & n3587 ;
  assign n3630 = n3628 & n3629 ;
  assign n3631 = ~n3542 & n3587 ;
  assign n3632 = ( n3491 & ~n3541 ) | ( n3491 & n3545 ) | ( ~n3541 & n3545 ) ;
  assign n3633 = ( n3540 & ~n3541 ) | ( n3540 & n3632 ) | ( ~n3541 & n3632 ) ;
  assign n3634 = ( n3541 & ~n3587 ) | ( n3541 & n3633 ) | ( ~n3587 & n3633 ) ;
  assign n3635 = ( n2814 & n3631 ) | ( n2814 & n3634 ) | ( n3631 & n3634 ) ;
  assign n3636 = ( n3628 & n3629 ) | ( n3628 & ~n3635 ) | ( n3629 & ~n3635 ) ;
  assign n3637 = ( n3587 & n3628 ) | ( n3587 & ~n3631 ) | ( n3628 & ~n3631 ) ;
  assign n3638 = ( n3630 & n3635 ) | ( n3630 & ~n3637 ) | ( n3635 & ~n3637 ) ;
  assign n3639 = ( ~n3630 & n3636 ) | ( ~n3630 & n3638 ) | ( n3636 & n3638 ) ;
  assign n3640 = ~n3630 & n3637 ;
  assign n3641 = ( n2814 & n3635 ) | ( n2814 & n3640 ) | ( n3635 & n3640 ) ;
  assign n3642 = ( n943 & n2457 ) | ( n943 & ~n2458 ) | ( n2457 & ~n2458 ) ;
  assign n3643 = ( n943 & n2539 ) | ( n943 & n2540 ) | ( n2539 & n2540 ) ;
  assign n3644 = ( ~n863 & n3642 ) | ( ~n863 & n3643 ) | ( n3642 & n3643 ) ;
  assign n3645 = ( n3642 & n3643 ) | ( n3642 & ~n3644 ) | ( n3643 & ~n3644 ) ;
  assign n3646 = ( n863 & n3644 ) | ( n863 & ~n3645 ) | ( n3644 & ~n3645 ) ;
  assign n3647 = n2418 & n2667 ;
  assign n3648 = n2322 & ~n2790 ;
  assign n3649 = n3647 | n3648 ;
  assign n3650 = n2316 & n2834 ;
  assign n3651 = n2324 & ~n2831 ;
  assign n3652 = ( ~n3649 & n3650 ) | ( ~n3649 & n3651 ) | ( n3650 & n3651 ) ;
  assign n3653 = ( ~n943 & n3649 ) | ( ~n943 & n3652 ) | ( n3649 & n3652 ) ;
  assign n3654 = ( n3649 & n3652 ) | ( n3649 & ~n3653 ) | ( n3652 & ~n3653 ) ;
  assign n3655 = ( n943 & n3653 ) | ( n943 & ~n3654 ) | ( n3653 & ~n3654 ) ;
  assign n3656 = ( n2523 & n3562 ) | ( n2523 & n3594 ) | ( n3562 & n3594 ) ;
  assign n3657 = ( ~n3646 & n3655 ) | ( ~n3646 & n3656 ) | ( n3655 & n3656 ) ;
  assign n3658 = ( n3646 & n3655 ) | ( n3646 & n3656 ) | ( n3655 & n3656 ) ;
  assign n3659 = ( n3646 & n3657 ) | ( n3646 & ~n3658 ) | ( n3657 & ~n3658 ) ;
  assign n3660 = ( ~n3609 & n3612 ) | ( ~n3609 & n3659 ) | ( n3612 & n3659 ) ;
  assign n3661 = ( n3612 & n3659 ) | ( n3612 & ~n3660 ) | ( n3659 & ~n3660 ) ;
  assign n3662 = ( n3609 & n3660 ) | ( n3609 & ~n3661 ) | ( n3660 & ~n3661 ) ;
  assign n3663 = n286 | n312 ;
  assign n3664 = ( n56 & n106 ) | ( n56 & n154 ) | ( n106 & n154 ) ;
  assign n3665 = ( n104 & n115 ) | ( n104 & n202 ) | ( n115 & n202 ) ;
  assign n3666 = ( n428 & ~n3664 ) | ( n428 & n3665 ) | ( ~n3664 & n3665 ) ;
  assign n3667 = n3664 | n3666 ;
  assign n3668 = ( n112 & ~n352 ) | ( n112 & n670 ) | ( ~n352 & n670 ) ;
  assign n3669 = n352 | n3668 ;
  assign n3670 = ( n3663 & ~n3667 ) | ( n3663 & n3669 ) | ( ~n3667 & n3669 ) ;
  assign n3671 = n2903 | n3667 ;
  assign n3672 = ( ~n128 & n305 ) | ( ~n128 & n341 ) | ( n305 & n341 ) ;
  assign n3673 = ( n128 & ~n2903 ) | ( n128 & n3672 ) | ( ~n2903 & n3672 ) ;
  assign n3674 = ( ~n3670 & n3671 ) | ( ~n3670 & n3673 ) | ( n3671 & n3673 ) ;
  assign n3675 = n2592 | n3670 ;
  assign n3676 = ( n263 & n2118 ) | ( n263 & ~n2592 ) | ( n2118 & ~n2592 ) ;
  assign n3677 = ( ~n3674 & n3675 ) | ( ~n3674 & n3676 ) | ( n3675 & n3676 ) ;
  assign n3678 = n3674 | n3677 ;
  assign n3679 = ( n3626 & n3662 ) | ( n3626 & n3678 ) | ( n3662 & n3678 ) ;
  assign n3680 = ( n3626 & ~n3662 ) | ( n3626 & n3678 ) | ( ~n3662 & n3678 ) ;
  assign n3681 = ( n3662 & ~n3679 ) | ( n3662 & n3680 ) | ( ~n3679 & n3680 ) ;
  assign n3682 = ( n3630 & ~n3641 ) | ( n3630 & n3681 ) | ( ~n3641 & n3681 ) ;
  assign n3683 = ( n3630 & n3681 ) | ( n3630 & ~n3682 ) | ( n3681 & ~n3682 ) ;
  assign n3684 = ( n3641 & n3682 ) | ( n3641 & ~n3683 ) | ( n3682 & ~n3683 ) ;
  assign n3685 = n943 & n2667 ;
  assign n3686 = n2418 & ~n2790 ;
  assign n3687 = n2316 & n2974 ;
  assign n3688 = n2322 & ~n2831 ;
  assign n3689 = ( ~n3686 & n3687 ) | ( ~n3686 & n3688 ) | ( n3687 & n3688 ) ;
  assign n3690 = ( ~n943 & n3686 ) | ( ~n943 & n3689 ) | ( n3686 & n3689 ) ;
  assign n3691 = ( n3686 & n3689 ) | ( n3686 & ~n3690 ) | ( n3689 & ~n3690 ) ;
  assign n3692 = ( n943 & n3690 ) | ( n943 & ~n3691 ) | ( n3690 & ~n3691 ) ;
  assign n3693 = ( n3644 & ~n3685 ) | ( n3644 & n3692 ) | ( ~n3685 & n3692 ) ;
  assign n3694 = ( n3644 & n3685 ) | ( n3644 & n3692 ) | ( n3685 & n3692 ) ;
  assign n3695 = ( n3685 & n3693 ) | ( n3685 & ~n3694 ) | ( n3693 & ~n3694 ) ;
  assign n3696 = ( ~n3657 & n3660 ) | ( ~n3657 & n3695 ) | ( n3660 & n3695 ) ;
  assign n3697 = ( n3660 & n3695 ) | ( n3660 & ~n3696 ) | ( n3695 & ~n3696 ) ;
  assign n3698 = ( n3657 & n3696 ) | ( n3657 & ~n3697 ) | ( n3696 & ~n3697 ) ;
  assign n3699 = n1575 | n2526 ;
  assign n3700 = n356 | n410 ;
  assign n3701 = n328 | n611 ;
  assign n3702 = n796 | n3701 ;
  assign n3703 = ( n128 & ~n3700 ) | ( n128 & n3702 ) | ( ~n3700 & n3702 ) ;
  assign n3704 = n3700 | n3703 ;
  assign n3705 = n167 | n1417 ;
  assign n3706 = ( ~n3699 & n3704 ) | ( ~n3699 & n3705 ) | ( n3704 & n3705 ) ;
  assign n3707 = n3699 | n3706 ;
  assign n3708 = ( n288 & ~n856 ) | ( n288 & n3707 ) | ( ~n856 & n3707 ) ;
  assign n3709 = n741 | n3708 ;
  assign n3710 = ( n856 & n1236 ) | ( n856 & ~n3709 ) | ( n1236 & ~n3709 ) ;
  assign n3711 = n3709 | n3710 ;
  assign n3712 = ( n3679 & n3698 ) | ( n3679 & n3711 ) | ( n3698 & n3711 ) ;
  assign n3713 = ( n3679 & ~n3698 ) | ( n3679 & n3711 ) | ( ~n3698 & n3711 ) ;
  assign n3714 = ( n3698 & ~n3712 ) | ( n3698 & n3713 ) | ( ~n3712 & n3713 ) ;
  assign n3715 = n3630 & n3681 ;
  assign n3716 = n3714 & n3715 ;
  assign n3717 = ~n3630 & n3681 ;
  assign n3718 = ( n3587 & ~n3629 ) | ( n3587 & n3634 ) | ( ~n3629 & n3634 ) ;
  assign n3719 = ( n3628 & ~n3629 ) | ( n3628 & n3718 ) | ( ~n3629 & n3718 ) ;
  assign n3720 = ( n3629 & ~n3681 ) | ( n3629 & n3719 ) | ( ~n3681 & n3719 ) ;
  assign n3721 = ( n2814 & n3717 ) | ( n2814 & n3720 ) | ( n3717 & n3720 ) ;
  assign n3722 = ( n3714 & n3715 ) | ( n3714 & ~n3721 ) | ( n3715 & ~n3721 ) ;
  assign n3723 = ( n3681 & n3714 ) | ( n3681 & ~n3717 ) | ( n3714 & ~n3717 ) ;
  assign n3724 = ( n3716 & n3721 ) | ( n3716 & ~n3723 ) | ( n3721 & ~n3723 ) ;
  assign n3725 = ( ~n3716 & n3722 ) | ( ~n3716 & n3724 ) | ( n3722 & n3724 ) ;
  assign n3726 = ~n3716 & n3723 ;
  assign n3727 = ( n2814 & n3721 ) | ( n2814 & n3726 ) | ( n3721 & n3726 ) ;
  assign n3728 = n2316 & ~n3045 ;
  assign n3729 = ( n2418 & ~n2831 ) | ( n2418 & n3728 ) | ( ~n2831 & n3728 ) ;
  assign n3730 = ~n2667 & n2790 ;
  assign n3731 = n2667 & ~n2790 ;
  assign n3732 = ( n943 & n3730 ) | ( n943 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3733 = n3729 | n3732 ;
  assign n3734 = ( n3729 & n3732 ) | ( n3729 & ~n3733 ) | ( n3732 & ~n3733 ) ;
  assign n3735 = n3733 & ~n3734 ;
  assign n3736 = ( ~n3693 & n3696 ) | ( ~n3693 & n3735 ) | ( n3696 & n3735 ) ;
  assign n3737 = ( n3696 & n3735 ) | ( n3696 & ~n3736 ) | ( n3735 & ~n3736 ) ;
  assign n3738 = ( n3693 & n3736 ) | ( n3693 & ~n3737 ) | ( n3736 & ~n3737 ) ;
  assign n3739 = ( n80 & n126 ) | ( n80 & n206 ) | ( n126 & n206 ) ;
  assign n3740 = n520 | n3739 ;
  assign n3741 = n336 | n3740 ;
  assign n3742 = n1584 | n1685 ;
  assign n3743 = n726 | n2562 ;
  assign n3744 = ( ~n56 & n165 ) | ( ~n56 & n237 ) | ( n165 & n237 ) ;
  assign n3745 = ( n565 & n610 ) | ( n565 & ~n3744 ) | ( n610 & ~n3744 ) ;
  assign n3746 = n3744 | n3745 ;
  assign n3747 = n302 | n3621 ;
  assign n3748 = n3746 | n3747 ;
  assign n3749 = ( ~n1685 & n3743 ) | ( ~n1685 & n3748 ) | ( n3743 & n3748 ) ;
  assign n3750 = ( ~n3741 & n3742 ) | ( ~n3741 & n3749 ) | ( n3742 & n3749 ) ;
  assign n3751 = n3741 | n3750 ;
  assign n3752 = ( n3712 & n3738 ) | ( n3712 & n3751 ) | ( n3738 & n3751 ) ;
  assign n3753 = ( n3712 & ~n3738 ) | ( n3712 & n3751 ) | ( ~n3738 & n3751 ) ;
  assign n3754 = ( n3738 & ~n3752 ) | ( n3738 & n3753 ) | ( ~n3752 & n3753 ) ;
  assign n3755 = ( n3716 & ~n3727 ) | ( n3716 & n3754 ) | ( ~n3727 & n3754 ) ;
  assign n3756 = ( n3716 & n3754 ) | ( n3716 & ~n3755 ) | ( n3754 & ~n3755 ) ;
  assign n3757 = ( n3727 & n3755 ) | ( n3727 & ~n3756 ) | ( n3755 & ~n3756 ) ;
  assign n3758 = n3716 & n3754 ;
  assign n3759 = ~n3716 & n3754 ;
  assign n3760 = ( n3681 & ~n3715 ) | ( n3681 & n3720 ) | ( ~n3715 & n3720 ) ;
  assign n3761 = ( n3714 & ~n3715 ) | ( n3714 & n3760 ) | ( ~n3715 & n3760 ) ;
  assign n3762 = ( n3715 & ~n3754 ) | ( n3715 & n3761 ) | ( ~n3754 & n3761 ) ;
  assign n3763 = ( n2814 & n3759 ) | ( n2814 & n3762 ) | ( n3759 & n3762 ) ;
  assign n3764 = n1749 | n2587 ;
  assign n3765 = n171 | n411 ;
  assign n3766 = ( n331 & ~n468 ) | ( n331 & n765 ) | ( ~n468 & n765 ) ;
  assign n3767 = n468 | n3766 ;
  assign n3768 = ( n1883 & ~n3765 ) | ( n1883 & n3767 ) | ( ~n3765 & n3767 ) ;
  assign n3769 = n3765 | n3768 ;
  assign n3770 = ( ~n2587 & n3667 ) | ( ~n2587 & n3769 ) | ( n3667 & n3769 ) ;
  assign n3771 = ( ~n2697 & n3764 ) | ( ~n2697 & n3770 ) | ( n3764 & n3770 ) ;
  assign n3772 = n2697 | n3771 ;
  assign n3773 = ~n2667 & n2831 ;
  assign n3774 = n2667 & ~n2831 ;
  assign n3775 = ( n943 & n3773 ) | ( n943 & n3774 ) | ( n3773 & n3774 ) ;
  assign n3776 = n943 | n3729 ;
  assign n3777 = ( ~n3729 & n3730 ) | ( ~n3729 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3778 = n2667 | n2790 ;
  assign n3779 = ( n943 & n3777 ) | ( n943 & ~n3778 ) | ( n3777 & ~n3778 ) ;
  assign n3780 = ( ~n943 & n3776 ) | ( ~n943 & n3779 ) | ( n3776 & n3779 ) ;
  assign n3781 = ( ~n3736 & n3775 ) | ( ~n3736 & n3780 ) | ( n3775 & n3780 ) ;
  assign n3782 = ( n3775 & n3780 ) | ( n3775 & ~n3781 ) | ( n3780 & ~n3781 ) ;
  assign n3783 = ( n3736 & n3781 ) | ( n3736 & ~n3782 ) | ( n3781 & ~n3782 ) ;
  assign n3784 = ( n3752 & n3772 ) | ( n3752 & n3783 ) | ( n3772 & n3783 ) ;
  assign n3785 = ( n3752 & ~n3772 ) | ( n3752 & n3783 ) | ( ~n3772 & n3783 ) ;
  assign n3786 = ( n3772 & ~n3784 ) | ( n3772 & n3785 ) | ( ~n3784 & n3785 ) ;
  assign n3787 = ( ~n3758 & n3763 ) | ( ~n3758 & n3786 ) | ( n3763 & n3786 ) ;
  assign n3788 = ( n3763 & n3786 ) | ( n3763 & ~n3787 ) | ( n3786 & ~n3787 ) ;
  assign n3789 = ( n3758 & n3787 ) | ( n3758 & ~n3788 ) | ( n3787 & ~n3788 ) ;
  assign n3790 = n3754 | n3786 ;
  assign n3791 = n3716 & n3786 ;
  assign n3792 = ( n3762 & n3790 ) | ( n3762 & ~n3791 ) | ( n3790 & ~n3791 ) ;
  assign n3793 = ( x22 & x23 ) | ( x22 & ~n3792 ) | ( x23 & ~n3792 ) ;
  assign n3794 = n3758 & n3786 ;
  assign n3795 = n137 | n184 ;
  assign n3796 = ( n458 & n524 ) | ( n458 & ~n3795 ) | ( n524 & ~n3795 ) ;
  assign n3797 = n3795 | n3796 ;
  assign n3798 = n286 | n2190 ;
  assign n3799 = ( n364 & n436 ) | ( n364 & ~n502 ) | ( n436 & ~n502 ) ;
  assign n3800 = n502 | n3799 ;
  assign n3801 = ( ~n3797 & n3798 ) | ( ~n3797 & n3800 ) | ( n3798 & n3800 ) ;
  assign n3802 = n3797 | n3801 ;
  assign n3803 = ( n646 & ~n672 ) | ( n646 & n2364 ) | ( ~n672 & n2364 ) ;
  assign n3804 = ( n672 & ~n3802 ) | ( n672 & n3803 ) | ( ~n3802 & n3803 ) ;
  assign n3805 = n3802 | n3804 ;
  assign n3806 = n3784 & n3805 ;
  assign n3807 = n3784 | n3805 ;
  assign n3808 = ( n3794 & ~n3806 ) | ( n3794 & n3807 ) | ( ~n3806 & n3807 ) ;
  assign n3809 = n3794 & n3805 ;
  assign n3810 = n3808 & ~n3809 ;
  assign n3811 = ( ~n2812 & n3793 ) | ( ~n2812 & n3810 ) | ( n3793 & n3810 ) ;
  assign n3812 = ( n3793 & n3810 ) | ( n3793 & ~n3811 ) | ( n3810 & ~n3811 ) ;
  assign n3813 = ( n2812 & n3811 ) | ( n2812 & ~n3812 ) | ( n3811 & ~n3812 ) ;
  assign n3814 = ( n3792 & n3808 ) | ( n3792 & ~n3809 ) | ( n3808 & ~n3809 ) ;
  assign n3815 = n217 | n717 ;
  assign n3816 = n228 | n410 ;
  assign n3817 = ( ~n717 & n785 ) | ( ~n717 & n3816 ) | ( n785 & n3816 ) ;
  assign n3818 = ( ~n217 & n351 ) | ( ~n217 & n2113 ) | ( n351 & n2113 ) ;
  assign n3819 = ( n3815 & ~n3817 ) | ( n3815 & n3818 ) | ( ~n3817 & n3818 ) ;
  assign n3820 = ( n380 & n458 ) | ( n380 & ~n569 ) | ( n458 & ~n569 ) ;
  assign n3821 = n569 | n3820 ;
  assign n3822 = ( n3817 & ~n3819 ) | ( n3817 & n3821 ) | ( ~n3819 & n3821 ) ;
  assign n3823 = n3819 | n3822 ;
  assign n3824 = ( n681 & n2578 ) | ( n681 & ~n3823 ) | ( n2578 & ~n3823 ) ;
  assign n3825 = n3823 | n3824 ;
  assign n3826 = ( ~n3806 & n3809 ) | ( ~n3806 & n3825 ) | ( n3809 & n3825 ) ;
  assign n3827 = ( n3809 & n3825 ) | ( n3809 & ~n3826 ) | ( n3825 & ~n3826 ) ;
  assign n3828 = ( n3806 & n3826 ) | ( n3806 & ~n3827 ) | ( n3826 & ~n3827 ) ;
  assign n3829 = n3814 | n3828 ;
  assign n3830 = ( n2814 & n3814 ) | ( n2814 & ~n3828 ) | ( n3814 & ~n3828 ) ;
  assign n3831 = n2814 & ~n3828 ;
  assign n3832 = ( n3829 & ~n3830 ) | ( n3829 & n3831 ) | ( ~n3830 & n3831 ) ;
  assign n3833 = n3809 & n3825 ;
  assign n3834 = n3806 & n3825 ;
  assign n3835 = n207 | n800 ;
  assign n3836 = ( n134 & n206 ) | ( n134 & n378 ) | ( n206 & n378 ) ;
  assign n3837 = ( n57 & n80 ) | ( n57 & n126 ) | ( n80 & n126 ) ;
  assign n3838 = ( n765 & ~n3836 ) | ( n765 & n3837 ) | ( ~n3836 & n3837 ) ;
  assign n3839 = ( n142 & n3836 ) | ( n142 & ~n3838 ) | ( n3836 & ~n3838 ) ;
  assign n3840 = n3838 | n3839 ;
  assign n3841 = ( n3213 & n3835 ) | ( n3213 & ~n3840 ) | ( n3835 & ~n3840 ) ;
  assign n3842 = ( n2271 & n3840 ) | ( n2271 & ~n3841 ) | ( n3840 & ~n3841 ) ;
  assign n3843 = n3841 | n3842 ;
  assign n3844 = n415 | n3741 ;
  assign n3845 = n3843 | n3844 ;
  assign n3846 = ( ~n3833 & n3834 ) | ( ~n3833 & n3845 ) | ( n3834 & n3845 ) ;
  assign n3847 = ( n3834 & n3845 ) | ( n3834 & ~n3846 ) | ( n3845 & ~n3846 ) ;
  assign n3848 = ( n3833 & n3846 ) | ( n3833 & ~n3847 ) | ( n3846 & ~n3847 ) ;
  assign n3849 = n3829 | n3848 ;
  assign n3850 = ( n2814 & n3829 ) | ( n2814 & ~n3848 ) | ( n3829 & ~n3848 ) ;
  assign n3851 = n2814 & ~n3848 ;
  assign n3852 = ( n3849 & ~n3850 ) | ( n3849 & n3851 ) | ( ~n3850 & n3851 ) ;
  assign n3853 = n3833 & n3845 ;
  assign n3854 = n3834 & n3845 ;
  assign n3855 = n145 | n2693 ;
  assign n3856 = n3357 | n3855 ;
  assign n3857 = ( n229 & ~n887 ) | ( n229 & n3211 ) | ( ~n887 & n3211 ) ;
  assign n3858 = n887 | n3857 ;
  assign n3859 = ( n158 & ~n3856 ) | ( n158 & n3858 ) | ( ~n3856 & n3858 ) ;
  assign n3860 = n3856 | n3859 ;
  assign n3861 = ( n723 & n3413 ) | ( n723 & ~n3860 ) | ( n3413 & ~n3860 ) ;
  assign n3862 = n3860 | n3861 ;
  assign n3863 = ( ~n3853 & n3854 ) | ( ~n3853 & n3862 ) | ( n3854 & n3862 ) ;
  assign n3864 = ( n3854 & n3862 ) | ( n3854 & ~n3863 ) | ( n3862 & ~n3863 ) ;
  assign n3865 = ( n3853 & n3863 ) | ( n3853 & ~n3864 ) | ( n3863 & ~n3864 ) ;
  assign n3866 = n3849 | n3865 ;
  assign n3867 = ( n2814 & n3849 ) | ( n2814 & ~n3865 ) | ( n3849 & ~n3865 ) ;
  assign n3868 = n2814 & ~n3865 ;
  assign n3869 = ( n3866 & ~n3867 ) | ( n3866 & n3868 ) | ( ~n3867 & n3868 ) ;
  assign n3870 = n2814 & n3866 ;
  assign n3871 = n3854 & n3862 ;
  assign n3872 = n106 | n2656 ;
  assign n3873 = ( n183 & n918 ) | ( n183 & ~n3872 ) | ( n918 & ~n3872 ) ;
  assign n3874 = n3872 | n3873 ;
  assign n3875 = ( n3853 & n3871 ) | ( n3853 & n3874 ) | ( n3871 & n3874 ) ;
  assign n3876 = ( ~n3853 & n3871 ) | ( ~n3853 & n3874 ) | ( n3871 & n3874 ) ;
  assign n3877 = ( n3853 & ~n3875 ) | ( n3853 & n3876 ) | ( ~n3875 & n3876 ) ;
  assign n3878 = n3870 | n3877 ;
  assign n3879 = ( n3870 & n3877 ) | ( n3870 & ~n3878 ) | ( n3877 & ~n3878 ) ;
  assign n3880 = n3878 & ~n3879 ;
  assign n3881 = ( n2814 & n3870 ) | ( n2814 & n3877 ) | ( n3870 & n3877 ) ;
  assign n3882 = n160 | n918 ;
  assign n3883 = ( ~n3875 & n3881 ) | ( ~n3875 & n3882 ) | ( n3881 & n3882 ) ;
  assign n3884 = ( n3881 & n3882 ) | ( n3881 & ~n3883 ) | ( n3882 & ~n3883 ) ;
  assign n3885 = ( n3875 & n3883 ) | ( n3875 & ~n3884 ) | ( n3883 & ~n3884 ) ;
  assign n3886 = n3875 & n3882 ;
  assign n3887 = x22 | n45 ;
  assign n3888 = ( n3881 & ~n3886 ) | ( n3881 & n3887 ) | ( ~n3886 & n3887 ) ;
  assign n3889 = n3875 | n3882 ;
  assign n3890 = ( n2814 & n3881 ) | ( n2814 & n3889 ) | ( n3881 & n3889 ) ;
  assign n3891 = n3886 | n3890 ;
  assign n3892 = ( n3886 & n3888 ) | ( n3886 & ~n3891 ) | ( n3888 & ~n3891 ) ;
  assign n3893 = ( n2814 & n3870 ) | ( n2814 & ~n3892 ) | ( n3870 & ~n3892 ) ;
  assign y0 = n2811 ;
  assign y1 = n2919 ;
  assign y2 = n3003 ;
  assign y3 = n3085 ;
  assign y4 = n3159 ;
  assign y5 = n3230 ;
  assign y6 = n3307 ;
  assign y7 = n3368 ;
  assign y8 = n3437 ;
  assign y9 = n3494 ;
  assign y10 = n3550 ;
  assign y11 = n3590 ;
  assign y12 = n3639 ;
  assign y13 = n3684 ;
  assign y14 = n3725 ;
  assign y15 = n3757 ;
  assign y16 = n3789 ;
  assign y17 = n3813 ;
  assign y18 = n3832 ;
  assign y19 = n3852 ;
  assign y20 = n3869 ;
  assign y21 = n3880 ;
  assign y22 = n3885 ;
  assign y23 = ~n3892 ;
  assign y24 = n3893 ;
endmodule
