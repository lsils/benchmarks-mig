module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , x544 , x545 , x546 , x547 , x548 , x549 , x550 , x551 , x552 , x553 , x554 , x555 , x556 , x557 , x558 , x559 , x560 , x561 , x562 , x563 , x564 , x565 , x566 , x567 , x568 , x569 , x570 , x571 , x572 , x573 , x574 , x575 , x576 , x577 , x578 , x579 , x580 , x581 , x582 , x583 , x584 , x585 , x586 , x587 , x588 , x589 , x590 , x591 , x592 , x593 , x594 , x595 , x596 , x597 , x598 , x599 , x600 , x601 , x602 , x603 , x604 , x605 , x606 , x607 , x608 , x609 , x610 , x611 , x612 , x613 , x614 , x615 , x616 , x617 , x618 , x619 , x620 , x621 , x622 , x623 , x624 , x625 , x626 , x627 , x628 , x629 , x630 , x631 , x632 , x633 , x634 , x635 , x636 , x637 , x638 , x639 , x640 , x641 , x642 , x643 , x644 , x645 , x646 , x647 , x648 , x649 , x650 , x651 , x652 , x653 , x654 , x655 , x656 , x657 , x658 , x659 , x660 , x661 , x662 , x663 , x664 , x665 , x666 , x667 , x668 , x669 , x670 , x671 , x672 , x673 , x674 , x675 , x676 , x677 , x678 , x679 , x680 , x681 , x682 , x683 , x684 , x685 , x686 , x687 , x688 , x689 , x690 , x691 , x692 , x693 , x694 , x695 , x696 , x697 , x698 , x699 , x700 , x701 , x702 , x703 , x704 , x705 , x706 , x707 , x708 , x709 , x710 , x711 , x712 , x713 , x714 , x715 , x716 , x717 , x718 , x719 , x720 , x721 , x722 , x723 , x724 , x725 , x726 , x727 , x728 , x729 , x730 , x731 , x732 , x733 , x734 , x735 , x736 , x737 , x738 , x739 , x740 , x741 , x742 , x743 , x744 , x745 , x746 , x747 , x748 , x749 , x750 , x751 , x752 , x753 , x754 , x755 , x756 , x757 , x758 , x759 , x760 , x761 , x762 , x763 , x764 , x765 , x766 , x767 , x768 , x769 , x770 , x771 , x772 , x773 , x774 , x775 , x776 , x777 , x778 , x779 , x780 , x781 , x782 , x783 , x784 , x785 , x786 , x787 , x788 , x789 , x790 , x791 , x792 , x793 , x794 , x795 , x796 , x797 , x798 , x799 , x800 , x801 , x802 , x803 , x804 , x805 , x806 , x807 , x808 , x809 , x810 , x811 , x812 , x813 , x814 , x815 , x816 , x817 , x818 , x819 , x820 , x821 , x822 , x823 , x824 , x825 , x826 , x827 , x828 , x829 , x830 , x831 , x832 , x833 , x834 , x835 , x836 , x837 , x838 , x839 , x840 , x841 , x842 , x843 , x844 , x845 , x846 , x847 , x848 , x849 , x850 , x851 , x852 , x853 , x854 , x855 , x856 , x857 , x858 , x859 , x860 , x861 , x862 , x863 , x864 , x865 , x866 , x867 , x868 , x869 , x870 , x871 , x872 , x873 , x874 , x875 , x876 , x877 , x878 , x879 , x880 , x881 , x882 , x883 , x884 , x885 , x886 , x887 , x888 , x889 , x890 , x891 , x892 , x893 , x894 , x895 , x896 , x897 , x898 , x899 , x900 , x901 , x902 , x903 , x904 , x905 , x906 , x907 , x908 , x909 , x910 , x911 , x912 , x913 , x914 , x915 , x916 , x917 , x918 , x919 , x920 , x921 , x922 , x923 , x924 , x925 , x926 , x927 , x928 , x929 , x930 , x931 , x932 , x933 , x934 , x935 , x936 , x937 , x938 , x939 , x940 , x941 , x942 , x943 , x944 , x945 , x946 , x947 , x948 , x949 , x950 , x951 , x952 , x953 , x954 , x955 , x956 , x957 , x958 , x959 , x960 , x961 , x962 , x963 , x964 , x965 , x966 , x967 , x968 , x969 , x970 , x971 , x972 , x973 , x974 , x975 , x976 , x977 , x978 , x979 , x980 , x981 , x982 , x983 , x984 , x985 , x986 , x987 , x988 , x989 , x990 , x991 , x992 , x993 , x994 , x995 , x996 , x997 , x998 , x999 , x1000 ;
  output y0 ;
  wire n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 ;
  assign n1002 = ( x460 & x461 ) | ( x460 & x462 ) | ( x461 & x462 ) ;
  assign n1003 = ( x457 & x458 ) | ( x457 & x459 ) | ( x458 & x459 ) ;
  assign n1004 = ( ~x460 & x461 ) | ( ~x460 & x462 ) | ( x461 & x462 ) ;
  assign n1005 = ( x460 & ~n1002 ) | ( x460 & n1004 ) | ( ~n1002 & n1004 ) ;
  assign n1006 = ( ~x457 & x458 ) | ( ~x457 & x459 ) | ( x458 & x459 ) ;
  assign n1007 = ( x457 & ~n1003 ) | ( x457 & n1006 ) | ( ~n1003 & n1006 ) ;
  assign n1008 = n1005 & n1007 ;
  assign n1009 = ( n1002 & n1003 ) | ( n1002 & n1008 ) | ( n1003 & n1008 ) ;
  assign n1010 = ( x451 & x452 ) | ( x451 & x453 ) | ( x452 & x453 ) ;
  assign n1011 = ( x454 & x455 ) | ( x454 & x456 ) | ( x455 & x456 ) ;
  assign n1012 = ( ~x454 & x455 ) | ( ~x454 & x456 ) | ( x455 & x456 ) ;
  assign n1013 = ( x454 & ~n1011 ) | ( x454 & n1012 ) | ( ~n1011 & n1012 ) ;
  assign n1014 = ( ~x451 & x452 ) | ( ~x451 & x453 ) | ( x452 & x453 ) ;
  assign n1015 = ( x451 & ~n1010 ) | ( x451 & n1014 ) | ( ~n1010 & n1014 ) ;
  assign n1016 = n1013 & n1015 ;
  assign n1017 = ( n1010 & n1011 ) | ( n1010 & n1016 ) | ( n1011 & n1016 ) ;
  assign n1018 = ( ~n1002 & n1003 ) | ( ~n1002 & n1008 ) | ( n1003 & n1008 ) ;
  assign n1019 = ( n1002 & ~n1009 ) | ( n1002 & n1018 ) | ( ~n1009 & n1018 ) ;
  assign n1020 = ( ~n1010 & n1011 ) | ( ~n1010 & n1016 ) | ( n1011 & n1016 ) ;
  assign n1021 = ( n1010 & ~n1017 ) | ( n1010 & n1020 ) | ( ~n1017 & n1020 ) ;
  assign n1022 = n1005 | n1007 ;
  assign n1023 = ~n1008 & n1022 ;
  assign n1024 = n1013 | n1015 ;
  assign n1025 = ~n1016 & n1024 ;
  assign n1026 = n1023 & n1025 ;
  assign n1027 = ( n1019 & n1021 ) | ( n1019 & n1026 ) | ( n1021 & n1026 ) ;
  assign n1028 = ( n1009 & n1017 ) | ( n1009 & n1027 ) | ( n1017 & n1027 ) ;
  assign n1029 = ( x448 & x449 ) | ( x448 & x450 ) | ( x449 & x450 ) ;
  assign n1030 = ( x445 & x446 ) | ( x445 & x447 ) | ( x446 & x447 ) ;
  assign n1031 = ( ~x448 & x449 ) | ( ~x448 & x450 ) | ( x449 & x450 ) ;
  assign n1032 = ( x448 & ~n1029 ) | ( x448 & n1031 ) | ( ~n1029 & n1031 ) ;
  assign n1033 = ( ~x445 & x446 ) | ( ~x445 & x447 ) | ( x446 & x447 ) ;
  assign n1034 = ( x445 & ~n1030 ) | ( x445 & n1033 ) | ( ~n1030 & n1033 ) ;
  assign n1035 = n1032 & n1034 ;
  assign n1036 = ( n1029 & n1030 ) | ( n1029 & n1035 ) | ( n1030 & n1035 ) ;
  assign n1037 = ( x439 & x440 ) | ( x439 & x441 ) | ( x440 & x441 ) ;
  assign n1038 = ( x442 & x443 ) | ( x442 & x444 ) | ( x443 & x444 ) ;
  assign n1039 = ( ~x442 & x443 ) | ( ~x442 & x444 ) | ( x443 & x444 ) ;
  assign n1040 = ( x442 & ~n1038 ) | ( x442 & n1039 ) | ( ~n1038 & n1039 ) ;
  assign n1041 = ( ~x439 & x440 ) | ( ~x439 & x441 ) | ( x440 & x441 ) ;
  assign n1042 = ( x439 & ~n1037 ) | ( x439 & n1041 ) | ( ~n1037 & n1041 ) ;
  assign n1043 = n1040 & n1042 ;
  assign n1044 = ( n1037 & n1038 ) | ( n1037 & n1043 ) | ( n1038 & n1043 ) ;
  assign n1045 = ( ~n1029 & n1030 ) | ( ~n1029 & n1035 ) | ( n1030 & n1035 ) ;
  assign n1046 = ( n1029 & ~n1036 ) | ( n1029 & n1045 ) | ( ~n1036 & n1045 ) ;
  assign n1047 = ( ~n1037 & n1038 ) | ( ~n1037 & n1043 ) | ( n1038 & n1043 ) ;
  assign n1048 = ( n1037 & ~n1044 ) | ( n1037 & n1047 ) | ( ~n1044 & n1047 ) ;
  assign n1049 = n1040 | n1042 ;
  assign n1050 = ~n1043 & n1049 ;
  assign n1051 = ( n1032 & n1034 ) | ( n1032 & n1050 ) | ( n1034 & n1050 ) ;
  assign n1052 = ~n1035 & n1051 ;
  assign n1053 = ( n1046 & n1048 ) | ( n1046 & n1052 ) | ( n1048 & n1052 ) ;
  assign n1054 = ( n1036 & n1044 ) | ( n1036 & n1053 ) | ( n1044 & n1053 ) ;
  assign n1055 = ( ~n1036 & n1044 ) | ( ~n1036 & n1053 ) | ( n1044 & n1053 ) ;
  assign n1056 = ( n1036 & ~n1054 ) | ( n1036 & n1055 ) | ( ~n1054 & n1055 ) ;
  assign n1057 = ( ~n1009 & n1017 ) | ( ~n1009 & n1027 ) | ( n1017 & n1027 ) ;
  assign n1058 = ( n1009 & ~n1028 ) | ( n1009 & n1057 ) | ( ~n1028 & n1057 ) ;
  assign n1059 = ( ~n1019 & n1021 ) | ( ~n1019 & n1026 ) | ( n1021 & n1026 ) ;
  assign n1060 = ( n1019 & ~n1027 ) | ( n1019 & n1059 ) | ( ~n1027 & n1059 ) ;
  assign n1061 = ( ~n1046 & n1048 ) | ( ~n1046 & n1052 ) | ( n1048 & n1052 ) ;
  assign n1062 = ( n1046 & ~n1053 ) | ( n1046 & n1061 ) | ( ~n1053 & n1061 ) ;
  assign n1063 = ( ~n1032 & n1034 ) | ( ~n1032 & n1050 ) | ( n1034 & n1050 ) ;
  assign n1064 = ( n1032 & ~n1051 ) | ( n1032 & n1063 ) | ( ~n1051 & n1063 ) ;
  assign n1065 = ( n1023 & n1025 ) | ( n1023 & n1064 ) | ( n1025 & n1064 ) ;
  assign n1066 = ~n1026 & n1065 ;
  assign n1067 = ( n1060 & n1062 ) | ( n1060 & n1066 ) | ( n1062 & n1066 ) ;
  assign n1068 = ( n1056 & n1058 ) | ( n1056 & n1067 ) | ( n1058 & n1067 ) ;
  assign n1069 = ( n1028 & n1054 ) | ( n1028 & n1068 ) | ( n1054 & n1068 ) ;
  assign n1070 = ( x436 & x437 ) | ( x436 & x438 ) | ( x437 & x438 ) ;
  assign n1071 = ( x433 & x434 ) | ( x433 & x435 ) | ( x434 & x435 ) ;
  assign n1072 = ( ~x436 & x437 ) | ( ~x436 & x438 ) | ( x437 & x438 ) ;
  assign n1073 = ( x436 & ~n1070 ) | ( x436 & n1072 ) | ( ~n1070 & n1072 ) ;
  assign n1074 = ( ~x433 & x434 ) | ( ~x433 & x435 ) | ( x434 & x435 ) ;
  assign n1075 = ( x433 & ~n1071 ) | ( x433 & n1074 ) | ( ~n1071 & n1074 ) ;
  assign n1076 = n1073 & n1075 ;
  assign n1077 = ( n1070 & n1071 ) | ( n1070 & n1076 ) | ( n1071 & n1076 ) ;
  assign n1078 = ( x427 & x428 ) | ( x427 & x429 ) | ( x428 & x429 ) ;
  assign n1079 = ( x430 & x431 ) | ( x430 & x432 ) | ( x431 & x432 ) ;
  assign n1080 = ( ~x430 & x431 ) | ( ~x430 & x432 ) | ( x431 & x432 ) ;
  assign n1081 = ( x430 & ~n1079 ) | ( x430 & n1080 ) | ( ~n1079 & n1080 ) ;
  assign n1082 = ( ~x427 & x428 ) | ( ~x427 & x429 ) | ( x428 & x429 ) ;
  assign n1083 = ( x427 & ~n1078 ) | ( x427 & n1082 ) | ( ~n1078 & n1082 ) ;
  assign n1084 = n1081 & n1083 ;
  assign n1085 = ( n1078 & n1079 ) | ( n1078 & n1084 ) | ( n1079 & n1084 ) ;
  assign n1086 = ( ~n1070 & n1071 ) | ( ~n1070 & n1076 ) | ( n1071 & n1076 ) ;
  assign n1087 = ( n1070 & ~n1077 ) | ( n1070 & n1086 ) | ( ~n1077 & n1086 ) ;
  assign n1088 = ( ~n1078 & n1079 ) | ( ~n1078 & n1084 ) | ( n1079 & n1084 ) ;
  assign n1089 = ( n1078 & ~n1085 ) | ( n1078 & n1088 ) | ( ~n1085 & n1088 ) ;
  assign n1090 = n1073 | n1075 ;
  assign n1091 = ~n1076 & n1090 ;
  assign n1092 = n1081 | n1083 ;
  assign n1093 = ~n1084 & n1092 ;
  assign n1094 = n1091 & n1093 ;
  assign n1095 = ( n1087 & n1089 ) | ( n1087 & n1094 ) | ( n1089 & n1094 ) ;
  assign n1096 = ( n1077 & n1085 ) | ( n1077 & n1095 ) | ( n1085 & n1095 ) ;
  assign n1097 = ( x424 & x425 ) | ( x424 & x426 ) | ( x425 & x426 ) ;
  assign n1098 = ( x421 & x422 ) | ( x421 & x423 ) | ( x422 & x423 ) ;
  assign n1099 = ( ~x424 & x425 ) | ( ~x424 & x426 ) | ( x425 & x426 ) ;
  assign n1100 = ( x424 & ~n1097 ) | ( x424 & n1099 ) | ( ~n1097 & n1099 ) ;
  assign n1101 = ( ~x421 & x422 ) | ( ~x421 & x423 ) | ( x422 & x423 ) ;
  assign n1102 = ( x421 & ~n1098 ) | ( x421 & n1101 ) | ( ~n1098 & n1101 ) ;
  assign n1103 = n1100 & n1102 ;
  assign n1104 = ( n1097 & n1098 ) | ( n1097 & n1103 ) | ( n1098 & n1103 ) ;
  assign n1105 = ( x415 & x416 ) | ( x415 & x417 ) | ( x416 & x417 ) ;
  assign n1106 = ( x418 & x419 ) | ( x418 & x420 ) | ( x419 & x420 ) ;
  assign n1107 = ( ~x418 & x419 ) | ( ~x418 & x420 ) | ( x419 & x420 ) ;
  assign n1108 = ( x418 & ~n1106 ) | ( x418 & n1107 ) | ( ~n1106 & n1107 ) ;
  assign n1109 = ( ~x415 & x416 ) | ( ~x415 & x417 ) | ( x416 & x417 ) ;
  assign n1110 = ( x415 & ~n1105 ) | ( x415 & n1109 ) | ( ~n1105 & n1109 ) ;
  assign n1111 = n1108 & n1110 ;
  assign n1112 = ( n1105 & n1106 ) | ( n1105 & n1111 ) | ( n1106 & n1111 ) ;
  assign n1113 = ( ~n1097 & n1098 ) | ( ~n1097 & n1103 ) | ( n1098 & n1103 ) ;
  assign n1114 = ( n1097 & ~n1104 ) | ( n1097 & n1113 ) | ( ~n1104 & n1113 ) ;
  assign n1115 = ( ~n1105 & n1106 ) | ( ~n1105 & n1111 ) | ( n1106 & n1111 ) ;
  assign n1116 = ( n1105 & ~n1112 ) | ( n1105 & n1115 ) | ( ~n1112 & n1115 ) ;
  assign n1117 = n1108 | n1110 ;
  assign n1118 = ~n1111 & n1117 ;
  assign n1119 = ( n1100 & n1102 ) | ( n1100 & n1118 ) | ( n1102 & n1118 ) ;
  assign n1120 = ~n1103 & n1119 ;
  assign n1121 = ( n1114 & n1116 ) | ( n1114 & n1120 ) | ( n1116 & n1120 ) ;
  assign n1122 = ( n1104 & n1112 ) | ( n1104 & n1121 ) | ( n1112 & n1121 ) ;
  assign n1123 = ( ~n1104 & n1112 ) | ( ~n1104 & n1121 ) | ( n1112 & n1121 ) ;
  assign n1124 = ( n1104 & ~n1122 ) | ( n1104 & n1123 ) | ( ~n1122 & n1123 ) ;
  assign n1125 = ( ~n1077 & n1085 ) | ( ~n1077 & n1095 ) | ( n1085 & n1095 ) ;
  assign n1126 = ( n1077 & ~n1096 ) | ( n1077 & n1125 ) | ( ~n1096 & n1125 ) ;
  assign n1127 = ( ~n1087 & n1089 ) | ( ~n1087 & n1094 ) | ( n1089 & n1094 ) ;
  assign n1128 = ( n1087 & ~n1095 ) | ( n1087 & n1127 ) | ( ~n1095 & n1127 ) ;
  assign n1129 = ( ~n1114 & n1116 ) | ( ~n1114 & n1120 ) | ( n1116 & n1120 ) ;
  assign n1130 = ( n1114 & ~n1121 ) | ( n1114 & n1129 ) | ( ~n1121 & n1129 ) ;
  assign n1131 = ( ~n1100 & n1102 ) | ( ~n1100 & n1118 ) | ( n1102 & n1118 ) ;
  assign n1132 = ( n1100 & ~n1119 ) | ( n1100 & n1131 ) | ( ~n1119 & n1131 ) ;
  assign n1133 = ( n1091 & n1093 ) | ( n1091 & n1132 ) | ( n1093 & n1132 ) ;
  assign n1134 = ~n1094 & n1133 ;
  assign n1135 = ( n1128 & n1130 ) | ( n1128 & n1134 ) | ( n1130 & n1134 ) ;
  assign n1136 = ( n1124 & n1126 ) | ( n1124 & n1135 ) | ( n1126 & n1135 ) ;
  assign n1137 = ( n1096 & n1122 ) | ( n1096 & n1136 ) | ( n1122 & n1136 ) ;
  assign n1138 = ( ~n1028 & n1054 ) | ( ~n1028 & n1068 ) | ( n1054 & n1068 ) ;
  assign n1139 = ( n1028 & ~n1069 ) | ( n1028 & n1138 ) | ( ~n1069 & n1138 ) ;
  assign n1140 = ( ~n1096 & n1122 ) | ( ~n1096 & n1136 ) | ( n1122 & n1136 ) ;
  assign n1141 = ( n1096 & ~n1137 ) | ( n1096 & n1140 ) | ( ~n1137 & n1140 ) ;
  assign n1142 = ( ~n1124 & n1126 ) | ( ~n1124 & n1135 ) | ( n1126 & n1135 ) ;
  assign n1143 = ( n1124 & ~n1136 ) | ( n1124 & n1142 ) | ( ~n1136 & n1142 ) ;
  assign n1144 = ( ~n1056 & n1058 ) | ( ~n1056 & n1067 ) | ( n1058 & n1067 ) ;
  assign n1145 = ( n1056 & ~n1068 ) | ( n1056 & n1144 ) | ( ~n1068 & n1144 ) ;
  assign n1146 = ( n1060 & n1062 ) | ( n1060 & ~n1066 ) | ( n1062 & ~n1066 ) ;
  assign n1147 = ( n1066 & ~n1067 ) | ( n1066 & n1146 ) | ( ~n1067 & n1146 ) ;
  assign n1148 = ( n1128 & n1130 ) | ( n1128 & ~n1134 ) | ( n1130 & ~n1134 ) ;
  assign n1149 = ( n1134 & ~n1135 ) | ( n1134 & n1148 ) | ( ~n1135 & n1148 ) ;
  assign n1150 = ( ~n1023 & n1025 ) | ( ~n1023 & n1064 ) | ( n1025 & n1064 ) ;
  assign n1151 = ( n1023 & ~n1065 ) | ( n1023 & n1150 ) | ( ~n1065 & n1150 ) ;
  assign n1152 = ( ~n1091 & n1093 ) | ( ~n1091 & n1132 ) | ( n1093 & n1132 ) ;
  assign n1153 = ( n1091 & ~n1133 ) | ( n1091 & n1152 ) | ( ~n1133 & n1152 ) ;
  assign n1154 = n1151 & n1153 ;
  assign n1155 = ( n1147 & n1149 ) | ( n1147 & n1154 ) | ( n1149 & n1154 ) ;
  assign n1156 = ( n1143 & n1145 ) | ( n1143 & n1155 ) | ( n1145 & n1155 ) ;
  assign n1157 = ( n1139 & n1141 ) | ( n1139 & n1156 ) | ( n1141 & n1156 ) ;
  assign n1158 = ( n1069 & n1137 ) | ( n1069 & n1157 ) | ( n1137 & n1157 ) ;
  assign n1159 = ( x412 & x413 ) | ( x412 & x414 ) | ( x413 & x414 ) ;
  assign n1160 = ( x409 & x410 ) | ( x409 & x411 ) | ( x410 & x411 ) ;
  assign n1161 = ( ~x412 & x413 ) | ( ~x412 & x414 ) | ( x413 & x414 ) ;
  assign n1162 = ( x412 & ~n1159 ) | ( x412 & n1161 ) | ( ~n1159 & n1161 ) ;
  assign n1163 = ( ~x409 & x410 ) | ( ~x409 & x411 ) | ( x410 & x411 ) ;
  assign n1164 = ( x409 & ~n1160 ) | ( x409 & n1163 ) | ( ~n1160 & n1163 ) ;
  assign n1165 = n1162 & n1164 ;
  assign n1166 = ( n1159 & n1160 ) | ( n1159 & n1165 ) | ( n1160 & n1165 ) ;
  assign n1167 = ( x403 & x404 ) | ( x403 & x405 ) | ( x404 & x405 ) ;
  assign n1168 = ( x406 & x407 ) | ( x406 & x408 ) | ( x407 & x408 ) ;
  assign n1169 = ( ~x406 & x407 ) | ( ~x406 & x408 ) | ( x407 & x408 ) ;
  assign n1170 = ( x406 & ~n1168 ) | ( x406 & n1169 ) | ( ~n1168 & n1169 ) ;
  assign n1171 = ( ~x403 & x404 ) | ( ~x403 & x405 ) | ( x404 & x405 ) ;
  assign n1172 = ( x403 & ~n1167 ) | ( x403 & n1171 ) | ( ~n1167 & n1171 ) ;
  assign n1173 = n1170 & n1172 ;
  assign n1174 = ( n1167 & n1168 ) | ( n1167 & n1173 ) | ( n1168 & n1173 ) ;
  assign n1175 = ( ~n1159 & n1160 ) | ( ~n1159 & n1165 ) | ( n1160 & n1165 ) ;
  assign n1176 = ( n1159 & ~n1166 ) | ( n1159 & n1175 ) | ( ~n1166 & n1175 ) ;
  assign n1177 = ( ~n1167 & n1168 ) | ( ~n1167 & n1173 ) | ( n1168 & n1173 ) ;
  assign n1178 = ( n1167 & ~n1174 ) | ( n1167 & n1177 ) | ( ~n1174 & n1177 ) ;
  assign n1179 = n1162 | n1164 ;
  assign n1180 = ~n1165 & n1179 ;
  assign n1181 = n1170 | n1172 ;
  assign n1182 = ~n1173 & n1181 ;
  assign n1183 = n1180 & n1182 ;
  assign n1184 = ( n1176 & n1178 ) | ( n1176 & n1183 ) | ( n1178 & n1183 ) ;
  assign n1185 = ( n1166 & n1174 ) | ( n1166 & n1184 ) | ( n1174 & n1184 ) ;
  assign n1186 = ( x400 & x401 ) | ( x400 & x402 ) | ( x401 & x402 ) ;
  assign n1187 = ( x397 & x398 ) | ( x397 & x399 ) | ( x398 & x399 ) ;
  assign n1188 = ( ~x400 & x401 ) | ( ~x400 & x402 ) | ( x401 & x402 ) ;
  assign n1189 = ( x400 & ~n1186 ) | ( x400 & n1188 ) | ( ~n1186 & n1188 ) ;
  assign n1190 = ( ~x397 & x398 ) | ( ~x397 & x399 ) | ( x398 & x399 ) ;
  assign n1191 = ( x397 & ~n1187 ) | ( x397 & n1190 ) | ( ~n1187 & n1190 ) ;
  assign n1192 = n1189 & n1191 ;
  assign n1193 = ( n1186 & n1187 ) | ( n1186 & n1192 ) | ( n1187 & n1192 ) ;
  assign n1194 = ( x391 & x392 ) | ( x391 & x393 ) | ( x392 & x393 ) ;
  assign n1195 = ( x394 & x395 ) | ( x394 & x396 ) | ( x395 & x396 ) ;
  assign n1196 = ( ~x394 & x395 ) | ( ~x394 & x396 ) | ( x395 & x396 ) ;
  assign n1197 = ( x394 & ~n1195 ) | ( x394 & n1196 ) | ( ~n1195 & n1196 ) ;
  assign n1198 = ( ~x391 & x392 ) | ( ~x391 & x393 ) | ( x392 & x393 ) ;
  assign n1199 = ( x391 & ~n1194 ) | ( x391 & n1198 ) | ( ~n1194 & n1198 ) ;
  assign n1200 = n1197 & n1199 ;
  assign n1201 = ( n1194 & n1195 ) | ( n1194 & n1200 ) | ( n1195 & n1200 ) ;
  assign n1202 = ( ~n1186 & n1187 ) | ( ~n1186 & n1192 ) | ( n1187 & n1192 ) ;
  assign n1203 = ( n1186 & ~n1193 ) | ( n1186 & n1202 ) | ( ~n1193 & n1202 ) ;
  assign n1204 = ( ~n1194 & n1195 ) | ( ~n1194 & n1200 ) | ( n1195 & n1200 ) ;
  assign n1205 = ( n1194 & ~n1201 ) | ( n1194 & n1204 ) | ( ~n1201 & n1204 ) ;
  assign n1206 = n1197 | n1199 ;
  assign n1207 = ~n1200 & n1206 ;
  assign n1208 = ( n1189 & n1191 ) | ( n1189 & n1207 ) | ( n1191 & n1207 ) ;
  assign n1209 = ~n1192 & n1208 ;
  assign n1210 = ( n1203 & n1205 ) | ( n1203 & n1209 ) | ( n1205 & n1209 ) ;
  assign n1211 = ( n1193 & n1201 ) | ( n1193 & n1210 ) | ( n1201 & n1210 ) ;
  assign n1212 = ( ~n1193 & n1201 ) | ( ~n1193 & n1210 ) | ( n1201 & n1210 ) ;
  assign n1213 = ( n1193 & ~n1211 ) | ( n1193 & n1212 ) | ( ~n1211 & n1212 ) ;
  assign n1214 = ( ~n1166 & n1174 ) | ( ~n1166 & n1184 ) | ( n1174 & n1184 ) ;
  assign n1215 = ( n1166 & ~n1185 ) | ( n1166 & n1214 ) | ( ~n1185 & n1214 ) ;
  assign n1216 = ( ~n1176 & n1178 ) | ( ~n1176 & n1183 ) | ( n1178 & n1183 ) ;
  assign n1217 = ( n1176 & ~n1184 ) | ( n1176 & n1216 ) | ( ~n1184 & n1216 ) ;
  assign n1218 = ( ~n1203 & n1205 ) | ( ~n1203 & n1209 ) | ( n1205 & n1209 ) ;
  assign n1219 = ( n1203 & ~n1210 ) | ( n1203 & n1218 ) | ( ~n1210 & n1218 ) ;
  assign n1220 = ( ~n1189 & n1191 ) | ( ~n1189 & n1207 ) | ( n1191 & n1207 ) ;
  assign n1221 = ( n1189 & ~n1208 ) | ( n1189 & n1220 ) | ( ~n1208 & n1220 ) ;
  assign n1222 = ( n1180 & n1182 ) | ( n1180 & n1221 ) | ( n1182 & n1221 ) ;
  assign n1223 = ~n1183 & n1222 ;
  assign n1224 = ( n1217 & n1219 ) | ( n1217 & n1223 ) | ( n1219 & n1223 ) ;
  assign n1225 = ( n1213 & n1215 ) | ( n1213 & n1224 ) | ( n1215 & n1224 ) ;
  assign n1226 = ( n1185 & n1211 ) | ( n1185 & n1225 ) | ( n1211 & n1225 ) ;
  assign n1227 = ( x388 & x389 ) | ( x388 & x390 ) | ( x389 & x390 ) ;
  assign n1228 = ( x385 & x386 ) | ( x385 & x387 ) | ( x386 & x387 ) ;
  assign n1229 = ( ~x388 & x389 ) | ( ~x388 & x390 ) | ( x389 & x390 ) ;
  assign n1230 = ( x388 & ~n1227 ) | ( x388 & n1229 ) | ( ~n1227 & n1229 ) ;
  assign n1231 = ( ~x385 & x386 ) | ( ~x385 & x387 ) | ( x386 & x387 ) ;
  assign n1232 = ( x385 & ~n1228 ) | ( x385 & n1231 ) | ( ~n1228 & n1231 ) ;
  assign n1233 = n1230 & n1232 ;
  assign n1234 = ( n1227 & n1228 ) | ( n1227 & n1233 ) | ( n1228 & n1233 ) ;
  assign n1235 = ( x379 & x380 ) | ( x379 & x381 ) | ( x380 & x381 ) ;
  assign n1236 = ( x382 & x383 ) | ( x382 & x384 ) | ( x383 & x384 ) ;
  assign n1237 = ( ~x382 & x383 ) | ( ~x382 & x384 ) | ( x383 & x384 ) ;
  assign n1238 = ( x382 & ~n1236 ) | ( x382 & n1237 ) | ( ~n1236 & n1237 ) ;
  assign n1239 = ( ~x379 & x380 ) | ( ~x379 & x381 ) | ( x380 & x381 ) ;
  assign n1240 = ( x379 & ~n1235 ) | ( x379 & n1239 ) | ( ~n1235 & n1239 ) ;
  assign n1241 = n1238 & n1240 ;
  assign n1242 = ( n1235 & n1236 ) | ( n1235 & n1241 ) | ( n1236 & n1241 ) ;
  assign n1243 = ( ~n1227 & n1228 ) | ( ~n1227 & n1233 ) | ( n1228 & n1233 ) ;
  assign n1244 = ( n1227 & ~n1234 ) | ( n1227 & n1243 ) | ( ~n1234 & n1243 ) ;
  assign n1245 = ( ~n1235 & n1236 ) | ( ~n1235 & n1241 ) | ( n1236 & n1241 ) ;
  assign n1246 = ( n1235 & ~n1242 ) | ( n1235 & n1245 ) | ( ~n1242 & n1245 ) ;
  assign n1247 = n1230 | n1232 ;
  assign n1248 = ~n1233 & n1247 ;
  assign n1249 = n1238 | n1240 ;
  assign n1250 = ~n1241 & n1249 ;
  assign n1251 = n1248 & n1250 ;
  assign n1252 = ( n1244 & n1246 ) | ( n1244 & n1251 ) | ( n1246 & n1251 ) ;
  assign n1253 = ( n1234 & n1242 ) | ( n1234 & n1252 ) | ( n1242 & n1252 ) ;
  assign n1254 = ( x376 & x377 ) | ( x376 & x378 ) | ( x377 & x378 ) ;
  assign n1255 = ( x373 & x374 ) | ( x373 & x375 ) | ( x374 & x375 ) ;
  assign n1256 = ( ~x376 & x377 ) | ( ~x376 & x378 ) | ( x377 & x378 ) ;
  assign n1257 = ( x376 & ~n1254 ) | ( x376 & n1256 ) | ( ~n1254 & n1256 ) ;
  assign n1258 = ( ~x373 & x374 ) | ( ~x373 & x375 ) | ( x374 & x375 ) ;
  assign n1259 = ( x373 & ~n1255 ) | ( x373 & n1258 ) | ( ~n1255 & n1258 ) ;
  assign n1260 = n1257 & n1259 ;
  assign n1261 = ( n1254 & n1255 ) | ( n1254 & n1260 ) | ( n1255 & n1260 ) ;
  assign n1262 = ( x367 & x368 ) | ( x367 & x369 ) | ( x368 & x369 ) ;
  assign n1263 = ( x370 & x371 ) | ( x370 & x372 ) | ( x371 & x372 ) ;
  assign n1264 = ( ~x370 & x371 ) | ( ~x370 & x372 ) | ( x371 & x372 ) ;
  assign n1265 = ( x370 & ~n1263 ) | ( x370 & n1264 ) | ( ~n1263 & n1264 ) ;
  assign n1266 = ( ~x367 & x368 ) | ( ~x367 & x369 ) | ( x368 & x369 ) ;
  assign n1267 = ( x367 & ~n1262 ) | ( x367 & n1266 ) | ( ~n1262 & n1266 ) ;
  assign n1268 = n1265 & n1267 ;
  assign n1269 = ( n1262 & n1263 ) | ( n1262 & n1268 ) | ( n1263 & n1268 ) ;
  assign n1270 = ( ~n1254 & n1255 ) | ( ~n1254 & n1260 ) | ( n1255 & n1260 ) ;
  assign n1271 = ( n1254 & ~n1261 ) | ( n1254 & n1270 ) | ( ~n1261 & n1270 ) ;
  assign n1272 = ( ~n1262 & n1263 ) | ( ~n1262 & n1268 ) | ( n1263 & n1268 ) ;
  assign n1273 = ( n1262 & ~n1269 ) | ( n1262 & n1272 ) | ( ~n1269 & n1272 ) ;
  assign n1274 = n1265 | n1267 ;
  assign n1275 = ~n1268 & n1274 ;
  assign n1276 = ( n1257 & n1259 ) | ( n1257 & n1275 ) | ( n1259 & n1275 ) ;
  assign n1277 = ~n1260 & n1276 ;
  assign n1278 = ( n1271 & n1273 ) | ( n1271 & n1277 ) | ( n1273 & n1277 ) ;
  assign n1279 = ( n1261 & n1269 ) | ( n1261 & n1278 ) | ( n1269 & n1278 ) ;
  assign n1280 = ( ~n1261 & n1269 ) | ( ~n1261 & n1278 ) | ( n1269 & n1278 ) ;
  assign n1281 = ( n1261 & ~n1279 ) | ( n1261 & n1280 ) | ( ~n1279 & n1280 ) ;
  assign n1282 = ( ~n1234 & n1242 ) | ( ~n1234 & n1252 ) | ( n1242 & n1252 ) ;
  assign n1283 = ( n1234 & ~n1253 ) | ( n1234 & n1282 ) | ( ~n1253 & n1282 ) ;
  assign n1284 = ( ~n1244 & n1246 ) | ( ~n1244 & n1251 ) | ( n1246 & n1251 ) ;
  assign n1285 = ( n1244 & ~n1252 ) | ( n1244 & n1284 ) | ( ~n1252 & n1284 ) ;
  assign n1286 = ( ~n1271 & n1273 ) | ( ~n1271 & n1277 ) | ( n1273 & n1277 ) ;
  assign n1287 = ( n1271 & ~n1278 ) | ( n1271 & n1286 ) | ( ~n1278 & n1286 ) ;
  assign n1288 = ( ~n1257 & n1259 ) | ( ~n1257 & n1275 ) | ( n1259 & n1275 ) ;
  assign n1289 = ( n1257 & ~n1276 ) | ( n1257 & n1288 ) | ( ~n1276 & n1288 ) ;
  assign n1290 = ( n1248 & n1250 ) | ( n1248 & n1289 ) | ( n1250 & n1289 ) ;
  assign n1291 = ~n1251 & n1290 ;
  assign n1292 = ( n1285 & n1287 ) | ( n1285 & n1291 ) | ( n1287 & n1291 ) ;
  assign n1293 = ( n1281 & n1283 ) | ( n1281 & n1292 ) | ( n1283 & n1292 ) ;
  assign n1294 = ( n1253 & n1279 ) | ( n1253 & n1293 ) | ( n1279 & n1293 ) ;
  assign n1295 = ( ~n1185 & n1211 ) | ( ~n1185 & n1225 ) | ( n1211 & n1225 ) ;
  assign n1296 = ( n1185 & ~n1226 ) | ( n1185 & n1295 ) | ( ~n1226 & n1295 ) ;
  assign n1297 = ( ~n1253 & n1279 ) | ( ~n1253 & n1293 ) | ( n1279 & n1293 ) ;
  assign n1298 = ( n1253 & ~n1294 ) | ( n1253 & n1297 ) | ( ~n1294 & n1297 ) ;
  assign n1299 = ( ~n1281 & n1283 ) | ( ~n1281 & n1292 ) | ( n1283 & n1292 ) ;
  assign n1300 = ( n1281 & ~n1293 ) | ( n1281 & n1299 ) | ( ~n1293 & n1299 ) ;
  assign n1301 = ( ~n1213 & n1215 ) | ( ~n1213 & n1224 ) | ( n1215 & n1224 ) ;
  assign n1302 = ( n1213 & ~n1225 ) | ( n1213 & n1301 ) | ( ~n1225 & n1301 ) ;
  assign n1303 = ( n1217 & n1219 ) | ( n1217 & ~n1223 ) | ( n1219 & ~n1223 ) ;
  assign n1304 = ( n1223 & ~n1224 ) | ( n1223 & n1303 ) | ( ~n1224 & n1303 ) ;
  assign n1305 = ( n1285 & n1287 ) | ( n1285 & ~n1291 ) | ( n1287 & ~n1291 ) ;
  assign n1306 = ( n1291 & ~n1292 ) | ( n1291 & n1305 ) | ( ~n1292 & n1305 ) ;
  assign n1307 = ( ~n1180 & n1182 ) | ( ~n1180 & n1221 ) | ( n1182 & n1221 ) ;
  assign n1308 = ( n1180 & ~n1222 ) | ( n1180 & n1307 ) | ( ~n1222 & n1307 ) ;
  assign n1309 = ( ~n1248 & n1250 ) | ( ~n1248 & n1289 ) | ( n1250 & n1289 ) ;
  assign n1310 = ( n1248 & ~n1290 ) | ( n1248 & n1309 ) | ( ~n1290 & n1309 ) ;
  assign n1311 = n1308 & n1310 ;
  assign n1312 = ( n1304 & n1306 ) | ( n1304 & n1311 ) | ( n1306 & n1311 ) ;
  assign n1313 = ( n1300 & n1302 ) | ( n1300 & n1312 ) | ( n1302 & n1312 ) ;
  assign n1314 = ( n1296 & n1298 ) | ( n1296 & n1313 ) | ( n1298 & n1313 ) ;
  assign n1315 = ( n1226 & n1294 ) | ( n1226 & n1314 ) | ( n1294 & n1314 ) ;
  assign n1316 = ( ~n1226 & n1294 ) | ( ~n1226 & n1314 ) | ( n1294 & n1314 ) ;
  assign n1317 = ( n1226 & ~n1315 ) | ( n1226 & n1316 ) | ( ~n1315 & n1316 ) ;
  assign n1318 = ( ~n1069 & n1137 ) | ( ~n1069 & n1157 ) | ( n1137 & n1157 ) ;
  assign n1319 = ( n1069 & ~n1158 ) | ( n1069 & n1318 ) | ( ~n1158 & n1318 ) ;
  assign n1320 = ( ~n1139 & n1141 ) | ( ~n1139 & n1156 ) | ( n1141 & n1156 ) ;
  assign n1321 = ( n1139 & ~n1157 ) | ( n1139 & n1320 ) | ( ~n1157 & n1320 ) ;
  assign n1322 = ( ~n1296 & n1298 ) | ( ~n1296 & n1313 ) | ( n1298 & n1313 ) ;
  assign n1323 = ( n1296 & ~n1314 ) | ( n1296 & n1322 ) | ( ~n1314 & n1322 ) ;
  assign n1324 = ( ~n1300 & n1302 ) | ( ~n1300 & n1312 ) | ( n1302 & n1312 ) ;
  assign n1325 = ( n1300 & ~n1313 ) | ( n1300 & n1324 ) | ( ~n1313 & n1324 ) ;
  assign n1326 = ( ~n1143 & n1145 ) | ( ~n1143 & n1155 ) | ( n1145 & n1155 ) ;
  assign n1327 = ( n1143 & ~n1156 ) | ( n1143 & n1326 ) | ( ~n1156 & n1326 ) ;
  assign n1328 = ( ~n1147 & n1149 ) | ( ~n1147 & n1154 ) | ( n1149 & n1154 ) ;
  assign n1329 = ( n1147 & ~n1155 ) | ( n1147 & n1328 ) | ( ~n1155 & n1328 ) ;
  assign n1330 = ( ~n1304 & n1306 ) | ( ~n1304 & n1311 ) | ( n1306 & n1311 ) ;
  assign n1331 = ( n1304 & ~n1312 ) | ( n1304 & n1330 ) | ( ~n1312 & n1330 ) ;
  assign n1332 = n1308 | n1310 ;
  assign n1333 = ~n1311 & n1332 ;
  assign n1334 = ( n1151 & n1153 ) | ( n1151 & n1333 ) | ( n1153 & n1333 ) ;
  assign n1335 = ~n1154 & n1334 ;
  assign n1336 = ( n1329 & n1331 ) | ( n1329 & n1335 ) | ( n1331 & n1335 ) ;
  assign n1337 = ( n1325 & n1327 ) | ( n1325 & n1336 ) | ( n1327 & n1336 ) ;
  assign n1338 = ( n1321 & n1323 ) | ( n1321 & n1337 ) | ( n1323 & n1337 ) ;
  assign n1339 = ( n1317 & n1319 ) | ( n1317 & n1338 ) | ( n1319 & n1338 ) ;
  assign n1340 = ( n1158 & n1315 ) | ( n1158 & n1339 ) | ( n1315 & n1339 ) ;
  assign n1341 = ( x364 & x365 ) | ( x364 & x366 ) | ( x365 & x366 ) ;
  assign n1342 = ( x361 & x362 ) | ( x361 & x363 ) | ( x362 & x363 ) ;
  assign n1343 = ( ~x364 & x365 ) | ( ~x364 & x366 ) | ( x365 & x366 ) ;
  assign n1344 = ( x364 & ~n1341 ) | ( x364 & n1343 ) | ( ~n1341 & n1343 ) ;
  assign n1345 = ( ~x361 & x362 ) | ( ~x361 & x363 ) | ( x362 & x363 ) ;
  assign n1346 = ( x361 & ~n1342 ) | ( x361 & n1345 ) | ( ~n1342 & n1345 ) ;
  assign n1347 = n1344 & n1346 ;
  assign n1348 = ( n1341 & n1342 ) | ( n1341 & n1347 ) | ( n1342 & n1347 ) ;
  assign n1349 = ( x355 & x356 ) | ( x355 & x357 ) | ( x356 & x357 ) ;
  assign n1350 = ( x358 & x359 ) | ( x358 & x360 ) | ( x359 & x360 ) ;
  assign n1351 = ( ~x358 & x359 ) | ( ~x358 & x360 ) | ( x359 & x360 ) ;
  assign n1352 = ( x358 & ~n1350 ) | ( x358 & n1351 ) | ( ~n1350 & n1351 ) ;
  assign n1353 = ( ~x355 & x356 ) | ( ~x355 & x357 ) | ( x356 & x357 ) ;
  assign n1354 = ( x355 & ~n1349 ) | ( x355 & n1353 ) | ( ~n1349 & n1353 ) ;
  assign n1355 = n1352 & n1354 ;
  assign n1356 = ( n1349 & n1350 ) | ( n1349 & n1355 ) | ( n1350 & n1355 ) ;
  assign n1357 = ( ~n1341 & n1342 ) | ( ~n1341 & n1347 ) | ( n1342 & n1347 ) ;
  assign n1358 = ( n1341 & ~n1348 ) | ( n1341 & n1357 ) | ( ~n1348 & n1357 ) ;
  assign n1359 = ( ~n1349 & n1350 ) | ( ~n1349 & n1355 ) | ( n1350 & n1355 ) ;
  assign n1360 = ( n1349 & ~n1356 ) | ( n1349 & n1359 ) | ( ~n1356 & n1359 ) ;
  assign n1361 = n1344 | n1346 ;
  assign n1362 = ~n1347 & n1361 ;
  assign n1363 = n1352 | n1354 ;
  assign n1364 = ~n1355 & n1363 ;
  assign n1365 = n1362 & n1364 ;
  assign n1366 = ( n1358 & n1360 ) | ( n1358 & n1365 ) | ( n1360 & n1365 ) ;
  assign n1367 = ( n1348 & n1356 ) | ( n1348 & n1366 ) | ( n1356 & n1366 ) ;
  assign n1368 = ( x352 & x353 ) | ( x352 & x354 ) | ( x353 & x354 ) ;
  assign n1369 = ( x349 & x350 ) | ( x349 & x351 ) | ( x350 & x351 ) ;
  assign n1370 = ( ~x352 & x353 ) | ( ~x352 & x354 ) | ( x353 & x354 ) ;
  assign n1371 = ( x352 & ~n1368 ) | ( x352 & n1370 ) | ( ~n1368 & n1370 ) ;
  assign n1372 = ( ~x349 & x350 ) | ( ~x349 & x351 ) | ( x350 & x351 ) ;
  assign n1373 = ( x349 & ~n1369 ) | ( x349 & n1372 ) | ( ~n1369 & n1372 ) ;
  assign n1374 = n1371 & n1373 ;
  assign n1375 = ( n1368 & n1369 ) | ( n1368 & n1374 ) | ( n1369 & n1374 ) ;
  assign n1376 = ( x343 & x344 ) | ( x343 & x345 ) | ( x344 & x345 ) ;
  assign n1377 = ( x346 & x347 ) | ( x346 & x348 ) | ( x347 & x348 ) ;
  assign n1378 = ( ~x346 & x347 ) | ( ~x346 & x348 ) | ( x347 & x348 ) ;
  assign n1379 = ( x346 & ~n1377 ) | ( x346 & n1378 ) | ( ~n1377 & n1378 ) ;
  assign n1380 = ( ~x343 & x344 ) | ( ~x343 & x345 ) | ( x344 & x345 ) ;
  assign n1381 = ( x343 & ~n1376 ) | ( x343 & n1380 ) | ( ~n1376 & n1380 ) ;
  assign n1382 = n1379 & n1381 ;
  assign n1383 = ( n1376 & n1377 ) | ( n1376 & n1382 ) | ( n1377 & n1382 ) ;
  assign n1384 = ( ~n1368 & n1369 ) | ( ~n1368 & n1374 ) | ( n1369 & n1374 ) ;
  assign n1385 = ( n1368 & ~n1375 ) | ( n1368 & n1384 ) | ( ~n1375 & n1384 ) ;
  assign n1386 = ( ~n1376 & n1377 ) | ( ~n1376 & n1382 ) | ( n1377 & n1382 ) ;
  assign n1387 = ( n1376 & ~n1383 ) | ( n1376 & n1386 ) | ( ~n1383 & n1386 ) ;
  assign n1388 = n1379 | n1381 ;
  assign n1389 = ~n1382 & n1388 ;
  assign n1390 = ( n1371 & n1373 ) | ( n1371 & n1389 ) | ( n1373 & n1389 ) ;
  assign n1391 = ~n1374 & n1390 ;
  assign n1392 = ( n1385 & n1387 ) | ( n1385 & n1391 ) | ( n1387 & n1391 ) ;
  assign n1393 = ( n1375 & n1383 ) | ( n1375 & n1392 ) | ( n1383 & n1392 ) ;
  assign n1394 = ( ~n1375 & n1383 ) | ( ~n1375 & n1392 ) | ( n1383 & n1392 ) ;
  assign n1395 = ( n1375 & ~n1393 ) | ( n1375 & n1394 ) | ( ~n1393 & n1394 ) ;
  assign n1396 = ( ~n1348 & n1356 ) | ( ~n1348 & n1366 ) | ( n1356 & n1366 ) ;
  assign n1397 = ( n1348 & ~n1367 ) | ( n1348 & n1396 ) | ( ~n1367 & n1396 ) ;
  assign n1398 = ( ~n1358 & n1360 ) | ( ~n1358 & n1365 ) | ( n1360 & n1365 ) ;
  assign n1399 = ( n1358 & ~n1366 ) | ( n1358 & n1398 ) | ( ~n1366 & n1398 ) ;
  assign n1400 = ( ~n1385 & n1387 ) | ( ~n1385 & n1391 ) | ( n1387 & n1391 ) ;
  assign n1401 = ( n1385 & ~n1392 ) | ( n1385 & n1400 ) | ( ~n1392 & n1400 ) ;
  assign n1402 = ( ~n1371 & n1373 ) | ( ~n1371 & n1389 ) | ( n1373 & n1389 ) ;
  assign n1403 = ( n1371 & ~n1390 ) | ( n1371 & n1402 ) | ( ~n1390 & n1402 ) ;
  assign n1404 = ( n1362 & n1364 ) | ( n1362 & n1403 ) | ( n1364 & n1403 ) ;
  assign n1405 = ~n1365 & n1404 ;
  assign n1406 = ( n1399 & n1401 ) | ( n1399 & n1405 ) | ( n1401 & n1405 ) ;
  assign n1407 = ( n1395 & n1397 ) | ( n1395 & n1406 ) | ( n1397 & n1406 ) ;
  assign n1408 = ( n1367 & n1393 ) | ( n1367 & n1407 ) | ( n1393 & n1407 ) ;
  assign n1409 = ( x340 & x341 ) | ( x340 & x342 ) | ( x341 & x342 ) ;
  assign n1410 = ( x337 & x338 ) | ( x337 & x339 ) | ( x338 & x339 ) ;
  assign n1411 = ( ~x340 & x341 ) | ( ~x340 & x342 ) | ( x341 & x342 ) ;
  assign n1412 = ( x340 & ~n1409 ) | ( x340 & n1411 ) | ( ~n1409 & n1411 ) ;
  assign n1413 = ( ~x337 & x338 ) | ( ~x337 & x339 ) | ( x338 & x339 ) ;
  assign n1414 = ( x337 & ~n1410 ) | ( x337 & n1413 ) | ( ~n1410 & n1413 ) ;
  assign n1415 = n1412 & n1414 ;
  assign n1416 = ( n1409 & n1410 ) | ( n1409 & n1415 ) | ( n1410 & n1415 ) ;
  assign n1417 = ( x331 & x332 ) | ( x331 & x333 ) | ( x332 & x333 ) ;
  assign n1418 = ( x334 & x335 ) | ( x334 & x336 ) | ( x335 & x336 ) ;
  assign n1419 = ( ~x334 & x335 ) | ( ~x334 & x336 ) | ( x335 & x336 ) ;
  assign n1420 = ( x334 & ~n1418 ) | ( x334 & n1419 ) | ( ~n1418 & n1419 ) ;
  assign n1421 = ( ~x331 & x332 ) | ( ~x331 & x333 ) | ( x332 & x333 ) ;
  assign n1422 = ( x331 & ~n1417 ) | ( x331 & n1421 ) | ( ~n1417 & n1421 ) ;
  assign n1423 = n1420 & n1422 ;
  assign n1424 = ( n1417 & n1418 ) | ( n1417 & n1423 ) | ( n1418 & n1423 ) ;
  assign n1425 = ( ~n1409 & n1410 ) | ( ~n1409 & n1415 ) | ( n1410 & n1415 ) ;
  assign n1426 = ( n1409 & ~n1416 ) | ( n1409 & n1425 ) | ( ~n1416 & n1425 ) ;
  assign n1427 = ( ~n1417 & n1418 ) | ( ~n1417 & n1423 ) | ( n1418 & n1423 ) ;
  assign n1428 = ( n1417 & ~n1424 ) | ( n1417 & n1427 ) | ( ~n1424 & n1427 ) ;
  assign n1429 = n1412 | n1414 ;
  assign n1430 = ~n1415 & n1429 ;
  assign n1431 = n1420 | n1422 ;
  assign n1432 = ~n1423 & n1431 ;
  assign n1433 = n1430 & n1432 ;
  assign n1434 = ( n1426 & n1428 ) | ( n1426 & n1433 ) | ( n1428 & n1433 ) ;
  assign n1435 = ( n1416 & n1424 ) | ( n1416 & n1434 ) | ( n1424 & n1434 ) ;
  assign n1436 = ( x328 & x329 ) | ( x328 & x330 ) | ( x329 & x330 ) ;
  assign n1437 = ( x325 & x326 ) | ( x325 & x327 ) | ( x326 & x327 ) ;
  assign n1438 = ( ~x328 & x329 ) | ( ~x328 & x330 ) | ( x329 & x330 ) ;
  assign n1439 = ( x328 & ~n1436 ) | ( x328 & n1438 ) | ( ~n1436 & n1438 ) ;
  assign n1440 = ( ~x325 & x326 ) | ( ~x325 & x327 ) | ( x326 & x327 ) ;
  assign n1441 = ( x325 & ~n1437 ) | ( x325 & n1440 ) | ( ~n1437 & n1440 ) ;
  assign n1442 = n1439 & n1441 ;
  assign n1443 = ( n1436 & n1437 ) | ( n1436 & n1442 ) | ( n1437 & n1442 ) ;
  assign n1444 = ( x319 & x320 ) | ( x319 & x321 ) | ( x320 & x321 ) ;
  assign n1445 = ( x322 & x323 ) | ( x322 & x324 ) | ( x323 & x324 ) ;
  assign n1446 = ( ~x322 & x323 ) | ( ~x322 & x324 ) | ( x323 & x324 ) ;
  assign n1447 = ( x322 & ~n1445 ) | ( x322 & n1446 ) | ( ~n1445 & n1446 ) ;
  assign n1448 = ( ~x319 & x320 ) | ( ~x319 & x321 ) | ( x320 & x321 ) ;
  assign n1449 = ( x319 & ~n1444 ) | ( x319 & n1448 ) | ( ~n1444 & n1448 ) ;
  assign n1450 = n1447 & n1449 ;
  assign n1451 = ( n1444 & n1445 ) | ( n1444 & n1450 ) | ( n1445 & n1450 ) ;
  assign n1452 = ( ~n1436 & n1437 ) | ( ~n1436 & n1442 ) | ( n1437 & n1442 ) ;
  assign n1453 = ( n1436 & ~n1443 ) | ( n1436 & n1452 ) | ( ~n1443 & n1452 ) ;
  assign n1454 = ( ~n1444 & n1445 ) | ( ~n1444 & n1450 ) | ( n1445 & n1450 ) ;
  assign n1455 = ( n1444 & ~n1451 ) | ( n1444 & n1454 ) | ( ~n1451 & n1454 ) ;
  assign n1456 = n1447 | n1449 ;
  assign n1457 = ~n1450 & n1456 ;
  assign n1458 = ( n1439 & n1441 ) | ( n1439 & n1457 ) | ( n1441 & n1457 ) ;
  assign n1459 = ~n1442 & n1458 ;
  assign n1460 = ( n1453 & n1455 ) | ( n1453 & n1459 ) | ( n1455 & n1459 ) ;
  assign n1461 = ( n1443 & n1451 ) | ( n1443 & n1460 ) | ( n1451 & n1460 ) ;
  assign n1462 = ( ~n1443 & n1451 ) | ( ~n1443 & n1460 ) | ( n1451 & n1460 ) ;
  assign n1463 = ( n1443 & ~n1461 ) | ( n1443 & n1462 ) | ( ~n1461 & n1462 ) ;
  assign n1464 = ( ~n1416 & n1424 ) | ( ~n1416 & n1434 ) | ( n1424 & n1434 ) ;
  assign n1465 = ( n1416 & ~n1435 ) | ( n1416 & n1464 ) | ( ~n1435 & n1464 ) ;
  assign n1466 = ( ~n1426 & n1428 ) | ( ~n1426 & n1433 ) | ( n1428 & n1433 ) ;
  assign n1467 = ( n1426 & ~n1434 ) | ( n1426 & n1466 ) | ( ~n1434 & n1466 ) ;
  assign n1468 = ( ~n1453 & n1455 ) | ( ~n1453 & n1459 ) | ( n1455 & n1459 ) ;
  assign n1469 = ( n1453 & ~n1460 ) | ( n1453 & n1468 ) | ( ~n1460 & n1468 ) ;
  assign n1470 = ( ~n1439 & n1441 ) | ( ~n1439 & n1457 ) | ( n1441 & n1457 ) ;
  assign n1471 = ( n1439 & ~n1458 ) | ( n1439 & n1470 ) | ( ~n1458 & n1470 ) ;
  assign n1472 = ( n1430 & n1432 ) | ( n1430 & n1471 ) | ( n1432 & n1471 ) ;
  assign n1473 = ~n1433 & n1472 ;
  assign n1474 = ( n1467 & n1469 ) | ( n1467 & n1473 ) | ( n1469 & n1473 ) ;
  assign n1475 = ( n1463 & n1465 ) | ( n1463 & n1474 ) | ( n1465 & n1474 ) ;
  assign n1476 = ( n1435 & n1461 ) | ( n1435 & n1475 ) | ( n1461 & n1475 ) ;
  assign n1477 = ( ~n1367 & n1393 ) | ( ~n1367 & n1407 ) | ( n1393 & n1407 ) ;
  assign n1478 = ( n1367 & ~n1408 ) | ( n1367 & n1477 ) | ( ~n1408 & n1477 ) ;
  assign n1479 = ( ~n1435 & n1461 ) | ( ~n1435 & n1475 ) | ( n1461 & n1475 ) ;
  assign n1480 = ( n1435 & ~n1476 ) | ( n1435 & n1479 ) | ( ~n1476 & n1479 ) ;
  assign n1481 = ( ~n1463 & n1465 ) | ( ~n1463 & n1474 ) | ( n1465 & n1474 ) ;
  assign n1482 = ( n1463 & ~n1475 ) | ( n1463 & n1481 ) | ( ~n1475 & n1481 ) ;
  assign n1483 = ( ~n1395 & n1397 ) | ( ~n1395 & n1406 ) | ( n1397 & n1406 ) ;
  assign n1484 = ( n1395 & ~n1407 ) | ( n1395 & n1483 ) | ( ~n1407 & n1483 ) ;
  assign n1485 = ( n1399 & n1401 ) | ( n1399 & ~n1405 ) | ( n1401 & ~n1405 ) ;
  assign n1486 = ( n1405 & ~n1406 ) | ( n1405 & n1485 ) | ( ~n1406 & n1485 ) ;
  assign n1487 = ( n1467 & n1469 ) | ( n1467 & ~n1473 ) | ( n1469 & ~n1473 ) ;
  assign n1488 = ( n1473 & ~n1474 ) | ( n1473 & n1487 ) | ( ~n1474 & n1487 ) ;
  assign n1489 = ( ~n1362 & n1364 ) | ( ~n1362 & n1403 ) | ( n1364 & n1403 ) ;
  assign n1490 = ( n1362 & ~n1404 ) | ( n1362 & n1489 ) | ( ~n1404 & n1489 ) ;
  assign n1491 = ( ~n1430 & n1432 ) | ( ~n1430 & n1471 ) | ( n1432 & n1471 ) ;
  assign n1492 = ( n1430 & ~n1472 ) | ( n1430 & n1491 ) | ( ~n1472 & n1491 ) ;
  assign n1493 = n1490 & n1492 ;
  assign n1494 = ( n1486 & n1488 ) | ( n1486 & n1493 ) | ( n1488 & n1493 ) ;
  assign n1495 = ( n1482 & n1484 ) | ( n1482 & n1494 ) | ( n1484 & n1494 ) ;
  assign n1496 = ( n1478 & n1480 ) | ( n1478 & n1495 ) | ( n1480 & n1495 ) ;
  assign n1497 = ( n1408 & n1476 ) | ( n1408 & n1496 ) | ( n1476 & n1496 ) ;
  assign n1498 = ( x316 & x317 ) | ( x316 & x318 ) | ( x317 & x318 ) ;
  assign n1499 = ( x313 & x314 ) | ( x313 & x315 ) | ( x314 & x315 ) ;
  assign n1500 = ( ~x316 & x317 ) | ( ~x316 & x318 ) | ( x317 & x318 ) ;
  assign n1501 = ( x316 & ~n1498 ) | ( x316 & n1500 ) | ( ~n1498 & n1500 ) ;
  assign n1502 = ( ~x313 & x314 ) | ( ~x313 & x315 ) | ( x314 & x315 ) ;
  assign n1503 = ( x313 & ~n1499 ) | ( x313 & n1502 ) | ( ~n1499 & n1502 ) ;
  assign n1504 = n1501 & n1503 ;
  assign n1505 = ( n1498 & n1499 ) | ( n1498 & n1504 ) | ( n1499 & n1504 ) ;
  assign n1506 = ( x307 & x308 ) | ( x307 & x309 ) | ( x308 & x309 ) ;
  assign n1507 = ( x310 & x311 ) | ( x310 & x312 ) | ( x311 & x312 ) ;
  assign n1508 = ( ~x310 & x311 ) | ( ~x310 & x312 ) | ( x311 & x312 ) ;
  assign n1509 = ( x310 & ~n1507 ) | ( x310 & n1508 ) | ( ~n1507 & n1508 ) ;
  assign n1510 = ( ~x307 & x308 ) | ( ~x307 & x309 ) | ( x308 & x309 ) ;
  assign n1511 = ( x307 & ~n1506 ) | ( x307 & n1510 ) | ( ~n1506 & n1510 ) ;
  assign n1512 = n1509 & n1511 ;
  assign n1513 = ( n1506 & n1507 ) | ( n1506 & n1512 ) | ( n1507 & n1512 ) ;
  assign n1514 = ( ~n1498 & n1499 ) | ( ~n1498 & n1504 ) | ( n1499 & n1504 ) ;
  assign n1515 = ( n1498 & ~n1505 ) | ( n1498 & n1514 ) | ( ~n1505 & n1514 ) ;
  assign n1516 = ( ~n1506 & n1507 ) | ( ~n1506 & n1512 ) | ( n1507 & n1512 ) ;
  assign n1517 = ( n1506 & ~n1513 ) | ( n1506 & n1516 ) | ( ~n1513 & n1516 ) ;
  assign n1518 = n1501 | n1503 ;
  assign n1519 = ~n1504 & n1518 ;
  assign n1520 = n1509 | n1511 ;
  assign n1521 = ~n1512 & n1520 ;
  assign n1522 = n1519 & n1521 ;
  assign n1523 = ( n1515 & n1517 ) | ( n1515 & n1522 ) | ( n1517 & n1522 ) ;
  assign n1524 = ( n1505 & n1513 ) | ( n1505 & n1523 ) | ( n1513 & n1523 ) ;
  assign n1525 = ( x304 & x305 ) | ( x304 & x306 ) | ( x305 & x306 ) ;
  assign n1526 = ( x301 & x302 ) | ( x301 & x303 ) | ( x302 & x303 ) ;
  assign n1527 = ( ~x304 & x305 ) | ( ~x304 & x306 ) | ( x305 & x306 ) ;
  assign n1528 = ( x304 & ~n1525 ) | ( x304 & n1527 ) | ( ~n1525 & n1527 ) ;
  assign n1529 = ( ~x301 & x302 ) | ( ~x301 & x303 ) | ( x302 & x303 ) ;
  assign n1530 = ( x301 & ~n1526 ) | ( x301 & n1529 ) | ( ~n1526 & n1529 ) ;
  assign n1531 = n1528 & n1530 ;
  assign n1532 = ( n1525 & n1526 ) | ( n1525 & n1531 ) | ( n1526 & n1531 ) ;
  assign n1533 = ( x295 & x296 ) | ( x295 & x297 ) | ( x296 & x297 ) ;
  assign n1534 = ( x298 & x299 ) | ( x298 & x300 ) | ( x299 & x300 ) ;
  assign n1535 = ( ~x298 & x299 ) | ( ~x298 & x300 ) | ( x299 & x300 ) ;
  assign n1536 = ( x298 & ~n1534 ) | ( x298 & n1535 ) | ( ~n1534 & n1535 ) ;
  assign n1537 = ( ~x295 & x296 ) | ( ~x295 & x297 ) | ( x296 & x297 ) ;
  assign n1538 = ( x295 & ~n1533 ) | ( x295 & n1537 ) | ( ~n1533 & n1537 ) ;
  assign n1539 = n1536 & n1538 ;
  assign n1540 = ( n1533 & n1534 ) | ( n1533 & n1539 ) | ( n1534 & n1539 ) ;
  assign n1541 = ( ~n1525 & n1526 ) | ( ~n1525 & n1531 ) | ( n1526 & n1531 ) ;
  assign n1542 = ( n1525 & ~n1532 ) | ( n1525 & n1541 ) | ( ~n1532 & n1541 ) ;
  assign n1543 = ( ~n1533 & n1534 ) | ( ~n1533 & n1539 ) | ( n1534 & n1539 ) ;
  assign n1544 = ( n1533 & ~n1540 ) | ( n1533 & n1543 ) | ( ~n1540 & n1543 ) ;
  assign n1545 = n1536 | n1538 ;
  assign n1546 = ~n1539 & n1545 ;
  assign n1547 = ( n1528 & n1530 ) | ( n1528 & n1546 ) | ( n1530 & n1546 ) ;
  assign n1548 = ~n1531 & n1547 ;
  assign n1549 = ( n1542 & n1544 ) | ( n1542 & n1548 ) | ( n1544 & n1548 ) ;
  assign n1550 = ( n1532 & n1540 ) | ( n1532 & n1549 ) | ( n1540 & n1549 ) ;
  assign n1551 = ( ~n1532 & n1540 ) | ( ~n1532 & n1549 ) | ( n1540 & n1549 ) ;
  assign n1552 = ( n1532 & ~n1550 ) | ( n1532 & n1551 ) | ( ~n1550 & n1551 ) ;
  assign n1553 = ( ~n1505 & n1513 ) | ( ~n1505 & n1523 ) | ( n1513 & n1523 ) ;
  assign n1554 = ( n1505 & ~n1524 ) | ( n1505 & n1553 ) | ( ~n1524 & n1553 ) ;
  assign n1555 = ( ~n1515 & n1517 ) | ( ~n1515 & n1522 ) | ( n1517 & n1522 ) ;
  assign n1556 = ( n1515 & ~n1523 ) | ( n1515 & n1555 ) | ( ~n1523 & n1555 ) ;
  assign n1557 = ( ~n1542 & n1544 ) | ( ~n1542 & n1548 ) | ( n1544 & n1548 ) ;
  assign n1558 = ( n1542 & ~n1549 ) | ( n1542 & n1557 ) | ( ~n1549 & n1557 ) ;
  assign n1559 = ( ~n1528 & n1530 ) | ( ~n1528 & n1546 ) | ( n1530 & n1546 ) ;
  assign n1560 = ( n1528 & ~n1547 ) | ( n1528 & n1559 ) | ( ~n1547 & n1559 ) ;
  assign n1561 = ( n1519 & n1521 ) | ( n1519 & n1560 ) | ( n1521 & n1560 ) ;
  assign n1562 = ~n1522 & n1561 ;
  assign n1563 = ( n1556 & n1558 ) | ( n1556 & n1562 ) | ( n1558 & n1562 ) ;
  assign n1564 = ( n1552 & n1554 ) | ( n1552 & n1563 ) | ( n1554 & n1563 ) ;
  assign n1565 = ( n1524 & n1550 ) | ( n1524 & n1564 ) | ( n1550 & n1564 ) ;
  assign n1566 = ( x292 & x293 ) | ( x292 & x294 ) | ( x293 & x294 ) ;
  assign n1567 = ( x289 & x290 ) | ( x289 & x291 ) | ( x290 & x291 ) ;
  assign n1568 = ( ~x292 & x293 ) | ( ~x292 & x294 ) | ( x293 & x294 ) ;
  assign n1569 = ( x292 & ~n1566 ) | ( x292 & n1568 ) | ( ~n1566 & n1568 ) ;
  assign n1570 = ( ~x289 & x290 ) | ( ~x289 & x291 ) | ( x290 & x291 ) ;
  assign n1571 = ( x289 & ~n1567 ) | ( x289 & n1570 ) | ( ~n1567 & n1570 ) ;
  assign n1572 = n1569 & n1571 ;
  assign n1573 = ( n1566 & n1567 ) | ( n1566 & n1572 ) | ( n1567 & n1572 ) ;
  assign n1574 = ( x283 & x284 ) | ( x283 & x285 ) | ( x284 & x285 ) ;
  assign n1575 = ( x286 & x287 ) | ( x286 & x288 ) | ( x287 & x288 ) ;
  assign n1576 = ( ~x286 & x287 ) | ( ~x286 & x288 ) | ( x287 & x288 ) ;
  assign n1577 = ( x286 & ~n1575 ) | ( x286 & n1576 ) | ( ~n1575 & n1576 ) ;
  assign n1578 = ( ~x283 & x284 ) | ( ~x283 & x285 ) | ( x284 & x285 ) ;
  assign n1579 = ( x283 & ~n1574 ) | ( x283 & n1578 ) | ( ~n1574 & n1578 ) ;
  assign n1580 = n1577 & n1579 ;
  assign n1581 = ( n1574 & n1575 ) | ( n1574 & n1580 ) | ( n1575 & n1580 ) ;
  assign n1582 = ( ~n1566 & n1567 ) | ( ~n1566 & n1572 ) | ( n1567 & n1572 ) ;
  assign n1583 = ( n1566 & ~n1573 ) | ( n1566 & n1582 ) | ( ~n1573 & n1582 ) ;
  assign n1584 = ( ~n1574 & n1575 ) | ( ~n1574 & n1580 ) | ( n1575 & n1580 ) ;
  assign n1585 = ( n1574 & ~n1581 ) | ( n1574 & n1584 ) | ( ~n1581 & n1584 ) ;
  assign n1586 = n1569 | n1571 ;
  assign n1587 = ~n1572 & n1586 ;
  assign n1588 = n1577 | n1579 ;
  assign n1589 = ~n1580 & n1588 ;
  assign n1590 = n1587 & n1589 ;
  assign n1591 = ( n1583 & n1585 ) | ( n1583 & n1590 ) | ( n1585 & n1590 ) ;
  assign n1592 = ( n1573 & n1581 ) | ( n1573 & n1591 ) | ( n1581 & n1591 ) ;
  assign n1593 = ( x280 & x281 ) | ( x280 & x282 ) | ( x281 & x282 ) ;
  assign n1594 = ( x277 & x278 ) | ( x277 & x279 ) | ( x278 & x279 ) ;
  assign n1595 = ( ~x280 & x281 ) | ( ~x280 & x282 ) | ( x281 & x282 ) ;
  assign n1596 = ( x280 & ~n1593 ) | ( x280 & n1595 ) | ( ~n1593 & n1595 ) ;
  assign n1597 = ( ~x277 & x278 ) | ( ~x277 & x279 ) | ( x278 & x279 ) ;
  assign n1598 = ( x277 & ~n1594 ) | ( x277 & n1597 ) | ( ~n1594 & n1597 ) ;
  assign n1599 = n1596 & n1598 ;
  assign n1600 = ( n1593 & n1594 ) | ( n1593 & n1599 ) | ( n1594 & n1599 ) ;
  assign n1601 = ( x271 & x272 ) | ( x271 & x273 ) | ( x272 & x273 ) ;
  assign n1602 = ( x274 & x275 ) | ( x274 & x276 ) | ( x275 & x276 ) ;
  assign n1603 = ( ~x274 & x275 ) | ( ~x274 & x276 ) | ( x275 & x276 ) ;
  assign n1604 = ( x274 & ~n1602 ) | ( x274 & n1603 ) | ( ~n1602 & n1603 ) ;
  assign n1605 = ( ~x271 & x272 ) | ( ~x271 & x273 ) | ( x272 & x273 ) ;
  assign n1606 = ( x271 & ~n1601 ) | ( x271 & n1605 ) | ( ~n1601 & n1605 ) ;
  assign n1607 = n1604 & n1606 ;
  assign n1608 = ( n1601 & n1602 ) | ( n1601 & n1607 ) | ( n1602 & n1607 ) ;
  assign n1609 = ( ~n1593 & n1594 ) | ( ~n1593 & n1599 ) | ( n1594 & n1599 ) ;
  assign n1610 = ( n1593 & ~n1600 ) | ( n1593 & n1609 ) | ( ~n1600 & n1609 ) ;
  assign n1611 = ( ~n1601 & n1602 ) | ( ~n1601 & n1607 ) | ( n1602 & n1607 ) ;
  assign n1612 = ( n1601 & ~n1608 ) | ( n1601 & n1611 ) | ( ~n1608 & n1611 ) ;
  assign n1613 = n1604 | n1606 ;
  assign n1614 = ~n1607 & n1613 ;
  assign n1615 = ( n1596 & n1598 ) | ( n1596 & n1614 ) | ( n1598 & n1614 ) ;
  assign n1616 = ~n1599 & n1615 ;
  assign n1617 = ( n1610 & n1612 ) | ( n1610 & n1616 ) | ( n1612 & n1616 ) ;
  assign n1618 = ( n1600 & n1608 ) | ( n1600 & n1617 ) | ( n1608 & n1617 ) ;
  assign n1619 = ( ~n1600 & n1608 ) | ( ~n1600 & n1617 ) | ( n1608 & n1617 ) ;
  assign n1620 = ( n1600 & ~n1618 ) | ( n1600 & n1619 ) | ( ~n1618 & n1619 ) ;
  assign n1621 = ( ~n1573 & n1581 ) | ( ~n1573 & n1591 ) | ( n1581 & n1591 ) ;
  assign n1622 = ( n1573 & ~n1592 ) | ( n1573 & n1621 ) | ( ~n1592 & n1621 ) ;
  assign n1623 = ( ~n1583 & n1585 ) | ( ~n1583 & n1590 ) | ( n1585 & n1590 ) ;
  assign n1624 = ( n1583 & ~n1591 ) | ( n1583 & n1623 ) | ( ~n1591 & n1623 ) ;
  assign n1625 = ( ~n1610 & n1612 ) | ( ~n1610 & n1616 ) | ( n1612 & n1616 ) ;
  assign n1626 = ( n1610 & ~n1617 ) | ( n1610 & n1625 ) | ( ~n1617 & n1625 ) ;
  assign n1627 = ( ~n1596 & n1598 ) | ( ~n1596 & n1614 ) | ( n1598 & n1614 ) ;
  assign n1628 = ( n1596 & ~n1615 ) | ( n1596 & n1627 ) | ( ~n1615 & n1627 ) ;
  assign n1629 = ( n1587 & n1589 ) | ( n1587 & n1628 ) | ( n1589 & n1628 ) ;
  assign n1630 = ~n1590 & n1629 ;
  assign n1631 = ( n1624 & n1626 ) | ( n1624 & n1630 ) | ( n1626 & n1630 ) ;
  assign n1632 = ( n1620 & n1622 ) | ( n1620 & n1631 ) | ( n1622 & n1631 ) ;
  assign n1633 = ( n1592 & n1618 ) | ( n1592 & n1632 ) | ( n1618 & n1632 ) ;
  assign n1634 = ( ~n1524 & n1550 ) | ( ~n1524 & n1564 ) | ( n1550 & n1564 ) ;
  assign n1635 = ( n1524 & ~n1565 ) | ( n1524 & n1634 ) | ( ~n1565 & n1634 ) ;
  assign n1636 = ( ~n1592 & n1618 ) | ( ~n1592 & n1632 ) | ( n1618 & n1632 ) ;
  assign n1637 = ( n1592 & ~n1633 ) | ( n1592 & n1636 ) | ( ~n1633 & n1636 ) ;
  assign n1638 = ( ~n1620 & n1622 ) | ( ~n1620 & n1631 ) | ( n1622 & n1631 ) ;
  assign n1639 = ( n1620 & ~n1632 ) | ( n1620 & n1638 ) | ( ~n1632 & n1638 ) ;
  assign n1640 = ( ~n1552 & n1554 ) | ( ~n1552 & n1563 ) | ( n1554 & n1563 ) ;
  assign n1641 = ( n1552 & ~n1564 ) | ( n1552 & n1640 ) | ( ~n1564 & n1640 ) ;
  assign n1642 = ( n1556 & n1558 ) | ( n1556 & ~n1562 ) | ( n1558 & ~n1562 ) ;
  assign n1643 = ( n1562 & ~n1563 ) | ( n1562 & n1642 ) | ( ~n1563 & n1642 ) ;
  assign n1644 = ( n1624 & n1626 ) | ( n1624 & ~n1630 ) | ( n1626 & ~n1630 ) ;
  assign n1645 = ( n1630 & ~n1631 ) | ( n1630 & n1644 ) | ( ~n1631 & n1644 ) ;
  assign n1646 = ( ~n1519 & n1521 ) | ( ~n1519 & n1560 ) | ( n1521 & n1560 ) ;
  assign n1647 = ( n1519 & ~n1561 ) | ( n1519 & n1646 ) | ( ~n1561 & n1646 ) ;
  assign n1648 = ( ~n1587 & n1589 ) | ( ~n1587 & n1628 ) | ( n1589 & n1628 ) ;
  assign n1649 = ( n1587 & ~n1629 ) | ( n1587 & n1648 ) | ( ~n1629 & n1648 ) ;
  assign n1650 = n1647 & n1649 ;
  assign n1651 = ( n1643 & n1645 ) | ( n1643 & n1650 ) | ( n1645 & n1650 ) ;
  assign n1652 = ( n1639 & n1641 ) | ( n1639 & n1651 ) | ( n1641 & n1651 ) ;
  assign n1653 = ( n1635 & n1637 ) | ( n1635 & n1652 ) | ( n1637 & n1652 ) ;
  assign n1654 = ( n1565 & n1633 ) | ( n1565 & n1653 ) | ( n1633 & n1653 ) ;
  assign n1655 = ( ~n1565 & n1633 ) | ( ~n1565 & n1653 ) | ( n1633 & n1653 ) ;
  assign n1656 = ( n1565 & ~n1654 ) | ( n1565 & n1655 ) | ( ~n1654 & n1655 ) ;
  assign n1657 = ( ~n1408 & n1476 ) | ( ~n1408 & n1496 ) | ( n1476 & n1496 ) ;
  assign n1658 = ( n1408 & ~n1497 ) | ( n1408 & n1657 ) | ( ~n1497 & n1657 ) ;
  assign n1659 = ( ~n1478 & n1480 ) | ( ~n1478 & n1495 ) | ( n1480 & n1495 ) ;
  assign n1660 = ( n1478 & ~n1496 ) | ( n1478 & n1659 ) | ( ~n1496 & n1659 ) ;
  assign n1661 = ( ~n1635 & n1637 ) | ( ~n1635 & n1652 ) | ( n1637 & n1652 ) ;
  assign n1662 = ( n1635 & ~n1653 ) | ( n1635 & n1661 ) | ( ~n1653 & n1661 ) ;
  assign n1663 = ( ~n1639 & n1641 ) | ( ~n1639 & n1651 ) | ( n1641 & n1651 ) ;
  assign n1664 = ( n1639 & ~n1652 ) | ( n1639 & n1663 ) | ( ~n1652 & n1663 ) ;
  assign n1665 = ( ~n1482 & n1484 ) | ( ~n1482 & n1494 ) | ( n1484 & n1494 ) ;
  assign n1666 = ( n1482 & ~n1495 ) | ( n1482 & n1665 ) | ( ~n1495 & n1665 ) ;
  assign n1667 = ( ~n1486 & n1488 ) | ( ~n1486 & n1493 ) | ( n1488 & n1493 ) ;
  assign n1668 = ( n1486 & ~n1494 ) | ( n1486 & n1667 ) | ( ~n1494 & n1667 ) ;
  assign n1669 = ( ~n1643 & n1645 ) | ( ~n1643 & n1650 ) | ( n1645 & n1650 ) ;
  assign n1670 = ( n1643 & ~n1651 ) | ( n1643 & n1669 ) | ( ~n1651 & n1669 ) ;
  assign n1671 = n1647 | n1649 ;
  assign n1672 = ~n1650 & n1671 ;
  assign n1673 = ( n1490 & n1492 ) | ( n1490 & n1672 ) | ( n1492 & n1672 ) ;
  assign n1674 = ~n1493 & n1673 ;
  assign n1675 = ( n1668 & n1670 ) | ( n1668 & n1674 ) | ( n1670 & n1674 ) ;
  assign n1676 = ( n1664 & n1666 ) | ( n1664 & n1675 ) | ( n1666 & n1675 ) ;
  assign n1677 = ( n1660 & n1662 ) | ( n1660 & n1676 ) | ( n1662 & n1676 ) ;
  assign n1678 = ( n1656 & n1658 ) | ( n1656 & n1677 ) | ( n1658 & n1677 ) ;
  assign n1679 = ( n1497 & n1654 ) | ( n1497 & n1678 ) | ( n1654 & n1678 ) ;
  assign n1680 = ( ~n1158 & n1315 ) | ( ~n1158 & n1339 ) | ( n1315 & n1339 ) ;
  assign n1681 = ( n1158 & ~n1340 ) | ( n1158 & n1680 ) | ( ~n1340 & n1680 ) ;
  assign n1682 = ( ~n1497 & n1654 ) | ( ~n1497 & n1678 ) | ( n1654 & n1678 ) ;
  assign n1683 = ( n1497 & ~n1679 ) | ( n1497 & n1682 ) | ( ~n1679 & n1682 ) ;
  assign n1684 = ( ~n1656 & n1658 ) | ( ~n1656 & n1677 ) | ( n1658 & n1677 ) ;
  assign n1685 = ( n1656 & ~n1678 ) | ( n1656 & n1684 ) | ( ~n1678 & n1684 ) ;
  assign n1686 = ( ~n1317 & n1319 ) | ( ~n1317 & n1338 ) | ( n1319 & n1338 ) ;
  assign n1687 = ( n1317 & ~n1339 ) | ( n1317 & n1686 ) | ( ~n1339 & n1686 ) ;
  assign n1688 = ( ~n1321 & n1323 ) | ( ~n1321 & n1337 ) | ( n1323 & n1337 ) ;
  assign n1689 = ( n1321 & ~n1338 ) | ( n1321 & n1688 ) | ( ~n1338 & n1688 ) ;
  assign n1690 = ( ~n1660 & n1662 ) | ( ~n1660 & n1676 ) | ( n1662 & n1676 ) ;
  assign n1691 = ( n1660 & ~n1677 ) | ( n1660 & n1690 ) | ( ~n1677 & n1690 ) ;
  assign n1692 = ( ~n1664 & n1666 ) | ( ~n1664 & n1675 ) | ( n1666 & n1675 ) ;
  assign n1693 = ( n1664 & ~n1676 ) | ( n1664 & n1692 ) | ( ~n1676 & n1692 ) ;
  assign n1694 = ( ~n1325 & n1327 ) | ( ~n1325 & n1336 ) | ( n1327 & n1336 ) ;
  assign n1695 = ( n1325 & ~n1337 ) | ( n1325 & n1694 ) | ( ~n1337 & n1694 ) ;
  assign n1696 = ( ~n1151 & n1153 ) | ( ~n1151 & n1333 ) | ( n1153 & n1333 ) ;
  assign n1697 = ( n1151 & ~n1334 ) | ( n1151 & n1696 ) | ( ~n1334 & n1696 ) ;
  assign n1698 = ( ~n1490 & n1492 ) | ( ~n1490 & n1672 ) | ( n1492 & n1672 ) ;
  assign n1699 = ( n1490 & ~n1673 ) | ( n1490 & n1698 ) | ( ~n1673 & n1698 ) ;
  assign n1700 = n1697 & n1699 ;
  assign n1701 = ( n1329 & n1331 ) | ( n1329 & ~n1335 ) | ( n1331 & ~n1335 ) ;
  assign n1702 = ( n1335 & ~n1336 ) | ( n1335 & n1701 ) | ( ~n1336 & n1701 ) ;
  assign n1703 = ( n1668 & n1670 ) | ( n1668 & ~n1674 ) | ( n1670 & ~n1674 ) ;
  assign n1704 = ( n1674 & ~n1675 ) | ( n1674 & n1703 ) | ( ~n1675 & n1703 ) ;
  assign n1705 = ( n1700 & n1702 ) | ( n1700 & n1704 ) | ( n1702 & n1704 ) ;
  assign n1706 = ( n1693 & n1695 ) | ( n1693 & n1705 ) | ( n1695 & n1705 ) ;
  assign n1707 = ( n1689 & n1691 ) | ( n1689 & n1706 ) | ( n1691 & n1706 ) ;
  assign n1708 = ( n1685 & n1687 ) | ( n1685 & n1707 ) | ( n1687 & n1707 ) ;
  assign n1709 = ( n1681 & n1683 ) | ( n1681 & n1708 ) | ( n1683 & n1708 ) ;
  assign n1710 = ( n1340 & n1679 ) | ( n1340 & n1709 ) | ( n1679 & n1709 ) ;
  assign n1711 = ( x268 & x269 ) | ( x268 & x270 ) | ( x269 & x270 ) ;
  assign n1712 = ( x265 & x266 ) | ( x265 & x267 ) | ( x266 & x267 ) ;
  assign n1713 = ( ~x268 & x269 ) | ( ~x268 & x270 ) | ( x269 & x270 ) ;
  assign n1714 = ( x268 & ~n1711 ) | ( x268 & n1713 ) | ( ~n1711 & n1713 ) ;
  assign n1715 = ( ~x265 & x266 ) | ( ~x265 & x267 ) | ( x266 & x267 ) ;
  assign n1716 = ( x265 & ~n1712 ) | ( x265 & n1715 ) | ( ~n1712 & n1715 ) ;
  assign n1717 = n1714 & n1716 ;
  assign n1718 = ( n1711 & n1712 ) | ( n1711 & n1717 ) | ( n1712 & n1717 ) ;
  assign n1719 = ( x259 & x260 ) | ( x259 & x261 ) | ( x260 & x261 ) ;
  assign n1720 = ( x262 & x263 ) | ( x262 & x264 ) | ( x263 & x264 ) ;
  assign n1721 = ( ~x262 & x263 ) | ( ~x262 & x264 ) | ( x263 & x264 ) ;
  assign n1722 = ( x262 & ~n1720 ) | ( x262 & n1721 ) | ( ~n1720 & n1721 ) ;
  assign n1723 = ( ~x259 & x260 ) | ( ~x259 & x261 ) | ( x260 & x261 ) ;
  assign n1724 = ( x259 & ~n1719 ) | ( x259 & n1723 ) | ( ~n1719 & n1723 ) ;
  assign n1725 = n1722 & n1724 ;
  assign n1726 = ( n1719 & n1720 ) | ( n1719 & n1725 ) | ( n1720 & n1725 ) ;
  assign n1727 = ( ~n1711 & n1712 ) | ( ~n1711 & n1717 ) | ( n1712 & n1717 ) ;
  assign n1728 = ( n1711 & ~n1718 ) | ( n1711 & n1727 ) | ( ~n1718 & n1727 ) ;
  assign n1729 = ( ~n1719 & n1720 ) | ( ~n1719 & n1725 ) | ( n1720 & n1725 ) ;
  assign n1730 = ( n1719 & ~n1726 ) | ( n1719 & n1729 ) | ( ~n1726 & n1729 ) ;
  assign n1731 = n1714 | n1716 ;
  assign n1732 = ~n1717 & n1731 ;
  assign n1733 = n1722 | n1724 ;
  assign n1734 = ~n1725 & n1733 ;
  assign n1735 = n1732 & n1734 ;
  assign n1736 = ( n1728 & n1730 ) | ( n1728 & n1735 ) | ( n1730 & n1735 ) ;
  assign n1737 = ( n1718 & n1726 ) | ( n1718 & n1736 ) | ( n1726 & n1736 ) ;
  assign n1738 = ( x256 & x257 ) | ( x256 & x258 ) | ( x257 & x258 ) ;
  assign n1739 = ( x253 & x254 ) | ( x253 & x255 ) | ( x254 & x255 ) ;
  assign n1740 = ( ~x256 & x257 ) | ( ~x256 & x258 ) | ( x257 & x258 ) ;
  assign n1741 = ( x256 & ~n1738 ) | ( x256 & n1740 ) | ( ~n1738 & n1740 ) ;
  assign n1742 = ( ~x253 & x254 ) | ( ~x253 & x255 ) | ( x254 & x255 ) ;
  assign n1743 = ( x253 & ~n1739 ) | ( x253 & n1742 ) | ( ~n1739 & n1742 ) ;
  assign n1744 = n1741 & n1743 ;
  assign n1745 = ( n1738 & n1739 ) | ( n1738 & n1744 ) | ( n1739 & n1744 ) ;
  assign n1746 = ( x247 & x248 ) | ( x247 & x249 ) | ( x248 & x249 ) ;
  assign n1747 = ( x250 & x251 ) | ( x250 & x252 ) | ( x251 & x252 ) ;
  assign n1748 = ( ~x250 & x251 ) | ( ~x250 & x252 ) | ( x251 & x252 ) ;
  assign n1749 = ( x250 & ~n1747 ) | ( x250 & n1748 ) | ( ~n1747 & n1748 ) ;
  assign n1750 = ( ~x247 & x248 ) | ( ~x247 & x249 ) | ( x248 & x249 ) ;
  assign n1751 = ( x247 & ~n1746 ) | ( x247 & n1750 ) | ( ~n1746 & n1750 ) ;
  assign n1752 = n1749 & n1751 ;
  assign n1753 = ( n1746 & n1747 ) | ( n1746 & n1752 ) | ( n1747 & n1752 ) ;
  assign n1754 = ( ~n1738 & n1739 ) | ( ~n1738 & n1744 ) | ( n1739 & n1744 ) ;
  assign n1755 = ( n1738 & ~n1745 ) | ( n1738 & n1754 ) | ( ~n1745 & n1754 ) ;
  assign n1756 = ( ~n1746 & n1747 ) | ( ~n1746 & n1752 ) | ( n1747 & n1752 ) ;
  assign n1757 = ( n1746 & ~n1753 ) | ( n1746 & n1756 ) | ( ~n1753 & n1756 ) ;
  assign n1758 = n1749 | n1751 ;
  assign n1759 = ~n1752 & n1758 ;
  assign n1760 = ( n1741 & n1743 ) | ( n1741 & n1759 ) | ( n1743 & n1759 ) ;
  assign n1761 = ~n1744 & n1760 ;
  assign n1762 = ( n1755 & n1757 ) | ( n1755 & n1761 ) | ( n1757 & n1761 ) ;
  assign n1763 = ( n1745 & n1753 ) | ( n1745 & n1762 ) | ( n1753 & n1762 ) ;
  assign n1764 = ( ~n1745 & n1753 ) | ( ~n1745 & n1762 ) | ( n1753 & n1762 ) ;
  assign n1765 = ( n1745 & ~n1763 ) | ( n1745 & n1764 ) | ( ~n1763 & n1764 ) ;
  assign n1766 = ( ~n1718 & n1726 ) | ( ~n1718 & n1736 ) | ( n1726 & n1736 ) ;
  assign n1767 = ( n1718 & ~n1737 ) | ( n1718 & n1766 ) | ( ~n1737 & n1766 ) ;
  assign n1768 = ( ~n1728 & n1730 ) | ( ~n1728 & n1735 ) | ( n1730 & n1735 ) ;
  assign n1769 = ( n1728 & ~n1736 ) | ( n1728 & n1768 ) | ( ~n1736 & n1768 ) ;
  assign n1770 = ( ~n1755 & n1757 ) | ( ~n1755 & n1761 ) | ( n1757 & n1761 ) ;
  assign n1771 = ( n1755 & ~n1762 ) | ( n1755 & n1770 ) | ( ~n1762 & n1770 ) ;
  assign n1772 = ( ~n1741 & n1743 ) | ( ~n1741 & n1759 ) | ( n1743 & n1759 ) ;
  assign n1773 = ( n1741 & ~n1760 ) | ( n1741 & n1772 ) | ( ~n1760 & n1772 ) ;
  assign n1774 = ( n1732 & n1734 ) | ( n1732 & n1773 ) | ( n1734 & n1773 ) ;
  assign n1775 = ~n1735 & n1774 ;
  assign n1776 = ( n1769 & n1771 ) | ( n1769 & n1775 ) | ( n1771 & n1775 ) ;
  assign n1777 = ( n1765 & n1767 ) | ( n1765 & n1776 ) | ( n1767 & n1776 ) ;
  assign n1778 = ( n1737 & n1763 ) | ( n1737 & n1777 ) | ( n1763 & n1777 ) ;
  assign n1779 = ( x244 & x245 ) | ( x244 & x246 ) | ( x245 & x246 ) ;
  assign n1780 = ( x241 & x242 ) | ( x241 & x243 ) | ( x242 & x243 ) ;
  assign n1781 = ( ~x244 & x245 ) | ( ~x244 & x246 ) | ( x245 & x246 ) ;
  assign n1782 = ( x244 & ~n1779 ) | ( x244 & n1781 ) | ( ~n1779 & n1781 ) ;
  assign n1783 = ( ~x241 & x242 ) | ( ~x241 & x243 ) | ( x242 & x243 ) ;
  assign n1784 = ( x241 & ~n1780 ) | ( x241 & n1783 ) | ( ~n1780 & n1783 ) ;
  assign n1785 = n1782 & n1784 ;
  assign n1786 = ( n1779 & n1780 ) | ( n1779 & n1785 ) | ( n1780 & n1785 ) ;
  assign n1787 = ( x235 & x236 ) | ( x235 & x237 ) | ( x236 & x237 ) ;
  assign n1788 = ( x238 & x239 ) | ( x238 & x240 ) | ( x239 & x240 ) ;
  assign n1789 = ( ~x238 & x239 ) | ( ~x238 & x240 ) | ( x239 & x240 ) ;
  assign n1790 = ( x238 & ~n1788 ) | ( x238 & n1789 ) | ( ~n1788 & n1789 ) ;
  assign n1791 = ( ~x235 & x236 ) | ( ~x235 & x237 ) | ( x236 & x237 ) ;
  assign n1792 = ( x235 & ~n1787 ) | ( x235 & n1791 ) | ( ~n1787 & n1791 ) ;
  assign n1793 = n1790 & n1792 ;
  assign n1794 = ( n1787 & n1788 ) | ( n1787 & n1793 ) | ( n1788 & n1793 ) ;
  assign n1795 = ( ~n1779 & n1780 ) | ( ~n1779 & n1785 ) | ( n1780 & n1785 ) ;
  assign n1796 = ( n1779 & ~n1786 ) | ( n1779 & n1795 ) | ( ~n1786 & n1795 ) ;
  assign n1797 = ( ~n1787 & n1788 ) | ( ~n1787 & n1793 ) | ( n1788 & n1793 ) ;
  assign n1798 = ( n1787 & ~n1794 ) | ( n1787 & n1797 ) | ( ~n1794 & n1797 ) ;
  assign n1799 = n1782 | n1784 ;
  assign n1800 = ~n1785 & n1799 ;
  assign n1801 = n1790 | n1792 ;
  assign n1802 = ~n1793 & n1801 ;
  assign n1803 = n1800 & n1802 ;
  assign n1804 = ( n1796 & n1798 ) | ( n1796 & n1803 ) | ( n1798 & n1803 ) ;
  assign n1805 = ( n1786 & n1794 ) | ( n1786 & n1804 ) | ( n1794 & n1804 ) ;
  assign n1806 = ( x232 & x233 ) | ( x232 & x234 ) | ( x233 & x234 ) ;
  assign n1807 = ( x229 & x230 ) | ( x229 & x231 ) | ( x230 & x231 ) ;
  assign n1808 = ( ~x232 & x233 ) | ( ~x232 & x234 ) | ( x233 & x234 ) ;
  assign n1809 = ( x232 & ~n1806 ) | ( x232 & n1808 ) | ( ~n1806 & n1808 ) ;
  assign n1810 = ( ~x229 & x230 ) | ( ~x229 & x231 ) | ( x230 & x231 ) ;
  assign n1811 = ( x229 & ~n1807 ) | ( x229 & n1810 ) | ( ~n1807 & n1810 ) ;
  assign n1812 = n1809 & n1811 ;
  assign n1813 = ( n1806 & n1807 ) | ( n1806 & n1812 ) | ( n1807 & n1812 ) ;
  assign n1814 = ( x223 & x224 ) | ( x223 & x225 ) | ( x224 & x225 ) ;
  assign n1815 = ( x226 & x227 ) | ( x226 & x228 ) | ( x227 & x228 ) ;
  assign n1816 = ( ~x226 & x227 ) | ( ~x226 & x228 ) | ( x227 & x228 ) ;
  assign n1817 = ( x226 & ~n1815 ) | ( x226 & n1816 ) | ( ~n1815 & n1816 ) ;
  assign n1818 = ( ~x223 & x224 ) | ( ~x223 & x225 ) | ( x224 & x225 ) ;
  assign n1819 = ( x223 & ~n1814 ) | ( x223 & n1818 ) | ( ~n1814 & n1818 ) ;
  assign n1820 = n1817 & n1819 ;
  assign n1821 = ( n1814 & n1815 ) | ( n1814 & n1820 ) | ( n1815 & n1820 ) ;
  assign n1822 = ( ~n1806 & n1807 ) | ( ~n1806 & n1812 ) | ( n1807 & n1812 ) ;
  assign n1823 = ( n1806 & ~n1813 ) | ( n1806 & n1822 ) | ( ~n1813 & n1822 ) ;
  assign n1824 = ( ~n1814 & n1815 ) | ( ~n1814 & n1820 ) | ( n1815 & n1820 ) ;
  assign n1825 = ( n1814 & ~n1821 ) | ( n1814 & n1824 ) | ( ~n1821 & n1824 ) ;
  assign n1826 = n1817 | n1819 ;
  assign n1827 = ~n1820 & n1826 ;
  assign n1828 = ( n1809 & n1811 ) | ( n1809 & n1827 ) | ( n1811 & n1827 ) ;
  assign n1829 = ~n1812 & n1828 ;
  assign n1830 = ( n1823 & n1825 ) | ( n1823 & n1829 ) | ( n1825 & n1829 ) ;
  assign n1831 = ( n1813 & n1821 ) | ( n1813 & n1830 ) | ( n1821 & n1830 ) ;
  assign n1832 = ( ~n1813 & n1821 ) | ( ~n1813 & n1830 ) | ( n1821 & n1830 ) ;
  assign n1833 = ( n1813 & ~n1831 ) | ( n1813 & n1832 ) | ( ~n1831 & n1832 ) ;
  assign n1834 = ( ~n1786 & n1794 ) | ( ~n1786 & n1804 ) | ( n1794 & n1804 ) ;
  assign n1835 = ( n1786 & ~n1805 ) | ( n1786 & n1834 ) | ( ~n1805 & n1834 ) ;
  assign n1836 = ( ~n1796 & n1798 ) | ( ~n1796 & n1803 ) | ( n1798 & n1803 ) ;
  assign n1837 = ( n1796 & ~n1804 ) | ( n1796 & n1836 ) | ( ~n1804 & n1836 ) ;
  assign n1838 = ( ~n1823 & n1825 ) | ( ~n1823 & n1829 ) | ( n1825 & n1829 ) ;
  assign n1839 = ( n1823 & ~n1830 ) | ( n1823 & n1838 ) | ( ~n1830 & n1838 ) ;
  assign n1840 = ( ~n1809 & n1811 ) | ( ~n1809 & n1827 ) | ( n1811 & n1827 ) ;
  assign n1841 = ( n1809 & ~n1828 ) | ( n1809 & n1840 ) | ( ~n1828 & n1840 ) ;
  assign n1842 = ( n1800 & n1802 ) | ( n1800 & n1841 ) | ( n1802 & n1841 ) ;
  assign n1843 = ~n1803 & n1842 ;
  assign n1844 = ( n1837 & n1839 ) | ( n1837 & n1843 ) | ( n1839 & n1843 ) ;
  assign n1845 = ( n1833 & n1835 ) | ( n1833 & n1844 ) | ( n1835 & n1844 ) ;
  assign n1846 = ( n1805 & n1831 ) | ( n1805 & n1845 ) | ( n1831 & n1845 ) ;
  assign n1847 = ( ~n1737 & n1763 ) | ( ~n1737 & n1777 ) | ( n1763 & n1777 ) ;
  assign n1848 = ( n1737 & ~n1778 ) | ( n1737 & n1847 ) | ( ~n1778 & n1847 ) ;
  assign n1849 = ( ~n1805 & n1831 ) | ( ~n1805 & n1845 ) | ( n1831 & n1845 ) ;
  assign n1850 = ( n1805 & ~n1846 ) | ( n1805 & n1849 ) | ( ~n1846 & n1849 ) ;
  assign n1851 = ( ~n1833 & n1835 ) | ( ~n1833 & n1844 ) | ( n1835 & n1844 ) ;
  assign n1852 = ( n1833 & ~n1845 ) | ( n1833 & n1851 ) | ( ~n1845 & n1851 ) ;
  assign n1853 = ( ~n1765 & n1767 ) | ( ~n1765 & n1776 ) | ( n1767 & n1776 ) ;
  assign n1854 = ( n1765 & ~n1777 ) | ( n1765 & n1853 ) | ( ~n1777 & n1853 ) ;
  assign n1855 = ( n1769 & n1771 ) | ( n1769 & ~n1775 ) | ( n1771 & ~n1775 ) ;
  assign n1856 = ( n1775 & ~n1776 ) | ( n1775 & n1855 ) | ( ~n1776 & n1855 ) ;
  assign n1857 = ( n1837 & n1839 ) | ( n1837 & ~n1843 ) | ( n1839 & ~n1843 ) ;
  assign n1858 = ( n1843 & ~n1844 ) | ( n1843 & n1857 ) | ( ~n1844 & n1857 ) ;
  assign n1859 = ( ~n1732 & n1734 ) | ( ~n1732 & n1773 ) | ( n1734 & n1773 ) ;
  assign n1860 = ( n1732 & ~n1774 ) | ( n1732 & n1859 ) | ( ~n1774 & n1859 ) ;
  assign n1861 = ( ~n1800 & n1802 ) | ( ~n1800 & n1841 ) | ( n1802 & n1841 ) ;
  assign n1862 = ( n1800 & ~n1842 ) | ( n1800 & n1861 ) | ( ~n1842 & n1861 ) ;
  assign n1863 = n1860 & n1862 ;
  assign n1864 = ( n1856 & n1858 ) | ( n1856 & n1863 ) | ( n1858 & n1863 ) ;
  assign n1865 = ( n1852 & n1854 ) | ( n1852 & n1864 ) | ( n1854 & n1864 ) ;
  assign n1866 = ( n1848 & n1850 ) | ( n1848 & n1865 ) | ( n1850 & n1865 ) ;
  assign n1867 = ( n1778 & n1846 ) | ( n1778 & n1866 ) | ( n1846 & n1866 ) ;
  assign n1868 = ( x220 & x221 ) | ( x220 & x222 ) | ( x221 & x222 ) ;
  assign n1869 = ( x217 & x218 ) | ( x217 & x219 ) | ( x218 & x219 ) ;
  assign n1870 = ( ~x220 & x221 ) | ( ~x220 & x222 ) | ( x221 & x222 ) ;
  assign n1871 = ( x220 & ~n1868 ) | ( x220 & n1870 ) | ( ~n1868 & n1870 ) ;
  assign n1872 = ( ~x217 & x218 ) | ( ~x217 & x219 ) | ( x218 & x219 ) ;
  assign n1873 = ( x217 & ~n1869 ) | ( x217 & n1872 ) | ( ~n1869 & n1872 ) ;
  assign n1874 = n1871 & n1873 ;
  assign n1875 = ( n1868 & n1869 ) | ( n1868 & n1874 ) | ( n1869 & n1874 ) ;
  assign n1876 = ( x211 & x212 ) | ( x211 & x213 ) | ( x212 & x213 ) ;
  assign n1877 = ( x214 & x215 ) | ( x214 & x216 ) | ( x215 & x216 ) ;
  assign n1878 = ( ~x214 & x215 ) | ( ~x214 & x216 ) | ( x215 & x216 ) ;
  assign n1879 = ( x214 & ~n1877 ) | ( x214 & n1878 ) | ( ~n1877 & n1878 ) ;
  assign n1880 = ( ~x211 & x212 ) | ( ~x211 & x213 ) | ( x212 & x213 ) ;
  assign n1881 = ( x211 & ~n1876 ) | ( x211 & n1880 ) | ( ~n1876 & n1880 ) ;
  assign n1882 = n1879 & n1881 ;
  assign n1883 = ( n1876 & n1877 ) | ( n1876 & n1882 ) | ( n1877 & n1882 ) ;
  assign n1884 = ( ~n1868 & n1869 ) | ( ~n1868 & n1874 ) | ( n1869 & n1874 ) ;
  assign n1885 = ( n1868 & ~n1875 ) | ( n1868 & n1884 ) | ( ~n1875 & n1884 ) ;
  assign n1886 = ( ~n1876 & n1877 ) | ( ~n1876 & n1882 ) | ( n1877 & n1882 ) ;
  assign n1887 = ( n1876 & ~n1883 ) | ( n1876 & n1886 ) | ( ~n1883 & n1886 ) ;
  assign n1888 = n1871 | n1873 ;
  assign n1889 = ~n1874 & n1888 ;
  assign n1890 = n1879 | n1881 ;
  assign n1891 = ~n1882 & n1890 ;
  assign n1892 = n1889 & n1891 ;
  assign n1893 = ( n1885 & n1887 ) | ( n1885 & n1892 ) | ( n1887 & n1892 ) ;
  assign n1894 = ( n1875 & n1883 ) | ( n1875 & n1893 ) | ( n1883 & n1893 ) ;
  assign n1895 = ( x208 & x209 ) | ( x208 & x210 ) | ( x209 & x210 ) ;
  assign n1896 = ( x205 & x206 ) | ( x205 & x207 ) | ( x206 & x207 ) ;
  assign n1897 = ( ~x208 & x209 ) | ( ~x208 & x210 ) | ( x209 & x210 ) ;
  assign n1898 = ( x208 & ~n1895 ) | ( x208 & n1897 ) | ( ~n1895 & n1897 ) ;
  assign n1899 = ( ~x205 & x206 ) | ( ~x205 & x207 ) | ( x206 & x207 ) ;
  assign n1900 = ( x205 & ~n1896 ) | ( x205 & n1899 ) | ( ~n1896 & n1899 ) ;
  assign n1901 = n1898 & n1900 ;
  assign n1902 = ( n1895 & n1896 ) | ( n1895 & n1901 ) | ( n1896 & n1901 ) ;
  assign n1903 = ( x199 & x200 ) | ( x199 & x201 ) | ( x200 & x201 ) ;
  assign n1904 = ( x202 & x203 ) | ( x202 & x204 ) | ( x203 & x204 ) ;
  assign n1905 = ( ~x202 & x203 ) | ( ~x202 & x204 ) | ( x203 & x204 ) ;
  assign n1906 = ( x202 & ~n1904 ) | ( x202 & n1905 ) | ( ~n1904 & n1905 ) ;
  assign n1907 = ( ~x199 & x200 ) | ( ~x199 & x201 ) | ( x200 & x201 ) ;
  assign n1908 = ( x199 & ~n1903 ) | ( x199 & n1907 ) | ( ~n1903 & n1907 ) ;
  assign n1909 = n1906 & n1908 ;
  assign n1910 = ( n1903 & n1904 ) | ( n1903 & n1909 ) | ( n1904 & n1909 ) ;
  assign n1911 = ( ~n1895 & n1896 ) | ( ~n1895 & n1901 ) | ( n1896 & n1901 ) ;
  assign n1912 = ( n1895 & ~n1902 ) | ( n1895 & n1911 ) | ( ~n1902 & n1911 ) ;
  assign n1913 = ( ~n1903 & n1904 ) | ( ~n1903 & n1909 ) | ( n1904 & n1909 ) ;
  assign n1914 = ( n1903 & ~n1910 ) | ( n1903 & n1913 ) | ( ~n1910 & n1913 ) ;
  assign n1915 = n1906 | n1908 ;
  assign n1916 = ~n1909 & n1915 ;
  assign n1917 = ( n1898 & n1900 ) | ( n1898 & n1916 ) | ( n1900 & n1916 ) ;
  assign n1918 = ~n1901 & n1917 ;
  assign n1919 = ( n1912 & n1914 ) | ( n1912 & n1918 ) | ( n1914 & n1918 ) ;
  assign n1920 = ( n1902 & n1910 ) | ( n1902 & n1919 ) | ( n1910 & n1919 ) ;
  assign n1921 = ( ~n1902 & n1910 ) | ( ~n1902 & n1919 ) | ( n1910 & n1919 ) ;
  assign n1922 = ( n1902 & ~n1920 ) | ( n1902 & n1921 ) | ( ~n1920 & n1921 ) ;
  assign n1923 = ( ~n1875 & n1883 ) | ( ~n1875 & n1893 ) | ( n1883 & n1893 ) ;
  assign n1924 = ( n1875 & ~n1894 ) | ( n1875 & n1923 ) | ( ~n1894 & n1923 ) ;
  assign n1925 = ( ~n1885 & n1887 ) | ( ~n1885 & n1892 ) | ( n1887 & n1892 ) ;
  assign n1926 = ( n1885 & ~n1893 ) | ( n1885 & n1925 ) | ( ~n1893 & n1925 ) ;
  assign n1927 = ( ~n1912 & n1914 ) | ( ~n1912 & n1918 ) | ( n1914 & n1918 ) ;
  assign n1928 = ( n1912 & ~n1919 ) | ( n1912 & n1927 ) | ( ~n1919 & n1927 ) ;
  assign n1929 = ( ~n1898 & n1900 ) | ( ~n1898 & n1916 ) | ( n1900 & n1916 ) ;
  assign n1930 = ( n1898 & ~n1917 ) | ( n1898 & n1929 ) | ( ~n1917 & n1929 ) ;
  assign n1931 = ( n1889 & n1891 ) | ( n1889 & n1930 ) | ( n1891 & n1930 ) ;
  assign n1932 = ~n1892 & n1931 ;
  assign n1933 = ( n1926 & n1928 ) | ( n1926 & n1932 ) | ( n1928 & n1932 ) ;
  assign n1934 = ( n1922 & n1924 ) | ( n1922 & n1933 ) | ( n1924 & n1933 ) ;
  assign n1935 = ( n1894 & n1920 ) | ( n1894 & n1934 ) | ( n1920 & n1934 ) ;
  assign n1936 = ( x196 & x197 ) | ( x196 & x198 ) | ( x197 & x198 ) ;
  assign n1937 = ( x193 & x194 ) | ( x193 & x195 ) | ( x194 & x195 ) ;
  assign n1938 = ( ~x196 & x197 ) | ( ~x196 & x198 ) | ( x197 & x198 ) ;
  assign n1939 = ( x196 & ~n1936 ) | ( x196 & n1938 ) | ( ~n1936 & n1938 ) ;
  assign n1940 = ( ~x193 & x194 ) | ( ~x193 & x195 ) | ( x194 & x195 ) ;
  assign n1941 = ( x193 & ~n1937 ) | ( x193 & n1940 ) | ( ~n1937 & n1940 ) ;
  assign n1942 = n1939 & n1941 ;
  assign n1943 = ( n1936 & n1937 ) | ( n1936 & n1942 ) | ( n1937 & n1942 ) ;
  assign n1944 = ( x187 & x188 ) | ( x187 & x189 ) | ( x188 & x189 ) ;
  assign n1945 = ( x190 & x191 ) | ( x190 & x192 ) | ( x191 & x192 ) ;
  assign n1946 = ( ~x190 & x191 ) | ( ~x190 & x192 ) | ( x191 & x192 ) ;
  assign n1947 = ( x190 & ~n1945 ) | ( x190 & n1946 ) | ( ~n1945 & n1946 ) ;
  assign n1948 = ( ~x187 & x188 ) | ( ~x187 & x189 ) | ( x188 & x189 ) ;
  assign n1949 = ( x187 & ~n1944 ) | ( x187 & n1948 ) | ( ~n1944 & n1948 ) ;
  assign n1950 = n1947 & n1949 ;
  assign n1951 = ( n1944 & n1945 ) | ( n1944 & n1950 ) | ( n1945 & n1950 ) ;
  assign n1952 = ( ~n1936 & n1937 ) | ( ~n1936 & n1942 ) | ( n1937 & n1942 ) ;
  assign n1953 = ( n1936 & ~n1943 ) | ( n1936 & n1952 ) | ( ~n1943 & n1952 ) ;
  assign n1954 = ( ~n1944 & n1945 ) | ( ~n1944 & n1950 ) | ( n1945 & n1950 ) ;
  assign n1955 = ( n1944 & ~n1951 ) | ( n1944 & n1954 ) | ( ~n1951 & n1954 ) ;
  assign n1956 = n1939 | n1941 ;
  assign n1957 = ~n1942 & n1956 ;
  assign n1958 = n1947 | n1949 ;
  assign n1959 = ~n1950 & n1958 ;
  assign n1960 = n1957 & n1959 ;
  assign n1961 = ( n1953 & n1955 ) | ( n1953 & n1960 ) | ( n1955 & n1960 ) ;
  assign n1962 = ( n1943 & n1951 ) | ( n1943 & n1961 ) | ( n1951 & n1961 ) ;
  assign n1963 = ( x184 & x185 ) | ( x184 & x186 ) | ( x185 & x186 ) ;
  assign n1964 = ( x181 & x182 ) | ( x181 & x183 ) | ( x182 & x183 ) ;
  assign n1965 = ( ~x184 & x185 ) | ( ~x184 & x186 ) | ( x185 & x186 ) ;
  assign n1966 = ( x184 & ~n1963 ) | ( x184 & n1965 ) | ( ~n1963 & n1965 ) ;
  assign n1967 = ( ~x181 & x182 ) | ( ~x181 & x183 ) | ( x182 & x183 ) ;
  assign n1968 = ( x181 & ~n1964 ) | ( x181 & n1967 ) | ( ~n1964 & n1967 ) ;
  assign n1969 = n1966 & n1968 ;
  assign n1970 = ( n1963 & n1964 ) | ( n1963 & n1969 ) | ( n1964 & n1969 ) ;
  assign n1971 = ( x175 & x176 ) | ( x175 & x177 ) | ( x176 & x177 ) ;
  assign n1972 = ( x178 & x179 ) | ( x178 & x180 ) | ( x179 & x180 ) ;
  assign n1973 = ( ~x178 & x179 ) | ( ~x178 & x180 ) | ( x179 & x180 ) ;
  assign n1974 = ( x178 & ~n1972 ) | ( x178 & n1973 ) | ( ~n1972 & n1973 ) ;
  assign n1975 = ( ~x175 & x176 ) | ( ~x175 & x177 ) | ( x176 & x177 ) ;
  assign n1976 = ( x175 & ~n1971 ) | ( x175 & n1975 ) | ( ~n1971 & n1975 ) ;
  assign n1977 = n1974 & n1976 ;
  assign n1978 = ( n1971 & n1972 ) | ( n1971 & n1977 ) | ( n1972 & n1977 ) ;
  assign n1979 = ( ~n1963 & n1964 ) | ( ~n1963 & n1969 ) | ( n1964 & n1969 ) ;
  assign n1980 = ( n1963 & ~n1970 ) | ( n1963 & n1979 ) | ( ~n1970 & n1979 ) ;
  assign n1981 = ( ~n1971 & n1972 ) | ( ~n1971 & n1977 ) | ( n1972 & n1977 ) ;
  assign n1982 = ( n1971 & ~n1978 ) | ( n1971 & n1981 ) | ( ~n1978 & n1981 ) ;
  assign n1983 = n1974 | n1976 ;
  assign n1984 = ~n1977 & n1983 ;
  assign n1985 = ( n1966 & n1968 ) | ( n1966 & n1984 ) | ( n1968 & n1984 ) ;
  assign n1986 = ~n1969 & n1985 ;
  assign n1987 = ( n1980 & n1982 ) | ( n1980 & n1986 ) | ( n1982 & n1986 ) ;
  assign n1988 = ( n1970 & n1978 ) | ( n1970 & n1987 ) | ( n1978 & n1987 ) ;
  assign n1989 = ( ~n1970 & n1978 ) | ( ~n1970 & n1987 ) | ( n1978 & n1987 ) ;
  assign n1990 = ( n1970 & ~n1988 ) | ( n1970 & n1989 ) | ( ~n1988 & n1989 ) ;
  assign n1991 = ( ~n1943 & n1951 ) | ( ~n1943 & n1961 ) | ( n1951 & n1961 ) ;
  assign n1992 = ( n1943 & ~n1962 ) | ( n1943 & n1991 ) | ( ~n1962 & n1991 ) ;
  assign n1993 = ( ~n1953 & n1955 ) | ( ~n1953 & n1960 ) | ( n1955 & n1960 ) ;
  assign n1994 = ( n1953 & ~n1961 ) | ( n1953 & n1993 ) | ( ~n1961 & n1993 ) ;
  assign n1995 = ( ~n1980 & n1982 ) | ( ~n1980 & n1986 ) | ( n1982 & n1986 ) ;
  assign n1996 = ( n1980 & ~n1987 ) | ( n1980 & n1995 ) | ( ~n1987 & n1995 ) ;
  assign n1997 = ( ~n1966 & n1968 ) | ( ~n1966 & n1984 ) | ( n1968 & n1984 ) ;
  assign n1998 = ( n1966 & ~n1985 ) | ( n1966 & n1997 ) | ( ~n1985 & n1997 ) ;
  assign n1999 = ( n1957 & n1959 ) | ( n1957 & n1998 ) | ( n1959 & n1998 ) ;
  assign n2000 = ~n1960 & n1999 ;
  assign n2001 = ( n1994 & n1996 ) | ( n1994 & n2000 ) | ( n1996 & n2000 ) ;
  assign n2002 = ( n1990 & n1992 ) | ( n1990 & n2001 ) | ( n1992 & n2001 ) ;
  assign n2003 = ( n1962 & n1988 ) | ( n1962 & n2002 ) | ( n1988 & n2002 ) ;
  assign n2004 = ( ~n1894 & n1920 ) | ( ~n1894 & n1934 ) | ( n1920 & n1934 ) ;
  assign n2005 = ( n1894 & ~n1935 ) | ( n1894 & n2004 ) | ( ~n1935 & n2004 ) ;
  assign n2006 = ( ~n1962 & n1988 ) | ( ~n1962 & n2002 ) | ( n1988 & n2002 ) ;
  assign n2007 = ( n1962 & ~n2003 ) | ( n1962 & n2006 ) | ( ~n2003 & n2006 ) ;
  assign n2008 = ( ~n1990 & n1992 ) | ( ~n1990 & n2001 ) | ( n1992 & n2001 ) ;
  assign n2009 = ( n1990 & ~n2002 ) | ( n1990 & n2008 ) | ( ~n2002 & n2008 ) ;
  assign n2010 = ( ~n1922 & n1924 ) | ( ~n1922 & n1933 ) | ( n1924 & n1933 ) ;
  assign n2011 = ( n1922 & ~n1934 ) | ( n1922 & n2010 ) | ( ~n1934 & n2010 ) ;
  assign n2012 = ( n1926 & n1928 ) | ( n1926 & ~n1932 ) | ( n1928 & ~n1932 ) ;
  assign n2013 = ( n1932 & ~n1933 ) | ( n1932 & n2012 ) | ( ~n1933 & n2012 ) ;
  assign n2014 = ( n1994 & n1996 ) | ( n1994 & ~n2000 ) | ( n1996 & ~n2000 ) ;
  assign n2015 = ( n2000 & ~n2001 ) | ( n2000 & n2014 ) | ( ~n2001 & n2014 ) ;
  assign n2016 = ( ~n1889 & n1891 ) | ( ~n1889 & n1930 ) | ( n1891 & n1930 ) ;
  assign n2017 = ( n1889 & ~n1931 ) | ( n1889 & n2016 ) | ( ~n1931 & n2016 ) ;
  assign n2018 = ( ~n1957 & n1959 ) | ( ~n1957 & n1998 ) | ( n1959 & n1998 ) ;
  assign n2019 = ( n1957 & ~n1999 ) | ( n1957 & n2018 ) | ( ~n1999 & n2018 ) ;
  assign n2020 = n2017 & n2019 ;
  assign n2021 = ( n2013 & n2015 ) | ( n2013 & n2020 ) | ( n2015 & n2020 ) ;
  assign n2022 = ( n2009 & n2011 ) | ( n2009 & n2021 ) | ( n2011 & n2021 ) ;
  assign n2023 = ( n2005 & n2007 ) | ( n2005 & n2022 ) | ( n2007 & n2022 ) ;
  assign n2024 = ( n1935 & n2003 ) | ( n1935 & n2023 ) | ( n2003 & n2023 ) ;
  assign n2025 = ( ~n1935 & n2003 ) | ( ~n1935 & n2023 ) | ( n2003 & n2023 ) ;
  assign n2026 = ( n1935 & ~n2024 ) | ( n1935 & n2025 ) | ( ~n2024 & n2025 ) ;
  assign n2027 = ( ~n1778 & n1846 ) | ( ~n1778 & n1866 ) | ( n1846 & n1866 ) ;
  assign n2028 = ( n1778 & ~n1867 ) | ( n1778 & n2027 ) | ( ~n1867 & n2027 ) ;
  assign n2029 = ( ~n1848 & n1850 ) | ( ~n1848 & n1865 ) | ( n1850 & n1865 ) ;
  assign n2030 = ( n1848 & ~n1866 ) | ( n1848 & n2029 ) | ( ~n1866 & n2029 ) ;
  assign n2031 = ( ~n2005 & n2007 ) | ( ~n2005 & n2022 ) | ( n2007 & n2022 ) ;
  assign n2032 = ( n2005 & ~n2023 ) | ( n2005 & n2031 ) | ( ~n2023 & n2031 ) ;
  assign n2033 = ( ~n2009 & n2011 ) | ( ~n2009 & n2021 ) | ( n2011 & n2021 ) ;
  assign n2034 = ( n2009 & ~n2022 ) | ( n2009 & n2033 ) | ( ~n2022 & n2033 ) ;
  assign n2035 = ( ~n1852 & n1854 ) | ( ~n1852 & n1864 ) | ( n1854 & n1864 ) ;
  assign n2036 = ( n1852 & ~n1865 ) | ( n1852 & n2035 ) | ( ~n1865 & n2035 ) ;
  assign n2037 = ( ~n1856 & n1858 ) | ( ~n1856 & n1863 ) | ( n1858 & n1863 ) ;
  assign n2038 = ( n1856 & ~n1864 ) | ( n1856 & n2037 ) | ( ~n1864 & n2037 ) ;
  assign n2039 = ( ~n2013 & n2015 ) | ( ~n2013 & n2020 ) | ( n2015 & n2020 ) ;
  assign n2040 = ( n2013 & ~n2021 ) | ( n2013 & n2039 ) | ( ~n2021 & n2039 ) ;
  assign n2041 = n2017 | n2019 ;
  assign n2042 = ~n2020 & n2041 ;
  assign n2043 = ( n1860 & n1862 ) | ( n1860 & n2042 ) | ( n1862 & n2042 ) ;
  assign n2044 = ~n1863 & n2043 ;
  assign n2045 = ( n2038 & n2040 ) | ( n2038 & n2044 ) | ( n2040 & n2044 ) ;
  assign n2046 = ( n2034 & n2036 ) | ( n2034 & n2045 ) | ( n2036 & n2045 ) ;
  assign n2047 = ( n2030 & n2032 ) | ( n2030 & n2046 ) | ( n2032 & n2046 ) ;
  assign n2048 = ( n2026 & n2028 ) | ( n2026 & n2047 ) | ( n2028 & n2047 ) ;
  assign n2049 = ( n1867 & n2024 ) | ( n1867 & n2048 ) | ( n2024 & n2048 ) ;
  assign n2050 = ( x172 & x173 ) | ( x172 & x174 ) | ( x173 & x174 ) ;
  assign n2051 = ( x169 & x170 ) | ( x169 & x171 ) | ( x170 & x171 ) ;
  assign n2052 = ( ~x172 & x173 ) | ( ~x172 & x174 ) | ( x173 & x174 ) ;
  assign n2053 = ( x172 & ~n2050 ) | ( x172 & n2052 ) | ( ~n2050 & n2052 ) ;
  assign n2054 = ( ~x169 & x170 ) | ( ~x169 & x171 ) | ( x170 & x171 ) ;
  assign n2055 = ( x169 & ~n2051 ) | ( x169 & n2054 ) | ( ~n2051 & n2054 ) ;
  assign n2056 = n2053 & n2055 ;
  assign n2057 = ( n2050 & n2051 ) | ( n2050 & n2056 ) | ( n2051 & n2056 ) ;
  assign n2058 = ( x163 & x164 ) | ( x163 & x165 ) | ( x164 & x165 ) ;
  assign n2059 = ( x166 & x167 ) | ( x166 & x168 ) | ( x167 & x168 ) ;
  assign n2060 = ( ~x166 & x167 ) | ( ~x166 & x168 ) | ( x167 & x168 ) ;
  assign n2061 = ( x166 & ~n2059 ) | ( x166 & n2060 ) | ( ~n2059 & n2060 ) ;
  assign n2062 = ( ~x163 & x164 ) | ( ~x163 & x165 ) | ( x164 & x165 ) ;
  assign n2063 = ( x163 & ~n2058 ) | ( x163 & n2062 ) | ( ~n2058 & n2062 ) ;
  assign n2064 = n2061 & n2063 ;
  assign n2065 = ( n2058 & n2059 ) | ( n2058 & n2064 ) | ( n2059 & n2064 ) ;
  assign n2066 = ( ~n2050 & n2051 ) | ( ~n2050 & n2056 ) | ( n2051 & n2056 ) ;
  assign n2067 = ( n2050 & ~n2057 ) | ( n2050 & n2066 ) | ( ~n2057 & n2066 ) ;
  assign n2068 = ( ~n2058 & n2059 ) | ( ~n2058 & n2064 ) | ( n2059 & n2064 ) ;
  assign n2069 = ( n2058 & ~n2065 ) | ( n2058 & n2068 ) | ( ~n2065 & n2068 ) ;
  assign n2070 = n2053 | n2055 ;
  assign n2071 = ~n2056 & n2070 ;
  assign n2072 = n2061 | n2063 ;
  assign n2073 = ~n2064 & n2072 ;
  assign n2074 = n2071 & n2073 ;
  assign n2075 = ( n2067 & n2069 ) | ( n2067 & n2074 ) | ( n2069 & n2074 ) ;
  assign n2076 = ( n2057 & n2065 ) | ( n2057 & n2075 ) | ( n2065 & n2075 ) ;
  assign n2077 = ( x160 & x161 ) | ( x160 & x162 ) | ( x161 & x162 ) ;
  assign n2078 = ( x157 & x158 ) | ( x157 & x159 ) | ( x158 & x159 ) ;
  assign n2079 = ( ~x160 & x161 ) | ( ~x160 & x162 ) | ( x161 & x162 ) ;
  assign n2080 = ( x160 & ~n2077 ) | ( x160 & n2079 ) | ( ~n2077 & n2079 ) ;
  assign n2081 = ( ~x157 & x158 ) | ( ~x157 & x159 ) | ( x158 & x159 ) ;
  assign n2082 = ( x157 & ~n2078 ) | ( x157 & n2081 ) | ( ~n2078 & n2081 ) ;
  assign n2083 = n2080 & n2082 ;
  assign n2084 = ( n2077 & n2078 ) | ( n2077 & n2083 ) | ( n2078 & n2083 ) ;
  assign n2085 = ( x151 & x152 ) | ( x151 & x153 ) | ( x152 & x153 ) ;
  assign n2086 = ( x154 & x155 ) | ( x154 & x156 ) | ( x155 & x156 ) ;
  assign n2087 = ( ~x154 & x155 ) | ( ~x154 & x156 ) | ( x155 & x156 ) ;
  assign n2088 = ( x154 & ~n2086 ) | ( x154 & n2087 ) | ( ~n2086 & n2087 ) ;
  assign n2089 = ( ~x151 & x152 ) | ( ~x151 & x153 ) | ( x152 & x153 ) ;
  assign n2090 = ( x151 & ~n2085 ) | ( x151 & n2089 ) | ( ~n2085 & n2089 ) ;
  assign n2091 = n2088 & n2090 ;
  assign n2092 = ( n2085 & n2086 ) | ( n2085 & n2091 ) | ( n2086 & n2091 ) ;
  assign n2093 = ( ~n2077 & n2078 ) | ( ~n2077 & n2083 ) | ( n2078 & n2083 ) ;
  assign n2094 = ( n2077 & ~n2084 ) | ( n2077 & n2093 ) | ( ~n2084 & n2093 ) ;
  assign n2095 = ( ~n2085 & n2086 ) | ( ~n2085 & n2091 ) | ( n2086 & n2091 ) ;
  assign n2096 = ( n2085 & ~n2092 ) | ( n2085 & n2095 ) | ( ~n2092 & n2095 ) ;
  assign n2097 = n2088 | n2090 ;
  assign n2098 = ~n2091 & n2097 ;
  assign n2099 = ( n2080 & n2082 ) | ( n2080 & n2098 ) | ( n2082 & n2098 ) ;
  assign n2100 = ~n2083 & n2099 ;
  assign n2101 = ( n2094 & n2096 ) | ( n2094 & n2100 ) | ( n2096 & n2100 ) ;
  assign n2102 = ( n2084 & n2092 ) | ( n2084 & n2101 ) | ( n2092 & n2101 ) ;
  assign n2103 = ( ~n2084 & n2092 ) | ( ~n2084 & n2101 ) | ( n2092 & n2101 ) ;
  assign n2104 = ( n2084 & ~n2102 ) | ( n2084 & n2103 ) | ( ~n2102 & n2103 ) ;
  assign n2105 = ( ~n2057 & n2065 ) | ( ~n2057 & n2075 ) | ( n2065 & n2075 ) ;
  assign n2106 = ( n2057 & ~n2076 ) | ( n2057 & n2105 ) | ( ~n2076 & n2105 ) ;
  assign n2107 = ( ~n2067 & n2069 ) | ( ~n2067 & n2074 ) | ( n2069 & n2074 ) ;
  assign n2108 = ( n2067 & ~n2075 ) | ( n2067 & n2107 ) | ( ~n2075 & n2107 ) ;
  assign n2109 = ( ~n2094 & n2096 ) | ( ~n2094 & n2100 ) | ( n2096 & n2100 ) ;
  assign n2110 = ( n2094 & ~n2101 ) | ( n2094 & n2109 ) | ( ~n2101 & n2109 ) ;
  assign n2111 = ( ~n2080 & n2082 ) | ( ~n2080 & n2098 ) | ( n2082 & n2098 ) ;
  assign n2112 = ( n2080 & ~n2099 ) | ( n2080 & n2111 ) | ( ~n2099 & n2111 ) ;
  assign n2113 = ( n2071 & n2073 ) | ( n2071 & n2112 ) | ( n2073 & n2112 ) ;
  assign n2114 = ~n2074 & n2113 ;
  assign n2115 = ( n2108 & n2110 ) | ( n2108 & n2114 ) | ( n2110 & n2114 ) ;
  assign n2116 = ( n2104 & n2106 ) | ( n2104 & n2115 ) | ( n2106 & n2115 ) ;
  assign n2117 = ( n2076 & n2102 ) | ( n2076 & n2116 ) | ( n2102 & n2116 ) ;
  assign n2118 = ( x148 & x149 ) | ( x148 & x150 ) | ( x149 & x150 ) ;
  assign n2119 = ( x145 & x146 ) | ( x145 & x147 ) | ( x146 & x147 ) ;
  assign n2120 = ( ~x148 & x149 ) | ( ~x148 & x150 ) | ( x149 & x150 ) ;
  assign n2121 = ( x148 & ~n2118 ) | ( x148 & n2120 ) | ( ~n2118 & n2120 ) ;
  assign n2122 = ( ~x145 & x146 ) | ( ~x145 & x147 ) | ( x146 & x147 ) ;
  assign n2123 = ( x145 & ~n2119 ) | ( x145 & n2122 ) | ( ~n2119 & n2122 ) ;
  assign n2124 = n2121 & n2123 ;
  assign n2125 = ( n2118 & n2119 ) | ( n2118 & n2124 ) | ( n2119 & n2124 ) ;
  assign n2126 = ( x139 & x140 ) | ( x139 & x141 ) | ( x140 & x141 ) ;
  assign n2127 = ( x142 & x143 ) | ( x142 & x144 ) | ( x143 & x144 ) ;
  assign n2128 = ( ~x142 & x143 ) | ( ~x142 & x144 ) | ( x143 & x144 ) ;
  assign n2129 = ( x142 & ~n2127 ) | ( x142 & n2128 ) | ( ~n2127 & n2128 ) ;
  assign n2130 = ( ~x139 & x140 ) | ( ~x139 & x141 ) | ( x140 & x141 ) ;
  assign n2131 = ( x139 & ~n2126 ) | ( x139 & n2130 ) | ( ~n2126 & n2130 ) ;
  assign n2132 = n2129 & n2131 ;
  assign n2133 = ( n2126 & n2127 ) | ( n2126 & n2132 ) | ( n2127 & n2132 ) ;
  assign n2134 = ( ~n2118 & n2119 ) | ( ~n2118 & n2124 ) | ( n2119 & n2124 ) ;
  assign n2135 = ( n2118 & ~n2125 ) | ( n2118 & n2134 ) | ( ~n2125 & n2134 ) ;
  assign n2136 = ( ~n2126 & n2127 ) | ( ~n2126 & n2132 ) | ( n2127 & n2132 ) ;
  assign n2137 = ( n2126 & ~n2133 ) | ( n2126 & n2136 ) | ( ~n2133 & n2136 ) ;
  assign n2138 = n2121 | n2123 ;
  assign n2139 = ~n2124 & n2138 ;
  assign n2140 = n2129 | n2131 ;
  assign n2141 = ~n2132 & n2140 ;
  assign n2142 = n2139 & n2141 ;
  assign n2143 = ( n2135 & n2137 ) | ( n2135 & n2142 ) | ( n2137 & n2142 ) ;
  assign n2144 = ( n2125 & n2133 ) | ( n2125 & n2143 ) | ( n2133 & n2143 ) ;
  assign n2145 = ( x136 & x137 ) | ( x136 & x138 ) | ( x137 & x138 ) ;
  assign n2146 = ( x133 & x134 ) | ( x133 & x135 ) | ( x134 & x135 ) ;
  assign n2147 = ( ~x136 & x137 ) | ( ~x136 & x138 ) | ( x137 & x138 ) ;
  assign n2148 = ( x136 & ~n2145 ) | ( x136 & n2147 ) | ( ~n2145 & n2147 ) ;
  assign n2149 = ( ~x133 & x134 ) | ( ~x133 & x135 ) | ( x134 & x135 ) ;
  assign n2150 = ( x133 & ~n2146 ) | ( x133 & n2149 ) | ( ~n2146 & n2149 ) ;
  assign n2151 = n2148 & n2150 ;
  assign n2152 = ( n2145 & n2146 ) | ( n2145 & n2151 ) | ( n2146 & n2151 ) ;
  assign n2153 = ( x127 & x128 ) | ( x127 & x129 ) | ( x128 & x129 ) ;
  assign n2154 = ( x130 & x131 ) | ( x130 & x132 ) | ( x131 & x132 ) ;
  assign n2155 = ( ~x130 & x131 ) | ( ~x130 & x132 ) | ( x131 & x132 ) ;
  assign n2156 = ( x130 & ~n2154 ) | ( x130 & n2155 ) | ( ~n2154 & n2155 ) ;
  assign n2157 = ( ~x127 & x128 ) | ( ~x127 & x129 ) | ( x128 & x129 ) ;
  assign n2158 = ( x127 & ~n2153 ) | ( x127 & n2157 ) | ( ~n2153 & n2157 ) ;
  assign n2159 = n2156 & n2158 ;
  assign n2160 = ( n2153 & n2154 ) | ( n2153 & n2159 ) | ( n2154 & n2159 ) ;
  assign n2161 = ( ~n2145 & n2146 ) | ( ~n2145 & n2151 ) | ( n2146 & n2151 ) ;
  assign n2162 = ( n2145 & ~n2152 ) | ( n2145 & n2161 ) | ( ~n2152 & n2161 ) ;
  assign n2163 = ( ~n2153 & n2154 ) | ( ~n2153 & n2159 ) | ( n2154 & n2159 ) ;
  assign n2164 = ( n2153 & ~n2160 ) | ( n2153 & n2163 ) | ( ~n2160 & n2163 ) ;
  assign n2165 = n2156 | n2158 ;
  assign n2166 = ~n2159 & n2165 ;
  assign n2167 = ( n2148 & n2150 ) | ( n2148 & n2166 ) | ( n2150 & n2166 ) ;
  assign n2168 = ~n2151 & n2167 ;
  assign n2169 = ( n2162 & n2164 ) | ( n2162 & n2168 ) | ( n2164 & n2168 ) ;
  assign n2170 = ( n2152 & n2160 ) | ( n2152 & n2169 ) | ( n2160 & n2169 ) ;
  assign n2171 = ( ~n2152 & n2160 ) | ( ~n2152 & n2169 ) | ( n2160 & n2169 ) ;
  assign n2172 = ( n2152 & ~n2170 ) | ( n2152 & n2171 ) | ( ~n2170 & n2171 ) ;
  assign n2173 = ( ~n2125 & n2133 ) | ( ~n2125 & n2143 ) | ( n2133 & n2143 ) ;
  assign n2174 = ( n2125 & ~n2144 ) | ( n2125 & n2173 ) | ( ~n2144 & n2173 ) ;
  assign n2175 = ( ~n2135 & n2137 ) | ( ~n2135 & n2142 ) | ( n2137 & n2142 ) ;
  assign n2176 = ( n2135 & ~n2143 ) | ( n2135 & n2175 ) | ( ~n2143 & n2175 ) ;
  assign n2177 = ( ~n2162 & n2164 ) | ( ~n2162 & n2168 ) | ( n2164 & n2168 ) ;
  assign n2178 = ( n2162 & ~n2169 ) | ( n2162 & n2177 ) | ( ~n2169 & n2177 ) ;
  assign n2179 = ( ~n2148 & n2150 ) | ( ~n2148 & n2166 ) | ( n2150 & n2166 ) ;
  assign n2180 = ( n2148 & ~n2167 ) | ( n2148 & n2179 ) | ( ~n2167 & n2179 ) ;
  assign n2181 = ( n2139 & n2141 ) | ( n2139 & n2180 ) | ( n2141 & n2180 ) ;
  assign n2182 = ~n2142 & n2181 ;
  assign n2183 = ( n2176 & n2178 ) | ( n2176 & n2182 ) | ( n2178 & n2182 ) ;
  assign n2184 = ( n2172 & n2174 ) | ( n2172 & n2183 ) | ( n2174 & n2183 ) ;
  assign n2185 = ( n2144 & n2170 ) | ( n2144 & n2184 ) | ( n2170 & n2184 ) ;
  assign n2186 = ( ~n2076 & n2102 ) | ( ~n2076 & n2116 ) | ( n2102 & n2116 ) ;
  assign n2187 = ( n2076 & ~n2117 ) | ( n2076 & n2186 ) | ( ~n2117 & n2186 ) ;
  assign n2188 = ( ~n2144 & n2170 ) | ( ~n2144 & n2184 ) | ( n2170 & n2184 ) ;
  assign n2189 = ( n2144 & ~n2185 ) | ( n2144 & n2188 ) | ( ~n2185 & n2188 ) ;
  assign n2190 = ( ~n2172 & n2174 ) | ( ~n2172 & n2183 ) | ( n2174 & n2183 ) ;
  assign n2191 = ( n2172 & ~n2184 ) | ( n2172 & n2190 ) | ( ~n2184 & n2190 ) ;
  assign n2192 = ( ~n2104 & n2106 ) | ( ~n2104 & n2115 ) | ( n2106 & n2115 ) ;
  assign n2193 = ( n2104 & ~n2116 ) | ( n2104 & n2192 ) | ( ~n2116 & n2192 ) ;
  assign n2194 = ( n2108 & n2110 ) | ( n2108 & ~n2114 ) | ( n2110 & ~n2114 ) ;
  assign n2195 = ( n2114 & ~n2115 ) | ( n2114 & n2194 ) | ( ~n2115 & n2194 ) ;
  assign n2196 = ( n2176 & n2178 ) | ( n2176 & ~n2182 ) | ( n2178 & ~n2182 ) ;
  assign n2197 = ( n2182 & ~n2183 ) | ( n2182 & n2196 ) | ( ~n2183 & n2196 ) ;
  assign n2198 = ( ~n2071 & n2073 ) | ( ~n2071 & n2112 ) | ( n2073 & n2112 ) ;
  assign n2199 = ( n2071 & ~n2113 ) | ( n2071 & n2198 ) | ( ~n2113 & n2198 ) ;
  assign n2200 = ( ~n2139 & n2141 ) | ( ~n2139 & n2180 ) | ( n2141 & n2180 ) ;
  assign n2201 = ( n2139 & ~n2181 ) | ( n2139 & n2200 ) | ( ~n2181 & n2200 ) ;
  assign n2202 = n2199 & n2201 ;
  assign n2203 = ( n2195 & n2197 ) | ( n2195 & n2202 ) | ( n2197 & n2202 ) ;
  assign n2204 = ( n2191 & n2193 ) | ( n2191 & n2203 ) | ( n2193 & n2203 ) ;
  assign n2205 = ( n2187 & n2189 ) | ( n2187 & n2204 ) | ( n2189 & n2204 ) ;
  assign n2206 = ( n2117 & n2185 ) | ( n2117 & n2205 ) | ( n2185 & n2205 ) ;
  assign n2207 = ( x124 & x125 ) | ( x124 & x126 ) | ( x125 & x126 ) ;
  assign n2208 = ( x121 & x122 ) | ( x121 & x123 ) | ( x122 & x123 ) ;
  assign n2209 = ( ~x124 & x125 ) | ( ~x124 & x126 ) | ( x125 & x126 ) ;
  assign n2210 = ( x124 & ~n2207 ) | ( x124 & n2209 ) | ( ~n2207 & n2209 ) ;
  assign n2211 = ( ~x121 & x122 ) | ( ~x121 & x123 ) | ( x122 & x123 ) ;
  assign n2212 = ( x121 & ~n2208 ) | ( x121 & n2211 ) | ( ~n2208 & n2211 ) ;
  assign n2213 = n2210 & n2212 ;
  assign n2214 = ( n2207 & n2208 ) | ( n2207 & n2213 ) | ( n2208 & n2213 ) ;
  assign n2215 = ( x115 & x116 ) | ( x115 & x117 ) | ( x116 & x117 ) ;
  assign n2216 = ( x118 & x119 ) | ( x118 & x120 ) | ( x119 & x120 ) ;
  assign n2217 = ( ~x118 & x119 ) | ( ~x118 & x120 ) | ( x119 & x120 ) ;
  assign n2218 = ( x118 & ~n2216 ) | ( x118 & n2217 ) | ( ~n2216 & n2217 ) ;
  assign n2219 = ( ~x115 & x116 ) | ( ~x115 & x117 ) | ( x116 & x117 ) ;
  assign n2220 = ( x115 & ~n2215 ) | ( x115 & n2219 ) | ( ~n2215 & n2219 ) ;
  assign n2221 = n2218 & n2220 ;
  assign n2222 = ( n2215 & n2216 ) | ( n2215 & n2221 ) | ( n2216 & n2221 ) ;
  assign n2223 = ( ~n2207 & n2208 ) | ( ~n2207 & n2213 ) | ( n2208 & n2213 ) ;
  assign n2224 = ( n2207 & ~n2214 ) | ( n2207 & n2223 ) | ( ~n2214 & n2223 ) ;
  assign n2225 = ( ~n2215 & n2216 ) | ( ~n2215 & n2221 ) | ( n2216 & n2221 ) ;
  assign n2226 = ( n2215 & ~n2222 ) | ( n2215 & n2225 ) | ( ~n2222 & n2225 ) ;
  assign n2227 = n2210 | n2212 ;
  assign n2228 = ~n2213 & n2227 ;
  assign n2229 = n2218 | n2220 ;
  assign n2230 = ~n2221 & n2229 ;
  assign n2231 = n2228 & n2230 ;
  assign n2232 = ( n2224 & n2226 ) | ( n2224 & n2231 ) | ( n2226 & n2231 ) ;
  assign n2233 = ( n2214 & n2222 ) | ( n2214 & n2232 ) | ( n2222 & n2232 ) ;
  assign n2234 = ( x112 & x113 ) | ( x112 & x114 ) | ( x113 & x114 ) ;
  assign n2235 = ( x109 & x110 ) | ( x109 & x111 ) | ( x110 & x111 ) ;
  assign n2236 = ( ~x112 & x113 ) | ( ~x112 & x114 ) | ( x113 & x114 ) ;
  assign n2237 = ( x112 & ~n2234 ) | ( x112 & n2236 ) | ( ~n2234 & n2236 ) ;
  assign n2238 = ( ~x109 & x110 ) | ( ~x109 & x111 ) | ( x110 & x111 ) ;
  assign n2239 = ( x109 & ~n2235 ) | ( x109 & n2238 ) | ( ~n2235 & n2238 ) ;
  assign n2240 = n2237 & n2239 ;
  assign n2241 = ( n2234 & n2235 ) | ( n2234 & n2240 ) | ( n2235 & n2240 ) ;
  assign n2242 = ( x103 & x104 ) | ( x103 & x105 ) | ( x104 & x105 ) ;
  assign n2243 = ( x106 & x107 ) | ( x106 & x108 ) | ( x107 & x108 ) ;
  assign n2244 = ( ~x106 & x107 ) | ( ~x106 & x108 ) | ( x107 & x108 ) ;
  assign n2245 = ( x106 & ~n2243 ) | ( x106 & n2244 ) | ( ~n2243 & n2244 ) ;
  assign n2246 = ( ~x103 & x104 ) | ( ~x103 & x105 ) | ( x104 & x105 ) ;
  assign n2247 = ( x103 & ~n2242 ) | ( x103 & n2246 ) | ( ~n2242 & n2246 ) ;
  assign n2248 = n2245 & n2247 ;
  assign n2249 = ( n2242 & n2243 ) | ( n2242 & n2248 ) | ( n2243 & n2248 ) ;
  assign n2250 = ( ~n2234 & n2235 ) | ( ~n2234 & n2240 ) | ( n2235 & n2240 ) ;
  assign n2251 = ( n2234 & ~n2241 ) | ( n2234 & n2250 ) | ( ~n2241 & n2250 ) ;
  assign n2252 = ( ~n2242 & n2243 ) | ( ~n2242 & n2248 ) | ( n2243 & n2248 ) ;
  assign n2253 = ( n2242 & ~n2249 ) | ( n2242 & n2252 ) | ( ~n2249 & n2252 ) ;
  assign n2254 = n2245 | n2247 ;
  assign n2255 = ~n2248 & n2254 ;
  assign n2256 = ( n2237 & n2239 ) | ( n2237 & n2255 ) | ( n2239 & n2255 ) ;
  assign n2257 = ~n2240 & n2256 ;
  assign n2258 = ( n2251 & n2253 ) | ( n2251 & n2257 ) | ( n2253 & n2257 ) ;
  assign n2259 = ( n2241 & n2249 ) | ( n2241 & n2258 ) | ( n2249 & n2258 ) ;
  assign n2260 = ( ~n2241 & n2249 ) | ( ~n2241 & n2258 ) | ( n2249 & n2258 ) ;
  assign n2261 = ( n2241 & ~n2259 ) | ( n2241 & n2260 ) | ( ~n2259 & n2260 ) ;
  assign n2262 = ( ~n2214 & n2222 ) | ( ~n2214 & n2232 ) | ( n2222 & n2232 ) ;
  assign n2263 = ( n2214 & ~n2233 ) | ( n2214 & n2262 ) | ( ~n2233 & n2262 ) ;
  assign n2264 = ( ~n2224 & n2226 ) | ( ~n2224 & n2231 ) | ( n2226 & n2231 ) ;
  assign n2265 = ( n2224 & ~n2232 ) | ( n2224 & n2264 ) | ( ~n2232 & n2264 ) ;
  assign n2266 = ( ~n2251 & n2253 ) | ( ~n2251 & n2257 ) | ( n2253 & n2257 ) ;
  assign n2267 = ( n2251 & ~n2258 ) | ( n2251 & n2266 ) | ( ~n2258 & n2266 ) ;
  assign n2268 = ( ~n2237 & n2239 ) | ( ~n2237 & n2255 ) | ( n2239 & n2255 ) ;
  assign n2269 = ( n2237 & ~n2256 ) | ( n2237 & n2268 ) | ( ~n2256 & n2268 ) ;
  assign n2270 = ( n2228 & n2230 ) | ( n2228 & n2269 ) | ( n2230 & n2269 ) ;
  assign n2271 = ~n2231 & n2270 ;
  assign n2272 = ( n2265 & n2267 ) | ( n2265 & n2271 ) | ( n2267 & n2271 ) ;
  assign n2273 = ( n2261 & n2263 ) | ( n2261 & n2272 ) | ( n2263 & n2272 ) ;
  assign n2274 = ( n2233 & n2259 ) | ( n2233 & n2273 ) | ( n2259 & n2273 ) ;
  assign n2275 = ( x100 & x101 ) | ( x100 & x102 ) | ( x101 & x102 ) ;
  assign n2276 = ( x97 & x98 ) | ( x97 & x99 ) | ( x98 & x99 ) ;
  assign n2277 = ( ~x100 & x101 ) | ( ~x100 & x102 ) | ( x101 & x102 ) ;
  assign n2278 = ( x100 & ~n2275 ) | ( x100 & n2277 ) | ( ~n2275 & n2277 ) ;
  assign n2279 = ( ~x97 & x98 ) | ( ~x97 & x99 ) | ( x98 & x99 ) ;
  assign n2280 = ( x97 & ~n2276 ) | ( x97 & n2279 ) | ( ~n2276 & n2279 ) ;
  assign n2281 = n2278 & n2280 ;
  assign n2282 = ( n2275 & n2276 ) | ( n2275 & n2281 ) | ( n2276 & n2281 ) ;
  assign n2283 = ( x91 & x92 ) | ( x91 & x93 ) | ( x92 & x93 ) ;
  assign n2284 = ( x94 & x95 ) | ( x94 & x96 ) | ( x95 & x96 ) ;
  assign n2285 = ( ~x94 & x95 ) | ( ~x94 & x96 ) | ( x95 & x96 ) ;
  assign n2286 = ( x94 & ~n2284 ) | ( x94 & n2285 ) | ( ~n2284 & n2285 ) ;
  assign n2287 = ( ~x91 & x92 ) | ( ~x91 & x93 ) | ( x92 & x93 ) ;
  assign n2288 = ( x91 & ~n2283 ) | ( x91 & n2287 ) | ( ~n2283 & n2287 ) ;
  assign n2289 = n2286 & n2288 ;
  assign n2290 = ( n2283 & n2284 ) | ( n2283 & n2289 ) | ( n2284 & n2289 ) ;
  assign n2291 = ( ~n2275 & n2276 ) | ( ~n2275 & n2281 ) | ( n2276 & n2281 ) ;
  assign n2292 = ( n2275 & ~n2282 ) | ( n2275 & n2291 ) | ( ~n2282 & n2291 ) ;
  assign n2293 = ( ~n2283 & n2284 ) | ( ~n2283 & n2289 ) | ( n2284 & n2289 ) ;
  assign n2294 = ( n2283 & ~n2290 ) | ( n2283 & n2293 ) | ( ~n2290 & n2293 ) ;
  assign n2295 = n2278 | n2280 ;
  assign n2296 = ~n2281 & n2295 ;
  assign n2297 = n2286 | n2288 ;
  assign n2298 = ~n2289 & n2297 ;
  assign n2299 = n2296 & n2298 ;
  assign n2300 = ( n2292 & n2294 ) | ( n2292 & n2299 ) | ( n2294 & n2299 ) ;
  assign n2301 = ( n2282 & n2290 ) | ( n2282 & n2300 ) | ( n2290 & n2300 ) ;
  assign n2302 = ( x88 & x89 ) | ( x88 & x90 ) | ( x89 & x90 ) ;
  assign n2303 = ( x85 & x86 ) | ( x85 & x87 ) | ( x86 & x87 ) ;
  assign n2304 = ( ~x88 & x89 ) | ( ~x88 & x90 ) | ( x89 & x90 ) ;
  assign n2305 = ( x88 & ~n2302 ) | ( x88 & n2304 ) | ( ~n2302 & n2304 ) ;
  assign n2306 = ( ~x85 & x86 ) | ( ~x85 & x87 ) | ( x86 & x87 ) ;
  assign n2307 = ( x85 & ~n2303 ) | ( x85 & n2306 ) | ( ~n2303 & n2306 ) ;
  assign n2308 = n2305 & n2307 ;
  assign n2309 = ( n2302 & n2303 ) | ( n2302 & n2308 ) | ( n2303 & n2308 ) ;
  assign n2310 = ( x79 & x80 ) | ( x79 & x81 ) | ( x80 & x81 ) ;
  assign n2311 = ( x82 & x83 ) | ( x82 & x84 ) | ( x83 & x84 ) ;
  assign n2312 = ( ~x82 & x83 ) | ( ~x82 & x84 ) | ( x83 & x84 ) ;
  assign n2313 = ( x82 & ~n2311 ) | ( x82 & n2312 ) | ( ~n2311 & n2312 ) ;
  assign n2314 = ( ~x79 & x80 ) | ( ~x79 & x81 ) | ( x80 & x81 ) ;
  assign n2315 = ( x79 & ~n2310 ) | ( x79 & n2314 ) | ( ~n2310 & n2314 ) ;
  assign n2316 = n2313 & n2315 ;
  assign n2317 = ( n2310 & n2311 ) | ( n2310 & n2316 ) | ( n2311 & n2316 ) ;
  assign n2318 = ( ~n2302 & n2303 ) | ( ~n2302 & n2308 ) | ( n2303 & n2308 ) ;
  assign n2319 = ( n2302 & ~n2309 ) | ( n2302 & n2318 ) | ( ~n2309 & n2318 ) ;
  assign n2320 = ( ~n2310 & n2311 ) | ( ~n2310 & n2316 ) | ( n2311 & n2316 ) ;
  assign n2321 = ( n2310 & ~n2317 ) | ( n2310 & n2320 ) | ( ~n2317 & n2320 ) ;
  assign n2322 = n2313 | n2315 ;
  assign n2323 = ~n2316 & n2322 ;
  assign n2324 = ( n2305 & n2307 ) | ( n2305 & n2323 ) | ( n2307 & n2323 ) ;
  assign n2325 = ~n2308 & n2324 ;
  assign n2326 = ( n2319 & n2321 ) | ( n2319 & n2325 ) | ( n2321 & n2325 ) ;
  assign n2327 = ( n2309 & n2317 ) | ( n2309 & n2326 ) | ( n2317 & n2326 ) ;
  assign n2328 = ( ~n2309 & n2317 ) | ( ~n2309 & n2326 ) | ( n2317 & n2326 ) ;
  assign n2329 = ( n2309 & ~n2327 ) | ( n2309 & n2328 ) | ( ~n2327 & n2328 ) ;
  assign n2330 = ( ~n2282 & n2290 ) | ( ~n2282 & n2300 ) | ( n2290 & n2300 ) ;
  assign n2331 = ( n2282 & ~n2301 ) | ( n2282 & n2330 ) | ( ~n2301 & n2330 ) ;
  assign n2332 = ( ~n2292 & n2294 ) | ( ~n2292 & n2299 ) | ( n2294 & n2299 ) ;
  assign n2333 = ( n2292 & ~n2300 ) | ( n2292 & n2332 ) | ( ~n2300 & n2332 ) ;
  assign n2334 = ( ~n2319 & n2321 ) | ( ~n2319 & n2325 ) | ( n2321 & n2325 ) ;
  assign n2335 = ( n2319 & ~n2326 ) | ( n2319 & n2334 ) | ( ~n2326 & n2334 ) ;
  assign n2336 = ( ~n2305 & n2307 ) | ( ~n2305 & n2323 ) | ( n2307 & n2323 ) ;
  assign n2337 = ( n2305 & ~n2324 ) | ( n2305 & n2336 ) | ( ~n2324 & n2336 ) ;
  assign n2338 = ( n2296 & n2298 ) | ( n2296 & n2337 ) | ( n2298 & n2337 ) ;
  assign n2339 = ~n2299 & n2338 ;
  assign n2340 = ( n2333 & n2335 ) | ( n2333 & n2339 ) | ( n2335 & n2339 ) ;
  assign n2341 = ( n2329 & n2331 ) | ( n2329 & n2340 ) | ( n2331 & n2340 ) ;
  assign n2342 = ( n2301 & n2327 ) | ( n2301 & n2341 ) | ( n2327 & n2341 ) ;
  assign n2343 = ( ~n2233 & n2259 ) | ( ~n2233 & n2273 ) | ( n2259 & n2273 ) ;
  assign n2344 = ( n2233 & ~n2274 ) | ( n2233 & n2343 ) | ( ~n2274 & n2343 ) ;
  assign n2345 = ( ~n2301 & n2327 ) | ( ~n2301 & n2341 ) | ( n2327 & n2341 ) ;
  assign n2346 = ( n2301 & ~n2342 ) | ( n2301 & n2345 ) | ( ~n2342 & n2345 ) ;
  assign n2347 = ( ~n2329 & n2331 ) | ( ~n2329 & n2340 ) | ( n2331 & n2340 ) ;
  assign n2348 = ( n2329 & ~n2341 ) | ( n2329 & n2347 ) | ( ~n2341 & n2347 ) ;
  assign n2349 = ( ~n2261 & n2263 ) | ( ~n2261 & n2272 ) | ( n2263 & n2272 ) ;
  assign n2350 = ( n2261 & ~n2273 ) | ( n2261 & n2349 ) | ( ~n2273 & n2349 ) ;
  assign n2351 = ( n2265 & n2267 ) | ( n2265 & ~n2271 ) | ( n2267 & ~n2271 ) ;
  assign n2352 = ( n2271 & ~n2272 ) | ( n2271 & n2351 ) | ( ~n2272 & n2351 ) ;
  assign n2353 = ( n2333 & n2335 ) | ( n2333 & ~n2339 ) | ( n2335 & ~n2339 ) ;
  assign n2354 = ( n2339 & ~n2340 ) | ( n2339 & n2353 ) | ( ~n2340 & n2353 ) ;
  assign n2355 = ( ~n2228 & n2230 ) | ( ~n2228 & n2269 ) | ( n2230 & n2269 ) ;
  assign n2356 = ( n2228 & ~n2270 ) | ( n2228 & n2355 ) | ( ~n2270 & n2355 ) ;
  assign n2357 = ( ~n2296 & n2298 ) | ( ~n2296 & n2337 ) | ( n2298 & n2337 ) ;
  assign n2358 = ( n2296 & ~n2338 ) | ( n2296 & n2357 ) | ( ~n2338 & n2357 ) ;
  assign n2359 = n2356 & n2358 ;
  assign n2360 = ( n2352 & n2354 ) | ( n2352 & n2359 ) | ( n2354 & n2359 ) ;
  assign n2361 = ( n2348 & n2350 ) | ( n2348 & n2360 ) | ( n2350 & n2360 ) ;
  assign n2362 = ( n2344 & n2346 ) | ( n2344 & n2361 ) | ( n2346 & n2361 ) ;
  assign n2363 = ( n2274 & n2342 ) | ( n2274 & n2362 ) | ( n2342 & n2362 ) ;
  assign n2364 = ( ~n2274 & n2342 ) | ( ~n2274 & n2362 ) | ( n2342 & n2362 ) ;
  assign n2365 = ( n2274 & ~n2363 ) | ( n2274 & n2364 ) | ( ~n2363 & n2364 ) ;
  assign n2366 = ( ~n2117 & n2185 ) | ( ~n2117 & n2205 ) | ( n2185 & n2205 ) ;
  assign n2367 = ( n2117 & ~n2206 ) | ( n2117 & n2366 ) | ( ~n2206 & n2366 ) ;
  assign n2368 = ( ~n2187 & n2189 ) | ( ~n2187 & n2204 ) | ( n2189 & n2204 ) ;
  assign n2369 = ( n2187 & ~n2205 ) | ( n2187 & n2368 ) | ( ~n2205 & n2368 ) ;
  assign n2370 = ( ~n2344 & n2346 ) | ( ~n2344 & n2361 ) | ( n2346 & n2361 ) ;
  assign n2371 = ( n2344 & ~n2362 ) | ( n2344 & n2370 ) | ( ~n2362 & n2370 ) ;
  assign n2372 = ( ~n2348 & n2350 ) | ( ~n2348 & n2360 ) | ( n2350 & n2360 ) ;
  assign n2373 = ( n2348 & ~n2361 ) | ( n2348 & n2372 ) | ( ~n2361 & n2372 ) ;
  assign n2374 = ( ~n2191 & n2193 ) | ( ~n2191 & n2203 ) | ( n2193 & n2203 ) ;
  assign n2375 = ( n2191 & ~n2204 ) | ( n2191 & n2374 ) | ( ~n2204 & n2374 ) ;
  assign n2376 = ( ~n2195 & n2197 ) | ( ~n2195 & n2202 ) | ( n2197 & n2202 ) ;
  assign n2377 = ( n2195 & ~n2203 ) | ( n2195 & n2376 ) | ( ~n2203 & n2376 ) ;
  assign n2378 = ( ~n2352 & n2354 ) | ( ~n2352 & n2359 ) | ( n2354 & n2359 ) ;
  assign n2379 = ( n2352 & ~n2360 ) | ( n2352 & n2378 ) | ( ~n2360 & n2378 ) ;
  assign n2380 = n2356 | n2358 ;
  assign n2381 = ~n2359 & n2380 ;
  assign n2382 = ( n2199 & n2201 ) | ( n2199 & n2381 ) | ( n2201 & n2381 ) ;
  assign n2383 = ~n2202 & n2382 ;
  assign n2384 = ( n2377 & n2379 ) | ( n2377 & n2383 ) | ( n2379 & n2383 ) ;
  assign n2385 = ( n2373 & n2375 ) | ( n2373 & n2384 ) | ( n2375 & n2384 ) ;
  assign n2386 = ( n2369 & n2371 ) | ( n2369 & n2385 ) | ( n2371 & n2385 ) ;
  assign n2387 = ( n2365 & n2367 ) | ( n2365 & n2386 ) | ( n2367 & n2386 ) ;
  assign n2388 = ( n2206 & n2363 ) | ( n2206 & n2387 ) | ( n2363 & n2387 ) ;
  assign n2389 = ( ~n1867 & n2024 ) | ( ~n1867 & n2048 ) | ( n2024 & n2048 ) ;
  assign n2390 = ( n1867 & ~n2049 ) | ( n1867 & n2389 ) | ( ~n2049 & n2389 ) ;
  assign n2391 = ( ~n2206 & n2363 ) | ( ~n2206 & n2387 ) | ( n2363 & n2387 ) ;
  assign n2392 = ( n2206 & ~n2388 ) | ( n2206 & n2391 ) | ( ~n2388 & n2391 ) ;
  assign n2393 = ( ~n2365 & n2367 ) | ( ~n2365 & n2386 ) | ( n2367 & n2386 ) ;
  assign n2394 = ( n2365 & ~n2387 ) | ( n2365 & n2393 ) | ( ~n2387 & n2393 ) ;
  assign n2395 = ( ~n2026 & n2028 ) | ( ~n2026 & n2047 ) | ( n2028 & n2047 ) ;
  assign n2396 = ( n2026 & ~n2048 ) | ( n2026 & n2395 ) | ( ~n2048 & n2395 ) ;
  assign n2397 = ( ~n2030 & n2032 ) | ( ~n2030 & n2046 ) | ( n2032 & n2046 ) ;
  assign n2398 = ( n2030 & ~n2047 ) | ( n2030 & n2397 ) | ( ~n2047 & n2397 ) ;
  assign n2399 = ( ~n2369 & n2371 ) | ( ~n2369 & n2385 ) | ( n2371 & n2385 ) ;
  assign n2400 = ( n2369 & ~n2386 ) | ( n2369 & n2399 ) | ( ~n2386 & n2399 ) ;
  assign n2401 = ( ~n2373 & n2375 ) | ( ~n2373 & n2384 ) | ( n2375 & n2384 ) ;
  assign n2402 = ( n2373 & ~n2385 ) | ( n2373 & n2401 ) | ( ~n2385 & n2401 ) ;
  assign n2403 = ( ~n2034 & n2036 ) | ( ~n2034 & n2045 ) | ( n2036 & n2045 ) ;
  assign n2404 = ( n2034 & ~n2046 ) | ( n2034 & n2403 ) | ( ~n2046 & n2403 ) ;
  assign n2405 = ( ~n1860 & n1862 ) | ( ~n1860 & n2042 ) | ( n1862 & n2042 ) ;
  assign n2406 = ( n1860 & ~n2043 ) | ( n1860 & n2405 ) | ( ~n2043 & n2405 ) ;
  assign n2407 = ( ~n2199 & n2201 ) | ( ~n2199 & n2381 ) | ( n2201 & n2381 ) ;
  assign n2408 = ( n2199 & ~n2382 ) | ( n2199 & n2407 ) | ( ~n2382 & n2407 ) ;
  assign n2409 = n2406 & n2408 ;
  assign n2410 = ( n2038 & n2040 ) | ( n2038 & ~n2044 ) | ( n2040 & ~n2044 ) ;
  assign n2411 = ( n2044 & ~n2045 ) | ( n2044 & n2410 ) | ( ~n2045 & n2410 ) ;
  assign n2412 = ( n2377 & n2379 ) | ( n2377 & ~n2383 ) | ( n2379 & ~n2383 ) ;
  assign n2413 = ( n2383 & ~n2384 ) | ( n2383 & n2412 ) | ( ~n2384 & n2412 ) ;
  assign n2414 = ( n2409 & n2411 ) | ( n2409 & n2413 ) | ( n2411 & n2413 ) ;
  assign n2415 = ( n2402 & n2404 ) | ( n2402 & n2414 ) | ( n2404 & n2414 ) ;
  assign n2416 = ( n2398 & n2400 ) | ( n2398 & n2415 ) | ( n2400 & n2415 ) ;
  assign n2417 = ( n2394 & n2396 ) | ( n2394 & n2416 ) | ( n2396 & n2416 ) ;
  assign n2418 = ( n2390 & n2392 ) | ( n2390 & n2417 ) | ( n2392 & n2417 ) ;
  assign n2419 = ( n2049 & n2388 ) | ( n2049 & n2418 ) | ( n2388 & n2418 ) ;
  assign n2420 = ( ~n2049 & n2388 ) | ( ~n2049 & n2418 ) | ( n2388 & n2418 ) ;
  assign n2421 = ( n2049 & ~n2419 ) | ( n2049 & n2420 ) | ( ~n2419 & n2420 ) ;
  assign n2422 = ( ~n1340 & n1679 ) | ( ~n1340 & n1709 ) | ( n1679 & n1709 ) ;
  assign n2423 = ( n1340 & ~n1710 ) | ( n1340 & n2422 ) | ( ~n1710 & n2422 ) ;
  assign n2424 = ( ~n1681 & n1683 ) | ( ~n1681 & n1708 ) | ( n1683 & n1708 ) ;
  assign n2425 = ( n1681 & ~n1709 ) | ( n1681 & n2424 ) | ( ~n1709 & n2424 ) ;
  assign n2426 = ( ~n2390 & n2392 ) | ( ~n2390 & n2417 ) | ( n2392 & n2417 ) ;
  assign n2427 = ( n2390 & ~n2418 ) | ( n2390 & n2426 ) | ( ~n2418 & n2426 ) ;
  assign n2428 = ( ~n2394 & n2396 ) | ( ~n2394 & n2416 ) | ( n2396 & n2416 ) ;
  assign n2429 = ( n2394 & ~n2417 ) | ( n2394 & n2428 ) | ( ~n2417 & n2428 ) ;
  assign n2430 = ( ~n1685 & n1687 ) | ( ~n1685 & n1707 ) | ( n1687 & n1707 ) ;
  assign n2431 = ( n1685 & ~n1708 ) | ( n1685 & n2430 ) | ( ~n1708 & n2430 ) ;
  assign n2432 = ( ~n1689 & n1691 ) | ( ~n1689 & n1706 ) | ( n1691 & n1706 ) ;
  assign n2433 = ( n1689 & ~n1707 ) | ( n1689 & n2432 ) | ( ~n1707 & n2432 ) ;
  assign n2434 = ( ~n2398 & n2400 ) | ( ~n2398 & n2415 ) | ( n2400 & n2415 ) ;
  assign n2435 = ( n2398 & ~n2416 ) | ( n2398 & n2434 ) | ( ~n2416 & n2434 ) ;
  assign n2436 = ( ~n2402 & n2404 ) | ( ~n2402 & n2414 ) | ( n2404 & n2414 ) ;
  assign n2437 = ( n2402 & ~n2415 ) | ( n2402 & n2436 ) | ( ~n2415 & n2436 ) ;
  assign n2438 = ( ~n1693 & n1695 ) | ( ~n1693 & n1705 ) | ( n1695 & n1705 ) ;
  assign n2439 = ( n1693 & ~n1706 ) | ( n1693 & n2438 ) | ( ~n1706 & n2438 ) ;
  assign n2440 = ( ~n1700 & n1702 ) | ( ~n1700 & n1704 ) | ( n1702 & n1704 ) ;
  assign n2441 = ( n1700 & ~n1705 ) | ( n1700 & n2440 ) | ( ~n1705 & n2440 ) ;
  assign n2442 = ( ~n2409 & n2411 ) | ( ~n2409 & n2413 ) | ( n2411 & n2413 ) ;
  assign n2443 = ( n2409 & ~n2414 ) | ( n2409 & n2442 ) | ( ~n2414 & n2442 ) ;
  assign n2444 = n1697 | n1699 ;
  assign n2445 = ~n1700 & n2444 ;
  assign n2446 = n2406 | n2408 ;
  assign n2447 = ~n2409 & n2446 ;
  assign n2448 = n2445 & n2447 ;
  assign n2449 = ( n2441 & n2443 ) | ( n2441 & n2448 ) | ( n2443 & n2448 ) ;
  assign n2450 = ( n2437 & n2439 ) | ( n2437 & n2449 ) | ( n2439 & n2449 ) ;
  assign n2451 = ( n2433 & n2435 ) | ( n2433 & n2450 ) | ( n2435 & n2450 ) ;
  assign n2452 = ( n2429 & n2431 ) | ( n2429 & n2451 ) | ( n2431 & n2451 ) ;
  assign n2453 = ( n2425 & n2427 ) | ( n2425 & n2452 ) | ( n2427 & n2452 ) ;
  assign n2454 = ( n2421 & n2423 ) | ( n2421 & n2453 ) | ( n2423 & n2453 ) ;
  assign n2455 = ( n1710 & n2419 ) | ( n1710 & n2454 ) | ( n2419 & n2454 ) ;
  assign n2456 = ( ~n1710 & n2419 ) | ( ~n1710 & n2454 ) | ( n2419 & n2454 ) ;
  assign n2457 = ( n1710 & ~n2455 ) | ( n1710 & n2456 ) | ( ~n2455 & n2456 ) ;
  assign n2458 = ( x28 & x29 ) | ( x28 & x30 ) | ( x29 & x30 ) ;
  assign n2459 = ( x25 & x26 ) | ( x25 & x27 ) | ( x26 & x27 ) ;
  assign n2460 = ( ~x28 & x29 ) | ( ~x28 & x30 ) | ( x29 & x30 ) ;
  assign n2461 = ( x28 & ~n2458 ) | ( x28 & n2460 ) | ( ~n2458 & n2460 ) ;
  assign n2462 = ( ~x25 & x26 ) | ( ~x25 & x27 ) | ( x26 & x27 ) ;
  assign n2463 = ( x25 & ~n2459 ) | ( x25 & n2462 ) | ( ~n2459 & n2462 ) ;
  assign n2464 = n2461 & n2463 ;
  assign n2465 = ( n2458 & n2459 ) | ( n2458 & n2464 ) | ( n2459 & n2464 ) ;
  assign n2466 = ( x19 & x20 ) | ( x19 & x21 ) | ( x20 & x21 ) ;
  assign n2467 = ( x22 & x23 ) | ( x22 & x24 ) | ( x23 & x24 ) ;
  assign n2468 = ( ~x22 & x23 ) | ( ~x22 & x24 ) | ( x23 & x24 ) ;
  assign n2469 = ( x22 & ~n2467 ) | ( x22 & n2468 ) | ( ~n2467 & n2468 ) ;
  assign n2470 = ( ~x19 & x20 ) | ( ~x19 & x21 ) | ( x20 & x21 ) ;
  assign n2471 = ( x19 & ~n2466 ) | ( x19 & n2470 ) | ( ~n2466 & n2470 ) ;
  assign n2472 = n2469 & n2471 ;
  assign n2473 = ( n2466 & n2467 ) | ( n2466 & n2472 ) | ( n2467 & n2472 ) ;
  assign n2474 = ( ~n2458 & n2459 ) | ( ~n2458 & n2464 ) | ( n2459 & n2464 ) ;
  assign n2475 = ( n2458 & ~n2465 ) | ( n2458 & n2474 ) | ( ~n2465 & n2474 ) ;
  assign n2476 = ( ~n2466 & n2467 ) | ( ~n2466 & n2472 ) | ( n2467 & n2472 ) ;
  assign n2477 = ( n2466 & ~n2473 ) | ( n2466 & n2476 ) | ( ~n2473 & n2476 ) ;
  assign n2478 = n2461 | n2463 ;
  assign n2479 = ~n2464 & n2478 ;
  assign n2480 = n2469 | n2471 ;
  assign n2481 = ~n2472 & n2480 ;
  assign n2482 = n2479 & n2481 ;
  assign n2483 = ( n2475 & n2477 ) | ( n2475 & n2482 ) | ( n2477 & n2482 ) ;
  assign n2484 = ( n2465 & n2473 ) | ( n2465 & n2483 ) | ( n2473 & n2483 ) ;
  assign n2485 = ( x16 & x17 ) | ( x16 & x18 ) | ( x17 & x18 ) ;
  assign n2486 = ( x13 & x14 ) | ( x13 & x15 ) | ( x14 & x15 ) ;
  assign n2487 = ( ~x16 & x17 ) | ( ~x16 & x18 ) | ( x17 & x18 ) ;
  assign n2488 = ( x16 & ~n2485 ) | ( x16 & n2487 ) | ( ~n2485 & n2487 ) ;
  assign n2489 = ( ~x13 & x14 ) | ( ~x13 & x15 ) | ( x14 & x15 ) ;
  assign n2490 = ( x13 & ~n2486 ) | ( x13 & n2489 ) | ( ~n2486 & n2489 ) ;
  assign n2491 = n2488 & n2490 ;
  assign n2492 = ( n2485 & n2486 ) | ( n2485 & n2491 ) | ( n2486 & n2491 ) ;
  assign n2493 = ( x7 & x8 ) | ( x7 & x9 ) | ( x8 & x9 ) ;
  assign n2494 = ( x10 & x11 ) | ( x10 & x12 ) | ( x11 & x12 ) ;
  assign n2495 = ( ~x10 & x11 ) | ( ~x10 & x12 ) | ( x11 & x12 ) ;
  assign n2496 = ( x10 & ~n2494 ) | ( x10 & n2495 ) | ( ~n2494 & n2495 ) ;
  assign n2497 = ( ~x7 & x8 ) | ( ~x7 & x9 ) | ( x8 & x9 ) ;
  assign n2498 = ( x7 & ~n2493 ) | ( x7 & n2497 ) | ( ~n2493 & n2497 ) ;
  assign n2499 = n2496 & n2498 ;
  assign n2500 = ( n2493 & n2494 ) | ( n2493 & n2499 ) | ( n2494 & n2499 ) ;
  assign n2501 = ( ~n2485 & n2486 ) | ( ~n2485 & n2491 ) | ( n2486 & n2491 ) ;
  assign n2502 = ( n2485 & ~n2492 ) | ( n2485 & n2501 ) | ( ~n2492 & n2501 ) ;
  assign n2503 = ( ~n2493 & n2494 ) | ( ~n2493 & n2499 ) | ( n2494 & n2499 ) ;
  assign n2504 = ( n2493 & ~n2500 ) | ( n2493 & n2503 ) | ( ~n2500 & n2503 ) ;
  assign n2505 = n2496 | n2498 ;
  assign n2506 = ~n2499 & n2505 ;
  assign n2507 = ( n2488 & n2490 ) | ( n2488 & n2506 ) | ( n2490 & n2506 ) ;
  assign n2508 = ~n2491 & n2507 ;
  assign n2509 = ( n2502 & n2504 ) | ( n2502 & n2508 ) | ( n2504 & n2508 ) ;
  assign n2510 = ( n2492 & n2500 ) | ( n2492 & n2509 ) | ( n2500 & n2509 ) ;
  assign n2511 = ( ~n2492 & n2500 ) | ( ~n2492 & n2509 ) | ( n2500 & n2509 ) ;
  assign n2512 = ( n2492 & ~n2510 ) | ( n2492 & n2511 ) | ( ~n2510 & n2511 ) ;
  assign n2513 = ( ~n2465 & n2473 ) | ( ~n2465 & n2483 ) | ( n2473 & n2483 ) ;
  assign n2514 = ( n2465 & ~n2484 ) | ( n2465 & n2513 ) | ( ~n2484 & n2513 ) ;
  assign n2515 = ( ~n2475 & n2477 ) | ( ~n2475 & n2482 ) | ( n2477 & n2482 ) ;
  assign n2516 = ( n2475 & ~n2483 ) | ( n2475 & n2515 ) | ( ~n2483 & n2515 ) ;
  assign n2517 = ( ~n2502 & n2504 ) | ( ~n2502 & n2508 ) | ( n2504 & n2508 ) ;
  assign n2518 = ( n2502 & ~n2509 ) | ( n2502 & n2517 ) | ( ~n2509 & n2517 ) ;
  assign n2519 = ( ~n2488 & n2490 ) | ( ~n2488 & n2506 ) | ( n2490 & n2506 ) ;
  assign n2520 = ( n2488 & ~n2507 ) | ( n2488 & n2519 ) | ( ~n2507 & n2519 ) ;
  assign n2521 = ( n2479 & n2481 ) | ( n2479 & n2520 ) | ( n2481 & n2520 ) ;
  assign n2522 = ~n2482 & n2521 ;
  assign n2523 = ( n2516 & n2518 ) | ( n2516 & n2522 ) | ( n2518 & n2522 ) ;
  assign n2524 = ( n2512 & n2514 ) | ( n2512 & n2523 ) | ( n2514 & n2523 ) ;
  assign n2525 = ( n2484 & n2510 ) | ( n2484 & n2524 ) | ( n2510 & n2524 ) ;
  assign n2526 = ( ~n2484 & n2510 ) | ( ~n2484 & n2524 ) | ( n2510 & n2524 ) ;
  assign n2527 = ( n2484 & ~n2525 ) | ( n2484 & n2526 ) | ( ~n2525 & n2526 ) ;
  assign n2528 = ( x0 & x1 ) | ( x0 & x2 ) | ( x1 & x2 ) ;
  assign n2529 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n2530 = ( ~x0 & x1 ) | ( ~x0 & x2 ) | ( x1 & x2 ) ;
  assign n2531 = ( x0 & ~n2528 ) | ( x0 & n2530 ) | ( ~n2528 & n2530 ) ;
  assign n2532 = ( ~x3 & x4 ) | ( ~x3 & x5 ) | ( x4 & x5 ) ;
  assign n2533 = ( x3 & ~n2529 ) | ( x3 & n2532 ) | ( ~n2529 & n2532 ) ;
  assign n2534 = ( x6 & n2531 ) | ( x6 & n2533 ) | ( n2531 & n2533 ) ;
  assign n2535 = ( n2528 & n2529 ) | ( n2528 & n2534 ) | ( n2529 & n2534 ) ;
  assign n2536 = ( ~n2528 & n2529 ) | ( ~n2528 & n2534 ) | ( n2529 & n2534 ) ;
  assign n2537 = ( n2528 & ~n2535 ) | ( n2528 & n2536 ) | ( ~n2535 & n2536 ) ;
  assign n2538 = ( x997 & x998 ) | ( x997 & x999 ) | ( x998 & x999 ) ;
  assign n2539 = ( ~x6 & n2531 ) | ( ~x6 & n2533 ) | ( n2531 & n2533 ) ;
  assign n2540 = ( x6 & ~n2534 ) | ( x6 & n2539 ) | ( ~n2534 & n2539 ) ;
  assign n2541 = ( ~x997 & x998 ) | ( ~x997 & x999 ) | ( x998 & x999 ) ;
  assign n2542 = ( x997 & ~n2538 ) | ( x997 & n2541 ) | ( ~n2538 & n2541 ) ;
  assign n2543 = n2540 & n2542 ;
  assign n2544 = ( n2537 & n2538 ) | ( n2537 & n2543 ) | ( n2538 & n2543 ) ;
  assign n2545 = ( x994 & x995 ) | ( x994 & x996 ) | ( x995 & x996 ) ;
  assign n2546 = ( x991 & x992 ) | ( x991 & x993 ) | ( x992 & x993 ) ;
  assign n2547 = ( ~x994 & x995 ) | ( ~x994 & x996 ) | ( x995 & x996 ) ;
  assign n2548 = ( x994 & ~n2545 ) | ( x994 & n2547 ) | ( ~n2545 & n2547 ) ;
  assign n2549 = ( x991 & x992 ) | ( x991 & ~x993 ) | ( x992 & ~x993 ) ;
  assign n2550 = ( x993 & ~n2546 ) | ( x993 & n2549 ) | ( ~n2546 & n2549 ) ;
  assign n2551 = n2548 & n2550 ;
  assign n2552 = ( n2545 & n2546 ) | ( n2545 & n2551 ) | ( n2546 & n2551 ) ;
  assign n2553 = ~n2535 & n2544 ;
  assign n2554 = ( n2544 & n2552 ) | ( n2544 & n2553 ) | ( n2552 & n2553 ) ;
  assign n2555 = n2548 | n2550 ;
  assign n2556 = ~n2551 & n2555 ;
  assign n2557 = ( ~x997 & x998 ) | ( ~x997 & n2540 ) | ( x998 & n2540 ) ;
  assign n2558 = ( x997 & x998 ) | ( x997 & n2540 ) | ( x998 & n2540 ) ;
  assign n2559 = ( x997 & n2557 ) | ( x997 & ~n2558 ) | ( n2557 & ~n2558 ) ;
  assign n2560 = ( x999 & ~n2556 ) | ( x999 & n2559 ) | ( ~n2556 & n2559 ) ;
  assign n2561 = ( x999 & n2556 ) | ( x999 & n2559 ) | ( n2556 & n2559 ) ;
  assign n2562 = ~n2560 & n2561 ;
  assign n2563 = ( ~n2537 & n2538 ) | ( ~n2537 & n2543 ) | ( n2538 & n2543 ) ;
  assign n2564 = ( n2537 & ~n2544 ) | ( n2537 & n2563 ) | ( ~n2544 & n2563 ) ;
  assign n2565 = ( ~n2545 & n2546 ) | ( ~n2545 & n2551 ) | ( n2546 & n2551 ) ;
  assign n2566 = ( n2545 & ~n2552 ) | ( n2545 & n2565 ) | ( ~n2552 & n2565 ) ;
  assign n2567 = ( n2562 & n2564 ) | ( n2562 & n2566 ) | ( n2564 & n2566 ) ;
  assign n2568 = ( n2544 & n2553 ) | ( n2544 & ~n2567 ) | ( n2553 & ~n2567 ) ;
  assign n2569 = n2535 | n2544 ;
  assign n2570 = ( n2552 & n2567 ) | ( n2552 & n2569 ) | ( n2567 & n2569 ) ;
  assign n2571 = ( ~n2554 & n2568 ) | ( ~n2554 & n2570 ) | ( n2568 & n2570 ) ;
  assign n2572 = ( ~n2512 & n2514 ) | ( ~n2512 & n2523 ) | ( n2514 & n2523 ) ;
  assign n2573 = ( n2512 & ~n2524 ) | ( n2512 & n2572 ) | ( ~n2524 & n2572 ) ;
  assign n2574 = ( ~n2544 & n2553 ) | ( ~n2544 & n2569 ) | ( n2553 & n2569 ) ;
  assign n2575 = ( n2552 & n2567 ) | ( n2552 & n2574 ) | ( n2567 & n2574 ) ;
  assign n2576 = ( ~n2552 & n2567 ) | ( ~n2552 & n2574 ) | ( n2567 & n2574 ) ;
  assign n2577 = ( n2552 & ~n2575 ) | ( n2552 & n2576 ) | ( ~n2575 & n2576 ) ;
  assign n2578 = ( ~n2479 & n2481 ) | ( ~n2479 & n2520 ) | ( n2481 & n2520 ) ;
  assign n2579 = ( n2479 & ~n2521 ) | ( n2479 & n2578 ) | ( ~n2521 & n2578 ) ;
  assign n2580 = ( n2556 & n2560 ) | ( n2556 & ~n2561 ) | ( n2560 & ~n2561 ) ;
  assign n2581 = n2579 & n2580 ;
  assign n2582 = ( n2516 & n2518 ) | ( n2516 & ~n2522 ) | ( n2518 & ~n2522 ) ;
  assign n2583 = ( n2522 & ~n2523 ) | ( n2522 & n2582 ) | ( ~n2523 & n2582 ) ;
  assign n2584 = ( ~n2562 & n2564 ) | ( ~n2562 & n2566 ) | ( n2564 & n2566 ) ;
  assign n2585 = ( n2562 & ~n2567 ) | ( n2562 & n2584 ) | ( ~n2567 & n2584 ) ;
  assign n2586 = ( n2581 & n2583 ) | ( n2581 & n2585 ) | ( n2583 & n2585 ) ;
  assign n2587 = ( n2573 & n2577 ) | ( n2573 & n2586 ) | ( n2577 & n2586 ) ;
  assign n2588 = ( n2527 & n2571 ) | ( n2527 & n2587 ) | ( n2571 & n2587 ) ;
  assign n2589 = n2570 & ~n2571 ;
  assign n2590 = ( n2525 & n2588 ) | ( n2525 & n2589 ) | ( n2588 & n2589 ) ;
  assign n2591 = ( x76 & x77 ) | ( x76 & x78 ) | ( x77 & x78 ) ;
  assign n2592 = ( x73 & x74 ) | ( x73 & x75 ) | ( x74 & x75 ) ;
  assign n2593 = ( ~x76 & x77 ) | ( ~x76 & x78 ) | ( x77 & x78 ) ;
  assign n2594 = ( x76 & ~n2591 ) | ( x76 & n2593 ) | ( ~n2591 & n2593 ) ;
  assign n2595 = ( ~x73 & x74 ) | ( ~x73 & x75 ) | ( x74 & x75 ) ;
  assign n2596 = ( x73 & ~n2592 ) | ( x73 & n2595 ) | ( ~n2592 & n2595 ) ;
  assign n2597 = n2594 & n2596 ;
  assign n2598 = ( n2591 & n2592 ) | ( n2591 & n2597 ) | ( n2592 & n2597 ) ;
  assign n2599 = ( x67 & x68 ) | ( x67 & x69 ) | ( x68 & x69 ) ;
  assign n2600 = ( x70 & x71 ) | ( x70 & x72 ) | ( x71 & x72 ) ;
  assign n2601 = ( ~x70 & x71 ) | ( ~x70 & x72 ) | ( x71 & x72 ) ;
  assign n2602 = ( x70 & ~n2600 ) | ( x70 & n2601 ) | ( ~n2600 & n2601 ) ;
  assign n2603 = ( ~x67 & x68 ) | ( ~x67 & x69 ) | ( x68 & x69 ) ;
  assign n2604 = ( x67 & ~n2599 ) | ( x67 & n2603 ) | ( ~n2599 & n2603 ) ;
  assign n2605 = n2602 & n2604 ;
  assign n2606 = ( n2599 & n2600 ) | ( n2599 & n2605 ) | ( n2600 & n2605 ) ;
  assign n2607 = ( ~n2591 & n2592 ) | ( ~n2591 & n2597 ) | ( n2592 & n2597 ) ;
  assign n2608 = ( n2591 & ~n2598 ) | ( n2591 & n2607 ) | ( ~n2598 & n2607 ) ;
  assign n2609 = ( ~n2599 & n2600 ) | ( ~n2599 & n2605 ) | ( n2600 & n2605 ) ;
  assign n2610 = ( n2599 & ~n2606 ) | ( n2599 & n2609 ) | ( ~n2606 & n2609 ) ;
  assign n2611 = n2594 | n2596 ;
  assign n2612 = ~n2597 & n2611 ;
  assign n2613 = n2602 | n2604 ;
  assign n2614 = ~n2605 & n2613 ;
  assign n2615 = n2612 & n2614 ;
  assign n2616 = ( n2608 & n2610 ) | ( n2608 & n2615 ) | ( n2610 & n2615 ) ;
  assign n2617 = ( n2598 & n2606 ) | ( n2598 & n2616 ) | ( n2606 & n2616 ) ;
  assign n2618 = ( x64 & x65 ) | ( x64 & x66 ) | ( x65 & x66 ) ;
  assign n2619 = ( x61 & x62 ) | ( x61 & x63 ) | ( x62 & x63 ) ;
  assign n2620 = ( ~x64 & x65 ) | ( ~x64 & x66 ) | ( x65 & x66 ) ;
  assign n2621 = ( x64 & ~n2618 ) | ( x64 & n2620 ) | ( ~n2618 & n2620 ) ;
  assign n2622 = ( ~x61 & x62 ) | ( ~x61 & x63 ) | ( x62 & x63 ) ;
  assign n2623 = ( x61 & ~n2619 ) | ( x61 & n2622 ) | ( ~n2619 & n2622 ) ;
  assign n2624 = n2621 & n2623 ;
  assign n2625 = ( n2618 & n2619 ) | ( n2618 & n2624 ) | ( n2619 & n2624 ) ;
  assign n2626 = ( x55 & x56 ) | ( x55 & x57 ) | ( x56 & x57 ) ;
  assign n2627 = ( x58 & x59 ) | ( x58 & x60 ) | ( x59 & x60 ) ;
  assign n2628 = ( ~x58 & x59 ) | ( ~x58 & x60 ) | ( x59 & x60 ) ;
  assign n2629 = ( x58 & ~n2627 ) | ( x58 & n2628 ) | ( ~n2627 & n2628 ) ;
  assign n2630 = ( ~x55 & x56 ) | ( ~x55 & x57 ) | ( x56 & x57 ) ;
  assign n2631 = ( x55 & ~n2626 ) | ( x55 & n2630 ) | ( ~n2626 & n2630 ) ;
  assign n2632 = n2629 & n2631 ;
  assign n2633 = ( n2626 & n2627 ) | ( n2626 & n2632 ) | ( n2627 & n2632 ) ;
  assign n2634 = ( ~n2618 & n2619 ) | ( ~n2618 & n2624 ) | ( n2619 & n2624 ) ;
  assign n2635 = ( n2618 & ~n2625 ) | ( n2618 & n2634 ) | ( ~n2625 & n2634 ) ;
  assign n2636 = ( ~n2626 & n2627 ) | ( ~n2626 & n2632 ) | ( n2627 & n2632 ) ;
  assign n2637 = ( n2626 & ~n2633 ) | ( n2626 & n2636 ) | ( ~n2633 & n2636 ) ;
  assign n2638 = n2629 | n2631 ;
  assign n2639 = ~n2632 & n2638 ;
  assign n2640 = ( n2621 & n2623 ) | ( n2621 & n2639 ) | ( n2623 & n2639 ) ;
  assign n2641 = ~n2624 & n2640 ;
  assign n2642 = ( n2635 & n2637 ) | ( n2635 & n2641 ) | ( n2637 & n2641 ) ;
  assign n2643 = ( n2625 & n2633 ) | ( n2625 & n2642 ) | ( n2633 & n2642 ) ;
  assign n2644 = ( ~n2625 & n2633 ) | ( ~n2625 & n2642 ) | ( n2633 & n2642 ) ;
  assign n2645 = ( n2625 & ~n2643 ) | ( n2625 & n2644 ) | ( ~n2643 & n2644 ) ;
  assign n2646 = ( ~n2598 & n2606 ) | ( ~n2598 & n2616 ) | ( n2606 & n2616 ) ;
  assign n2647 = ( n2598 & ~n2617 ) | ( n2598 & n2646 ) | ( ~n2617 & n2646 ) ;
  assign n2648 = ( ~n2608 & n2610 ) | ( ~n2608 & n2615 ) | ( n2610 & n2615 ) ;
  assign n2649 = ( n2608 & ~n2616 ) | ( n2608 & n2648 ) | ( ~n2616 & n2648 ) ;
  assign n2650 = ( ~n2635 & n2637 ) | ( ~n2635 & n2641 ) | ( n2637 & n2641 ) ;
  assign n2651 = ( n2635 & ~n2642 ) | ( n2635 & n2650 ) | ( ~n2642 & n2650 ) ;
  assign n2652 = ( ~n2621 & n2623 ) | ( ~n2621 & n2639 ) | ( n2623 & n2639 ) ;
  assign n2653 = ( n2621 & ~n2640 ) | ( n2621 & n2652 ) | ( ~n2640 & n2652 ) ;
  assign n2654 = ( n2612 & n2614 ) | ( n2612 & n2653 ) | ( n2614 & n2653 ) ;
  assign n2655 = ~n2615 & n2654 ;
  assign n2656 = ( n2649 & n2651 ) | ( n2649 & n2655 ) | ( n2651 & n2655 ) ;
  assign n2657 = ( n2645 & n2647 ) | ( n2645 & n2656 ) | ( n2647 & n2656 ) ;
  assign n2658 = ( n2617 & n2643 ) | ( n2617 & n2657 ) | ( n2643 & n2657 ) ;
  assign n2659 = ( x52 & x53 ) | ( x52 & x54 ) | ( x53 & x54 ) ;
  assign n2660 = ( x49 & x50 ) | ( x49 & x51 ) | ( x50 & x51 ) ;
  assign n2661 = ( ~x52 & x53 ) | ( ~x52 & x54 ) | ( x53 & x54 ) ;
  assign n2662 = ( x52 & ~n2659 ) | ( x52 & n2661 ) | ( ~n2659 & n2661 ) ;
  assign n2663 = ( ~x49 & x50 ) | ( ~x49 & x51 ) | ( x50 & x51 ) ;
  assign n2664 = ( x49 & ~n2660 ) | ( x49 & n2663 ) | ( ~n2660 & n2663 ) ;
  assign n2665 = n2662 & n2664 ;
  assign n2666 = ( n2659 & n2660 ) | ( n2659 & n2665 ) | ( n2660 & n2665 ) ;
  assign n2667 = ( x43 & x44 ) | ( x43 & x45 ) | ( x44 & x45 ) ;
  assign n2668 = ( x46 & x47 ) | ( x46 & x48 ) | ( x47 & x48 ) ;
  assign n2669 = ( ~x46 & x47 ) | ( ~x46 & x48 ) | ( x47 & x48 ) ;
  assign n2670 = ( x46 & ~n2668 ) | ( x46 & n2669 ) | ( ~n2668 & n2669 ) ;
  assign n2671 = ( ~x43 & x44 ) | ( ~x43 & x45 ) | ( x44 & x45 ) ;
  assign n2672 = ( x43 & ~n2667 ) | ( x43 & n2671 ) | ( ~n2667 & n2671 ) ;
  assign n2673 = n2670 & n2672 ;
  assign n2674 = ( n2667 & n2668 ) | ( n2667 & n2673 ) | ( n2668 & n2673 ) ;
  assign n2675 = ( ~n2659 & n2660 ) | ( ~n2659 & n2665 ) | ( n2660 & n2665 ) ;
  assign n2676 = ( n2659 & ~n2666 ) | ( n2659 & n2675 ) | ( ~n2666 & n2675 ) ;
  assign n2677 = ( ~n2667 & n2668 ) | ( ~n2667 & n2673 ) | ( n2668 & n2673 ) ;
  assign n2678 = ( n2667 & ~n2674 ) | ( n2667 & n2677 ) | ( ~n2674 & n2677 ) ;
  assign n2679 = n2662 | n2664 ;
  assign n2680 = ~n2665 & n2679 ;
  assign n2681 = n2670 | n2672 ;
  assign n2682 = ~n2673 & n2681 ;
  assign n2683 = n2680 & n2682 ;
  assign n2684 = ( n2676 & n2678 ) | ( n2676 & n2683 ) | ( n2678 & n2683 ) ;
  assign n2685 = ( n2666 & n2674 ) | ( n2666 & n2684 ) | ( n2674 & n2684 ) ;
  assign n2686 = ( x40 & x41 ) | ( x40 & x42 ) | ( x41 & x42 ) ;
  assign n2687 = ( x37 & x38 ) | ( x37 & x39 ) | ( x38 & x39 ) ;
  assign n2688 = ( ~x40 & x41 ) | ( ~x40 & x42 ) | ( x41 & x42 ) ;
  assign n2689 = ( x40 & ~n2686 ) | ( x40 & n2688 ) | ( ~n2686 & n2688 ) ;
  assign n2690 = ( ~x37 & x38 ) | ( ~x37 & x39 ) | ( x38 & x39 ) ;
  assign n2691 = ( x37 & ~n2687 ) | ( x37 & n2690 ) | ( ~n2687 & n2690 ) ;
  assign n2692 = n2689 & n2691 ;
  assign n2693 = ( n2686 & n2687 ) | ( n2686 & n2692 ) | ( n2687 & n2692 ) ;
  assign n2694 = ( x31 & x32 ) | ( x31 & x33 ) | ( x32 & x33 ) ;
  assign n2695 = ( x34 & x35 ) | ( x34 & x36 ) | ( x35 & x36 ) ;
  assign n2696 = ( ~x34 & x35 ) | ( ~x34 & x36 ) | ( x35 & x36 ) ;
  assign n2697 = ( x34 & ~n2695 ) | ( x34 & n2696 ) | ( ~n2695 & n2696 ) ;
  assign n2698 = ( ~x31 & x32 ) | ( ~x31 & x33 ) | ( x32 & x33 ) ;
  assign n2699 = ( x31 & ~n2694 ) | ( x31 & n2698 ) | ( ~n2694 & n2698 ) ;
  assign n2700 = n2697 & n2699 ;
  assign n2701 = ( n2694 & n2695 ) | ( n2694 & n2700 ) | ( n2695 & n2700 ) ;
  assign n2702 = ( ~n2686 & n2687 ) | ( ~n2686 & n2692 ) | ( n2687 & n2692 ) ;
  assign n2703 = ( n2686 & ~n2693 ) | ( n2686 & n2702 ) | ( ~n2693 & n2702 ) ;
  assign n2704 = ( ~n2694 & n2695 ) | ( ~n2694 & n2700 ) | ( n2695 & n2700 ) ;
  assign n2705 = ( n2694 & ~n2701 ) | ( n2694 & n2704 ) | ( ~n2701 & n2704 ) ;
  assign n2706 = n2697 | n2699 ;
  assign n2707 = ~n2700 & n2706 ;
  assign n2708 = ( n2689 & n2691 ) | ( n2689 & n2707 ) | ( n2691 & n2707 ) ;
  assign n2709 = ~n2692 & n2708 ;
  assign n2710 = ( n2703 & n2705 ) | ( n2703 & n2709 ) | ( n2705 & n2709 ) ;
  assign n2711 = ( n2693 & n2701 ) | ( n2693 & n2710 ) | ( n2701 & n2710 ) ;
  assign n2712 = ( ~n2693 & n2701 ) | ( ~n2693 & n2710 ) | ( n2701 & n2710 ) ;
  assign n2713 = ( n2693 & ~n2711 ) | ( n2693 & n2712 ) | ( ~n2711 & n2712 ) ;
  assign n2714 = ( ~n2666 & n2674 ) | ( ~n2666 & n2684 ) | ( n2674 & n2684 ) ;
  assign n2715 = ( n2666 & ~n2685 ) | ( n2666 & n2714 ) | ( ~n2685 & n2714 ) ;
  assign n2716 = ( ~n2676 & n2678 ) | ( ~n2676 & n2683 ) | ( n2678 & n2683 ) ;
  assign n2717 = ( n2676 & ~n2684 ) | ( n2676 & n2716 ) | ( ~n2684 & n2716 ) ;
  assign n2718 = ( ~n2703 & n2705 ) | ( ~n2703 & n2709 ) | ( n2705 & n2709 ) ;
  assign n2719 = ( n2703 & ~n2710 ) | ( n2703 & n2718 ) | ( ~n2710 & n2718 ) ;
  assign n2720 = ( ~n2689 & n2691 ) | ( ~n2689 & n2707 ) | ( n2691 & n2707 ) ;
  assign n2721 = ( n2689 & ~n2708 ) | ( n2689 & n2720 ) | ( ~n2708 & n2720 ) ;
  assign n2722 = ( n2680 & n2682 ) | ( n2680 & n2721 ) | ( n2682 & n2721 ) ;
  assign n2723 = ~n2683 & n2722 ;
  assign n2724 = ( n2717 & n2719 ) | ( n2717 & n2723 ) | ( n2719 & n2723 ) ;
  assign n2725 = ( n2713 & n2715 ) | ( n2713 & n2724 ) | ( n2715 & n2724 ) ;
  assign n2726 = ( n2685 & n2711 ) | ( n2685 & n2725 ) | ( n2711 & n2725 ) ;
  assign n2727 = ( ~n2617 & n2643 ) | ( ~n2617 & n2657 ) | ( n2643 & n2657 ) ;
  assign n2728 = ( n2617 & ~n2658 ) | ( n2617 & n2727 ) | ( ~n2658 & n2727 ) ;
  assign n2729 = ( ~n2685 & n2711 ) | ( ~n2685 & n2725 ) | ( n2711 & n2725 ) ;
  assign n2730 = ( n2685 & ~n2726 ) | ( n2685 & n2729 ) | ( ~n2726 & n2729 ) ;
  assign n2731 = ( ~n2713 & n2715 ) | ( ~n2713 & n2724 ) | ( n2715 & n2724 ) ;
  assign n2732 = ( n2713 & ~n2725 ) | ( n2713 & n2731 ) | ( ~n2725 & n2731 ) ;
  assign n2733 = ( ~n2645 & n2647 ) | ( ~n2645 & n2656 ) | ( n2647 & n2656 ) ;
  assign n2734 = ( n2645 & ~n2657 ) | ( n2645 & n2733 ) | ( ~n2657 & n2733 ) ;
  assign n2735 = ( ~n2612 & n2614 ) | ( ~n2612 & n2653 ) | ( n2614 & n2653 ) ;
  assign n2736 = ( n2612 & ~n2654 ) | ( n2612 & n2735 ) | ( ~n2654 & n2735 ) ;
  assign n2737 = ( ~n2680 & n2682 ) | ( ~n2680 & n2721 ) | ( n2682 & n2721 ) ;
  assign n2738 = ( n2680 & ~n2722 ) | ( n2680 & n2737 ) | ( ~n2722 & n2737 ) ;
  assign n2739 = n2736 & n2738 ;
  assign n2740 = ( n2649 & n2651 ) | ( n2649 & ~n2655 ) | ( n2651 & ~n2655 ) ;
  assign n2741 = ( n2655 & ~n2656 ) | ( n2655 & n2740 ) | ( ~n2656 & n2740 ) ;
  assign n2742 = ( n2717 & n2719 ) | ( n2717 & ~n2723 ) | ( n2719 & ~n2723 ) ;
  assign n2743 = ( n2723 & ~n2724 ) | ( n2723 & n2742 ) | ( ~n2724 & n2742 ) ;
  assign n2744 = ( n2739 & n2741 ) | ( n2739 & n2743 ) | ( n2741 & n2743 ) ;
  assign n2745 = ( n2732 & n2734 ) | ( n2732 & n2744 ) | ( n2734 & n2744 ) ;
  assign n2746 = ( n2728 & n2730 ) | ( n2728 & n2745 ) | ( n2730 & n2745 ) ;
  assign n2747 = ( n2658 & n2726 ) | ( n2658 & n2746 ) | ( n2726 & n2746 ) ;
  assign n2748 = ( ~n2525 & n2588 ) | ( ~n2525 & n2589 ) | ( n2588 & n2589 ) ;
  assign n2749 = ( n2525 & ~n2590 ) | ( n2525 & n2748 ) | ( ~n2590 & n2748 ) ;
  assign n2750 = ( ~n2658 & n2726 ) | ( ~n2658 & n2746 ) | ( n2726 & n2746 ) ;
  assign n2751 = ( n2658 & ~n2747 ) | ( n2658 & n2750 ) | ( ~n2747 & n2750 ) ;
  assign n2752 = ( ~n2728 & n2730 ) | ( ~n2728 & n2745 ) | ( n2730 & n2745 ) ;
  assign n2753 = ( n2728 & ~n2746 ) | ( n2728 & n2752 ) | ( ~n2746 & n2752 ) ;
  assign n2754 = ( ~n2527 & n2571 ) | ( ~n2527 & n2587 ) | ( n2571 & n2587 ) ;
  assign n2755 = ( n2527 & ~n2588 ) | ( n2527 & n2754 ) | ( ~n2588 & n2754 ) ;
  assign n2756 = ( ~n2573 & n2577 ) | ( ~n2573 & n2586 ) | ( n2577 & n2586 ) ;
  assign n2757 = ( n2573 & ~n2587 ) | ( n2573 & n2756 ) | ( ~n2587 & n2756 ) ;
  assign n2758 = ( ~n2732 & n2734 ) | ( ~n2732 & n2744 ) | ( n2734 & n2744 ) ;
  assign n2759 = ( n2732 & ~n2745 ) | ( n2732 & n2758 ) | ( ~n2745 & n2758 ) ;
  assign n2760 = ( ~n2739 & n2741 ) | ( ~n2739 & n2743 ) | ( n2741 & n2743 ) ;
  assign n2761 = ( n2739 & ~n2744 ) | ( n2739 & n2760 ) | ( ~n2744 & n2760 ) ;
  assign n2762 = ( ~n2581 & n2583 ) | ( ~n2581 & n2585 ) | ( n2583 & n2585 ) ;
  assign n2763 = ( n2581 & ~n2586 ) | ( n2581 & n2762 ) | ( ~n2586 & n2762 ) ;
  assign n2764 = n2736 | n2738 ;
  assign n2765 = ~n2739 & n2764 ;
  assign n2766 = n2579 | n2580 ;
  assign n2767 = ~n2581 & n2766 ;
  assign n2768 = n2765 & n2767 ;
  assign n2769 = ( n2761 & n2763 ) | ( n2761 & n2768 ) | ( n2763 & n2768 ) ;
  assign n2770 = ( n2757 & n2759 ) | ( n2757 & n2769 ) | ( n2759 & n2769 ) ;
  assign n2771 = ( n2753 & n2755 ) | ( n2753 & n2770 ) | ( n2755 & n2770 ) ;
  assign n2772 = ( n2749 & n2751 ) | ( n2749 & n2771 ) | ( n2751 & n2771 ) ;
  assign n2773 = ( n2590 & n2747 ) | ( n2590 & n2772 ) | ( n2747 & n2772 ) ;
  assign n2774 = ( ~n2590 & n2747 ) | ( ~n2590 & n2772 ) | ( n2747 & n2772 ) ;
  assign n2775 = ( n2590 & ~n2773 ) | ( n2590 & n2774 ) | ( ~n2773 & n2774 ) ;
  assign n2776 = ( x988 & x989 ) | ( x988 & x990 ) | ( x989 & x990 ) ;
  assign n2777 = ( x985 & x986 ) | ( x985 & x987 ) | ( x986 & x987 ) ;
  assign n2778 = ( ~x988 & x989 ) | ( ~x988 & x990 ) | ( x989 & x990 ) ;
  assign n2779 = ( x988 & ~n2776 ) | ( x988 & n2778 ) | ( ~n2776 & n2778 ) ;
  assign n2780 = ( ~x985 & x986 ) | ( ~x985 & x987 ) | ( x986 & x987 ) ;
  assign n2781 = ( x985 & ~n2777 ) | ( x985 & n2780 ) | ( ~n2777 & n2780 ) ;
  assign n2782 = n2779 & n2781 ;
  assign n2783 = ( n2776 & n2777 ) | ( n2776 & n2782 ) | ( n2777 & n2782 ) ;
  assign n2784 = ( x979 & x980 ) | ( x979 & x981 ) | ( x980 & x981 ) ;
  assign n2785 = ( x982 & x983 ) | ( x982 & x984 ) | ( x983 & x984 ) ;
  assign n2786 = ( ~x982 & x983 ) | ( ~x982 & x984 ) | ( x983 & x984 ) ;
  assign n2787 = ( x982 & ~n2785 ) | ( x982 & n2786 ) | ( ~n2785 & n2786 ) ;
  assign n2788 = ( ~x979 & x980 ) | ( ~x979 & x981 ) | ( x980 & x981 ) ;
  assign n2789 = ( x979 & ~n2784 ) | ( x979 & n2788 ) | ( ~n2784 & n2788 ) ;
  assign n2790 = n2787 & n2789 ;
  assign n2791 = ( n2784 & n2785 ) | ( n2784 & n2790 ) | ( n2785 & n2790 ) ;
  assign n2792 = ( ~n2776 & n2777 ) | ( ~n2776 & n2782 ) | ( n2777 & n2782 ) ;
  assign n2793 = ( n2776 & ~n2783 ) | ( n2776 & n2792 ) | ( ~n2783 & n2792 ) ;
  assign n2794 = ( ~n2784 & n2785 ) | ( ~n2784 & n2790 ) | ( n2785 & n2790 ) ;
  assign n2795 = ( n2784 & ~n2791 ) | ( n2784 & n2794 ) | ( ~n2791 & n2794 ) ;
  assign n2796 = n2779 | n2781 ;
  assign n2797 = ~n2782 & n2796 ;
  assign n2798 = n2787 | n2789 ;
  assign n2799 = ~n2790 & n2798 ;
  assign n2800 = n2797 & n2799 ;
  assign n2801 = ( n2793 & n2795 ) | ( n2793 & n2800 ) | ( n2795 & n2800 ) ;
  assign n2802 = ( n2783 & n2791 ) | ( n2783 & n2801 ) | ( n2791 & n2801 ) ;
  assign n2803 = ( x976 & x977 ) | ( x976 & x978 ) | ( x977 & x978 ) ;
  assign n2804 = ( x973 & x974 ) | ( x973 & x975 ) | ( x974 & x975 ) ;
  assign n2805 = ( ~x976 & x977 ) | ( ~x976 & x978 ) | ( x977 & x978 ) ;
  assign n2806 = ( x976 & ~n2803 ) | ( x976 & n2805 ) | ( ~n2803 & n2805 ) ;
  assign n2807 = ( ~x973 & x974 ) | ( ~x973 & x975 ) | ( x974 & x975 ) ;
  assign n2808 = ( x973 & ~n2804 ) | ( x973 & n2807 ) | ( ~n2804 & n2807 ) ;
  assign n2809 = n2806 & n2808 ;
  assign n2810 = ( n2803 & n2804 ) | ( n2803 & n2809 ) | ( n2804 & n2809 ) ;
  assign n2811 = ( x967 & x968 ) | ( x967 & x969 ) | ( x968 & x969 ) ;
  assign n2812 = ( x970 & x971 ) | ( x970 & x972 ) | ( x971 & x972 ) ;
  assign n2813 = ( ~x970 & x971 ) | ( ~x970 & x972 ) | ( x971 & x972 ) ;
  assign n2814 = ( x970 & ~n2812 ) | ( x970 & n2813 ) | ( ~n2812 & n2813 ) ;
  assign n2815 = ( ~x967 & x968 ) | ( ~x967 & x969 ) | ( x968 & x969 ) ;
  assign n2816 = ( x967 & ~n2811 ) | ( x967 & n2815 ) | ( ~n2811 & n2815 ) ;
  assign n2817 = n2814 & n2816 ;
  assign n2818 = ( n2811 & n2812 ) | ( n2811 & n2817 ) | ( n2812 & n2817 ) ;
  assign n2819 = ( ~n2803 & n2804 ) | ( ~n2803 & n2809 ) | ( n2804 & n2809 ) ;
  assign n2820 = ( n2803 & ~n2810 ) | ( n2803 & n2819 ) | ( ~n2810 & n2819 ) ;
  assign n2821 = ( ~n2811 & n2812 ) | ( ~n2811 & n2817 ) | ( n2812 & n2817 ) ;
  assign n2822 = ( n2811 & ~n2818 ) | ( n2811 & n2821 ) | ( ~n2818 & n2821 ) ;
  assign n2823 = n2814 | n2816 ;
  assign n2824 = ~n2817 & n2823 ;
  assign n2825 = ( n2806 & n2808 ) | ( n2806 & n2824 ) | ( n2808 & n2824 ) ;
  assign n2826 = ~n2809 & n2825 ;
  assign n2827 = ( n2820 & n2822 ) | ( n2820 & n2826 ) | ( n2822 & n2826 ) ;
  assign n2828 = ( n2810 & n2818 ) | ( n2810 & n2827 ) | ( n2818 & n2827 ) ;
  assign n2829 = ( ~n2810 & n2818 ) | ( ~n2810 & n2827 ) | ( n2818 & n2827 ) ;
  assign n2830 = ( n2810 & ~n2828 ) | ( n2810 & n2829 ) | ( ~n2828 & n2829 ) ;
  assign n2831 = ( ~n2783 & n2791 ) | ( ~n2783 & n2801 ) | ( n2791 & n2801 ) ;
  assign n2832 = ( n2783 & ~n2802 ) | ( n2783 & n2831 ) | ( ~n2802 & n2831 ) ;
  assign n2833 = ( ~n2793 & n2795 ) | ( ~n2793 & n2800 ) | ( n2795 & n2800 ) ;
  assign n2834 = ( n2793 & ~n2801 ) | ( n2793 & n2833 ) | ( ~n2801 & n2833 ) ;
  assign n2835 = ( ~n2820 & n2822 ) | ( ~n2820 & n2826 ) | ( n2822 & n2826 ) ;
  assign n2836 = ( n2820 & ~n2827 ) | ( n2820 & n2835 ) | ( ~n2827 & n2835 ) ;
  assign n2837 = ( ~n2806 & n2808 ) | ( ~n2806 & n2824 ) | ( n2808 & n2824 ) ;
  assign n2838 = ( n2806 & ~n2825 ) | ( n2806 & n2837 ) | ( ~n2825 & n2837 ) ;
  assign n2839 = ( n2797 & n2799 ) | ( n2797 & n2838 ) | ( n2799 & n2838 ) ;
  assign n2840 = ~n2800 & n2839 ;
  assign n2841 = ( n2834 & n2836 ) | ( n2834 & n2840 ) | ( n2836 & n2840 ) ;
  assign n2842 = ( n2830 & n2832 ) | ( n2830 & n2841 ) | ( n2832 & n2841 ) ;
  assign n2843 = ( n2802 & n2828 ) | ( n2802 & n2842 ) | ( n2828 & n2842 ) ;
  assign n2844 = ( x964 & x965 ) | ( x964 & x966 ) | ( x965 & x966 ) ;
  assign n2845 = ( x961 & x962 ) | ( x961 & x963 ) | ( x962 & x963 ) ;
  assign n2846 = ( ~x964 & x965 ) | ( ~x964 & x966 ) | ( x965 & x966 ) ;
  assign n2847 = ( x964 & ~n2844 ) | ( x964 & n2846 ) | ( ~n2844 & n2846 ) ;
  assign n2848 = ( ~x961 & x962 ) | ( ~x961 & x963 ) | ( x962 & x963 ) ;
  assign n2849 = ( x961 & ~n2845 ) | ( x961 & n2848 ) | ( ~n2845 & n2848 ) ;
  assign n2850 = n2847 & n2849 ;
  assign n2851 = ( n2844 & n2845 ) | ( n2844 & n2850 ) | ( n2845 & n2850 ) ;
  assign n2852 = ( x955 & x956 ) | ( x955 & x957 ) | ( x956 & x957 ) ;
  assign n2853 = ( x958 & x959 ) | ( x958 & x960 ) | ( x959 & x960 ) ;
  assign n2854 = ( ~x958 & x959 ) | ( ~x958 & x960 ) | ( x959 & x960 ) ;
  assign n2855 = ( x958 & ~n2853 ) | ( x958 & n2854 ) | ( ~n2853 & n2854 ) ;
  assign n2856 = ( ~x955 & x956 ) | ( ~x955 & x957 ) | ( x956 & x957 ) ;
  assign n2857 = ( x955 & ~n2852 ) | ( x955 & n2856 ) | ( ~n2852 & n2856 ) ;
  assign n2858 = n2855 & n2857 ;
  assign n2859 = ( n2852 & n2853 ) | ( n2852 & n2858 ) | ( n2853 & n2858 ) ;
  assign n2860 = ( ~n2844 & n2845 ) | ( ~n2844 & n2850 ) | ( n2845 & n2850 ) ;
  assign n2861 = ( n2844 & ~n2851 ) | ( n2844 & n2860 ) | ( ~n2851 & n2860 ) ;
  assign n2862 = ( ~n2852 & n2853 ) | ( ~n2852 & n2858 ) | ( n2853 & n2858 ) ;
  assign n2863 = ( n2852 & ~n2859 ) | ( n2852 & n2862 ) | ( ~n2859 & n2862 ) ;
  assign n2864 = n2847 | n2849 ;
  assign n2865 = ~n2850 & n2864 ;
  assign n2866 = n2855 | n2857 ;
  assign n2867 = ~n2858 & n2866 ;
  assign n2868 = n2865 & n2867 ;
  assign n2869 = ( n2861 & n2863 ) | ( n2861 & n2868 ) | ( n2863 & n2868 ) ;
  assign n2870 = ( n2851 & n2859 ) | ( n2851 & n2869 ) | ( n2859 & n2869 ) ;
  assign n2871 = ( x952 & x953 ) | ( x952 & x954 ) | ( x953 & x954 ) ;
  assign n2872 = ( x949 & x950 ) | ( x949 & x951 ) | ( x950 & x951 ) ;
  assign n2873 = ( ~x952 & x953 ) | ( ~x952 & x954 ) | ( x953 & x954 ) ;
  assign n2874 = ( x952 & ~n2871 ) | ( x952 & n2873 ) | ( ~n2871 & n2873 ) ;
  assign n2875 = ( ~x949 & x950 ) | ( ~x949 & x951 ) | ( x950 & x951 ) ;
  assign n2876 = ( x949 & ~n2872 ) | ( x949 & n2875 ) | ( ~n2872 & n2875 ) ;
  assign n2877 = n2874 & n2876 ;
  assign n2878 = ( n2871 & n2872 ) | ( n2871 & n2877 ) | ( n2872 & n2877 ) ;
  assign n2879 = ( x943 & x944 ) | ( x943 & x945 ) | ( x944 & x945 ) ;
  assign n2880 = ( x946 & x947 ) | ( x946 & x948 ) | ( x947 & x948 ) ;
  assign n2881 = ( ~x946 & x947 ) | ( ~x946 & x948 ) | ( x947 & x948 ) ;
  assign n2882 = ( x946 & ~n2880 ) | ( x946 & n2881 ) | ( ~n2880 & n2881 ) ;
  assign n2883 = ( ~x943 & x944 ) | ( ~x943 & x945 ) | ( x944 & x945 ) ;
  assign n2884 = ( x943 & ~n2879 ) | ( x943 & n2883 ) | ( ~n2879 & n2883 ) ;
  assign n2885 = n2882 & n2884 ;
  assign n2886 = ( n2879 & n2880 ) | ( n2879 & n2885 ) | ( n2880 & n2885 ) ;
  assign n2887 = ( ~n2871 & n2872 ) | ( ~n2871 & n2877 ) | ( n2872 & n2877 ) ;
  assign n2888 = ( n2871 & ~n2878 ) | ( n2871 & n2887 ) | ( ~n2878 & n2887 ) ;
  assign n2889 = ( ~n2879 & n2880 ) | ( ~n2879 & n2885 ) | ( n2880 & n2885 ) ;
  assign n2890 = ( n2879 & ~n2886 ) | ( n2879 & n2889 ) | ( ~n2886 & n2889 ) ;
  assign n2891 = n2882 | n2884 ;
  assign n2892 = ~n2885 & n2891 ;
  assign n2893 = ( n2874 & n2876 ) | ( n2874 & n2892 ) | ( n2876 & n2892 ) ;
  assign n2894 = ~n2877 & n2893 ;
  assign n2895 = ( n2888 & n2890 ) | ( n2888 & n2894 ) | ( n2890 & n2894 ) ;
  assign n2896 = ( n2878 & n2886 ) | ( n2878 & n2895 ) | ( n2886 & n2895 ) ;
  assign n2897 = ( ~n2878 & n2886 ) | ( ~n2878 & n2895 ) | ( n2886 & n2895 ) ;
  assign n2898 = ( n2878 & ~n2896 ) | ( n2878 & n2897 ) | ( ~n2896 & n2897 ) ;
  assign n2899 = ( ~n2851 & n2859 ) | ( ~n2851 & n2869 ) | ( n2859 & n2869 ) ;
  assign n2900 = ( n2851 & ~n2870 ) | ( n2851 & n2899 ) | ( ~n2870 & n2899 ) ;
  assign n2901 = ( ~n2861 & n2863 ) | ( ~n2861 & n2868 ) | ( n2863 & n2868 ) ;
  assign n2902 = ( n2861 & ~n2869 ) | ( n2861 & n2901 ) | ( ~n2869 & n2901 ) ;
  assign n2903 = ( ~n2888 & n2890 ) | ( ~n2888 & n2894 ) | ( n2890 & n2894 ) ;
  assign n2904 = ( n2888 & ~n2895 ) | ( n2888 & n2903 ) | ( ~n2895 & n2903 ) ;
  assign n2905 = ( ~n2874 & n2876 ) | ( ~n2874 & n2892 ) | ( n2876 & n2892 ) ;
  assign n2906 = ( n2874 & ~n2893 ) | ( n2874 & n2905 ) | ( ~n2893 & n2905 ) ;
  assign n2907 = ( n2865 & n2867 ) | ( n2865 & n2906 ) | ( n2867 & n2906 ) ;
  assign n2908 = ~n2868 & n2907 ;
  assign n2909 = ( n2902 & n2904 ) | ( n2902 & n2908 ) | ( n2904 & n2908 ) ;
  assign n2910 = ( n2898 & n2900 ) | ( n2898 & n2909 ) | ( n2900 & n2909 ) ;
  assign n2911 = ( n2870 & n2896 ) | ( n2870 & n2910 ) | ( n2896 & n2910 ) ;
  assign n2912 = ( ~n2802 & n2828 ) | ( ~n2802 & n2842 ) | ( n2828 & n2842 ) ;
  assign n2913 = ( n2802 & ~n2843 ) | ( n2802 & n2912 ) | ( ~n2843 & n2912 ) ;
  assign n2914 = ( ~n2870 & n2896 ) | ( ~n2870 & n2910 ) | ( n2896 & n2910 ) ;
  assign n2915 = ( n2870 & ~n2911 ) | ( n2870 & n2914 ) | ( ~n2911 & n2914 ) ;
  assign n2916 = ( ~n2898 & n2900 ) | ( ~n2898 & n2909 ) | ( n2900 & n2909 ) ;
  assign n2917 = ( n2898 & ~n2910 ) | ( n2898 & n2916 ) | ( ~n2910 & n2916 ) ;
  assign n2918 = ( ~n2830 & n2832 ) | ( ~n2830 & n2841 ) | ( n2832 & n2841 ) ;
  assign n2919 = ( n2830 & ~n2842 ) | ( n2830 & n2918 ) | ( ~n2842 & n2918 ) ;
  assign n2920 = ( ~n2797 & n2799 ) | ( ~n2797 & n2838 ) | ( n2799 & n2838 ) ;
  assign n2921 = ( n2797 & ~n2839 ) | ( n2797 & n2920 ) | ( ~n2839 & n2920 ) ;
  assign n2922 = ( ~n2865 & n2867 ) | ( ~n2865 & n2906 ) | ( n2867 & n2906 ) ;
  assign n2923 = ( n2865 & ~n2907 ) | ( n2865 & n2922 ) | ( ~n2907 & n2922 ) ;
  assign n2924 = n2921 & n2923 ;
  assign n2925 = ( n2834 & n2836 ) | ( n2834 & ~n2840 ) | ( n2836 & ~n2840 ) ;
  assign n2926 = ( n2840 & ~n2841 ) | ( n2840 & n2925 ) | ( ~n2841 & n2925 ) ;
  assign n2927 = ( n2902 & n2904 ) | ( n2902 & ~n2908 ) | ( n2904 & ~n2908 ) ;
  assign n2928 = ( n2908 & ~n2909 ) | ( n2908 & n2927 ) | ( ~n2909 & n2927 ) ;
  assign n2929 = ( n2924 & n2926 ) | ( n2924 & n2928 ) | ( n2926 & n2928 ) ;
  assign n2930 = ( n2917 & n2919 ) | ( n2917 & n2929 ) | ( n2919 & n2929 ) ;
  assign n2931 = ( n2913 & n2915 ) | ( n2913 & n2930 ) | ( n2915 & n2930 ) ;
  assign n2932 = ( n2843 & n2911 ) | ( n2843 & n2931 ) | ( n2911 & n2931 ) ;
  assign n2933 = ( ~n2843 & n2911 ) | ( ~n2843 & n2931 ) | ( n2911 & n2931 ) ;
  assign n2934 = ( n2843 & ~n2932 ) | ( n2843 & n2933 ) | ( ~n2932 & n2933 ) ;
  assign n2935 = ( ~n2749 & n2751 ) | ( ~n2749 & n2771 ) | ( n2751 & n2771 ) ;
  assign n2936 = ( n2749 & ~n2772 ) | ( n2749 & n2935 ) | ( ~n2772 & n2935 ) ;
  assign n2937 = ( ~n2753 & n2755 ) | ( ~n2753 & n2770 ) | ( n2755 & n2770 ) ;
  assign n2938 = ( n2753 & ~n2771 ) | ( n2753 & n2937 ) | ( ~n2771 & n2937 ) ;
  assign n2939 = ( ~n2913 & n2915 ) | ( ~n2913 & n2930 ) | ( n2915 & n2930 ) ;
  assign n2940 = ( n2913 & ~n2931 ) | ( n2913 & n2939 ) | ( ~n2931 & n2939 ) ;
  assign n2941 = ( ~n2917 & n2919 ) | ( ~n2917 & n2929 ) | ( n2919 & n2929 ) ;
  assign n2942 = ( n2917 & ~n2930 ) | ( n2917 & n2941 ) | ( ~n2930 & n2941 ) ;
  assign n2943 = ( ~n2757 & n2759 ) | ( ~n2757 & n2769 ) | ( n2759 & n2769 ) ;
  assign n2944 = ( n2757 & ~n2770 ) | ( n2757 & n2943 ) | ( ~n2770 & n2943 ) ;
  assign n2945 = n2921 | n2923 ;
  assign n2946 = ~n2924 & n2945 ;
  assign n2947 = ( n2765 & n2767 ) | ( n2765 & n2946 ) | ( n2767 & n2946 ) ;
  assign n2948 = ( n2765 & n2767 ) | ( n2765 & ~n2946 ) | ( n2767 & ~n2946 ) ;
  assign n2949 = n2947 & ~n2948 ;
  assign n2950 = ( ~n2761 & n2763 ) | ( ~n2761 & n2768 ) | ( n2763 & n2768 ) ;
  assign n2951 = ( n2761 & ~n2769 ) | ( n2761 & n2950 ) | ( ~n2769 & n2950 ) ;
  assign n2952 = ( ~n2924 & n2926 ) | ( ~n2924 & n2928 ) | ( n2926 & n2928 ) ;
  assign n2953 = ( n2924 & ~n2929 ) | ( n2924 & n2952 ) | ( ~n2929 & n2952 ) ;
  assign n2954 = ( n2949 & n2951 ) | ( n2949 & n2953 ) | ( n2951 & n2953 ) ;
  assign n2955 = ( n2942 & n2944 ) | ( n2942 & n2954 ) | ( n2944 & n2954 ) ;
  assign n2956 = ( n2938 & n2940 ) | ( n2938 & n2955 ) | ( n2940 & n2955 ) ;
  assign n2957 = ( n2934 & n2936 ) | ( n2934 & n2956 ) | ( n2936 & n2956 ) ;
  assign n2958 = ( n2775 & n2932 ) | ( n2775 & n2957 ) | ( n2932 & n2957 ) ;
  assign n2959 = ( x940 & x941 ) | ( x940 & x942 ) | ( x941 & x942 ) ;
  assign n2960 = ( x937 & x938 ) | ( x937 & x939 ) | ( x938 & x939 ) ;
  assign n2961 = ( ~x940 & x941 ) | ( ~x940 & x942 ) | ( x941 & x942 ) ;
  assign n2962 = ( x940 & ~n2959 ) | ( x940 & n2961 ) | ( ~n2959 & n2961 ) ;
  assign n2963 = ( ~x937 & x938 ) | ( ~x937 & x939 ) | ( x938 & x939 ) ;
  assign n2964 = ( x937 & ~n2960 ) | ( x937 & n2963 ) | ( ~n2960 & n2963 ) ;
  assign n2965 = n2962 & n2964 ;
  assign n2966 = ( n2959 & n2960 ) | ( n2959 & n2965 ) | ( n2960 & n2965 ) ;
  assign n2967 = ( x931 & x932 ) | ( x931 & x933 ) | ( x932 & x933 ) ;
  assign n2968 = ( x934 & x935 ) | ( x934 & x936 ) | ( x935 & x936 ) ;
  assign n2969 = ( ~x934 & x935 ) | ( ~x934 & x936 ) | ( x935 & x936 ) ;
  assign n2970 = ( x934 & ~n2968 ) | ( x934 & n2969 ) | ( ~n2968 & n2969 ) ;
  assign n2971 = ( ~x931 & x932 ) | ( ~x931 & x933 ) | ( x932 & x933 ) ;
  assign n2972 = ( x931 & ~n2967 ) | ( x931 & n2971 ) | ( ~n2967 & n2971 ) ;
  assign n2973 = n2970 & n2972 ;
  assign n2974 = ( n2967 & n2968 ) | ( n2967 & n2973 ) | ( n2968 & n2973 ) ;
  assign n2975 = ( ~n2959 & n2960 ) | ( ~n2959 & n2965 ) | ( n2960 & n2965 ) ;
  assign n2976 = ( n2959 & ~n2966 ) | ( n2959 & n2975 ) | ( ~n2966 & n2975 ) ;
  assign n2977 = ( ~n2967 & n2968 ) | ( ~n2967 & n2973 ) | ( n2968 & n2973 ) ;
  assign n2978 = ( n2967 & ~n2974 ) | ( n2967 & n2977 ) | ( ~n2974 & n2977 ) ;
  assign n2979 = n2962 | n2964 ;
  assign n2980 = ~n2965 & n2979 ;
  assign n2981 = n2970 | n2972 ;
  assign n2982 = ~n2973 & n2981 ;
  assign n2983 = n2980 & n2982 ;
  assign n2984 = ( n2976 & n2978 ) | ( n2976 & n2983 ) | ( n2978 & n2983 ) ;
  assign n2985 = ( n2966 & n2974 ) | ( n2966 & n2984 ) | ( n2974 & n2984 ) ;
  assign n2986 = ( x928 & x929 ) | ( x928 & x930 ) | ( x929 & x930 ) ;
  assign n2987 = ( x925 & x926 ) | ( x925 & x927 ) | ( x926 & x927 ) ;
  assign n2988 = ( ~x928 & x929 ) | ( ~x928 & x930 ) | ( x929 & x930 ) ;
  assign n2989 = ( x928 & ~n2986 ) | ( x928 & n2988 ) | ( ~n2986 & n2988 ) ;
  assign n2990 = ( ~x925 & x926 ) | ( ~x925 & x927 ) | ( x926 & x927 ) ;
  assign n2991 = ( x925 & ~n2987 ) | ( x925 & n2990 ) | ( ~n2987 & n2990 ) ;
  assign n2992 = n2989 & n2991 ;
  assign n2993 = ( n2986 & n2987 ) | ( n2986 & n2992 ) | ( n2987 & n2992 ) ;
  assign n2994 = ( x919 & x920 ) | ( x919 & x921 ) | ( x920 & x921 ) ;
  assign n2995 = ( x922 & x923 ) | ( x922 & x924 ) | ( x923 & x924 ) ;
  assign n2996 = ( ~x922 & x923 ) | ( ~x922 & x924 ) | ( x923 & x924 ) ;
  assign n2997 = ( x922 & ~n2995 ) | ( x922 & n2996 ) | ( ~n2995 & n2996 ) ;
  assign n2998 = ( ~x919 & x920 ) | ( ~x919 & x921 ) | ( x920 & x921 ) ;
  assign n2999 = ( x919 & ~n2994 ) | ( x919 & n2998 ) | ( ~n2994 & n2998 ) ;
  assign n3000 = n2997 & n2999 ;
  assign n3001 = ( n2994 & n2995 ) | ( n2994 & n3000 ) | ( n2995 & n3000 ) ;
  assign n3002 = ( ~n2986 & n2987 ) | ( ~n2986 & n2992 ) | ( n2987 & n2992 ) ;
  assign n3003 = ( n2986 & ~n2993 ) | ( n2986 & n3002 ) | ( ~n2993 & n3002 ) ;
  assign n3004 = ( ~n2994 & n2995 ) | ( ~n2994 & n3000 ) | ( n2995 & n3000 ) ;
  assign n3005 = ( n2994 & ~n3001 ) | ( n2994 & n3004 ) | ( ~n3001 & n3004 ) ;
  assign n3006 = n2997 | n2999 ;
  assign n3007 = ~n3000 & n3006 ;
  assign n3008 = ( n2989 & n2991 ) | ( n2989 & n3007 ) | ( n2991 & n3007 ) ;
  assign n3009 = ~n2992 & n3008 ;
  assign n3010 = ( n3003 & n3005 ) | ( n3003 & n3009 ) | ( n3005 & n3009 ) ;
  assign n3011 = ( n2993 & n3001 ) | ( n2993 & n3010 ) | ( n3001 & n3010 ) ;
  assign n3012 = ( ~n2993 & n3001 ) | ( ~n2993 & n3010 ) | ( n3001 & n3010 ) ;
  assign n3013 = ( n2993 & ~n3011 ) | ( n2993 & n3012 ) | ( ~n3011 & n3012 ) ;
  assign n3014 = ( ~n2966 & n2974 ) | ( ~n2966 & n2984 ) | ( n2974 & n2984 ) ;
  assign n3015 = ( n2966 & ~n2985 ) | ( n2966 & n3014 ) | ( ~n2985 & n3014 ) ;
  assign n3016 = ( ~n2976 & n2978 ) | ( ~n2976 & n2983 ) | ( n2978 & n2983 ) ;
  assign n3017 = ( n2976 & ~n2984 ) | ( n2976 & n3016 ) | ( ~n2984 & n3016 ) ;
  assign n3018 = ( ~n3003 & n3005 ) | ( ~n3003 & n3009 ) | ( n3005 & n3009 ) ;
  assign n3019 = ( n3003 & ~n3010 ) | ( n3003 & n3018 ) | ( ~n3010 & n3018 ) ;
  assign n3020 = ( ~n2989 & n2991 ) | ( ~n2989 & n3007 ) | ( n2991 & n3007 ) ;
  assign n3021 = ( n2989 & ~n3008 ) | ( n2989 & n3020 ) | ( ~n3008 & n3020 ) ;
  assign n3022 = ( n2980 & n2982 ) | ( n2980 & n3021 ) | ( n2982 & n3021 ) ;
  assign n3023 = ~n2983 & n3022 ;
  assign n3024 = ( n3017 & n3019 ) | ( n3017 & n3023 ) | ( n3019 & n3023 ) ;
  assign n3025 = ( n3013 & n3015 ) | ( n3013 & n3024 ) | ( n3015 & n3024 ) ;
  assign n3026 = ( n2985 & n3011 ) | ( n2985 & n3025 ) | ( n3011 & n3025 ) ;
  assign n3027 = ( x916 & x917 ) | ( x916 & x918 ) | ( x917 & x918 ) ;
  assign n3028 = ( x913 & x914 ) | ( x913 & x915 ) | ( x914 & x915 ) ;
  assign n3029 = ( ~x916 & x917 ) | ( ~x916 & x918 ) | ( x917 & x918 ) ;
  assign n3030 = ( x916 & ~n3027 ) | ( x916 & n3029 ) | ( ~n3027 & n3029 ) ;
  assign n3031 = ( ~x913 & x914 ) | ( ~x913 & x915 ) | ( x914 & x915 ) ;
  assign n3032 = ( x913 & ~n3028 ) | ( x913 & n3031 ) | ( ~n3028 & n3031 ) ;
  assign n3033 = n3030 & n3032 ;
  assign n3034 = ( n3027 & n3028 ) | ( n3027 & n3033 ) | ( n3028 & n3033 ) ;
  assign n3035 = ( x907 & x908 ) | ( x907 & x909 ) | ( x908 & x909 ) ;
  assign n3036 = ( x910 & x911 ) | ( x910 & x912 ) | ( x911 & x912 ) ;
  assign n3037 = ( ~x910 & x911 ) | ( ~x910 & x912 ) | ( x911 & x912 ) ;
  assign n3038 = ( x910 & ~n3036 ) | ( x910 & n3037 ) | ( ~n3036 & n3037 ) ;
  assign n3039 = ( ~x907 & x908 ) | ( ~x907 & x909 ) | ( x908 & x909 ) ;
  assign n3040 = ( x907 & ~n3035 ) | ( x907 & n3039 ) | ( ~n3035 & n3039 ) ;
  assign n3041 = n3038 & n3040 ;
  assign n3042 = ( n3035 & n3036 ) | ( n3035 & n3041 ) | ( n3036 & n3041 ) ;
  assign n3043 = ( ~n3027 & n3028 ) | ( ~n3027 & n3033 ) | ( n3028 & n3033 ) ;
  assign n3044 = ( n3027 & ~n3034 ) | ( n3027 & n3043 ) | ( ~n3034 & n3043 ) ;
  assign n3045 = ( ~n3035 & n3036 ) | ( ~n3035 & n3041 ) | ( n3036 & n3041 ) ;
  assign n3046 = ( n3035 & ~n3042 ) | ( n3035 & n3045 ) | ( ~n3042 & n3045 ) ;
  assign n3047 = n3030 | n3032 ;
  assign n3048 = ~n3033 & n3047 ;
  assign n3049 = n3038 | n3040 ;
  assign n3050 = ~n3041 & n3049 ;
  assign n3051 = n3048 & n3050 ;
  assign n3052 = ( n3044 & n3046 ) | ( n3044 & n3051 ) | ( n3046 & n3051 ) ;
  assign n3053 = ( n3034 & n3042 ) | ( n3034 & n3052 ) | ( n3042 & n3052 ) ;
  assign n3054 = ( x904 & x905 ) | ( x904 & x906 ) | ( x905 & x906 ) ;
  assign n3055 = ( x901 & x902 ) | ( x901 & x903 ) | ( x902 & x903 ) ;
  assign n3056 = ( ~x904 & x905 ) | ( ~x904 & x906 ) | ( x905 & x906 ) ;
  assign n3057 = ( x904 & ~n3054 ) | ( x904 & n3056 ) | ( ~n3054 & n3056 ) ;
  assign n3058 = ( ~x901 & x902 ) | ( ~x901 & x903 ) | ( x902 & x903 ) ;
  assign n3059 = ( x901 & ~n3055 ) | ( x901 & n3058 ) | ( ~n3055 & n3058 ) ;
  assign n3060 = n3057 & n3059 ;
  assign n3061 = ( n3054 & n3055 ) | ( n3054 & n3060 ) | ( n3055 & n3060 ) ;
  assign n3062 = ( x895 & x896 ) | ( x895 & x897 ) | ( x896 & x897 ) ;
  assign n3063 = ( x898 & x899 ) | ( x898 & x900 ) | ( x899 & x900 ) ;
  assign n3064 = ( ~x898 & x899 ) | ( ~x898 & x900 ) | ( x899 & x900 ) ;
  assign n3065 = ( x898 & ~n3063 ) | ( x898 & n3064 ) | ( ~n3063 & n3064 ) ;
  assign n3066 = ( ~x895 & x896 ) | ( ~x895 & x897 ) | ( x896 & x897 ) ;
  assign n3067 = ( x895 & ~n3062 ) | ( x895 & n3066 ) | ( ~n3062 & n3066 ) ;
  assign n3068 = n3065 & n3067 ;
  assign n3069 = ( n3062 & n3063 ) | ( n3062 & n3068 ) | ( n3063 & n3068 ) ;
  assign n3070 = ( ~n3054 & n3055 ) | ( ~n3054 & n3060 ) | ( n3055 & n3060 ) ;
  assign n3071 = ( n3054 & ~n3061 ) | ( n3054 & n3070 ) | ( ~n3061 & n3070 ) ;
  assign n3072 = ( ~n3062 & n3063 ) | ( ~n3062 & n3068 ) | ( n3063 & n3068 ) ;
  assign n3073 = ( n3062 & ~n3069 ) | ( n3062 & n3072 ) | ( ~n3069 & n3072 ) ;
  assign n3074 = n3065 | n3067 ;
  assign n3075 = ~n3068 & n3074 ;
  assign n3076 = ( n3057 & n3059 ) | ( n3057 & n3075 ) | ( n3059 & n3075 ) ;
  assign n3077 = ~n3060 & n3076 ;
  assign n3078 = ( n3071 & n3073 ) | ( n3071 & n3077 ) | ( n3073 & n3077 ) ;
  assign n3079 = ( n3061 & n3069 ) | ( n3061 & n3078 ) | ( n3069 & n3078 ) ;
  assign n3080 = ( ~n3061 & n3069 ) | ( ~n3061 & n3078 ) | ( n3069 & n3078 ) ;
  assign n3081 = ( n3061 & ~n3079 ) | ( n3061 & n3080 ) | ( ~n3079 & n3080 ) ;
  assign n3082 = ( ~n3034 & n3042 ) | ( ~n3034 & n3052 ) | ( n3042 & n3052 ) ;
  assign n3083 = ( n3034 & ~n3053 ) | ( n3034 & n3082 ) | ( ~n3053 & n3082 ) ;
  assign n3084 = ( ~n3044 & n3046 ) | ( ~n3044 & n3051 ) | ( n3046 & n3051 ) ;
  assign n3085 = ( n3044 & ~n3052 ) | ( n3044 & n3084 ) | ( ~n3052 & n3084 ) ;
  assign n3086 = ( ~n3071 & n3073 ) | ( ~n3071 & n3077 ) | ( n3073 & n3077 ) ;
  assign n3087 = ( n3071 & ~n3078 ) | ( n3071 & n3086 ) | ( ~n3078 & n3086 ) ;
  assign n3088 = ( ~n3057 & n3059 ) | ( ~n3057 & n3075 ) | ( n3059 & n3075 ) ;
  assign n3089 = ( n3057 & ~n3076 ) | ( n3057 & n3088 ) | ( ~n3076 & n3088 ) ;
  assign n3090 = ( n3048 & n3050 ) | ( n3048 & n3089 ) | ( n3050 & n3089 ) ;
  assign n3091 = ~n3051 & n3090 ;
  assign n3092 = ( n3085 & n3087 ) | ( n3085 & n3091 ) | ( n3087 & n3091 ) ;
  assign n3093 = ( n3081 & n3083 ) | ( n3081 & n3092 ) | ( n3083 & n3092 ) ;
  assign n3094 = ( n3053 & n3079 ) | ( n3053 & n3093 ) | ( n3079 & n3093 ) ;
  assign n3095 = ( ~n2985 & n3011 ) | ( ~n2985 & n3025 ) | ( n3011 & n3025 ) ;
  assign n3096 = ( n2985 & ~n3026 ) | ( n2985 & n3095 ) | ( ~n3026 & n3095 ) ;
  assign n3097 = ( ~n3053 & n3079 ) | ( ~n3053 & n3093 ) | ( n3079 & n3093 ) ;
  assign n3098 = ( n3053 & ~n3094 ) | ( n3053 & n3097 ) | ( ~n3094 & n3097 ) ;
  assign n3099 = ( ~n3081 & n3083 ) | ( ~n3081 & n3092 ) | ( n3083 & n3092 ) ;
  assign n3100 = ( n3081 & ~n3093 ) | ( n3081 & n3099 ) | ( ~n3093 & n3099 ) ;
  assign n3101 = ( ~n3013 & n3015 ) | ( ~n3013 & n3024 ) | ( n3015 & n3024 ) ;
  assign n3102 = ( n3013 & ~n3025 ) | ( n3013 & n3101 ) | ( ~n3025 & n3101 ) ;
  assign n3103 = ( n3017 & n3019 ) | ( n3017 & ~n3023 ) | ( n3019 & ~n3023 ) ;
  assign n3104 = ( n3023 & ~n3024 ) | ( n3023 & n3103 ) | ( ~n3024 & n3103 ) ;
  assign n3105 = ( n3085 & n3087 ) | ( n3085 & ~n3091 ) | ( n3087 & ~n3091 ) ;
  assign n3106 = ( n3091 & ~n3092 ) | ( n3091 & n3105 ) | ( ~n3092 & n3105 ) ;
  assign n3107 = ( ~n2980 & n2982 ) | ( ~n2980 & n3021 ) | ( n2982 & n3021 ) ;
  assign n3108 = ( n2980 & ~n3022 ) | ( n2980 & n3107 ) | ( ~n3022 & n3107 ) ;
  assign n3109 = ( ~n3048 & n3050 ) | ( ~n3048 & n3089 ) | ( n3050 & n3089 ) ;
  assign n3110 = ( n3048 & ~n3090 ) | ( n3048 & n3109 ) | ( ~n3090 & n3109 ) ;
  assign n3111 = n3108 & n3110 ;
  assign n3112 = ( n3104 & n3106 ) | ( n3104 & n3111 ) | ( n3106 & n3111 ) ;
  assign n3113 = ( n3100 & n3102 ) | ( n3100 & n3112 ) | ( n3102 & n3112 ) ;
  assign n3114 = ( n3096 & n3098 ) | ( n3096 & n3113 ) | ( n3098 & n3113 ) ;
  assign n3115 = ( n3026 & n3094 ) | ( n3026 & n3114 ) | ( n3094 & n3114 ) ;
  assign n3116 = ( x892 & x893 ) | ( x892 & x894 ) | ( x893 & x894 ) ;
  assign n3117 = ( x889 & x890 ) | ( x889 & x891 ) | ( x890 & x891 ) ;
  assign n3118 = ( ~x892 & x893 ) | ( ~x892 & x894 ) | ( x893 & x894 ) ;
  assign n3119 = ( x892 & ~n3116 ) | ( x892 & n3118 ) | ( ~n3116 & n3118 ) ;
  assign n3120 = ( ~x889 & x890 ) | ( ~x889 & x891 ) | ( x890 & x891 ) ;
  assign n3121 = ( x889 & ~n3117 ) | ( x889 & n3120 ) | ( ~n3117 & n3120 ) ;
  assign n3122 = n3119 & n3121 ;
  assign n3123 = ( n3116 & n3117 ) | ( n3116 & n3122 ) | ( n3117 & n3122 ) ;
  assign n3124 = ( x883 & x884 ) | ( x883 & x885 ) | ( x884 & x885 ) ;
  assign n3125 = ( x886 & x887 ) | ( x886 & x888 ) | ( x887 & x888 ) ;
  assign n3126 = ( ~x886 & x887 ) | ( ~x886 & x888 ) | ( x887 & x888 ) ;
  assign n3127 = ( x886 & ~n3125 ) | ( x886 & n3126 ) | ( ~n3125 & n3126 ) ;
  assign n3128 = ( ~x883 & x884 ) | ( ~x883 & x885 ) | ( x884 & x885 ) ;
  assign n3129 = ( x883 & ~n3124 ) | ( x883 & n3128 ) | ( ~n3124 & n3128 ) ;
  assign n3130 = n3127 & n3129 ;
  assign n3131 = ( n3124 & n3125 ) | ( n3124 & n3130 ) | ( n3125 & n3130 ) ;
  assign n3132 = ( ~n3116 & n3117 ) | ( ~n3116 & n3122 ) | ( n3117 & n3122 ) ;
  assign n3133 = ( n3116 & ~n3123 ) | ( n3116 & n3132 ) | ( ~n3123 & n3132 ) ;
  assign n3134 = ( ~n3124 & n3125 ) | ( ~n3124 & n3130 ) | ( n3125 & n3130 ) ;
  assign n3135 = ( n3124 & ~n3131 ) | ( n3124 & n3134 ) | ( ~n3131 & n3134 ) ;
  assign n3136 = n3119 | n3121 ;
  assign n3137 = ~n3122 & n3136 ;
  assign n3138 = n3127 | n3129 ;
  assign n3139 = ~n3130 & n3138 ;
  assign n3140 = n3137 & n3139 ;
  assign n3141 = ( n3133 & n3135 ) | ( n3133 & n3140 ) | ( n3135 & n3140 ) ;
  assign n3142 = ( n3123 & n3131 ) | ( n3123 & n3141 ) | ( n3131 & n3141 ) ;
  assign n3143 = ( x880 & x881 ) | ( x880 & x882 ) | ( x881 & x882 ) ;
  assign n3144 = ( x877 & x878 ) | ( x877 & x879 ) | ( x878 & x879 ) ;
  assign n3145 = ( ~x880 & x881 ) | ( ~x880 & x882 ) | ( x881 & x882 ) ;
  assign n3146 = ( x880 & ~n3143 ) | ( x880 & n3145 ) | ( ~n3143 & n3145 ) ;
  assign n3147 = ( ~x877 & x878 ) | ( ~x877 & x879 ) | ( x878 & x879 ) ;
  assign n3148 = ( x877 & ~n3144 ) | ( x877 & n3147 ) | ( ~n3144 & n3147 ) ;
  assign n3149 = n3146 & n3148 ;
  assign n3150 = ( n3143 & n3144 ) | ( n3143 & n3149 ) | ( n3144 & n3149 ) ;
  assign n3151 = ( x871 & x872 ) | ( x871 & x873 ) | ( x872 & x873 ) ;
  assign n3152 = ( x874 & x875 ) | ( x874 & x876 ) | ( x875 & x876 ) ;
  assign n3153 = ( ~x874 & x875 ) | ( ~x874 & x876 ) | ( x875 & x876 ) ;
  assign n3154 = ( x874 & ~n3152 ) | ( x874 & n3153 ) | ( ~n3152 & n3153 ) ;
  assign n3155 = ( ~x871 & x872 ) | ( ~x871 & x873 ) | ( x872 & x873 ) ;
  assign n3156 = ( x871 & ~n3151 ) | ( x871 & n3155 ) | ( ~n3151 & n3155 ) ;
  assign n3157 = n3154 & n3156 ;
  assign n3158 = ( n3151 & n3152 ) | ( n3151 & n3157 ) | ( n3152 & n3157 ) ;
  assign n3159 = ( ~n3143 & n3144 ) | ( ~n3143 & n3149 ) | ( n3144 & n3149 ) ;
  assign n3160 = ( n3143 & ~n3150 ) | ( n3143 & n3159 ) | ( ~n3150 & n3159 ) ;
  assign n3161 = ( ~n3151 & n3152 ) | ( ~n3151 & n3157 ) | ( n3152 & n3157 ) ;
  assign n3162 = ( n3151 & ~n3158 ) | ( n3151 & n3161 ) | ( ~n3158 & n3161 ) ;
  assign n3163 = n3154 | n3156 ;
  assign n3164 = ~n3157 & n3163 ;
  assign n3165 = ( n3146 & n3148 ) | ( n3146 & n3164 ) | ( n3148 & n3164 ) ;
  assign n3166 = ~n3149 & n3165 ;
  assign n3167 = ( n3160 & n3162 ) | ( n3160 & n3166 ) | ( n3162 & n3166 ) ;
  assign n3168 = ( n3150 & n3158 ) | ( n3150 & n3167 ) | ( n3158 & n3167 ) ;
  assign n3169 = ( ~n3150 & n3158 ) | ( ~n3150 & n3167 ) | ( n3158 & n3167 ) ;
  assign n3170 = ( n3150 & ~n3168 ) | ( n3150 & n3169 ) | ( ~n3168 & n3169 ) ;
  assign n3171 = ( ~n3123 & n3131 ) | ( ~n3123 & n3141 ) | ( n3131 & n3141 ) ;
  assign n3172 = ( n3123 & ~n3142 ) | ( n3123 & n3171 ) | ( ~n3142 & n3171 ) ;
  assign n3173 = ( ~n3133 & n3135 ) | ( ~n3133 & n3140 ) | ( n3135 & n3140 ) ;
  assign n3174 = ( n3133 & ~n3141 ) | ( n3133 & n3173 ) | ( ~n3141 & n3173 ) ;
  assign n3175 = ( ~n3160 & n3162 ) | ( ~n3160 & n3166 ) | ( n3162 & n3166 ) ;
  assign n3176 = ( n3160 & ~n3167 ) | ( n3160 & n3175 ) | ( ~n3167 & n3175 ) ;
  assign n3177 = ( ~n3146 & n3148 ) | ( ~n3146 & n3164 ) | ( n3148 & n3164 ) ;
  assign n3178 = ( n3146 & ~n3165 ) | ( n3146 & n3177 ) | ( ~n3165 & n3177 ) ;
  assign n3179 = ( n3137 & n3139 ) | ( n3137 & n3178 ) | ( n3139 & n3178 ) ;
  assign n3180 = ~n3140 & n3179 ;
  assign n3181 = ( n3174 & n3176 ) | ( n3174 & n3180 ) | ( n3176 & n3180 ) ;
  assign n3182 = ( n3170 & n3172 ) | ( n3170 & n3181 ) | ( n3172 & n3181 ) ;
  assign n3183 = ( n3142 & n3168 ) | ( n3142 & n3182 ) | ( n3168 & n3182 ) ;
  assign n3184 = ( x868 & x869 ) | ( x868 & x870 ) | ( x869 & x870 ) ;
  assign n3185 = ( x865 & x866 ) | ( x865 & x867 ) | ( x866 & x867 ) ;
  assign n3186 = ( ~x868 & x869 ) | ( ~x868 & x870 ) | ( x869 & x870 ) ;
  assign n3187 = ( x868 & ~n3184 ) | ( x868 & n3186 ) | ( ~n3184 & n3186 ) ;
  assign n3188 = ( ~x865 & x866 ) | ( ~x865 & x867 ) | ( x866 & x867 ) ;
  assign n3189 = ( x865 & ~n3185 ) | ( x865 & n3188 ) | ( ~n3185 & n3188 ) ;
  assign n3190 = n3187 & n3189 ;
  assign n3191 = ( n3184 & n3185 ) | ( n3184 & n3190 ) | ( n3185 & n3190 ) ;
  assign n3192 = ( x859 & x860 ) | ( x859 & x861 ) | ( x860 & x861 ) ;
  assign n3193 = ( x862 & x863 ) | ( x862 & x864 ) | ( x863 & x864 ) ;
  assign n3194 = ( ~x862 & x863 ) | ( ~x862 & x864 ) | ( x863 & x864 ) ;
  assign n3195 = ( x862 & ~n3193 ) | ( x862 & n3194 ) | ( ~n3193 & n3194 ) ;
  assign n3196 = ( ~x859 & x860 ) | ( ~x859 & x861 ) | ( x860 & x861 ) ;
  assign n3197 = ( x859 & ~n3192 ) | ( x859 & n3196 ) | ( ~n3192 & n3196 ) ;
  assign n3198 = n3195 & n3197 ;
  assign n3199 = ( n3192 & n3193 ) | ( n3192 & n3198 ) | ( n3193 & n3198 ) ;
  assign n3200 = ( ~n3184 & n3185 ) | ( ~n3184 & n3190 ) | ( n3185 & n3190 ) ;
  assign n3201 = ( n3184 & ~n3191 ) | ( n3184 & n3200 ) | ( ~n3191 & n3200 ) ;
  assign n3202 = ( ~n3192 & n3193 ) | ( ~n3192 & n3198 ) | ( n3193 & n3198 ) ;
  assign n3203 = ( n3192 & ~n3199 ) | ( n3192 & n3202 ) | ( ~n3199 & n3202 ) ;
  assign n3204 = n3187 | n3189 ;
  assign n3205 = ~n3190 & n3204 ;
  assign n3206 = n3195 | n3197 ;
  assign n3207 = ~n3198 & n3206 ;
  assign n3208 = n3205 & n3207 ;
  assign n3209 = ( n3201 & n3203 ) | ( n3201 & n3208 ) | ( n3203 & n3208 ) ;
  assign n3210 = ( n3191 & n3199 ) | ( n3191 & n3209 ) | ( n3199 & n3209 ) ;
  assign n3211 = ( x856 & x857 ) | ( x856 & x858 ) | ( x857 & x858 ) ;
  assign n3212 = ( x853 & x854 ) | ( x853 & x855 ) | ( x854 & x855 ) ;
  assign n3213 = ( ~x856 & x857 ) | ( ~x856 & x858 ) | ( x857 & x858 ) ;
  assign n3214 = ( x856 & ~n3211 ) | ( x856 & n3213 ) | ( ~n3211 & n3213 ) ;
  assign n3215 = ( ~x853 & x854 ) | ( ~x853 & x855 ) | ( x854 & x855 ) ;
  assign n3216 = ( x853 & ~n3212 ) | ( x853 & n3215 ) | ( ~n3212 & n3215 ) ;
  assign n3217 = n3214 & n3216 ;
  assign n3218 = ( n3211 & n3212 ) | ( n3211 & n3217 ) | ( n3212 & n3217 ) ;
  assign n3219 = ( x847 & x848 ) | ( x847 & x849 ) | ( x848 & x849 ) ;
  assign n3220 = ( x850 & x851 ) | ( x850 & x852 ) | ( x851 & x852 ) ;
  assign n3221 = ( ~x850 & x851 ) | ( ~x850 & x852 ) | ( x851 & x852 ) ;
  assign n3222 = ( x850 & ~n3220 ) | ( x850 & n3221 ) | ( ~n3220 & n3221 ) ;
  assign n3223 = ( ~x847 & x848 ) | ( ~x847 & x849 ) | ( x848 & x849 ) ;
  assign n3224 = ( x847 & ~n3219 ) | ( x847 & n3223 ) | ( ~n3219 & n3223 ) ;
  assign n3225 = n3222 & n3224 ;
  assign n3226 = ( n3219 & n3220 ) | ( n3219 & n3225 ) | ( n3220 & n3225 ) ;
  assign n3227 = ( ~n3211 & n3212 ) | ( ~n3211 & n3217 ) | ( n3212 & n3217 ) ;
  assign n3228 = ( n3211 & ~n3218 ) | ( n3211 & n3227 ) | ( ~n3218 & n3227 ) ;
  assign n3229 = ( ~n3219 & n3220 ) | ( ~n3219 & n3225 ) | ( n3220 & n3225 ) ;
  assign n3230 = ( n3219 & ~n3226 ) | ( n3219 & n3229 ) | ( ~n3226 & n3229 ) ;
  assign n3231 = n3222 | n3224 ;
  assign n3232 = ~n3225 & n3231 ;
  assign n3233 = ( n3214 & n3216 ) | ( n3214 & n3232 ) | ( n3216 & n3232 ) ;
  assign n3234 = ~n3217 & n3233 ;
  assign n3235 = ( n3228 & n3230 ) | ( n3228 & n3234 ) | ( n3230 & n3234 ) ;
  assign n3236 = ( n3218 & n3226 ) | ( n3218 & n3235 ) | ( n3226 & n3235 ) ;
  assign n3237 = ( ~n3218 & n3226 ) | ( ~n3218 & n3235 ) | ( n3226 & n3235 ) ;
  assign n3238 = ( n3218 & ~n3236 ) | ( n3218 & n3237 ) | ( ~n3236 & n3237 ) ;
  assign n3239 = ( ~n3191 & n3199 ) | ( ~n3191 & n3209 ) | ( n3199 & n3209 ) ;
  assign n3240 = ( n3191 & ~n3210 ) | ( n3191 & n3239 ) | ( ~n3210 & n3239 ) ;
  assign n3241 = ( ~n3201 & n3203 ) | ( ~n3201 & n3208 ) | ( n3203 & n3208 ) ;
  assign n3242 = ( n3201 & ~n3209 ) | ( n3201 & n3241 ) | ( ~n3209 & n3241 ) ;
  assign n3243 = ( ~n3228 & n3230 ) | ( ~n3228 & n3234 ) | ( n3230 & n3234 ) ;
  assign n3244 = ( n3228 & ~n3235 ) | ( n3228 & n3243 ) | ( ~n3235 & n3243 ) ;
  assign n3245 = ( ~n3214 & n3216 ) | ( ~n3214 & n3232 ) | ( n3216 & n3232 ) ;
  assign n3246 = ( n3214 & ~n3233 ) | ( n3214 & n3245 ) | ( ~n3233 & n3245 ) ;
  assign n3247 = ( n3205 & n3207 ) | ( n3205 & n3246 ) | ( n3207 & n3246 ) ;
  assign n3248 = ~n3208 & n3247 ;
  assign n3249 = ( n3242 & n3244 ) | ( n3242 & n3248 ) | ( n3244 & n3248 ) ;
  assign n3250 = ( n3238 & n3240 ) | ( n3238 & n3249 ) | ( n3240 & n3249 ) ;
  assign n3251 = ( n3210 & n3236 ) | ( n3210 & n3250 ) | ( n3236 & n3250 ) ;
  assign n3252 = ( ~n3142 & n3168 ) | ( ~n3142 & n3182 ) | ( n3168 & n3182 ) ;
  assign n3253 = ( n3142 & ~n3183 ) | ( n3142 & n3252 ) | ( ~n3183 & n3252 ) ;
  assign n3254 = ( ~n3210 & n3236 ) | ( ~n3210 & n3250 ) | ( n3236 & n3250 ) ;
  assign n3255 = ( n3210 & ~n3251 ) | ( n3210 & n3254 ) | ( ~n3251 & n3254 ) ;
  assign n3256 = ( ~n3238 & n3240 ) | ( ~n3238 & n3249 ) | ( n3240 & n3249 ) ;
  assign n3257 = ( n3238 & ~n3250 ) | ( n3238 & n3256 ) | ( ~n3250 & n3256 ) ;
  assign n3258 = ( ~n3170 & n3172 ) | ( ~n3170 & n3181 ) | ( n3172 & n3181 ) ;
  assign n3259 = ( n3170 & ~n3182 ) | ( n3170 & n3258 ) | ( ~n3182 & n3258 ) ;
  assign n3260 = ( n3174 & n3176 ) | ( n3174 & ~n3180 ) | ( n3176 & ~n3180 ) ;
  assign n3261 = ( n3180 & ~n3181 ) | ( n3180 & n3260 ) | ( ~n3181 & n3260 ) ;
  assign n3262 = ( n3242 & n3244 ) | ( n3242 & ~n3248 ) | ( n3244 & ~n3248 ) ;
  assign n3263 = ( n3248 & ~n3249 ) | ( n3248 & n3262 ) | ( ~n3249 & n3262 ) ;
  assign n3264 = ( ~n3137 & n3139 ) | ( ~n3137 & n3178 ) | ( n3139 & n3178 ) ;
  assign n3265 = ( n3137 & ~n3179 ) | ( n3137 & n3264 ) | ( ~n3179 & n3264 ) ;
  assign n3266 = ( ~n3205 & n3207 ) | ( ~n3205 & n3246 ) | ( n3207 & n3246 ) ;
  assign n3267 = ( n3205 & ~n3247 ) | ( n3205 & n3266 ) | ( ~n3247 & n3266 ) ;
  assign n3268 = n3265 & n3267 ;
  assign n3269 = ( n3261 & n3263 ) | ( n3261 & n3268 ) | ( n3263 & n3268 ) ;
  assign n3270 = ( n3257 & n3259 ) | ( n3257 & n3269 ) | ( n3259 & n3269 ) ;
  assign n3271 = ( n3253 & n3255 ) | ( n3253 & n3270 ) | ( n3255 & n3270 ) ;
  assign n3272 = ( n3183 & n3251 ) | ( n3183 & n3271 ) | ( n3251 & n3271 ) ;
  assign n3273 = ( ~n3183 & n3251 ) | ( ~n3183 & n3271 ) | ( n3251 & n3271 ) ;
  assign n3274 = ( n3183 & ~n3272 ) | ( n3183 & n3273 ) | ( ~n3272 & n3273 ) ;
  assign n3275 = ( ~n3026 & n3094 ) | ( ~n3026 & n3114 ) | ( n3094 & n3114 ) ;
  assign n3276 = ( n3026 & ~n3115 ) | ( n3026 & n3275 ) | ( ~n3115 & n3275 ) ;
  assign n3277 = ( ~n3096 & n3098 ) | ( ~n3096 & n3113 ) | ( n3098 & n3113 ) ;
  assign n3278 = ( n3096 & ~n3114 ) | ( n3096 & n3277 ) | ( ~n3114 & n3277 ) ;
  assign n3279 = ( ~n3253 & n3255 ) | ( ~n3253 & n3270 ) | ( n3255 & n3270 ) ;
  assign n3280 = ( n3253 & ~n3271 ) | ( n3253 & n3279 ) | ( ~n3271 & n3279 ) ;
  assign n3281 = ( ~n3257 & n3259 ) | ( ~n3257 & n3269 ) | ( n3259 & n3269 ) ;
  assign n3282 = ( n3257 & ~n3270 ) | ( n3257 & n3281 ) | ( ~n3270 & n3281 ) ;
  assign n3283 = ( ~n3100 & n3102 ) | ( ~n3100 & n3112 ) | ( n3102 & n3112 ) ;
  assign n3284 = ( n3100 & ~n3113 ) | ( n3100 & n3283 ) | ( ~n3113 & n3283 ) ;
  assign n3285 = ( ~n3104 & n3106 ) | ( ~n3104 & n3111 ) | ( n3106 & n3111 ) ;
  assign n3286 = ( n3104 & ~n3112 ) | ( n3104 & n3285 ) | ( ~n3112 & n3285 ) ;
  assign n3287 = ( ~n3261 & n3263 ) | ( ~n3261 & n3268 ) | ( n3263 & n3268 ) ;
  assign n3288 = ( n3261 & ~n3269 ) | ( n3261 & n3287 ) | ( ~n3269 & n3287 ) ;
  assign n3289 = n3265 | n3267 ;
  assign n3290 = ~n3268 & n3289 ;
  assign n3291 = ( n3108 & n3110 ) | ( n3108 & n3290 ) | ( n3110 & n3290 ) ;
  assign n3292 = ~n3111 & n3291 ;
  assign n3293 = ( n3286 & n3288 ) | ( n3286 & n3292 ) | ( n3288 & n3292 ) ;
  assign n3294 = ( n3282 & n3284 ) | ( n3282 & n3293 ) | ( n3284 & n3293 ) ;
  assign n3295 = ( n3278 & n3280 ) | ( n3278 & n3294 ) | ( n3280 & n3294 ) ;
  assign n3296 = ( n3274 & n3276 ) | ( n3274 & n3295 ) | ( n3276 & n3295 ) ;
  assign n3297 = ( n3115 & n3272 ) | ( n3115 & n3296 ) | ( n3272 & n3296 ) ;
  assign n3298 = n2773 & ~n3297 ;
  assign n3299 = ( n2773 & n2958 ) | ( n2773 & n3298 ) | ( n2958 & n3298 ) ;
  assign n3300 = ( ~n3115 & n3272 ) | ( ~n3115 & n3296 ) | ( n3272 & n3296 ) ;
  assign n3301 = ( n3115 & ~n3297 ) | ( n3115 & n3300 ) | ( ~n3297 & n3300 ) ;
  assign n3302 = ( ~n2775 & n2932 ) | ( ~n2775 & n2957 ) | ( n2932 & n2957 ) ;
  assign n3303 = ( n2775 & ~n2958 ) | ( n2775 & n3302 ) | ( ~n2958 & n3302 ) ;
  assign n3304 = ( ~n3274 & n3276 ) | ( ~n3274 & n3295 ) | ( n3276 & n3295 ) ;
  assign n3305 = ( n3274 & ~n3296 ) | ( n3274 & n3304 ) | ( ~n3296 & n3304 ) ;
  assign n3306 = ( ~n2934 & n2936 ) | ( ~n2934 & n2956 ) | ( n2936 & n2956 ) ;
  assign n3307 = ( n2934 & ~n2957 ) | ( n2934 & n3306 ) | ( ~n2957 & n3306 ) ;
  assign n3308 = ( ~n2938 & n2940 ) | ( ~n2938 & n2955 ) | ( n2940 & n2955 ) ;
  assign n3309 = ( n2938 & ~n2956 ) | ( n2938 & n3308 ) | ( ~n2956 & n3308 ) ;
  assign n3310 = ( ~n3278 & n3280 ) | ( ~n3278 & n3294 ) | ( n3280 & n3294 ) ;
  assign n3311 = ( n3278 & ~n3295 ) | ( n3278 & n3310 ) | ( ~n3295 & n3310 ) ;
  assign n3312 = ( ~n3282 & n3284 ) | ( ~n3282 & n3293 ) | ( n3284 & n3293 ) ;
  assign n3313 = ( n3282 & ~n3294 ) | ( n3282 & n3312 ) | ( ~n3294 & n3312 ) ;
  assign n3314 = ( ~n2942 & n2944 ) | ( ~n2942 & n2954 ) | ( n2944 & n2954 ) ;
  assign n3315 = ( n2942 & ~n2955 ) | ( n2942 & n3314 ) | ( ~n2955 & n3314 ) ;
  assign n3316 = ( ~n3108 & n3110 ) | ( ~n3108 & n3290 ) | ( n3110 & n3290 ) ;
  assign n3317 = ( n3108 & ~n3291 ) | ( n3108 & n3316 ) | ( ~n3291 & n3316 ) ;
  assign n3318 = ( n2946 & ~n2947 ) | ( n2946 & n2948 ) | ( ~n2947 & n2948 ) ;
  assign n3319 = n3317 & n3318 ;
  assign n3320 = ( ~n2949 & n2951 ) | ( ~n2949 & n2953 ) | ( n2951 & n2953 ) ;
  assign n3321 = ( n2949 & ~n2954 ) | ( n2949 & n3320 ) | ( ~n2954 & n3320 ) ;
  assign n3322 = ( n3286 & n3288 ) | ( n3286 & ~n3292 ) | ( n3288 & ~n3292 ) ;
  assign n3323 = ( n3292 & ~n3293 ) | ( n3292 & n3322 ) | ( ~n3293 & n3322 ) ;
  assign n3324 = ( n3319 & n3321 ) | ( n3319 & n3323 ) | ( n3321 & n3323 ) ;
  assign n3325 = ( n3313 & n3315 ) | ( n3313 & n3324 ) | ( n3315 & n3324 ) ;
  assign n3326 = ( n3309 & n3311 ) | ( n3309 & n3325 ) | ( n3311 & n3325 ) ;
  assign n3327 = ( n3305 & n3307 ) | ( n3305 & n3326 ) | ( n3307 & n3326 ) ;
  assign n3328 = ( n3301 & n3303 ) | ( n3301 & n3327 ) | ( n3303 & n3327 ) ;
  assign n3329 = ( n2773 & n3298 ) | ( n2773 & ~n3328 ) | ( n3298 & ~n3328 ) ;
  assign n3330 = n2773 | n3297 ;
  assign n3331 = ( n2958 & n3328 ) | ( n2958 & n3330 ) | ( n3328 & n3330 ) ;
  assign n3332 = ( ~n3299 & n3329 ) | ( ~n3299 & n3331 ) | ( n3329 & n3331 ) ;
  assign n3333 = ( ~n2421 & n2423 ) | ( ~n2421 & n2453 ) | ( n2423 & n2453 ) ;
  assign n3334 = ( n2421 & ~n2454 ) | ( n2421 & n3333 ) | ( ~n2454 & n3333 ) ;
  assign n3335 = ( ~n2773 & n3298 ) | ( ~n2773 & n3330 ) | ( n3298 & n3330 ) ;
  assign n3336 = ( n2958 & n3328 ) | ( n2958 & n3335 ) | ( n3328 & n3335 ) ;
  assign n3337 = ( ~n2958 & n3328 ) | ( ~n2958 & n3335 ) | ( n3328 & n3335 ) ;
  assign n3338 = ( n2958 & ~n3336 ) | ( n2958 & n3337 ) | ( ~n3336 & n3337 ) ;
  assign n3339 = ( ~n2425 & n2427 ) | ( ~n2425 & n2452 ) | ( n2427 & n2452 ) ;
  assign n3340 = ( n2425 & ~n2453 ) | ( n2425 & n3339 ) | ( ~n2453 & n3339 ) ;
  assign n3341 = ( ~n3301 & n3303 ) | ( ~n3301 & n3327 ) | ( n3303 & n3327 ) ;
  assign n3342 = ( n3301 & ~n3328 ) | ( n3301 & n3341 ) | ( ~n3328 & n3341 ) ;
  assign n3343 = ( ~n3305 & n3307 ) | ( ~n3305 & n3326 ) | ( n3307 & n3326 ) ;
  assign n3344 = ( n3305 & ~n3327 ) | ( n3305 & n3343 ) | ( ~n3327 & n3343 ) ;
  assign n3345 = ( ~n2429 & n2431 ) | ( ~n2429 & n2451 ) | ( n2431 & n2451 ) ;
  assign n3346 = ( n2429 & ~n2452 ) | ( n2429 & n3345 ) | ( ~n2452 & n3345 ) ;
  assign n3347 = ( ~n2433 & n2435 ) | ( ~n2433 & n2450 ) | ( n2435 & n2450 ) ;
  assign n3348 = ( n2433 & ~n2451 ) | ( n2433 & n3347 ) | ( ~n2451 & n3347 ) ;
  assign n3349 = ( ~n3309 & n3311 ) | ( ~n3309 & n3325 ) | ( n3311 & n3325 ) ;
  assign n3350 = ( n3309 & ~n3326 ) | ( n3309 & n3349 ) | ( ~n3326 & n3349 ) ;
  assign n3351 = ( ~n3313 & n3315 ) | ( ~n3313 & n3324 ) | ( n3315 & n3324 ) ;
  assign n3352 = ( n3313 & ~n3325 ) | ( n3313 & n3351 ) | ( ~n3325 & n3351 ) ;
  assign n3353 = ( ~n2437 & n2439 ) | ( ~n2437 & n2449 ) | ( n2439 & n2449 ) ;
  assign n3354 = ( n2437 & ~n2450 ) | ( n2437 & n3353 ) | ( ~n2450 & n3353 ) ;
  assign n3355 = ( ~n2441 & n2443 ) | ( ~n2441 & n2448 ) | ( n2443 & n2448 ) ;
  assign n3356 = ( n2441 & ~n2449 ) | ( n2441 & n3355 ) | ( ~n2449 & n3355 ) ;
  assign n3357 = ( ~n3319 & n3321 ) | ( ~n3319 & n3323 ) | ( n3321 & n3323 ) ;
  assign n3358 = ( n3319 & ~n3324 ) | ( n3319 & n3357 ) | ( ~n3324 & n3357 ) ;
  assign n3359 = n3317 | n3318 ;
  assign n3360 = ~n3319 & n3359 ;
  assign n3361 = ( n2445 & n2447 ) | ( n2445 & n3360 ) | ( n2447 & n3360 ) ;
  assign n3362 = ~n2448 & n3361 ;
  assign n3363 = ( n3356 & n3358 ) | ( n3356 & n3362 ) | ( n3358 & n3362 ) ;
  assign n3364 = ( n3352 & n3354 ) | ( n3352 & n3363 ) | ( n3354 & n3363 ) ;
  assign n3365 = ( n3348 & n3350 ) | ( n3348 & n3364 ) | ( n3350 & n3364 ) ;
  assign n3366 = ( n3344 & n3346 ) | ( n3344 & n3365 ) | ( n3346 & n3365 ) ;
  assign n3367 = ( n3340 & n3342 ) | ( n3340 & n3366 ) | ( n3342 & n3366 ) ;
  assign n3368 = ( n3334 & n3338 ) | ( n3334 & n3367 ) | ( n3338 & n3367 ) ;
  assign n3369 = ( n2457 & n3332 ) | ( n2457 & n3368 ) | ( n3332 & n3368 ) ;
  assign n3370 = n3331 & ~n3332 ;
  assign n3371 = ( n2455 & n3369 ) | ( n2455 & n3370 ) | ( n3369 & n3370 ) ;
  assign n3372 = ( x844 & x845 ) | ( x844 & x846 ) | ( x845 & x846 ) ;
  assign n3373 = ( x841 & x842 ) | ( x841 & x843 ) | ( x842 & x843 ) ;
  assign n3374 = ( ~x844 & x845 ) | ( ~x844 & x846 ) | ( x845 & x846 ) ;
  assign n3375 = ( x844 & ~n3372 ) | ( x844 & n3374 ) | ( ~n3372 & n3374 ) ;
  assign n3376 = ( ~x841 & x842 ) | ( ~x841 & x843 ) | ( x842 & x843 ) ;
  assign n3377 = ( x841 & ~n3373 ) | ( x841 & n3376 ) | ( ~n3373 & n3376 ) ;
  assign n3378 = n3375 & n3377 ;
  assign n3379 = ( n3372 & n3373 ) | ( n3372 & n3378 ) | ( n3373 & n3378 ) ;
  assign n3380 = ( x835 & x836 ) | ( x835 & x837 ) | ( x836 & x837 ) ;
  assign n3381 = ( x838 & x839 ) | ( x838 & x840 ) | ( x839 & x840 ) ;
  assign n3382 = ( ~x838 & x839 ) | ( ~x838 & x840 ) | ( x839 & x840 ) ;
  assign n3383 = ( x838 & ~n3381 ) | ( x838 & n3382 ) | ( ~n3381 & n3382 ) ;
  assign n3384 = ( ~x835 & x836 ) | ( ~x835 & x837 ) | ( x836 & x837 ) ;
  assign n3385 = ( x835 & ~n3380 ) | ( x835 & n3384 ) | ( ~n3380 & n3384 ) ;
  assign n3386 = n3383 & n3385 ;
  assign n3387 = ( n3380 & n3381 ) | ( n3380 & n3386 ) | ( n3381 & n3386 ) ;
  assign n3388 = ( ~n3372 & n3373 ) | ( ~n3372 & n3378 ) | ( n3373 & n3378 ) ;
  assign n3389 = ( n3372 & ~n3379 ) | ( n3372 & n3388 ) | ( ~n3379 & n3388 ) ;
  assign n3390 = ( ~n3380 & n3381 ) | ( ~n3380 & n3386 ) | ( n3381 & n3386 ) ;
  assign n3391 = ( n3380 & ~n3387 ) | ( n3380 & n3390 ) | ( ~n3387 & n3390 ) ;
  assign n3392 = n3375 | n3377 ;
  assign n3393 = ~n3378 & n3392 ;
  assign n3394 = n3383 | n3385 ;
  assign n3395 = ~n3386 & n3394 ;
  assign n3396 = n3393 & n3395 ;
  assign n3397 = ( n3389 & n3391 ) | ( n3389 & n3396 ) | ( n3391 & n3396 ) ;
  assign n3398 = ( n3379 & n3387 ) | ( n3379 & n3397 ) | ( n3387 & n3397 ) ;
  assign n3399 = ( x832 & x833 ) | ( x832 & x834 ) | ( x833 & x834 ) ;
  assign n3400 = ( x829 & x830 ) | ( x829 & x831 ) | ( x830 & x831 ) ;
  assign n3401 = ( ~x832 & x833 ) | ( ~x832 & x834 ) | ( x833 & x834 ) ;
  assign n3402 = ( x832 & ~n3399 ) | ( x832 & n3401 ) | ( ~n3399 & n3401 ) ;
  assign n3403 = ( ~x829 & x830 ) | ( ~x829 & x831 ) | ( x830 & x831 ) ;
  assign n3404 = ( x829 & ~n3400 ) | ( x829 & n3403 ) | ( ~n3400 & n3403 ) ;
  assign n3405 = n3402 & n3404 ;
  assign n3406 = ( n3399 & n3400 ) | ( n3399 & n3405 ) | ( n3400 & n3405 ) ;
  assign n3407 = ( x823 & x824 ) | ( x823 & x825 ) | ( x824 & x825 ) ;
  assign n3408 = ( x826 & x827 ) | ( x826 & x828 ) | ( x827 & x828 ) ;
  assign n3409 = ( ~x826 & x827 ) | ( ~x826 & x828 ) | ( x827 & x828 ) ;
  assign n3410 = ( x826 & ~n3408 ) | ( x826 & n3409 ) | ( ~n3408 & n3409 ) ;
  assign n3411 = ( ~x823 & x824 ) | ( ~x823 & x825 ) | ( x824 & x825 ) ;
  assign n3412 = ( x823 & ~n3407 ) | ( x823 & n3411 ) | ( ~n3407 & n3411 ) ;
  assign n3413 = n3410 & n3412 ;
  assign n3414 = ( n3407 & n3408 ) | ( n3407 & n3413 ) | ( n3408 & n3413 ) ;
  assign n3415 = ( ~n3399 & n3400 ) | ( ~n3399 & n3405 ) | ( n3400 & n3405 ) ;
  assign n3416 = ( n3399 & ~n3406 ) | ( n3399 & n3415 ) | ( ~n3406 & n3415 ) ;
  assign n3417 = ( ~n3407 & n3408 ) | ( ~n3407 & n3413 ) | ( n3408 & n3413 ) ;
  assign n3418 = ( n3407 & ~n3414 ) | ( n3407 & n3417 ) | ( ~n3414 & n3417 ) ;
  assign n3419 = n3410 | n3412 ;
  assign n3420 = ~n3413 & n3419 ;
  assign n3421 = ( n3402 & n3404 ) | ( n3402 & n3420 ) | ( n3404 & n3420 ) ;
  assign n3422 = ~n3405 & n3421 ;
  assign n3423 = ( n3416 & n3418 ) | ( n3416 & n3422 ) | ( n3418 & n3422 ) ;
  assign n3424 = ( n3406 & n3414 ) | ( n3406 & n3423 ) | ( n3414 & n3423 ) ;
  assign n3425 = ( ~n3406 & n3414 ) | ( ~n3406 & n3423 ) | ( n3414 & n3423 ) ;
  assign n3426 = ( n3406 & ~n3424 ) | ( n3406 & n3425 ) | ( ~n3424 & n3425 ) ;
  assign n3427 = ( ~n3379 & n3387 ) | ( ~n3379 & n3397 ) | ( n3387 & n3397 ) ;
  assign n3428 = ( n3379 & ~n3398 ) | ( n3379 & n3427 ) | ( ~n3398 & n3427 ) ;
  assign n3429 = ( ~n3389 & n3391 ) | ( ~n3389 & n3396 ) | ( n3391 & n3396 ) ;
  assign n3430 = ( n3389 & ~n3397 ) | ( n3389 & n3429 ) | ( ~n3397 & n3429 ) ;
  assign n3431 = ( ~n3416 & n3418 ) | ( ~n3416 & n3422 ) | ( n3418 & n3422 ) ;
  assign n3432 = ( n3416 & ~n3423 ) | ( n3416 & n3431 ) | ( ~n3423 & n3431 ) ;
  assign n3433 = ( ~n3402 & n3404 ) | ( ~n3402 & n3420 ) | ( n3404 & n3420 ) ;
  assign n3434 = ( n3402 & ~n3421 ) | ( n3402 & n3433 ) | ( ~n3421 & n3433 ) ;
  assign n3435 = ( n3393 & n3395 ) | ( n3393 & n3434 ) | ( n3395 & n3434 ) ;
  assign n3436 = ~n3396 & n3435 ;
  assign n3437 = ( n3430 & n3432 ) | ( n3430 & n3436 ) | ( n3432 & n3436 ) ;
  assign n3438 = ( n3426 & n3428 ) | ( n3426 & n3437 ) | ( n3428 & n3437 ) ;
  assign n3439 = ( n3398 & n3424 ) | ( n3398 & n3438 ) | ( n3424 & n3438 ) ;
  assign n3440 = ( x820 & x821 ) | ( x820 & x822 ) | ( x821 & x822 ) ;
  assign n3441 = ( x817 & x818 ) | ( x817 & x819 ) | ( x818 & x819 ) ;
  assign n3442 = ( ~x820 & x821 ) | ( ~x820 & x822 ) | ( x821 & x822 ) ;
  assign n3443 = ( x820 & ~n3440 ) | ( x820 & n3442 ) | ( ~n3440 & n3442 ) ;
  assign n3444 = ( ~x817 & x818 ) | ( ~x817 & x819 ) | ( x818 & x819 ) ;
  assign n3445 = ( x817 & ~n3441 ) | ( x817 & n3444 ) | ( ~n3441 & n3444 ) ;
  assign n3446 = n3443 & n3445 ;
  assign n3447 = ( n3440 & n3441 ) | ( n3440 & n3446 ) | ( n3441 & n3446 ) ;
  assign n3448 = ( x811 & x812 ) | ( x811 & x813 ) | ( x812 & x813 ) ;
  assign n3449 = ( x814 & x815 ) | ( x814 & x816 ) | ( x815 & x816 ) ;
  assign n3450 = ( ~x814 & x815 ) | ( ~x814 & x816 ) | ( x815 & x816 ) ;
  assign n3451 = ( x814 & ~n3449 ) | ( x814 & n3450 ) | ( ~n3449 & n3450 ) ;
  assign n3452 = ( ~x811 & x812 ) | ( ~x811 & x813 ) | ( x812 & x813 ) ;
  assign n3453 = ( x811 & ~n3448 ) | ( x811 & n3452 ) | ( ~n3448 & n3452 ) ;
  assign n3454 = n3451 & n3453 ;
  assign n3455 = ( n3448 & n3449 ) | ( n3448 & n3454 ) | ( n3449 & n3454 ) ;
  assign n3456 = ( ~n3440 & n3441 ) | ( ~n3440 & n3446 ) | ( n3441 & n3446 ) ;
  assign n3457 = ( n3440 & ~n3447 ) | ( n3440 & n3456 ) | ( ~n3447 & n3456 ) ;
  assign n3458 = ( ~n3448 & n3449 ) | ( ~n3448 & n3454 ) | ( n3449 & n3454 ) ;
  assign n3459 = ( n3448 & ~n3455 ) | ( n3448 & n3458 ) | ( ~n3455 & n3458 ) ;
  assign n3460 = n3443 | n3445 ;
  assign n3461 = ~n3446 & n3460 ;
  assign n3462 = n3451 | n3453 ;
  assign n3463 = ~n3454 & n3462 ;
  assign n3464 = n3461 & n3463 ;
  assign n3465 = ( n3457 & n3459 ) | ( n3457 & n3464 ) | ( n3459 & n3464 ) ;
  assign n3466 = ( n3447 & n3455 ) | ( n3447 & n3465 ) | ( n3455 & n3465 ) ;
  assign n3467 = ( x808 & x809 ) | ( x808 & x810 ) | ( x809 & x810 ) ;
  assign n3468 = ( x805 & x806 ) | ( x805 & x807 ) | ( x806 & x807 ) ;
  assign n3469 = ( ~x808 & x809 ) | ( ~x808 & x810 ) | ( x809 & x810 ) ;
  assign n3470 = ( x808 & ~n3467 ) | ( x808 & n3469 ) | ( ~n3467 & n3469 ) ;
  assign n3471 = ( ~x805 & x806 ) | ( ~x805 & x807 ) | ( x806 & x807 ) ;
  assign n3472 = ( x805 & ~n3468 ) | ( x805 & n3471 ) | ( ~n3468 & n3471 ) ;
  assign n3473 = n3470 & n3472 ;
  assign n3474 = ( n3467 & n3468 ) | ( n3467 & n3473 ) | ( n3468 & n3473 ) ;
  assign n3475 = ( x799 & x800 ) | ( x799 & x801 ) | ( x800 & x801 ) ;
  assign n3476 = ( x802 & x803 ) | ( x802 & x804 ) | ( x803 & x804 ) ;
  assign n3477 = ( ~x802 & x803 ) | ( ~x802 & x804 ) | ( x803 & x804 ) ;
  assign n3478 = ( x802 & ~n3476 ) | ( x802 & n3477 ) | ( ~n3476 & n3477 ) ;
  assign n3479 = ( ~x799 & x800 ) | ( ~x799 & x801 ) | ( x800 & x801 ) ;
  assign n3480 = ( x799 & ~n3475 ) | ( x799 & n3479 ) | ( ~n3475 & n3479 ) ;
  assign n3481 = n3478 & n3480 ;
  assign n3482 = ( n3475 & n3476 ) | ( n3475 & n3481 ) | ( n3476 & n3481 ) ;
  assign n3483 = ( ~n3467 & n3468 ) | ( ~n3467 & n3473 ) | ( n3468 & n3473 ) ;
  assign n3484 = ( n3467 & ~n3474 ) | ( n3467 & n3483 ) | ( ~n3474 & n3483 ) ;
  assign n3485 = ( ~n3475 & n3476 ) | ( ~n3475 & n3481 ) | ( n3476 & n3481 ) ;
  assign n3486 = ( n3475 & ~n3482 ) | ( n3475 & n3485 ) | ( ~n3482 & n3485 ) ;
  assign n3487 = n3478 | n3480 ;
  assign n3488 = ~n3481 & n3487 ;
  assign n3489 = ( n3470 & n3472 ) | ( n3470 & n3488 ) | ( n3472 & n3488 ) ;
  assign n3490 = ~n3473 & n3489 ;
  assign n3491 = ( n3484 & n3486 ) | ( n3484 & n3490 ) | ( n3486 & n3490 ) ;
  assign n3492 = ( n3474 & n3482 ) | ( n3474 & n3491 ) | ( n3482 & n3491 ) ;
  assign n3493 = ( ~n3474 & n3482 ) | ( ~n3474 & n3491 ) | ( n3482 & n3491 ) ;
  assign n3494 = ( n3474 & ~n3492 ) | ( n3474 & n3493 ) | ( ~n3492 & n3493 ) ;
  assign n3495 = ( ~n3447 & n3455 ) | ( ~n3447 & n3465 ) | ( n3455 & n3465 ) ;
  assign n3496 = ( n3447 & ~n3466 ) | ( n3447 & n3495 ) | ( ~n3466 & n3495 ) ;
  assign n3497 = ( ~n3457 & n3459 ) | ( ~n3457 & n3464 ) | ( n3459 & n3464 ) ;
  assign n3498 = ( n3457 & ~n3465 ) | ( n3457 & n3497 ) | ( ~n3465 & n3497 ) ;
  assign n3499 = ( ~n3484 & n3486 ) | ( ~n3484 & n3490 ) | ( n3486 & n3490 ) ;
  assign n3500 = ( n3484 & ~n3491 ) | ( n3484 & n3499 ) | ( ~n3491 & n3499 ) ;
  assign n3501 = ( ~n3470 & n3472 ) | ( ~n3470 & n3488 ) | ( n3472 & n3488 ) ;
  assign n3502 = ( n3470 & ~n3489 ) | ( n3470 & n3501 ) | ( ~n3489 & n3501 ) ;
  assign n3503 = ( n3461 & n3463 ) | ( n3461 & n3502 ) | ( n3463 & n3502 ) ;
  assign n3504 = ~n3464 & n3503 ;
  assign n3505 = ( n3498 & n3500 ) | ( n3498 & n3504 ) | ( n3500 & n3504 ) ;
  assign n3506 = ( n3494 & n3496 ) | ( n3494 & n3505 ) | ( n3496 & n3505 ) ;
  assign n3507 = ( n3466 & n3492 ) | ( n3466 & n3506 ) | ( n3492 & n3506 ) ;
  assign n3508 = ( ~n3398 & n3424 ) | ( ~n3398 & n3438 ) | ( n3424 & n3438 ) ;
  assign n3509 = ( n3398 & ~n3439 ) | ( n3398 & n3508 ) | ( ~n3439 & n3508 ) ;
  assign n3510 = ( ~n3466 & n3492 ) | ( ~n3466 & n3506 ) | ( n3492 & n3506 ) ;
  assign n3511 = ( n3466 & ~n3507 ) | ( n3466 & n3510 ) | ( ~n3507 & n3510 ) ;
  assign n3512 = ( ~n3494 & n3496 ) | ( ~n3494 & n3505 ) | ( n3496 & n3505 ) ;
  assign n3513 = ( n3494 & ~n3506 ) | ( n3494 & n3512 ) | ( ~n3506 & n3512 ) ;
  assign n3514 = ( ~n3426 & n3428 ) | ( ~n3426 & n3437 ) | ( n3428 & n3437 ) ;
  assign n3515 = ( n3426 & ~n3438 ) | ( n3426 & n3514 ) | ( ~n3438 & n3514 ) ;
  assign n3516 = ( n3430 & n3432 ) | ( n3430 & ~n3436 ) | ( n3432 & ~n3436 ) ;
  assign n3517 = ( n3436 & ~n3437 ) | ( n3436 & n3516 ) | ( ~n3437 & n3516 ) ;
  assign n3518 = ( n3498 & n3500 ) | ( n3498 & ~n3504 ) | ( n3500 & ~n3504 ) ;
  assign n3519 = ( n3504 & ~n3505 ) | ( n3504 & n3518 ) | ( ~n3505 & n3518 ) ;
  assign n3520 = ( ~n3393 & n3395 ) | ( ~n3393 & n3434 ) | ( n3395 & n3434 ) ;
  assign n3521 = ( n3393 & ~n3435 ) | ( n3393 & n3520 ) | ( ~n3435 & n3520 ) ;
  assign n3522 = ( ~n3461 & n3463 ) | ( ~n3461 & n3502 ) | ( n3463 & n3502 ) ;
  assign n3523 = ( n3461 & ~n3503 ) | ( n3461 & n3522 ) | ( ~n3503 & n3522 ) ;
  assign n3524 = n3521 & n3523 ;
  assign n3525 = ( n3517 & n3519 ) | ( n3517 & n3524 ) | ( n3519 & n3524 ) ;
  assign n3526 = ( n3513 & n3515 ) | ( n3513 & n3525 ) | ( n3515 & n3525 ) ;
  assign n3527 = ( n3509 & n3511 ) | ( n3509 & n3526 ) | ( n3511 & n3526 ) ;
  assign n3528 = ( n3439 & n3507 ) | ( n3439 & n3527 ) | ( n3507 & n3527 ) ;
  assign n3529 = ( x796 & x797 ) | ( x796 & x798 ) | ( x797 & x798 ) ;
  assign n3530 = ( x793 & x794 ) | ( x793 & x795 ) | ( x794 & x795 ) ;
  assign n3531 = ( ~x796 & x797 ) | ( ~x796 & x798 ) | ( x797 & x798 ) ;
  assign n3532 = ( x796 & ~n3529 ) | ( x796 & n3531 ) | ( ~n3529 & n3531 ) ;
  assign n3533 = ( ~x793 & x794 ) | ( ~x793 & x795 ) | ( x794 & x795 ) ;
  assign n3534 = ( x793 & ~n3530 ) | ( x793 & n3533 ) | ( ~n3530 & n3533 ) ;
  assign n3535 = n3532 & n3534 ;
  assign n3536 = ( n3529 & n3530 ) | ( n3529 & n3535 ) | ( n3530 & n3535 ) ;
  assign n3537 = ( x787 & x788 ) | ( x787 & x789 ) | ( x788 & x789 ) ;
  assign n3538 = ( x790 & x791 ) | ( x790 & x792 ) | ( x791 & x792 ) ;
  assign n3539 = ( ~x790 & x791 ) | ( ~x790 & x792 ) | ( x791 & x792 ) ;
  assign n3540 = ( x790 & ~n3538 ) | ( x790 & n3539 ) | ( ~n3538 & n3539 ) ;
  assign n3541 = ( ~x787 & x788 ) | ( ~x787 & x789 ) | ( x788 & x789 ) ;
  assign n3542 = ( x787 & ~n3537 ) | ( x787 & n3541 ) | ( ~n3537 & n3541 ) ;
  assign n3543 = n3540 & n3542 ;
  assign n3544 = ( n3537 & n3538 ) | ( n3537 & n3543 ) | ( n3538 & n3543 ) ;
  assign n3545 = ( ~n3529 & n3530 ) | ( ~n3529 & n3535 ) | ( n3530 & n3535 ) ;
  assign n3546 = ( n3529 & ~n3536 ) | ( n3529 & n3545 ) | ( ~n3536 & n3545 ) ;
  assign n3547 = ( ~n3537 & n3538 ) | ( ~n3537 & n3543 ) | ( n3538 & n3543 ) ;
  assign n3548 = ( n3537 & ~n3544 ) | ( n3537 & n3547 ) | ( ~n3544 & n3547 ) ;
  assign n3549 = n3532 | n3534 ;
  assign n3550 = ~n3535 & n3549 ;
  assign n3551 = n3540 | n3542 ;
  assign n3552 = ~n3543 & n3551 ;
  assign n3553 = n3550 & n3552 ;
  assign n3554 = ( n3546 & n3548 ) | ( n3546 & n3553 ) | ( n3548 & n3553 ) ;
  assign n3555 = ( n3536 & n3544 ) | ( n3536 & n3554 ) | ( n3544 & n3554 ) ;
  assign n3556 = ( x784 & x785 ) | ( x784 & x786 ) | ( x785 & x786 ) ;
  assign n3557 = ( x781 & x782 ) | ( x781 & x783 ) | ( x782 & x783 ) ;
  assign n3558 = ( ~x784 & x785 ) | ( ~x784 & x786 ) | ( x785 & x786 ) ;
  assign n3559 = ( x784 & ~n3556 ) | ( x784 & n3558 ) | ( ~n3556 & n3558 ) ;
  assign n3560 = ( ~x781 & x782 ) | ( ~x781 & x783 ) | ( x782 & x783 ) ;
  assign n3561 = ( x781 & ~n3557 ) | ( x781 & n3560 ) | ( ~n3557 & n3560 ) ;
  assign n3562 = n3559 & n3561 ;
  assign n3563 = ( n3556 & n3557 ) | ( n3556 & n3562 ) | ( n3557 & n3562 ) ;
  assign n3564 = ( x775 & x776 ) | ( x775 & x777 ) | ( x776 & x777 ) ;
  assign n3565 = ( x778 & x779 ) | ( x778 & x780 ) | ( x779 & x780 ) ;
  assign n3566 = ( ~x778 & x779 ) | ( ~x778 & x780 ) | ( x779 & x780 ) ;
  assign n3567 = ( x778 & ~n3565 ) | ( x778 & n3566 ) | ( ~n3565 & n3566 ) ;
  assign n3568 = ( ~x775 & x776 ) | ( ~x775 & x777 ) | ( x776 & x777 ) ;
  assign n3569 = ( x775 & ~n3564 ) | ( x775 & n3568 ) | ( ~n3564 & n3568 ) ;
  assign n3570 = n3567 & n3569 ;
  assign n3571 = ( n3564 & n3565 ) | ( n3564 & n3570 ) | ( n3565 & n3570 ) ;
  assign n3572 = ( ~n3556 & n3557 ) | ( ~n3556 & n3562 ) | ( n3557 & n3562 ) ;
  assign n3573 = ( n3556 & ~n3563 ) | ( n3556 & n3572 ) | ( ~n3563 & n3572 ) ;
  assign n3574 = ( ~n3564 & n3565 ) | ( ~n3564 & n3570 ) | ( n3565 & n3570 ) ;
  assign n3575 = ( n3564 & ~n3571 ) | ( n3564 & n3574 ) | ( ~n3571 & n3574 ) ;
  assign n3576 = n3567 | n3569 ;
  assign n3577 = ~n3570 & n3576 ;
  assign n3578 = ( n3559 & n3561 ) | ( n3559 & n3577 ) | ( n3561 & n3577 ) ;
  assign n3579 = ~n3562 & n3578 ;
  assign n3580 = ( n3573 & n3575 ) | ( n3573 & n3579 ) | ( n3575 & n3579 ) ;
  assign n3581 = ( n3563 & n3571 ) | ( n3563 & n3580 ) | ( n3571 & n3580 ) ;
  assign n3582 = ( ~n3563 & n3571 ) | ( ~n3563 & n3580 ) | ( n3571 & n3580 ) ;
  assign n3583 = ( n3563 & ~n3581 ) | ( n3563 & n3582 ) | ( ~n3581 & n3582 ) ;
  assign n3584 = ( ~n3536 & n3544 ) | ( ~n3536 & n3554 ) | ( n3544 & n3554 ) ;
  assign n3585 = ( n3536 & ~n3555 ) | ( n3536 & n3584 ) | ( ~n3555 & n3584 ) ;
  assign n3586 = ( ~n3546 & n3548 ) | ( ~n3546 & n3553 ) | ( n3548 & n3553 ) ;
  assign n3587 = ( n3546 & ~n3554 ) | ( n3546 & n3586 ) | ( ~n3554 & n3586 ) ;
  assign n3588 = ( ~n3573 & n3575 ) | ( ~n3573 & n3579 ) | ( n3575 & n3579 ) ;
  assign n3589 = ( n3573 & ~n3580 ) | ( n3573 & n3588 ) | ( ~n3580 & n3588 ) ;
  assign n3590 = ( ~n3559 & n3561 ) | ( ~n3559 & n3577 ) | ( n3561 & n3577 ) ;
  assign n3591 = ( n3559 & ~n3578 ) | ( n3559 & n3590 ) | ( ~n3578 & n3590 ) ;
  assign n3592 = ( n3550 & n3552 ) | ( n3550 & n3591 ) | ( n3552 & n3591 ) ;
  assign n3593 = ~n3553 & n3592 ;
  assign n3594 = ( n3587 & n3589 ) | ( n3587 & n3593 ) | ( n3589 & n3593 ) ;
  assign n3595 = ( n3583 & n3585 ) | ( n3583 & n3594 ) | ( n3585 & n3594 ) ;
  assign n3596 = ( n3555 & n3581 ) | ( n3555 & n3595 ) | ( n3581 & n3595 ) ;
  assign n3597 = ( x772 & x773 ) | ( x772 & x774 ) | ( x773 & x774 ) ;
  assign n3598 = ( x769 & x770 ) | ( x769 & x771 ) | ( x770 & x771 ) ;
  assign n3599 = ( ~x772 & x773 ) | ( ~x772 & x774 ) | ( x773 & x774 ) ;
  assign n3600 = ( x772 & ~n3597 ) | ( x772 & n3599 ) | ( ~n3597 & n3599 ) ;
  assign n3601 = ( ~x769 & x770 ) | ( ~x769 & x771 ) | ( x770 & x771 ) ;
  assign n3602 = ( x769 & ~n3598 ) | ( x769 & n3601 ) | ( ~n3598 & n3601 ) ;
  assign n3603 = n3600 & n3602 ;
  assign n3604 = ( n3597 & n3598 ) | ( n3597 & n3603 ) | ( n3598 & n3603 ) ;
  assign n3605 = ( x763 & x764 ) | ( x763 & x765 ) | ( x764 & x765 ) ;
  assign n3606 = ( x766 & x767 ) | ( x766 & x768 ) | ( x767 & x768 ) ;
  assign n3607 = ( ~x766 & x767 ) | ( ~x766 & x768 ) | ( x767 & x768 ) ;
  assign n3608 = ( x766 & ~n3606 ) | ( x766 & n3607 ) | ( ~n3606 & n3607 ) ;
  assign n3609 = ( ~x763 & x764 ) | ( ~x763 & x765 ) | ( x764 & x765 ) ;
  assign n3610 = ( x763 & ~n3605 ) | ( x763 & n3609 ) | ( ~n3605 & n3609 ) ;
  assign n3611 = n3608 & n3610 ;
  assign n3612 = ( n3605 & n3606 ) | ( n3605 & n3611 ) | ( n3606 & n3611 ) ;
  assign n3613 = ( ~n3597 & n3598 ) | ( ~n3597 & n3603 ) | ( n3598 & n3603 ) ;
  assign n3614 = ( n3597 & ~n3604 ) | ( n3597 & n3613 ) | ( ~n3604 & n3613 ) ;
  assign n3615 = ( ~n3605 & n3606 ) | ( ~n3605 & n3611 ) | ( n3606 & n3611 ) ;
  assign n3616 = ( n3605 & ~n3612 ) | ( n3605 & n3615 ) | ( ~n3612 & n3615 ) ;
  assign n3617 = n3600 | n3602 ;
  assign n3618 = ~n3603 & n3617 ;
  assign n3619 = n3608 | n3610 ;
  assign n3620 = ~n3611 & n3619 ;
  assign n3621 = n3618 & n3620 ;
  assign n3622 = ( n3614 & n3616 ) | ( n3614 & n3621 ) | ( n3616 & n3621 ) ;
  assign n3623 = ( n3604 & n3612 ) | ( n3604 & n3622 ) | ( n3612 & n3622 ) ;
  assign n3624 = ( x760 & x761 ) | ( x760 & x762 ) | ( x761 & x762 ) ;
  assign n3625 = ( x757 & x758 ) | ( x757 & x759 ) | ( x758 & x759 ) ;
  assign n3626 = ( ~x760 & x761 ) | ( ~x760 & x762 ) | ( x761 & x762 ) ;
  assign n3627 = ( x760 & ~n3624 ) | ( x760 & n3626 ) | ( ~n3624 & n3626 ) ;
  assign n3628 = ( ~x757 & x758 ) | ( ~x757 & x759 ) | ( x758 & x759 ) ;
  assign n3629 = ( x757 & ~n3625 ) | ( x757 & n3628 ) | ( ~n3625 & n3628 ) ;
  assign n3630 = n3627 & n3629 ;
  assign n3631 = ( n3624 & n3625 ) | ( n3624 & n3630 ) | ( n3625 & n3630 ) ;
  assign n3632 = ( x751 & x752 ) | ( x751 & x753 ) | ( x752 & x753 ) ;
  assign n3633 = ( x754 & x755 ) | ( x754 & x756 ) | ( x755 & x756 ) ;
  assign n3634 = ( ~x754 & x755 ) | ( ~x754 & x756 ) | ( x755 & x756 ) ;
  assign n3635 = ( x754 & ~n3633 ) | ( x754 & n3634 ) | ( ~n3633 & n3634 ) ;
  assign n3636 = ( ~x751 & x752 ) | ( ~x751 & x753 ) | ( x752 & x753 ) ;
  assign n3637 = ( x751 & ~n3632 ) | ( x751 & n3636 ) | ( ~n3632 & n3636 ) ;
  assign n3638 = n3635 & n3637 ;
  assign n3639 = ( n3632 & n3633 ) | ( n3632 & n3638 ) | ( n3633 & n3638 ) ;
  assign n3640 = ( ~n3624 & n3625 ) | ( ~n3624 & n3630 ) | ( n3625 & n3630 ) ;
  assign n3641 = ( n3624 & ~n3631 ) | ( n3624 & n3640 ) | ( ~n3631 & n3640 ) ;
  assign n3642 = ( ~n3632 & n3633 ) | ( ~n3632 & n3638 ) | ( n3633 & n3638 ) ;
  assign n3643 = ( n3632 & ~n3639 ) | ( n3632 & n3642 ) | ( ~n3639 & n3642 ) ;
  assign n3644 = n3635 | n3637 ;
  assign n3645 = ~n3638 & n3644 ;
  assign n3646 = ( n3627 & n3629 ) | ( n3627 & n3645 ) | ( n3629 & n3645 ) ;
  assign n3647 = ~n3630 & n3646 ;
  assign n3648 = ( n3641 & n3643 ) | ( n3641 & n3647 ) | ( n3643 & n3647 ) ;
  assign n3649 = ( n3631 & n3639 ) | ( n3631 & n3648 ) | ( n3639 & n3648 ) ;
  assign n3650 = ( ~n3631 & n3639 ) | ( ~n3631 & n3648 ) | ( n3639 & n3648 ) ;
  assign n3651 = ( n3631 & ~n3649 ) | ( n3631 & n3650 ) | ( ~n3649 & n3650 ) ;
  assign n3652 = ( ~n3604 & n3612 ) | ( ~n3604 & n3622 ) | ( n3612 & n3622 ) ;
  assign n3653 = ( n3604 & ~n3623 ) | ( n3604 & n3652 ) | ( ~n3623 & n3652 ) ;
  assign n3654 = ( ~n3614 & n3616 ) | ( ~n3614 & n3621 ) | ( n3616 & n3621 ) ;
  assign n3655 = ( n3614 & ~n3622 ) | ( n3614 & n3654 ) | ( ~n3622 & n3654 ) ;
  assign n3656 = ( ~n3641 & n3643 ) | ( ~n3641 & n3647 ) | ( n3643 & n3647 ) ;
  assign n3657 = ( n3641 & ~n3648 ) | ( n3641 & n3656 ) | ( ~n3648 & n3656 ) ;
  assign n3658 = ( ~n3627 & n3629 ) | ( ~n3627 & n3645 ) | ( n3629 & n3645 ) ;
  assign n3659 = ( n3627 & ~n3646 ) | ( n3627 & n3658 ) | ( ~n3646 & n3658 ) ;
  assign n3660 = ( n3618 & n3620 ) | ( n3618 & n3659 ) | ( n3620 & n3659 ) ;
  assign n3661 = ~n3621 & n3660 ;
  assign n3662 = ( n3655 & n3657 ) | ( n3655 & n3661 ) | ( n3657 & n3661 ) ;
  assign n3663 = ( n3651 & n3653 ) | ( n3651 & n3662 ) | ( n3653 & n3662 ) ;
  assign n3664 = ( n3623 & n3649 ) | ( n3623 & n3663 ) | ( n3649 & n3663 ) ;
  assign n3665 = ( ~n3555 & n3581 ) | ( ~n3555 & n3595 ) | ( n3581 & n3595 ) ;
  assign n3666 = ( n3555 & ~n3596 ) | ( n3555 & n3665 ) | ( ~n3596 & n3665 ) ;
  assign n3667 = ( ~n3623 & n3649 ) | ( ~n3623 & n3663 ) | ( n3649 & n3663 ) ;
  assign n3668 = ( n3623 & ~n3664 ) | ( n3623 & n3667 ) | ( ~n3664 & n3667 ) ;
  assign n3669 = ( ~n3651 & n3653 ) | ( ~n3651 & n3662 ) | ( n3653 & n3662 ) ;
  assign n3670 = ( n3651 & ~n3663 ) | ( n3651 & n3669 ) | ( ~n3663 & n3669 ) ;
  assign n3671 = ( ~n3583 & n3585 ) | ( ~n3583 & n3594 ) | ( n3585 & n3594 ) ;
  assign n3672 = ( n3583 & ~n3595 ) | ( n3583 & n3671 ) | ( ~n3595 & n3671 ) ;
  assign n3673 = ( n3587 & n3589 ) | ( n3587 & ~n3593 ) | ( n3589 & ~n3593 ) ;
  assign n3674 = ( n3593 & ~n3594 ) | ( n3593 & n3673 ) | ( ~n3594 & n3673 ) ;
  assign n3675 = ( n3655 & n3657 ) | ( n3655 & ~n3661 ) | ( n3657 & ~n3661 ) ;
  assign n3676 = ( n3661 & ~n3662 ) | ( n3661 & n3675 ) | ( ~n3662 & n3675 ) ;
  assign n3677 = ( ~n3550 & n3552 ) | ( ~n3550 & n3591 ) | ( n3552 & n3591 ) ;
  assign n3678 = ( n3550 & ~n3592 ) | ( n3550 & n3677 ) | ( ~n3592 & n3677 ) ;
  assign n3679 = ( ~n3618 & n3620 ) | ( ~n3618 & n3659 ) | ( n3620 & n3659 ) ;
  assign n3680 = ( n3618 & ~n3660 ) | ( n3618 & n3679 ) | ( ~n3660 & n3679 ) ;
  assign n3681 = n3678 & n3680 ;
  assign n3682 = ( n3674 & n3676 ) | ( n3674 & n3681 ) | ( n3676 & n3681 ) ;
  assign n3683 = ( n3670 & n3672 ) | ( n3670 & n3682 ) | ( n3672 & n3682 ) ;
  assign n3684 = ( n3666 & n3668 ) | ( n3666 & n3683 ) | ( n3668 & n3683 ) ;
  assign n3685 = ( n3596 & n3664 ) | ( n3596 & n3684 ) | ( n3664 & n3684 ) ;
  assign n3686 = ( ~n3596 & n3664 ) | ( ~n3596 & n3684 ) | ( n3664 & n3684 ) ;
  assign n3687 = ( n3596 & ~n3685 ) | ( n3596 & n3686 ) | ( ~n3685 & n3686 ) ;
  assign n3688 = ( ~n3439 & n3507 ) | ( ~n3439 & n3527 ) | ( n3507 & n3527 ) ;
  assign n3689 = ( n3439 & ~n3528 ) | ( n3439 & n3688 ) | ( ~n3528 & n3688 ) ;
  assign n3690 = ( ~n3509 & n3511 ) | ( ~n3509 & n3526 ) | ( n3511 & n3526 ) ;
  assign n3691 = ( n3509 & ~n3527 ) | ( n3509 & n3690 ) | ( ~n3527 & n3690 ) ;
  assign n3692 = ( ~n3666 & n3668 ) | ( ~n3666 & n3683 ) | ( n3668 & n3683 ) ;
  assign n3693 = ( n3666 & ~n3684 ) | ( n3666 & n3692 ) | ( ~n3684 & n3692 ) ;
  assign n3694 = ( ~n3670 & n3672 ) | ( ~n3670 & n3682 ) | ( n3672 & n3682 ) ;
  assign n3695 = ( n3670 & ~n3683 ) | ( n3670 & n3694 ) | ( ~n3683 & n3694 ) ;
  assign n3696 = ( ~n3513 & n3515 ) | ( ~n3513 & n3525 ) | ( n3515 & n3525 ) ;
  assign n3697 = ( n3513 & ~n3526 ) | ( n3513 & n3696 ) | ( ~n3526 & n3696 ) ;
  assign n3698 = ( ~n3517 & n3519 ) | ( ~n3517 & n3524 ) | ( n3519 & n3524 ) ;
  assign n3699 = ( n3517 & ~n3525 ) | ( n3517 & n3698 ) | ( ~n3525 & n3698 ) ;
  assign n3700 = ( ~n3674 & n3676 ) | ( ~n3674 & n3681 ) | ( n3676 & n3681 ) ;
  assign n3701 = ( n3674 & ~n3682 ) | ( n3674 & n3700 ) | ( ~n3682 & n3700 ) ;
  assign n3702 = n3678 | n3680 ;
  assign n3703 = ~n3681 & n3702 ;
  assign n3704 = ( n3521 & n3523 ) | ( n3521 & n3703 ) | ( n3523 & n3703 ) ;
  assign n3705 = ~n3524 & n3704 ;
  assign n3706 = ( n3699 & n3701 ) | ( n3699 & n3705 ) | ( n3701 & n3705 ) ;
  assign n3707 = ( n3695 & n3697 ) | ( n3695 & n3706 ) | ( n3697 & n3706 ) ;
  assign n3708 = ( n3691 & n3693 ) | ( n3691 & n3707 ) | ( n3693 & n3707 ) ;
  assign n3709 = ( n3687 & n3689 ) | ( n3687 & n3708 ) | ( n3689 & n3708 ) ;
  assign n3710 = ( n3528 & n3685 ) | ( n3528 & n3709 ) | ( n3685 & n3709 ) ;
  assign n3711 = ( x748 & x749 ) | ( x748 & x750 ) | ( x749 & x750 ) ;
  assign n3712 = ( x745 & x746 ) | ( x745 & x747 ) | ( x746 & x747 ) ;
  assign n3713 = ( ~x748 & x749 ) | ( ~x748 & x750 ) | ( x749 & x750 ) ;
  assign n3714 = ( x748 & ~n3711 ) | ( x748 & n3713 ) | ( ~n3711 & n3713 ) ;
  assign n3715 = ( ~x745 & x746 ) | ( ~x745 & x747 ) | ( x746 & x747 ) ;
  assign n3716 = ( x745 & ~n3712 ) | ( x745 & n3715 ) | ( ~n3712 & n3715 ) ;
  assign n3717 = n3714 & n3716 ;
  assign n3718 = ( n3711 & n3712 ) | ( n3711 & n3717 ) | ( n3712 & n3717 ) ;
  assign n3719 = ( x739 & x740 ) | ( x739 & x741 ) | ( x740 & x741 ) ;
  assign n3720 = ( x742 & x743 ) | ( x742 & x744 ) | ( x743 & x744 ) ;
  assign n3721 = ( ~x742 & x743 ) | ( ~x742 & x744 ) | ( x743 & x744 ) ;
  assign n3722 = ( x742 & ~n3720 ) | ( x742 & n3721 ) | ( ~n3720 & n3721 ) ;
  assign n3723 = ( ~x739 & x740 ) | ( ~x739 & x741 ) | ( x740 & x741 ) ;
  assign n3724 = ( x739 & ~n3719 ) | ( x739 & n3723 ) | ( ~n3719 & n3723 ) ;
  assign n3725 = n3722 & n3724 ;
  assign n3726 = ( n3719 & n3720 ) | ( n3719 & n3725 ) | ( n3720 & n3725 ) ;
  assign n3727 = ( ~n3711 & n3712 ) | ( ~n3711 & n3717 ) | ( n3712 & n3717 ) ;
  assign n3728 = ( n3711 & ~n3718 ) | ( n3711 & n3727 ) | ( ~n3718 & n3727 ) ;
  assign n3729 = ( ~n3719 & n3720 ) | ( ~n3719 & n3725 ) | ( n3720 & n3725 ) ;
  assign n3730 = ( n3719 & ~n3726 ) | ( n3719 & n3729 ) | ( ~n3726 & n3729 ) ;
  assign n3731 = n3714 | n3716 ;
  assign n3732 = ~n3717 & n3731 ;
  assign n3733 = n3722 | n3724 ;
  assign n3734 = ~n3725 & n3733 ;
  assign n3735 = n3732 & n3734 ;
  assign n3736 = ( n3728 & n3730 ) | ( n3728 & n3735 ) | ( n3730 & n3735 ) ;
  assign n3737 = ( n3718 & n3726 ) | ( n3718 & n3736 ) | ( n3726 & n3736 ) ;
  assign n3738 = ( x736 & x737 ) | ( x736 & x738 ) | ( x737 & x738 ) ;
  assign n3739 = ( x733 & x734 ) | ( x733 & x735 ) | ( x734 & x735 ) ;
  assign n3740 = ( ~x736 & x737 ) | ( ~x736 & x738 ) | ( x737 & x738 ) ;
  assign n3741 = ( x736 & ~n3738 ) | ( x736 & n3740 ) | ( ~n3738 & n3740 ) ;
  assign n3742 = ( ~x733 & x734 ) | ( ~x733 & x735 ) | ( x734 & x735 ) ;
  assign n3743 = ( x733 & ~n3739 ) | ( x733 & n3742 ) | ( ~n3739 & n3742 ) ;
  assign n3744 = n3741 & n3743 ;
  assign n3745 = ( n3738 & n3739 ) | ( n3738 & n3744 ) | ( n3739 & n3744 ) ;
  assign n3746 = ( x727 & x728 ) | ( x727 & x729 ) | ( x728 & x729 ) ;
  assign n3747 = ( x730 & x731 ) | ( x730 & x732 ) | ( x731 & x732 ) ;
  assign n3748 = ( ~x730 & x731 ) | ( ~x730 & x732 ) | ( x731 & x732 ) ;
  assign n3749 = ( x730 & ~n3747 ) | ( x730 & n3748 ) | ( ~n3747 & n3748 ) ;
  assign n3750 = ( ~x727 & x728 ) | ( ~x727 & x729 ) | ( x728 & x729 ) ;
  assign n3751 = ( x727 & ~n3746 ) | ( x727 & n3750 ) | ( ~n3746 & n3750 ) ;
  assign n3752 = n3749 & n3751 ;
  assign n3753 = ( n3746 & n3747 ) | ( n3746 & n3752 ) | ( n3747 & n3752 ) ;
  assign n3754 = ( ~n3738 & n3739 ) | ( ~n3738 & n3744 ) | ( n3739 & n3744 ) ;
  assign n3755 = ( n3738 & ~n3745 ) | ( n3738 & n3754 ) | ( ~n3745 & n3754 ) ;
  assign n3756 = ( ~n3746 & n3747 ) | ( ~n3746 & n3752 ) | ( n3747 & n3752 ) ;
  assign n3757 = ( n3746 & ~n3753 ) | ( n3746 & n3756 ) | ( ~n3753 & n3756 ) ;
  assign n3758 = n3749 | n3751 ;
  assign n3759 = ~n3752 & n3758 ;
  assign n3760 = ( n3741 & n3743 ) | ( n3741 & n3759 ) | ( n3743 & n3759 ) ;
  assign n3761 = ~n3744 & n3760 ;
  assign n3762 = ( n3755 & n3757 ) | ( n3755 & n3761 ) | ( n3757 & n3761 ) ;
  assign n3763 = ( n3745 & n3753 ) | ( n3745 & n3762 ) | ( n3753 & n3762 ) ;
  assign n3764 = ( ~n3745 & n3753 ) | ( ~n3745 & n3762 ) | ( n3753 & n3762 ) ;
  assign n3765 = ( n3745 & ~n3763 ) | ( n3745 & n3764 ) | ( ~n3763 & n3764 ) ;
  assign n3766 = ( ~n3718 & n3726 ) | ( ~n3718 & n3736 ) | ( n3726 & n3736 ) ;
  assign n3767 = ( n3718 & ~n3737 ) | ( n3718 & n3766 ) | ( ~n3737 & n3766 ) ;
  assign n3768 = ( ~n3728 & n3730 ) | ( ~n3728 & n3735 ) | ( n3730 & n3735 ) ;
  assign n3769 = ( n3728 & ~n3736 ) | ( n3728 & n3768 ) | ( ~n3736 & n3768 ) ;
  assign n3770 = ( ~n3755 & n3757 ) | ( ~n3755 & n3761 ) | ( n3757 & n3761 ) ;
  assign n3771 = ( n3755 & ~n3762 ) | ( n3755 & n3770 ) | ( ~n3762 & n3770 ) ;
  assign n3772 = ( ~n3741 & n3743 ) | ( ~n3741 & n3759 ) | ( n3743 & n3759 ) ;
  assign n3773 = ( n3741 & ~n3760 ) | ( n3741 & n3772 ) | ( ~n3760 & n3772 ) ;
  assign n3774 = ( n3732 & n3734 ) | ( n3732 & n3773 ) | ( n3734 & n3773 ) ;
  assign n3775 = ~n3735 & n3774 ;
  assign n3776 = ( n3769 & n3771 ) | ( n3769 & n3775 ) | ( n3771 & n3775 ) ;
  assign n3777 = ( n3765 & n3767 ) | ( n3765 & n3776 ) | ( n3767 & n3776 ) ;
  assign n3778 = ( n3737 & n3763 ) | ( n3737 & n3777 ) | ( n3763 & n3777 ) ;
  assign n3779 = ( x724 & x725 ) | ( x724 & x726 ) | ( x725 & x726 ) ;
  assign n3780 = ( x721 & x722 ) | ( x721 & x723 ) | ( x722 & x723 ) ;
  assign n3781 = ( ~x724 & x725 ) | ( ~x724 & x726 ) | ( x725 & x726 ) ;
  assign n3782 = ( x724 & ~n3779 ) | ( x724 & n3781 ) | ( ~n3779 & n3781 ) ;
  assign n3783 = ( ~x721 & x722 ) | ( ~x721 & x723 ) | ( x722 & x723 ) ;
  assign n3784 = ( x721 & ~n3780 ) | ( x721 & n3783 ) | ( ~n3780 & n3783 ) ;
  assign n3785 = n3782 & n3784 ;
  assign n3786 = ( n3779 & n3780 ) | ( n3779 & n3785 ) | ( n3780 & n3785 ) ;
  assign n3787 = ( x715 & x716 ) | ( x715 & x717 ) | ( x716 & x717 ) ;
  assign n3788 = ( x718 & x719 ) | ( x718 & x720 ) | ( x719 & x720 ) ;
  assign n3789 = ( ~x718 & x719 ) | ( ~x718 & x720 ) | ( x719 & x720 ) ;
  assign n3790 = ( x718 & ~n3788 ) | ( x718 & n3789 ) | ( ~n3788 & n3789 ) ;
  assign n3791 = ( ~x715 & x716 ) | ( ~x715 & x717 ) | ( x716 & x717 ) ;
  assign n3792 = ( x715 & ~n3787 ) | ( x715 & n3791 ) | ( ~n3787 & n3791 ) ;
  assign n3793 = n3790 & n3792 ;
  assign n3794 = ( n3787 & n3788 ) | ( n3787 & n3793 ) | ( n3788 & n3793 ) ;
  assign n3795 = ( ~n3779 & n3780 ) | ( ~n3779 & n3785 ) | ( n3780 & n3785 ) ;
  assign n3796 = ( n3779 & ~n3786 ) | ( n3779 & n3795 ) | ( ~n3786 & n3795 ) ;
  assign n3797 = ( ~n3787 & n3788 ) | ( ~n3787 & n3793 ) | ( n3788 & n3793 ) ;
  assign n3798 = ( n3787 & ~n3794 ) | ( n3787 & n3797 ) | ( ~n3794 & n3797 ) ;
  assign n3799 = n3782 | n3784 ;
  assign n3800 = ~n3785 & n3799 ;
  assign n3801 = n3790 | n3792 ;
  assign n3802 = ~n3793 & n3801 ;
  assign n3803 = n3800 & n3802 ;
  assign n3804 = ( n3796 & n3798 ) | ( n3796 & n3803 ) | ( n3798 & n3803 ) ;
  assign n3805 = ( n3786 & n3794 ) | ( n3786 & n3804 ) | ( n3794 & n3804 ) ;
  assign n3806 = ( x712 & x713 ) | ( x712 & x714 ) | ( x713 & x714 ) ;
  assign n3807 = ( x709 & x710 ) | ( x709 & x711 ) | ( x710 & x711 ) ;
  assign n3808 = ( ~x712 & x713 ) | ( ~x712 & x714 ) | ( x713 & x714 ) ;
  assign n3809 = ( x712 & ~n3806 ) | ( x712 & n3808 ) | ( ~n3806 & n3808 ) ;
  assign n3810 = ( ~x709 & x710 ) | ( ~x709 & x711 ) | ( x710 & x711 ) ;
  assign n3811 = ( x709 & ~n3807 ) | ( x709 & n3810 ) | ( ~n3807 & n3810 ) ;
  assign n3812 = n3809 & n3811 ;
  assign n3813 = ( n3806 & n3807 ) | ( n3806 & n3812 ) | ( n3807 & n3812 ) ;
  assign n3814 = ( x703 & x704 ) | ( x703 & x705 ) | ( x704 & x705 ) ;
  assign n3815 = ( x706 & x707 ) | ( x706 & x708 ) | ( x707 & x708 ) ;
  assign n3816 = ( ~x706 & x707 ) | ( ~x706 & x708 ) | ( x707 & x708 ) ;
  assign n3817 = ( x706 & ~n3815 ) | ( x706 & n3816 ) | ( ~n3815 & n3816 ) ;
  assign n3818 = ( ~x703 & x704 ) | ( ~x703 & x705 ) | ( x704 & x705 ) ;
  assign n3819 = ( x703 & ~n3814 ) | ( x703 & n3818 ) | ( ~n3814 & n3818 ) ;
  assign n3820 = n3817 & n3819 ;
  assign n3821 = ( n3814 & n3815 ) | ( n3814 & n3820 ) | ( n3815 & n3820 ) ;
  assign n3822 = ( ~n3806 & n3807 ) | ( ~n3806 & n3812 ) | ( n3807 & n3812 ) ;
  assign n3823 = ( n3806 & ~n3813 ) | ( n3806 & n3822 ) | ( ~n3813 & n3822 ) ;
  assign n3824 = ( ~n3814 & n3815 ) | ( ~n3814 & n3820 ) | ( n3815 & n3820 ) ;
  assign n3825 = ( n3814 & ~n3821 ) | ( n3814 & n3824 ) | ( ~n3821 & n3824 ) ;
  assign n3826 = n3817 | n3819 ;
  assign n3827 = ~n3820 & n3826 ;
  assign n3828 = ( n3809 & n3811 ) | ( n3809 & n3827 ) | ( n3811 & n3827 ) ;
  assign n3829 = ~n3812 & n3828 ;
  assign n3830 = ( n3823 & n3825 ) | ( n3823 & n3829 ) | ( n3825 & n3829 ) ;
  assign n3831 = ( n3813 & n3821 ) | ( n3813 & n3830 ) | ( n3821 & n3830 ) ;
  assign n3832 = ( ~n3813 & n3821 ) | ( ~n3813 & n3830 ) | ( n3821 & n3830 ) ;
  assign n3833 = ( n3813 & ~n3831 ) | ( n3813 & n3832 ) | ( ~n3831 & n3832 ) ;
  assign n3834 = ( ~n3786 & n3794 ) | ( ~n3786 & n3804 ) | ( n3794 & n3804 ) ;
  assign n3835 = ( n3786 & ~n3805 ) | ( n3786 & n3834 ) | ( ~n3805 & n3834 ) ;
  assign n3836 = ( ~n3796 & n3798 ) | ( ~n3796 & n3803 ) | ( n3798 & n3803 ) ;
  assign n3837 = ( n3796 & ~n3804 ) | ( n3796 & n3836 ) | ( ~n3804 & n3836 ) ;
  assign n3838 = ( ~n3823 & n3825 ) | ( ~n3823 & n3829 ) | ( n3825 & n3829 ) ;
  assign n3839 = ( n3823 & ~n3830 ) | ( n3823 & n3838 ) | ( ~n3830 & n3838 ) ;
  assign n3840 = ( ~n3809 & n3811 ) | ( ~n3809 & n3827 ) | ( n3811 & n3827 ) ;
  assign n3841 = ( n3809 & ~n3828 ) | ( n3809 & n3840 ) | ( ~n3828 & n3840 ) ;
  assign n3842 = ( n3800 & n3802 ) | ( n3800 & n3841 ) | ( n3802 & n3841 ) ;
  assign n3843 = ~n3803 & n3842 ;
  assign n3844 = ( n3837 & n3839 ) | ( n3837 & n3843 ) | ( n3839 & n3843 ) ;
  assign n3845 = ( n3833 & n3835 ) | ( n3833 & n3844 ) | ( n3835 & n3844 ) ;
  assign n3846 = ( n3805 & n3831 ) | ( n3805 & n3845 ) | ( n3831 & n3845 ) ;
  assign n3847 = ( ~n3737 & n3763 ) | ( ~n3737 & n3777 ) | ( n3763 & n3777 ) ;
  assign n3848 = ( n3737 & ~n3778 ) | ( n3737 & n3847 ) | ( ~n3778 & n3847 ) ;
  assign n3849 = ( ~n3805 & n3831 ) | ( ~n3805 & n3845 ) | ( n3831 & n3845 ) ;
  assign n3850 = ( n3805 & ~n3846 ) | ( n3805 & n3849 ) | ( ~n3846 & n3849 ) ;
  assign n3851 = ( ~n3833 & n3835 ) | ( ~n3833 & n3844 ) | ( n3835 & n3844 ) ;
  assign n3852 = ( n3833 & ~n3845 ) | ( n3833 & n3851 ) | ( ~n3845 & n3851 ) ;
  assign n3853 = ( ~n3765 & n3767 ) | ( ~n3765 & n3776 ) | ( n3767 & n3776 ) ;
  assign n3854 = ( n3765 & ~n3777 ) | ( n3765 & n3853 ) | ( ~n3777 & n3853 ) ;
  assign n3855 = ( n3769 & n3771 ) | ( n3769 & ~n3775 ) | ( n3771 & ~n3775 ) ;
  assign n3856 = ( n3775 & ~n3776 ) | ( n3775 & n3855 ) | ( ~n3776 & n3855 ) ;
  assign n3857 = ( n3837 & n3839 ) | ( n3837 & ~n3843 ) | ( n3839 & ~n3843 ) ;
  assign n3858 = ( n3843 & ~n3844 ) | ( n3843 & n3857 ) | ( ~n3844 & n3857 ) ;
  assign n3859 = ( ~n3732 & n3734 ) | ( ~n3732 & n3773 ) | ( n3734 & n3773 ) ;
  assign n3860 = ( n3732 & ~n3774 ) | ( n3732 & n3859 ) | ( ~n3774 & n3859 ) ;
  assign n3861 = ( ~n3800 & n3802 ) | ( ~n3800 & n3841 ) | ( n3802 & n3841 ) ;
  assign n3862 = ( n3800 & ~n3842 ) | ( n3800 & n3861 ) | ( ~n3842 & n3861 ) ;
  assign n3863 = n3860 & n3862 ;
  assign n3864 = ( n3856 & n3858 ) | ( n3856 & n3863 ) | ( n3858 & n3863 ) ;
  assign n3865 = ( n3852 & n3854 ) | ( n3852 & n3864 ) | ( n3854 & n3864 ) ;
  assign n3866 = ( n3848 & n3850 ) | ( n3848 & n3865 ) | ( n3850 & n3865 ) ;
  assign n3867 = ( n3778 & n3846 ) | ( n3778 & n3866 ) | ( n3846 & n3866 ) ;
  assign n3868 = ( x700 & x701 ) | ( x700 & x702 ) | ( x701 & x702 ) ;
  assign n3869 = ( x697 & x698 ) | ( x697 & x699 ) | ( x698 & x699 ) ;
  assign n3870 = ( ~x700 & x701 ) | ( ~x700 & x702 ) | ( x701 & x702 ) ;
  assign n3871 = ( x700 & ~n3868 ) | ( x700 & n3870 ) | ( ~n3868 & n3870 ) ;
  assign n3872 = ( ~x697 & x698 ) | ( ~x697 & x699 ) | ( x698 & x699 ) ;
  assign n3873 = ( x697 & ~n3869 ) | ( x697 & n3872 ) | ( ~n3869 & n3872 ) ;
  assign n3874 = n3871 & n3873 ;
  assign n3875 = ( n3868 & n3869 ) | ( n3868 & n3874 ) | ( n3869 & n3874 ) ;
  assign n3876 = ( x691 & x692 ) | ( x691 & x693 ) | ( x692 & x693 ) ;
  assign n3877 = ( x694 & x695 ) | ( x694 & x696 ) | ( x695 & x696 ) ;
  assign n3878 = ( ~x694 & x695 ) | ( ~x694 & x696 ) | ( x695 & x696 ) ;
  assign n3879 = ( x694 & ~n3877 ) | ( x694 & n3878 ) | ( ~n3877 & n3878 ) ;
  assign n3880 = ( ~x691 & x692 ) | ( ~x691 & x693 ) | ( x692 & x693 ) ;
  assign n3881 = ( x691 & ~n3876 ) | ( x691 & n3880 ) | ( ~n3876 & n3880 ) ;
  assign n3882 = n3879 & n3881 ;
  assign n3883 = ( n3876 & n3877 ) | ( n3876 & n3882 ) | ( n3877 & n3882 ) ;
  assign n3884 = ( ~n3868 & n3869 ) | ( ~n3868 & n3874 ) | ( n3869 & n3874 ) ;
  assign n3885 = ( n3868 & ~n3875 ) | ( n3868 & n3884 ) | ( ~n3875 & n3884 ) ;
  assign n3886 = ( ~n3876 & n3877 ) | ( ~n3876 & n3882 ) | ( n3877 & n3882 ) ;
  assign n3887 = ( n3876 & ~n3883 ) | ( n3876 & n3886 ) | ( ~n3883 & n3886 ) ;
  assign n3888 = n3871 | n3873 ;
  assign n3889 = ~n3874 & n3888 ;
  assign n3890 = n3879 | n3881 ;
  assign n3891 = ~n3882 & n3890 ;
  assign n3892 = n3889 & n3891 ;
  assign n3893 = ( n3885 & n3887 ) | ( n3885 & n3892 ) | ( n3887 & n3892 ) ;
  assign n3894 = ( n3875 & n3883 ) | ( n3875 & n3893 ) | ( n3883 & n3893 ) ;
  assign n3895 = ( x688 & x689 ) | ( x688 & x690 ) | ( x689 & x690 ) ;
  assign n3896 = ( x685 & x686 ) | ( x685 & x687 ) | ( x686 & x687 ) ;
  assign n3897 = ( ~x688 & x689 ) | ( ~x688 & x690 ) | ( x689 & x690 ) ;
  assign n3898 = ( x688 & ~n3895 ) | ( x688 & n3897 ) | ( ~n3895 & n3897 ) ;
  assign n3899 = ( ~x685 & x686 ) | ( ~x685 & x687 ) | ( x686 & x687 ) ;
  assign n3900 = ( x685 & ~n3896 ) | ( x685 & n3899 ) | ( ~n3896 & n3899 ) ;
  assign n3901 = n3898 & n3900 ;
  assign n3902 = ( n3895 & n3896 ) | ( n3895 & n3901 ) | ( n3896 & n3901 ) ;
  assign n3903 = ( x679 & x680 ) | ( x679 & x681 ) | ( x680 & x681 ) ;
  assign n3904 = ( x682 & x683 ) | ( x682 & x684 ) | ( x683 & x684 ) ;
  assign n3905 = ( ~x682 & x683 ) | ( ~x682 & x684 ) | ( x683 & x684 ) ;
  assign n3906 = ( x682 & ~n3904 ) | ( x682 & n3905 ) | ( ~n3904 & n3905 ) ;
  assign n3907 = ( ~x679 & x680 ) | ( ~x679 & x681 ) | ( x680 & x681 ) ;
  assign n3908 = ( x679 & ~n3903 ) | ( x679 & n3907 ) | ( ~n3903 & n3907 ) ;
  assign n3909 = n3906 & n3908 ;
  assign n3910 = ( n3903 & n3904 ) | ( n3903 & n3909 ) | ( n3904 & n3909 ) ;
  assign n3911 = ( ~n3895 & n3896 ) | ( ~n3895 & n3901 ) | ( n3896 & n3901 ) ;
  assign n3912 = ( n3895 & ~n3902 ) | ( n3895 & n3911 ) | ( ~n3902 & n3911 ) ;
  assign n3913 = ( ~n3903 & n3904 ) | ( ~n3903 & n3909 ) | ( n3904 & n3909 ) ;
  assign n3914 = ( n3903 & ~n3910 ) | ( n3903 & n3913 ) | ( ~n3910 & n3913 ) ;
  assign n3915 = n3906 | n3908 ;
  assign n3916 = ~n3909 & n3915 ;
  assign n3917 = ( n3898 & n3900 ) | ( n3898 & n3916 ) | ( n3900 & n3916 ) ;
  assign n3918 = ~n3901 & n3917 ;
  assign n3919 = ( n3912 & n3914 ) | ( n3912 & n3918 ) | ( n3914 & n3918 ) ;
  assign n3920 = ( n3902 & n3910 ) | ( n3902 & n3919 ) | ( n3910 & n3919 ) ;
  assign n3921 = ( ~n3902 & n3910 ) | ( ~n3902 & n3919 ) | ( n3910 & n3919 ) ;
  assign n3922 = ( n3902 & ~n3920 ) | ( n3902 & n3921 ) | ( ~n3920 & n3921 ) ;
  assign n3923 = ( ~n3875 & n3883 ) | ( ~n3875 & n3893 ) | ( n3883 & n3893 ) ;
  assign n3924 = ( n3875 & ~n3894 ) | ( n3875 & n3923 ) | ( ~n3894 & n3923 ) ;
  assign n3925 = ( ~n3885 & n3887 ) | ( ~n3885 & n3892 ) | ( n3887 & n3892 ) ;
  assign n3926 = ( n3885 & ~n3893 ) | ( n3885 & n3925 ) | ( ~n3893 & n3925 ) ;
  assign n3927 = ( ~n3912 & n3914 ) | ( ~n3912 & n3918 ) | ( n3914 & n3918 ) ;
  assign n3928 = ( n3912 & ~n3919 ) | ( n3912 & n3927 ) | ( ~n3919 & n3927 ) ;
  assign n3929 = ( ~n3898 & n3900 ) | ( ~n3898 & n3916 ) | ( n3900 & n3916 ) ;
  assign n3930 = ( n3898 & ~n3917 ) | ( n3898 & n3929 ) | ( ~n3917 & n3929 ) ;
  assign n3931 = ( n3889 & n3891 ) | ( n3889 & n3930 ) | ( n3891 & n3930 ) ;
  assign n3932 = ~n3892 & n3931 ;
  assign n3933 = ( n3926 & n3928 ) | ( n3926 & n3932 ) | ( n3928 & n3932 ) ;
  assign n3934 = ( n3922 & n3924 ) | ( n3922 & n3933 ) | ( n3924 & n3933 ) ;
  assign n3935 = ( n3894 & n3920 ) | ( n3894 & n3934 ) | ( n3920 & n3934 ) ;
  assign n3936 = ( x676 & x677 ) | ( x676 & x678 ) | ( x677 & x678 ) ;
  assign n3937 = ( x673 & x674 ) | ( x673 & x675 ) | ( x674 & x675 ) ;
  assign n3938 = ( ~x676 & x677 ) | ( ~x676 & x678 ) | ( x677 & x678 ) ;
  assign n3939 = ( x676 & ~n3936 ) | ( x676 & n3938 ) | ( ~n3936 & n3938 ) ;
  assign n3940 = ( ~x673 & x674 ) | ( ~x673 & x675 ) | ( x674 & x675 ) ;
  assign n3941 = ( x673 & ~n3937 ) | ( x673 & n3940 ) | ( ~n3937 & n3940 ) ;
  assign n3942 = n3939 & n3941 ;
  assign n3943 = ( n3936 & n3937 ) | ( n3936 & n3942 ) | ( n3937 & n3942 ) ;
  assign n3944 = ( x667 & x668 ) | ( x667 & x669 ) | ( x668 & x669 ) ;
  assign n3945 = ( x670 & x671 ) | ( x670 & x672 ) | ( x671 & x672 ) ;
  assign n3946 = ( ~x670 & x671 ) | ( ~x670 & x672 ) | ( x671 & x672 ) ;
  assign n3947 = ( x670 & ~n3945 ) | ( x670 & n3946 ) | ( ~n3945 & n3946 ) ;
  assign n3948 = ( ~x667 & x668 ) | ( ~x667 & x669 ) | ( x668 & x669 ) ;
  assign n3949 = ( x667 & ~n3944 ) | ( x667 & n3948 ) | ( ~n3944 & n3948 ) ;
  assign n3950 = n3947 & n3949 ;
  assign n3951 = ( n3944 & n3945 ) | ( n3944 & n3950 ) | ( n3945 & n3950 ) ;
  assign n3952 = ( ~n3936 & n3937 ) | ( ~n3936 & n3942 ) | ( n3937 & n3942 ) ;
  assign n3953 = ( n3936 & ~n3943 ) | ( n3936 & n3952 ) | ( ~n3943 & n3952 ) ;
  assign n3954 = ( ~n3944 & n3945 ) | ( ~n3944 & n3950 ) | ( n3945 & n3950 ) ;
  assign n3955 = ( n3944 & ~n3951 ) | ( n3944 & n3954 ) | ( ~n3951 & n3954 ) ;
  assign n3956 = n3939 | n3941 ;
  assign n3957 = ~n3942 & n3956 ;
  assign n3958 = n3947 | n3949 ;
  assign n3959 = ~n3950 & n3958 ;
  assign n3960 = n3957 & n3959 ;
  assign n3961 = ( n3953 & n3955 ) | ( n3953 & n3960 ) | ( n3955 & n3960 ) ;
  assign n3962 = ( n3943 & n3951 ) | ( n3943 & n3961 ) | ( n3951 & n3961 ) ;
  assign n3963 = ( x664 & x665 ) | ( x664 & x666 ) | ( x665 & x666 ) ;
  assign n3964 = ( x661 & x662 ) | ( x661 & x663 ) | ( x662 & x663 ) ;
  assign n3965 = ( ~x664 & x665 ) | ( ~x664 & x666 ) | ( x665 & x666 ) ;
  assign n3966 = ( x664 & ~n3963 ) | ( x664 & n3965 ) | ( ~n3963 & n3965 ) ;
  assign n3967 = ( ~x661 & x662 ) | ( ~x661 & x663 ) | ( x662 & x663 ) ;
  assign n3968 = ( x661 & ~n3964 ) | ( x661 & n3967 ) | ( ~n3964 & n3967 ) ;
  assign n3969 = n3966 & n3968 ;
  assign n3970 = ( n3963 & n3964 ) | ( n3963 & n3969 ) | ( n3964 & n3969 ) ;
  assign n3971 = ( x655 & x656 ) | ( x655 & x657 ) | ( x656 & x657 ) ;
  assign n3972 = ( x658 & x659 ) | ( x658 & x660 ) | ( x659 & x660 ) ;
  assign n3973 = ( ~x658 & x659 ) | ( ~x658 & x660 ) | ( x659 & x660 ) ;
  assign n3974 = ( x658 & ~n3972 ) | ( x658 & n3973 ) | ( ~n3972 & n3973 ) ;
  assign n3975 = ( ~x655 & x656 ) | ( ~x655 & x657 ) | ( x656 & x657 ) ;
  assign n3976 = ( x655 & ~n3971 ) | ( x655 & n3975 ) | ( ~n3971 & n3975 ) ;
  assign n3977 = n3974 & n3976 ;
  assign n3978 = ( n3971 & n3972 ) | ( n3971 & n3977 ) | ( n3972 & n3977 ) ;
  assign n3979 = ( ~n3963 & n3964 ) | ( ~n3963 & n3969 ) | ( n3964 & n3969 ) ;
  assign n3980 = ( n3963 & ~n3970 ) | ( n3963 & n3979 ) | ( ~n3970 & n3979 ) ;
  assign n3981 = ( ~n3971 & n3972 ) | ( ~n3971 & n3977 ) | ( n3972 & n3977 ) ;
  assign n3982 = ( n3971 & ~n3978 ) | ( n3971 & n3981 ) | ( ~n3978 & n3981 ) ;
  assign n3983 = n3974 | n3976 ;
  assign n3984 = ~n3977 & n3983 ;
  assign n3985 = ( n3966 & n3968 ) | ( n3966 & n3984 ) | ( n3968 & n3984 ) ;
  assign n3986 = ~n3969 & n3985 ;
  assign n3987 = ( n3980 & n3982 ) | ( n3980 & n3986 ) | ( n3982 & n3986 ) ;
  assign n3988 = ( n3970 & n3978 ) | ( n3970 & n3987 ) | ( n3978 & n3987 ) ;
  assign n3989 = ( ~n3970 & n3978 ) | ( ~n3970 & n3987 ) | ( n3978 & n3987 ) ;
  assign n3990 = ( n3970 & ~n3988 ) | ( n3970 & n3989 ) | ( ~n3988 & n3989 ) ;
  assign n3991 = ( ~n3943 & n3951 ) | ( ~n3943 & n3961 ) | ( n3951 & n3961 ) ;
  assign n3992 = ( n3943 & ~n3962 ) | ( n3943 & n3991 ) | ( ~n3962 & n3991 ) ;
  assign n3993 = ( ~n3953 & n3955 ) | ( ~n3953 & n3960 ) | ( n3955 & n3960 ) ;
  assign n3994 = ( n3953 & ~n3961 ) | ( n3953 & n3993 ) | ( ~n3961 & n3993 ) ;
  assign n3995 = ( ~n3980 & n3982 ) | ( ~n3980 & n3986 ) | ( n3982 & n3986 ) ;
  assign n3996 = ( n3980 & ~n3987 ) | ( n3980 & n3995 ) | ( ~n3987 & n3995 ) ;
  assign n3997 = ( ~n3966 & n3968 ) | ( ~n3966 & n3984 ) | ( n3968 & n3984 ) ;
  assign n3998 = ( n3966 & ~n3985 ) | ( n3966 & n3997 ) | ( ~n3985 & n3997 ) ;
  assign n3999 = ( n3957 & n3959 ) | ( n3957 & n3998 ) | ( n3959 & n3998 ) ;
  assign n4000 = ~n3960 & n3999 ;
  assign n4001 = ( n3994 & n3996 ) | ( n3994 & n4000 ) | ( n3996 & n4000 ) ;
  assign n4002 = ( n3990 & n3992 ) | ( n3990 & n4001 ) | ( n3992 & n4001 ) ;
  assign n4003 = ( n3962 & n3988 ) | ( n3962 & n4002 ) | ( n3988 & n4002 ) ;
  assign n4004 = ( ~n3894 & n3920 ) | ( ~n3894 & n3934 ) | ( n3920 & n3934 ) ;
  assign n4005 = ( n3894 & ~n3935 ) | ( n3894 & n4004 ) | ( ~n3935 & n4004 ) ;
  assign n4006 = ( ~n3962 & n3988 ) | ( ~n3962 & n4002 ) | ( n3988 & n4002 ) ;
  assign n4007 = ( n3962 & ~n4003 ) | ( n3962 & n4006 ) | ( ~n4003 & n4006 ) ;
  assign n4008 = ( ~n3990 & n3992 ) | ( ~n3990 & n4001 ) | ( n3992 & n4001 ) ;
  assign n4009 = ( n3990 & ~n4002 ) | ( n3990 & n4008 ) | ( ~n4002 & n4008 ) ;
  assign n4010 = ( ~n3922 & n3924 ) | ( ~n3922 & n3933 ) | ( n3924 & n3933 ) ;
  assign n4011 = ( n3922 & ~n3934 ) | ( n3922 & n4010 ) | ( ~n3934 & n4010 ) ;
  assign n4012 = ( n3926 & n3928 ) | ( n3926 & ~n3932 ) | ( n3928 & ~n3932 ) ;
  assign n4013 = ( n3932 & ~n3933 ) | ( n3932 & n4012 ) | ( ~n3933 & n4012 ) ;
  assign n4014 = ( n3994 & n3996 ) | ( n3994 & ~n4000 ) | ( n3996 & ~n4000 ) ;
  assign n4015 = ( n4000 & ~n4001 ) | ( n4000 & n4014 ) | ( ~n4001 & n4014 ) ;
  assign n4016 = ( ~n3889 & n3891 ) | ( ~n3889 & n3930 ) | ( n3891 & n3930 ) ;
  assign n4017 = ( n3889 & ~n3931 ) | ( n3889 & n4016 ) | ( ~n3931 & n4016 ) ;
  assign n4018 = ( ~n3957 & n3959 ) | ( ~n3957 & n3998 ) | ( n3959 & n3998 ) ;
  assign n4019 = ( n3957 & ~n3999 ) | ( n3957 & n4018 ) | ( ~n3999 & n4018 ) ;
  assign n4020 = n4017 & n4019 ;
  assign n4021 = ( n4013 & n4015 ) | ( n4013 & n4020 ) | ( n4015 & n4020 ) ;
  assign n4022 = ( n4009 & n4011 ) | ( n4009 & n4021 ) | ( n4011 & n4021 ) ;
  assign n4023 = ( n4005 & n4007 ) | ( n4005 & n4022 ) | ( n4007 & n4022 ) ;
  assign n4024 = ( n3935 & n4003 ) | ( n3935 & n4023 ) | ( n4003 & n4023 ) ;
  assign n4025 = ( ~n3935 & n4003 ) | ( ~n3935 & n4023 ) | ( n4003 & n4023 ) ;
  assign n4026 = ( n3935 & ~n4024 ) | ( n3935 & n4025 ) | ( ~n4024 & n4025 ) ;
  assign n4027 = ( ~n3778 & n3846 ) | ( ~n3778 & n3866 ) | ( n3846 & n3866 ) ;
  assign n4028 = ( n3778 & ~n3867 ) | ( n3778 & n4027 ) | ( ~n3867 & n4027 ) ;
  assign n4029 = ( ~n3848 & n3850 ) | ( ~n3848 & n3865 ) | ( n3850 & n3865 ) ;
  assign n4030 = ( n3848 & ~n3866 ) | ( n3848 & n4029 ) | ( ~n3866 & n4029 ) ;
  assign n4031 = ( ~n4005 & n4007 ) | ( ~n4005 & n4022 ) | ( n4007 & n4022 ) ;
  assign n4032 = ( n4005 & ~n4023 ) | ( n4005 & n4031 ) | ( ~n4023 & n4031 ) ;
  assign n4033 = ( ~n4009 & n4011 ) | ( ~n4009 & n4021 ) | ( n4011 & n4021 ) ;
  assign n4034 = ( n4009 & ~n4022 ) | ( n4009 & n4033 ) | ( ~n4022 & n4033 ) ;
  assign n4035 = ( ~n3852 & n3854 ) | ( ~n3852 & n3864 ) | ( n3854 & n3864 ) ;
  assign n4036 = ( n3852 & ~n3865 ) | ( n3852 & n4035 ) | ( ~n3865 & n4035 ) ;
  assign n4037 = ( ~n3856 & n3858 ) | ( ~n3856 & n3863 ) | ( n3858 & n3863 ) ;
  assign n4038 = ( n3856 & ~n3864 ) | ( n3856 & n4037 ) | ( ~n3864 & n4037 ) ;
  assign n4039 = ( ~n4013 & n4015 ) | ( ~n4013 & n4020 ) | ( n4015 & n4020 ) ;
  assign n4040 = ( n4013 & ~n4021 ) | ( n4013 & n4039 ) | ( ~n4021 & n4039 ) ;
  assign n4041 = n4017 | n4019 ;
  assign n4042 = ~n4020 & n4041 ;
  assign n4043 = ( n3860 & n3862 ) | ( n3860 & n4042 ) | ( n3862 & n4042 ) ;
  assign n4044 = ~n3863 & n4043 ;
  assign n4045 = ( n4038 & n4040 ) | ( n4038 & n4044 ) | ( n4040 & n4044 ) ;
  assign n4046 = ( n4034 & n4036 ) | ( n4034 & n4045 ) | ( n4036 & n4045 ) ;
  assign n4047 = ( n4030 & n4032 ) | ( n4030 & n4046 ) | ( n4032 & n4046 ) ;
  assign n4048 = ( n4026 & n4028 ) | ( n4026 & n4047 ) | ( n4028 & n4047 ) ;
  assign n4049 = ( n3867 & n4024 ) | ( n3867 & n4048 ) | ( n4024 & n4048 ) ;
  assign n4050 = ( ~n3528 & n3685 ) | ( ~n3528 & n3709 ) | ( n3685 & n3709 ) ;
  assign n4051 = ( n3528 & ~n3710 ) | ( n3528 & n4050 ) | ( ~n3710 & n4050 ) ;
  assign n4052 = ( ~n3867 & n4024 ) | ( ~n3867 & n4048 ) | ( n4024 & n4048 ) ;
  assign n4053 = ( n3867 & ~n4049 ) | ( n3867 & n4052 ) | ( ~n4049 & n4052 ) ;
  assign n4054 = ( ~n4026 & n4028 ) | ( ~n4026 & n4047 ) | ( n4028 & n4047 ) ;
  assign n4055 = ( n4026 & ~n4048 ) | ( n4026 & n4054 ) | ( ~n4048 & n4054 ) ;
  assign n4056 = ( ~n3687 & n3689 ) | ( ~n3687 & n3708 ) | ( n3689 & n3708 ) ;
  assign n4057 = ( n3687 & ~n3709 ) | ( n3687 & n4056 ) | ( ~n3709 & n4056 ) ;
  assign n4058 = ( ~n3691 & n3693 ) | ( ~n3691 & n3707 ) | ( n3693 & n3707 ) ;
  assign n4059 = ( n3691 & ~n3708 ) | ( n3691 & n4058 ) | ( ~n3708 & n4058 ) ;
  assign n4060 = ( ~n4030 & n4032 ) | ( ~n4030 & n4046 ) | ( n4032 & n4046 ) ;
  assign n4061 = ( n4030 & ~n4047 ) | ( n4030 & n4060 ) | ( ~n4047 & n4060 ) ;
  assign n4062 = ( ~n4034 & n4036 ) | ( ~n4034 & n4045 ) | ( n4036 & n4045 ) ;
  assign n4063 = ( n4034 & ~n4046 ) | ( n4034 & n4062 ) | ( ~n4046 & n4062 ) ;
  assign n4064 = ( ~n3695 & n3697 ) | ( ~n3695 & n3706 ) | ( n3697 & n3706 ) ;
  assign n4065 = ( n3695 & ~n3707 ) | ( n3695 & n4064 ) | ( ~n3707 & n4064 ) ;
  assign n4066 = ( n3699 & n3701 ) | ( n3699 & ~n3705 ) | ( n3701 & ~n3705 ) ;
  assign n4067 = ( n3705 & ~n3706 ) | ( n3705 & n4066 ) | ( ~n3706 & n4066 ) ;
  assign n4068 = ( n4038 & n4040 ) | ( n4038 & ~n4044 ) | ( n4040 & ~n4044 ) ;
  assign n4069 = ( n4044 & ~n4045 ) | ( n4044 & n4068 ) | ( ~n4045 & n4068 ) ;
  assign n4070 = ( ~n3521 & n3523 ) | ( ~n3521 & n3703 ) | ( n3523 & n3703 ) ;
  assign n4071 = ( n3521 & ~n3704 ) | ( n3521 & n4070 ) | ( ~n3704 & n4070 ) ;
  assign n4072 = ( ~n3860 & n3862 ) | ( ~n3860 & n4042 ) | ( n3862 & n4042 ) ;
  assign n4073 = ( n3860 & ~n4043 ) | ( n3860 & n4072 ) | ( ~n4043 & n4072 ) ;
  assign n4074 = n4071 & n4073 ;
  assign n4075 = ( n4067 & n4069 ) | ( n4067 & n4074 ) | ( n4069 & n4074 ) ;
  assign n4076 = ( n4063 & n4065 ) | ( n4063 & n4075 ) | ( n4065 & n4075 ) ;
  assign n4077 = ( n4059 & n4061 ) | ( n4059 & n4076 ) | ( n4061 & n4076 ) ;
  assign n4078 = ( n4055 & n4057 ) | ( n4055 & n4077 ) | ( n4057 & n4077 ) ;
  assign n4079 = ( n4051 & n4053 ) | ( n4051 & n4078 ) | ( n4053 & n4078 ) ;
  assign n4080 = ( n3710 & n4049 ) | ( n3710 & n4079 ) | ( n4049 & n4079 ) ;
  assign n4081 = ( x652 & x653 ) | ( x652 & x654 ) | ( x653 & x654 ) ;
  assign n4082 = ( x649 & x650 ) | ( x649 & x651 ) | ( x650 & x651 ) ;
  assign n4083 = ( ~x652 & x653 ) | ( ~x652 & x654 ) | ( x653 & x654 ) ;
  assign n4084 = ( x652 & ~n4081 ) | ( x652 & n4083 ) | ( ~n4081 & n4083 ) ;
  assign n4085 = ( ~x649 & x650 ) | ( ~x649 & x651 ) | ( x650 & x651 ) ;
  assign n4086 = ( x649 & ~n4082 ) | ( x649 & n4085 ) | ( ~n4082 & n4085 ) ;
  assign n4087 = n4084 & n4086 ;
  assign n4088 = ( n4081 & n4082 ) | ( n4081 & n4087 ) | ( n4082 & n4087 ) ;
  assign n4089 = ( x643 & x644 ) | ( x643 & x645 ) | ( x644 & x645 ) ;
  assign n4090 = ( x646 & x647 ) | ( x646 & x648 ) | ( x647 & x648 ) ;
  assign n4091 = ( ~x646 & x647 ) | ( ~x646 & x648 ) | ( x647 & x648 ) ;
  assign n4092 = ( x646 & ~n4090 ) | ( x646 & n4091 ) | ( ~n4090 & n4091 ) ;
  assign n4093 = ( ~x643 & x644 ) | ( ~x643 & x645 ) | ( x644 & x645 ) ;
  assign n4094 = ( x643 & ~n4089 ) | ( x643 & n4093 ) | ( ~n4089 & n4093 ) ;
  assign n4095 = n4092 & n4094 ;
  assign n4096 = ( n4089 & n4090 ) | ( n4089 & n4095 ) | ( n4090 & n4095 ) ;
  assign n4097 = ( ~n4081 & n4082 ) | ( ~n4081 & n4087 ) | ( n4082 & n4087 ) ;
  assign n4098 = ( n4081 & ~n4088 ) | ( n4081 & n4097 ) | ( ~n4088 & n4097 ) ;
  assign n4099 = ( ~n4089 & n4090 ) | ( ~n4089 & n4095 ) | ( n4090 & n4095 ) ;
  assign n4100 = ( n4089 & ~n4096 ) | ( n4089 & n4099 ) | ( ~n4096 & n4099 ) ;
  assign n4101 = n4084 | n4086 ;
  assign n4102 = ~n4087 & n4101 ;
  assign n4103 = n4092 | n4094 ;
  assign n4104 = ~n4095 & n4103 ;
  assign n4105 = n4102 & n4104 ;
  assign n4106 = ( n4098 & n4100 ) | ( n4098 & n4105 ) | ( n4100 & n4105 ) ;
  assign n4107 = ( n4088 & n4096 ) | ( n4088 & n4106 ) | ( n4096 & n4106 ) ;
  assign n4108 = ( x640 & x641 ) | ( x640 & x642 ) | ( x641 & x642 ) ;
  assign n4109 = ( x637 & x638 ) | ( x637 & x639 ) | ( x638 & x639 ) ;
  assign n4110 = ( ~x640 & x641 ) | ( ~x640 & x642 ) | ( x641 & x642 ) ;
  assign n4111 = ( x640 & ~n4108 ) | ( x640 & n4110 ) | ( ~n4108 & n4110 ) ;
  assign n4112 = ( ~x637 & x638 ) | ( ~x637 & x639 ) | ( x638 & x639 ) ;
  assign n4113 = ( x637 & ~n4109 ) | ( x637 & n4112 ) | ( ~n4109 & n4112 ) ;
  assign n4114 = n4111 & n4113 ;
  assign n4115 = ( n4108 & n4109 ) | ( n4108 & n4114 ) | ( n4109 & n4114 ) ;
  assign n4116 = ( x631 & x632 ) | ( x631 & x633 ) | ( x632 & x633 ) ;
  assign n4117 = ( x634 & x635 ) | ( x634 & x636 ) | ( x635 & x636 ) ;
  assign n4118 = ( ~x634 & x635 ) | ( ~x634 & x636 ) | ( x635 & x636 ) ;
  assign n4119 = ( x634 & ~n4117 ) | ( x634 & n4118 ) | ( ~n4117 & n4118 ) ;
  assign n4120 = ( ~x631 & x632 ) | ( ~x631 & x633 ) | ( x632 & x633 ) ;
  assign n4121 = ( x631 & ~n4116 ) | ( x631 & n4120 ) | ( ~n4116 & n4120 ) ;
  assign n4122 = n4119 & n4121 ;
  assign n4123 = ( n4116 & n4117 ) | ( n4116 & n4122 ) | ( n4117 & n4122 ) ;
  assign n4124 = ( ~n4108 & n4109 ) | ( ~n4108 & n4114 ) | ( n4109 & n4114 ) ;
  assign n4125 = ( n4108 & ~n4115 ) | ( n4108 & n4124 ) | ( ~n4115 & n4124 ) ;
  assign n4126 = ( ~n4116 & n4117 ) | ( ~n4116 & n4122 ) | ( n4117 & n4122 ) ;
  assign n4127 = ( n4116 & ~n4123 ) | ( n4116 & n4126 ) | ( ~n4123 & n4126 ) ;
  assign n4128 = n4119 | n4121 ;
  assign n4129 = ~n4122 & n4128 ;
  assign n4130 = ( n4111 & n4113 ) | ( n4111 & n4129 ) | ( n4113 & n4129 ) ;
  assign n4131 = ~n4114 & n4130 ;
  assign n4132 = ( n4125 & n4127 ) | ( n4125 & n4131 ) | ( n4127 & n4131 ) ;
  assign n4133 = ( n4115 & n4123 ) | ( n4115 & n4132 ) | ( n4123 & n4132 ) ;
  assign n4134 = ( ~n4115 & n4123 ) | ( ~n4115 & n4132 ) | ( n4123 & n4132 ) ;
  assign n4135 = ( n4115 & ~n4133 ) | ( n4115 & n4134 ) | ( ~n4133 & n4134 ) ;
  assign n4136 = ( ~n4088 & n4096 ) | ( ~n4088 & n4106 ) | ( n4096 & n4106 ) ;
  assign n4137 = ( n4088 & ~n4107 ) | ( n4088 & n4136 ) | ( ~n4107 & n4136 ) ;
  assign n4138 = ( ~n4098 & n4100 ) | ( ~n4098 & n4105 ) | ( n4100 & n4105 ) ;
  assign n4139 = ( n4098 & ~n4106 ) | ( n4098 & n4138 ) | ( ~n4106 & n4138 ) ;
  assign n4140 = ( ~n4125 & n4127 ) | ( ~n4125 & n4131 ) | ( n4127 & n4131 ) ;
  assign n4141 = ( n4125 & ~n4132 ) | ( n4125 & n4140 ) | ( ~n4132 & n4140 ) ;
  assign n4142 = ( ~n4111 & n4113 ) | ( ~n4111 & n4129 ) | ( n4113 & n4129 ) ;
  assign n4143 = ( n4111 & ~n4130 ) | ( n4111 & n4142 ) | ( ~n4130 & n4142 ) ;
  assign n4144 = ( n4102 & n4104 ) | ( n4102 & n4143 ) | ( n4104 & n4143 ) ;
  assign n4145 = ~n4105 & n4144 ;
  assign n4146 = ( n4139 & n4141 ) | ( n4139 & n4145 ) | ( n4141 & n4145 ) ;
  assign n4147 = ( n4135 & n4137 ) | ( n4135 & n4146 ) | ( n4137 & n4146 ) ;
  assign n4148 = ( n4107 & n4133 ) | ( n4107 & n4147 ) | ( n4133 & n4147 ) ;
  assign n4149 = ( x628 & x629 ) | ( x628 & x630 ) | ( x629 & x630 ) ;
  assign n4150 = ( x625 & x626 ) | ( x625 & x627 ) | ( x626 & x627 ) ;
  assign n4151 = ( ~x628 & x629 ) | ( ~x628 & x630 ) | ( x629 & x630 ) ;
  assign n4152 = ( x628 & ~n4149 ) | ( x628 & n4151 ) | ( ~n4149 & n4151 ) ;
  assign n4153 = ( ~x625 & x626 ) | ( ~x625 & x627 ) | ( x626 & x627 ) ;
  assign n4154 = ( x625 & ~n4150 ) | ( x625 & n4153 ) | ( ~n4150 & n4153 ) ;
  assign n4155 = n4152 & n4154 ;
  assign n4156 = ( n4149 & n4150 ) | ( n4149 & n4155 ) | ( n4150 & n4155 ) ;
  assign n4157 = ( x619 & x620 ) | ( x619 & x621 ) | ( x620 & x621 ) ;
  assign n4158 = ( x622 & x623 ) | ( x622 & x624 ) | ( x623 & x624 ) ;
  assign n4159 = ( ~x622 & x623 ) | ( ~x622 & x624 ) | ( x623 & x624 ) ;
  assign n4160 = ( x622 & ~n4158 ) | ( x622 & n4159 ) | ( ~n4158 & n4159 ) ;
  assign n4161 = ( ~x619 & x620 ) | ( ~x619 & x621 ) | ( x620 & x621 ) ;
  assign n4162 = ( x619 & ~n4157 ) | ( x619 & n4161 ) | ( ~n4157 & n4161 ) ;
  assign n4163 = n4160 & n4162 ;
  assign n4164 = ( n4157 & n4158 ) | ( n4157 & n4163 ) | ( n4158 & n4163 ) ;
  assign n4165 = ( ~n4149 & n4150 ) | ( ~n4149 & n4155 ) | ( n4150 & n4155 ) ;
  assign n4166 = ( n4149 & ~n4156 ) | ( n4149 & n4165 ) | ( ~n4156 & n4165 ) ;
  assign n4167 = ( ~n4157 & n4158 ) | ( ~n4157 & n4163 ) | ( n4158 & n4163 ) ;
  assign n4168 = ( n4157 & ~n4164 ) | ( n4157 & n4167 ) | ( ~n4164 & n4167 ) ;
  assign n4169 = n4152 | n4154 ;
  assign n4170 = ~n4155 & n4169 ;
  assign n4171 = n4160 | n4162 ;
  assign n4172 = ~n4163 & n4171 ;
  assign n4173 = n4170 & n4172 ;
  assign n4174 = ( n4166 & n4168 ) | ( n4166 & n4173 ) | ( n4168 & n4173 ) ;
  assign n4175 = ( n4156 & n4164 ) | ( n4156 & n4174 ) | ( n4164 & n4174 ) ;
  assign n4176 = ( x616 & x617 ) | ( x616 & x618 ) | ( x617 & x618 ) ;
  assign n4177 = ( x613 & x614 ) | ( x613 & x615 ) | ( x614 & x615 ) ;
  assign n4178 = ( ~x616 & x617 ) | ( ~x616 & x618 ) | ( x617 & x618 ) ;
  assign n4179 = ( x616 & ~n4176 ) | ( x616 & n4178 ) | ( ~n4176 & n4178 ) ;
  assign n4180 = ( ~x613 & x614 ) | ( ~x613 & x615 ) | ( x614 & x615 ) ;
  assign n4181 = ( x613 & ~n4177 ) | ( x613 & n4180 ) | ( ~n4177 & n4180 ) ;
  assign n4182 = n4179 & n4181 ;
  assign n4183 = ( n4176 & n4177 ) | ( n4176 & n4182 ) | ( n4177 & n4182 ) ;
  assign n4184 = ( x607 & x608 ) | ( x607 & x609 ) | ( x608 & x609 ) ;
  assign n4185 = ( x610 & x611 ) | ( x610 & x612 ) | ( x611 & x612 ) ;
  assign n4186 = ( ~x610 & x611 ) | ( ~x610 & x612 ) | ( x611 & x612 ) ;
  assign n4187 = ( x610 & ~n4185 ) | ( x610 & n4186 ) | ( ~n4185 & n4186 ) ;
  assign n4188 = ( ~x607 & x608 ) | ( ~x607 & x609 ) | ( x608 & x609 ) ;
  assign n4189 = ( x607 & ~n4184 ) | ( x607 & n4188 ) | ( ~n4184 & n4188 ) ;
  assign n4190 = n4187 & n4189 ;
  assign n4191 = ( n4184 & n4185 ) | ( n4184 & n4190 ) | ( n4185 & n4190 ) ;
  assign n4192 = ( ~n4176 & n4177 ) | ( ~n4176 & n4182 ) | ( n4177 & n4182 ) ;
  assign n4193 = ( n4176 & ~n4183 ) | ( n4176 & n4192 ) | ( ~n4183 & n4192 ) ;
  assign n4194 = ( ~n4184 & n4185 ) | ( ~n4184 & n4190 ) | ( n4185 & n4190 ) ;
  assign n4195 = ( n4184 & ~n4191 ) | ( n4184 & n4194 ) | ( ~n4191 & n4194 ) ;
  assign n4196 = n4187 | n4189 ;
  assign n4197 = ~n4190 & n4196 ;
  assign n4198 = ( n4179 & n4181 ) | ( n4179 & n4197 ) | ( n4181 & n4197 ) ;
  assign n4199 = ~n4182 & n4198 ;
  assign n4200 = ( n4193 & n4195 ) | ( n4193 & n4199 ) | ( n4195 & n4199 ) ;
  assign n4201 = ( n4183 & n4191 ) | ( n4183 & n4200 ) | ( n4191 & n4200 ) ;
  assign n4202 = ( ~n4183 & n4191 ) | ( ~n4183 & n4200 ) | ( n4191 & n4200 ) ;
  assign n4203 = ( n4183 & ~n4201 ) | ( n4183 & n4202 ) | ( ~n4201 & n4202 ) ;
  assign n4204 = ( ~n4156 & n4164 ) | ( ~n4156 & n4174 ) | ( n4164 & n4174 ) ;
  assign n4205 = ( n4156 & ~n4175 ) | ( n4156 & n4204 ) | ( ~n4175 & n4204 ) ;
  assign n4206 = ( ~n4166 & n4168 ) | ( ~n4166 & n4173 ) | ( n4168 & n4173 ) ;
  assign n4207 = ( n4166 & ~n4174 ) | ( n4166 & n4206 ) | ( ~n4174 & n4206 ) ;
  assign n4208 = ( ~n4193 & n4195 ) | ( ~n4193 & n4199 ) | ( n4195 & n4199 ) ;
  assign n4209 = ( n4193 & ~n4200 ) | ( n4193 & n4208 ) | ( ~n4200 & n4208 ) ;
  assign n4210 = ( ~n4179 & n4181 ) | ( ~n4179 & n4197 ) | ( n4181 & n4197 ) ;
  assign n4211 = ( n4179 & ~n4198 ) | ( n4179 & n4210 ) | ( ~n4198 & n4210 ) ;
  assign n4212 = ( n4170 & n4172 ) | ( n4170 & n4211 ) | ( n4172 & n4211 ) ;
  assign n4213 = ~n4173 & n4212 ;
  assign n4214 = ( n4207 & n4209 ) | ( n4207 & n4213 ) | ( n4209 & n4213 ) ;
  assign n4215 = ( n4203 & n4205 ) | ( n4203 & n4214 ) | ( n4205 & n4214 ) ;
  assign n4216 = ( n4175 & n4201 ) | ( n4175 & n4215 ) | ( n4201 & n4215 ) ;
  assign n4217 = ( ~n4107 & n4133 ) | ( ~n4107 & n4147 ) | ( n4133 & n4147 ) ;
  assign n4218 = ( n4107 & ~n4148 ) | ( n4107 & n4217 ) | ( ~n4148 & n4217 ) ;
  assign n4219 = ( ~n4175 & n4201 ) | ( ~n4175 & n4215 ) | ( n4201 & n4215 ) ;
  assign n4220 = ( n4175 & ~n4216 ) | ( n4175 & n4219 ) | ( ~n4216 & n4219 ) ;
  assign n4221 = ( ~n4203 & n4205 ) | ( ~n4203 & n4214 ) | ( n4205 & n4214 ) ;
  assign n4222 = ( n4203 & ~n4215 ) | ( n4203 & n4221 ) | ( ~n4215 & n4221 ) ;
  assign n4223 = ( ~n4135 & n4137 ) | ( ~n4135 & n4146 ) | ( n4137 & n4146 ) ;
  assign n4224 = ( n4135 & ~n4147 ) | ( n4135 & n4223 ) | ( ~n4147 & n4223 ) ;
  assign n4225 = ( n4139 & n4141 ) | ( n4139 & ~n4145 ) | ( n4141 & ~n4145 ) ;
  assign n4226 = ( n4145 & ~n4146 ) | ( n4145 & n4225 ) | ( ~n4146 & n4225 ) ;
  assign n4227 = ( n4207 & n4209 ) | ( n4207 & ~n4213 ) | ( n4209 & ~n4213 ) ;
  assign n4228 = ( n4213 & ~n4214 ) | ( n4213 & n4227 ) | ( ~n4214 & n4227 ) ;
  assign n4229 = ( ~n4102 & n4104 ) | ( ~n4102 & n4143 ) | ( n4104 & n4143 ) ;
  assign n4230 = ( n4102 & ~n4144 ) | ( n4102 & n4229 ) | ( ~n4144 & n4229 ) ;
  assign n4231 = ( ~n4170 & n4172 ) | ( ~n4170 & n4211 ) | ( n4172 & n4211 ) ;
  assign n4232 = ( n4170 & ~n4212 ) | ( n4170 & n4231 ) | ( ~n4212 & n4231 ) ;
  assign n4233 = n4230 & n4232 ;
  assign n4234 = ( n4226 & n4228 ) | ( n4226 & n4233 ) | ( n4228 & n4233 ) ;
  assign n4235 = ( n4222 & n4224 ) | ( n4222 & n4234 ) | ( n4224 & n4234 ) ;
  assign n4236 = ( n4218 & n4220 ) | ( n4218 & n4235 ) | ( n4220 & n4235 ) ;
  assign n4237 = ( n4148 & n4216 ) | ( n4148 & n4236 ) | ( n4216 & n4236 ) ;
  assign n4238 = ( x604 & x605 ) | ( x604 & x606 ) | ( x605 & x606 ) ;
  assign n4239 = ( x601 & x602 ) | ( x601 & x603 ) | ( x602 & x603 ) ;
  assign n4240 = ( ~x604 & x605 ) | ( ~x604 & x606 ) | ( x605 & x606 ) ;
  assign n4241 = ( x604 & ~n4238 ) | ( x604 & n4240 ) | ( ~n4238 & n4240 ) ;
  assign n4242 = ( ~x601 & x602 ) | ( ~x601 & x603 ) | ( x602 & x603 ) ;
  assign n4243 = ( x601 & ~n4239 ) | ( x601 & n4242 ) | ( ~n4239 & n4242 ) ;
  assign n4244 = n4241 & n4243 ;
  assign n4245 = ( n4238 & n4239 ) | ( n4238 & n4244 ) | ( n4239 & n4244 ) ;
  assign n4246 = ( x595 & x596 ) | ( x595 & x597 ) | ( x596 & x597 ) ;
  assign n4247 = ( x598 & x599 ) | ( x598 & x600 ) | ( x599 & x600 ) ;
  assign n4248 = ( ~x598 & x599 ) | ( ~x598 & x600 ) | ( x599 & x600 ) ;
  assign n4249 = ( x598 & ~n4247 ) | ( x598 & n4248 ) | ( ~n4247 & n4248 ) ;
  assign n4250 = ( ~x595 & x596 ) | ( ~x595 & x597 ) | ( x596 & x597 ) ;
  assign n4251 = ( x595 & ~n4246 ) | ( x595 & n4250 ) | ( ~n4246 & n4250 ) ;
  assign n4252 = n4249 & n4251 ;
  assign n4253 = ( n4246 & n4247 ) | ( n4246 & n4252 ) | ( n4247 & n4252 ) ;
  assign n4254 = ( ~n4238 & n4239 ) | ( ~n4238 & n4244 ) | ( n4239 & n4244 ) ;
  assign n4255 = ( n4238 & ~n4245 ) | ( n4238 & n4254 ) | ( ~n4245 & n4254 ) ;
  assign n4256 = ( ~n4246 & n4247 ) | ( ~n4246 & n4252 ) | ( n4247 & n4252 ) ;
  assign n4257 = ( n4246 & ~n4253 ) | ( n4246 & n4256 ) | ( ~n4253 & n4256 ) ;
  assign n4258 = n4241 | n4243 ;
  assign n4259 = ~n4244 & n4258 ;
  assign n4260 = n4249 | n4251 ;
  assign n4261 = ~n4252 & n4260 ;
  assign n4262 = n4259 & n4261 ;
  assign n4263 = ( n4255 & n4257 ) | ( n4255 & n4262 ) | ( n4257 & n4262 ) ;
  assign n4264 = ( n4245 & n4253 ) | ( n4245 & n4263 ) | ( n4253 & n4263 ) ;
  assign n4265 = ( x592 & x593 ) | ( x592 & x594 ) | ( x593 & x594 ) ;
  assign n4266 = ( x589 & x590 ) | ( x589 & x591 ) | ( x590 & x591 ) ;
  assign n4267 = ( ~x592 & x593 ) | ( ~x592 & x594 ) | ( x593 & x594 ) ;
  assign n4268 = ( x592 & ~n4265 ) | ( x592 & n4267 ) | ( ~n4265 & n4267 ) ;
  assign n4269 = ( ~x589 & x590 ) | ( ~x589 & x591 ) | ( x590 & x591 ) ;
  assign n4270 = ( x589 & ~n4266 ) | ( x589 & n4269 ) | ( ~n4266 & n4269 ) ;
  assign n4271 = n4268 & n4270 ;
  assign n4272 = ( n4265 & n4266 ) | ( n4265 & n4271 ) | ( n4266 & n4271 ) ;
  assign n4273 = ( x583 & x584 ) | ( x583 & x585 ) | ( x584 & x585 ) ;
  assign n4274 = ( x586 & x587 ) | ( x586 & x588 ) | ( x587 & x588 ) ;
  assign n4275 = ( ~x586 & x587 ) | ( ~x586 & x588 ) | ( x587 & x588 ) ;
  assign n4276 = ( x586 & ~n4274 ) | ( x586 & n4275 ) | ( ~n4274 & n4275 ) ;
  assign n4277 = ( ~x583 & x584 ) | ( ~x583 & x585 ) | ( x584 & x585 ) ;
  assign n4278 = ( x583 & ~n4273 ) | ( x583 & n4277 ) | ( ~n4273 & n4277 ) ;
  assign n4279 = n4276 & n4278 ;
  assign n4280 = ( n4273 & n4274 ) | ( n4273 & n4279 ) | ( n4274 & n4279 ) ;
  assign n4281 = ( ~n4265 & n4266 ) | ( ~n4265 & n4271 ) | ( n4266 & n4271 ) ;
  assign n4282 = ( n4265 & ~n4272 ) | ( n4265 & n4281 ) | ( ~n4272 & n4281 ) ;
  assign n4283 = ( ~n4273 & n4274 ) | ( ~n4273 & n4279 ) | ( n4274 & n4279 ) ;
  assign n4284 = ( n4273 & ~n4280 ) | ( n4273 & n4283 ) | ( ~n4280 & n4283 ) ;
  assign n4285 = n4276 | n4278 ;
  assign n4286 = ~n4279 & n4285 ;
  assign n4287 = ( n4268 & n4270 ) | ( n4268 & n4286 ) | ( n4270 & n4286 ) ;
  assign n4288 = ~n4271 & n4287 ;
  assign n4289 = ( n4282 & n4284 ) | ( n4282 & n4288 ) | ( n4284 & n4288 ) ;
  assign n4290 = ( n4272 & n4280 ) | ( n4272 & n4289 ) | ( n4280 & n4289 ) ;
  assign n4291 = ( ~n4272 & n4280 ) | ( ~n4272 & n4289 ) | ( n4280 & n4289 ) ;
  assign n4292 = ( n4272 & ~n4290 ) | ( n4272 & n4291 ) | ( ~n4290 & n4291 ) ;
  assign n4293 = ( ~n4245 & n4253 ) | ( ~n4245 & n4263 ) | ( n4253 & n4263 ) ;
  assign n4294 = ( n4245 & ~n4264 ) | ( n4245 & n4293 ) | ( ~n4264 & n4293 ) ;
  assign n4295 = ( ~n4255 & n4257 ) | ( ~n4255 & n4262 ) | ( n4257 & n4262 ) ;
  assign n4296 = ( n4255 & ~n4263 ) | ( n4255 & n4295 ) | ( ~n4263 & n4295 ) ;
  assign n4297 = ( ~n4282 & n4284 ) | ( ~n4282 & n4288 ) | ( n4284 & n4288 ) ;
  assign n4298 = ( n4282 & ~n4289 ) | ( n4282 & n4297 ) | ( ~n4289 & n4297 ) ;
  assign n4299 = ( ~n4268 & n4270 ) | ( ~n4268 & n4286 ) | ( n4270 & n4286 ) ;
  assign n4300 = ( n4268 & ~n4287 ) | ( n4268 & n4299 ) | ( ~n4287 & n4299 ) ;
  assign n4301 = ( n4259 & n4261 ) | ( n4259 & n4300 ) | ( n4261 & n4300 ) ;
  assign n4302 = ~n4262 & n4301 ;
  assign n4303 = ( n4296 & n4298 ) | ( n4296 & n4302 ) | ( n4298 & n4302 ) ;
  assign n4304 = ( n4292 & n4294 ) | ( n4292 & n4303 ) | ( n4294 & n4303 ) ;
  assign n4305 = ( n4264 & n4290 ) | ( n4264 & n4304 ) | ( n4290 & n4304 ) ;
  assign n4306 = ( x580 & x581 ) | ( x580 & x582 ) | ( x581 & x582 ) ;
  assign n4307 = ( x577 & x578 ) | ( x577 & x579 ) | ( x578 & x579 ) ;
  assign n4308 = ( ~x580 & x581 ) | ( ~x580 & x582 ) | ( x581 & x582 ) ;
  assign n4309 = ( x580 & ~n4306 ) | ( x580 & n4308 ) | ( ~n4306 & n4308 ) ;
  assign n4310 = ( ~x577 & x578 ) | ( ~x577 & x579 ) | ( x578 & x579 ) ;
  assign n4311 = ( x577 & ~n4307 ) | ( x577 & n4310 ) | ( ~n4307 & n4310 ) ;
  assign n4312 = n4309 & n4311 ;
  assign n4313 = ( n4306 & n4307 ) | ( n4306 & n4312 ) | ( n4307 & n4312 ) ;
  assign n4314 = ( x571 & x572 ) | ( x571 & x573 ) | ( x572 & x573 ) ;
  assign n4315 = ( x574 & x575 ) | ( x574 & x576 ) | ( x575 & x576 ) ;
  assign n4316 = ( ~x574 & x575 ) | ( ~x574 & x576 ) | ( x575 & x576 ) ;
  assign n4317 = ( x574 & ~n4315 ) | ( x574 & n4316 ) | ( ~n4315 & n4316 ) ;
  assign n4318 = ( ~x571 & x572 ) | ( ~x571 & x573 ) | ( x572 & x573 ) ;
  assign n4319 = ( x571 & ~n4314 ) | ( x571 & n4318 ) | ( ~n4314 & n4318 ) ;
  assign n4320 = n4317 & n4319 ;
  assign n4321 = ( n4314 & n4315 ) | ( n4314 & n4320 ) | ( n4315 & n4320 ) ;
  assign n4322 = ( ~n4306 & n4307 ) | ( ~n4306 & n4312 ) | ( n4307 & n4312 ) ;
  assign n4323 = ( n4306 & ~n4313 ) | ( n4306 & n4322 ) | ( ~n4313 & n4322 ) ;
  assign n4324 = ( ~n4314 & n4315 ) | ( ~n4314 & n4320 ) | ( n4315 & n4320 ) ;
  assign n4325 = ( n4314 & ~n4321 ) | ( n4314 & n4324 ) | ( ~n4321 & n4324 ) ;
  assign n4326 = n4309 | n4311 ;
  assign n4327 = ~n4312 & n4326 ;
  assign n4328 = n4317 | n4319 ;
  assign n4329 = ~n4320 & n4328 ;
  assign n4330 = n4327 & n4329 ;
  assign n4331 = ( n4323 & n4325 ) | ( n4323 & n4330 ) | ( n4325 & n4330 ) ;
  assign n4332 = ( n4313 & n4321 ) | ( n4313 & n4331 ) | ( n4321 & n4331 ) ;
  assign n4333 = ( x568 & x569 ) | ( x568 & x570 ) | ( x569 & x570 ) ;
  assign n4334 = ( x565 & x566 ) | ( x565 & x567 ) | ( x566 & x567 ) ;
  assign n4335 = ( ~x568 & x569 ) | ( ~x568 & x570 ) | ( x569 & x570 ) ;
  assign n4336 = ( x568 & ~n4333 ) | ( x568 & n4335 ) | ( ~n4333 & n4335 ) ;
  assign n4337 = ( ~x565 & x566 ) | ( ~x565 & x567 ) | ( x566 & x567 ) ;
  assign n4338 = ( x565 & ~n4334 ) | ( x565 & n4337 ) | ( ~n4334 & n4337 ) ;
  assign n4339 = n4336 & n4338 ;
  assign n4340 = ( n4333 & n4334 ) | ( n4333 & n4339 ) | ( n4334 & n4339 ) ;
  assign n4341 = ( x559 & x560 ) | ( x559 & x561 ) | ( x560 & x561 ) ;
  assign n4342 = ( x562 & x563 ) | ( x562 & x564 ) | ( x563 & x564 ) ;
  assign n4343 = ( ~x562 & x563 ) | ( ~x562 & x564 ) | ( x563 & x564 ) ;
  assign n4344 = ( x562 & ~n4342 ) | ( x562 & n4343 ) | ( ~n4342 & n4343 ) ;
  assign n4345 = ( ~x559 & x560 ) | ( ~x559 & x561 ) | ( x560 & x561 ) ;
  assign n4346 = ( x559 & ~n4341 ) | ( x559 & n4345 ) | ( ~n4341 & n4345 ) ;
  assign n4347 = n4344 & n4346 ;
  assign n4348 = ( n4341 & n4342 ) | ( n4341 & n4347 ) | ( n4342 & n4347 ) ;
  assign n4349 = ( ~n4333 & n4334 ) | ( ~n4333 & n4339 ) | ( n4334 & n4339 ) ;
  assign n4350 = ( n4333 & ~n4340 ) | ( n4333 & n4349 ) | ( ~n4340 & n4349 ) ;
  assign n4351 = ( ~n4341 & n4342 ) | ( ~n4341 & n4347 ) | ( n4342 & n4347 ) ;
  assign n4352 = ( n4341 & ~n4348 ) | ( n4341 & n4351 ) | ( ~n4348 & n4351 ) ;
  assign n4353 = n4344 | n4346 ;
  assign n4354 = ~n4347 & n4353 ;
  assign n4355 = ( n4336 & n4338 ) | ( n4336 & n4354 ) | ( n4338 & n4354 ) ;
  assign n4356 = ~n4339 & n4355 ;
  assign n4357 = ( n4350 & n4352 ) | ( n4350 & n4356 ) | ( n4352 & n4356 ) ;
  assign n4358 = ( n4340 & n4348 ) | ( n4340 & n4357 ) | ( n4348 & n4357 ) ;
  assign n4359 = ( ~n4340 & n4348 ) | ( ~n4340 & n4357 ) | ( n4348 & n4357 ) ;
  assign n4360 = ( n4340 & ~n4358 ) | ( n4340 & n4359 ) | ( ~n4358 & n4359 ) ;
  assign n4361 = ( ~n4313 & n4321 ) | ( ~n4313 & n4331 ) | ( n4321 & n4331 ) ;
  assign n4362 = ( n4313 & ~n4332 ) | ( n4313 & n4361 ) | ( ~n4332 & n4361 ) ;
  assign n4363 = ( ~n4323 & n4325 ) | ( ~n4323 & n4330 ) | ( n4325 & n4330 ) ;
  assign n4364 = ( n4323 & ~n4331 ) | ( n4323 & n4363 ) | ( ~n4331 & n4363 ) ;
  assign n4365 = ( ~n4350 & n4352 ) | ( ~n4350 & n4356 ) | ( n4352 & n4356 ) ;
  assign n4366 = ( n4350 & ~n4357 ) | ( n4350 & n4365 ) | ( ~n4357 & n4365 ) ;
  assign n4367 = ( ~n4336 & n4338 ) | ( ~n4336 & n4354 ) | ( n4338 & n4354 ) ;
  assign n4368 = ( n4336 & ~n4355 ) | ( n4336 & n4367 ) | ( ~n4355 & n4367 ) ;
  assign n4369 = ( n4327 & n4329 ) | ( n4327 & n4368 ) | ( n4329 & n4368 ) ;
  assign n4370 = ~n4330 & n4369 ;
  assign n4371 = ( n4364 & n4366 ) | ( n4364 & n4370 ) | ( n4366 & n4370 ) ;
  assign n4372 = ( n4360 & n4362 ) | ( n4360 & n4371 ) | ( n4362 & n4371 ) ;
  assign n4373 = ( n4332 & n4358 ) | ( n4332 & n4372 ) | ( n4358 & n4372 ) ;
  assign n4374 = ( ~n4264 & n4290 ) | ( ~n4264 & n4304 ) | ( n4290 & n4304 ) ;
  assign n4375 = ( n4264 & ~n4305 ) | ( n4264 & n4374 ) | ( ~n4305 & n4374 ) ;
  assign n4376 = ( ~n4332 & n4358 ) | ( ~n4332 & n4372 ) | ( n4358 & n4372 ) ;
  assign n4377 = ( n4332 & ~n4373 ) | ( n4332 & n4376 ) | ( ~n4373 & n4376 ) ;
  assign n4378 = ( ~n4360 & n4362 ) | ( ~n4360 & n4371 ) | ( n4362 & n4371 ) ;
  assign n4379 = ( n4360 & ~n4372 ) | ( n4360 & n4378 ) | ( ~n4372 & n4378 ) ;
  assign n4380 = ( ~n4292 & n4294 ) | ( ~n4292 & n4303 ) | ( n4294 & n4303 ) ;
  assign n4381 = ( n4292 & ~n4304 ) | ( n4292 & n4380 ) | ( ~n4304 & n4380 ) ;
  assign n4382 = ( n4296 & n4298 ) | ( n4296 & ~n4302 ) | ( n4298 & ~n4302 ) ;
  assign n4383 = ( n4302 & ~n4303 ) | ( n4302 & n4382 ) | ( ~n4303 & n4382 ) ;
  assign n4384 = ( n4364 & n4366 ) | ( n4364 & ~n4370 ) | ( n4366 & ~n4370 ) ;
  assign n4385 = ( n4370 & ~n4371 ) | ( n4370 & n4384 ) | ( ~n4371 & n4384 ) ;
  assign n4386 = ( ~n4259 & n4261 ) | ( ~n4259 & n4300 ) | ( n4261 & n4300 ) ;
  assign n4387 = ( n4259 & ~n4301 ) | ( n4259 & n4386 ) | ( ~n4301 & n4386 ) ;
  assign n4388 = ( ~n4327 & n4329 ) | ( ~n4327 & n4368 ) | ( n4329 & n4368 ) ;
  assign n4389 = ( n4327 & ~n4369 ) | ( n4327 & n4388 ) | ( ~n4369 & n4388 ) ;
  assign n4390 = n4387 & n4389 ;
  assign n4391 = ( n4383 & n4385 ) | ( n4383 & n4390 ) | ( n4385 & n4390 ) ;
  assign n4392 = ( n4379 & n4381 ) | ( n4379 & n4391 ) | ( n4381 & n4391 ) ;
  assign n4393 = ( n4375 & n4377 ) | ( n4375 & n4392 ) | ( n4377 & n4392 ) ;
  assign n4394 = ( n4305 & n4373 ) | ( n4305 & n4393 ) | ( n4373 & n4393 ) ;
  assign n4395 = ( ~n4305 & n4373 ) | ( ~n4305 & n4393 ) | ( n4373 & n4393 ) ;
  assign n4396 = ( n4305 & ~n4394 ) | ( n4305 & n4395 ) | ( ~n4394 & n4395 ) ;
  assign n4397 = ( ~n4148 & n4216 ) | ( ~n4148 & n4236 ) | ( n4216 & n4236 ) ;
  assign n4398 = ( n4148 & ~n4237 ) | ( n4148 & n4397 ) | ( ~n4237 & n4397 ) ;
  assign n4399 = ( ~n4218 & n4220 ) | ( ~n4218 & n4235 ) | ( n4220 & n4235 ) ;
  assign n4400 = ( n4218 & ~n4236 ) | ( n4218 & n4399 ) | ( ~n4236 & n4399 ) ;
  assign n4401 = ( ~n4375 & n4377 ) | ( ~n4375 & n4392 ) | ( n4377 & n4392 ) ;
  assign n4402 = ( n4375 & ~n4393 ) | ( n4375 & n4401 ) | ( ~n4393 & n4401 ) ;
  assign n4403 = ( ~n4379 & n4381 ) | ( ~n4379 & n4391 ) | ( n4381 & n4391 ) ;
  assign n4404 = ( n4379 & ~n4392 ) | ( n4379 & n4403 ) | ( ~n4392 & n4403 ) ;
  assign n4405 = ( ~n4222 & n4224 ) | ( ~n4222 & n4234 ) | ( n4224 & n4234 ) ;
  assign n4406 = ( n4222 & ~n4235 ) | ( n4222 & n4405 ) | ( ~n4235 & n4405 ) ;
  assign n4407 = ( ~n4226 & n4228 ) | ( ~n4226 & n4233 ) | ( n4228 & n4233 ) ;
  assign n4408 = ( n4226 & ~n4234 ) | ( n4226 & n4407 ) | ( ~n4234 & n4407 ) ;
  assign n4409 = ( ~n4383 & n4385 ) | ( ~n4383 & n4390 ) | ( n4385 & n4390 ) ;
  assign n4410 = ( n4383 & ~n4391 ) | ( n4383 & n4409 ) | ( ~n4391 & n4409 ) ;
  assign n4411 = n4387 | n4389 ;
  assign n4412 = ~n4390 & n4411 ;
  assign n4413 = ( n4230 & n4232 ) | ( n4230 & n4412 ) | ( n4232 & n4412 ) ;
  assign n4414 = ~n4233 & n4413 ;
  assign n4415 = ( n4408 & n4410 ) | ( n4408 & n4414 ) | ( n4410 & n4414 ) ;
  assign n4416 = ( n4404 & n4406 ) | ( n4404 & n4415 ) | ( n4406 & n4415 ) ;
  assign n4417 = ( n4400 & n4402 ) | ( n4400 & n4416 ) | ( n4402 & n4416 ) ;
  assign n4418 = ( n4396 & n4398 ) | ( n4396 & n4417 ) | ( n4398 & n4417 ) ;
  assign n4419 = ( n4237 & n4394 ) | ( n4237 & n4418 ) | ( n4394 & n4418 ) ;
  assign n4420 = ( x556 & x557 ) | ( x556 & x558 ) | ( x557 & x558 ) ;
  assign n4421 = ( x553 & x554 ) | ( x553 & x555 ) | ( x554 & x555 ) ;
  assign n4422 = ( ~x556 & x557 ) | ( ~x556 & x558 ) | ( x557 & x558 ) ;
  assign n4423 = ( x556 & ~n4420 ) | ( x556 & n4422 ) | ( ~n4420 & n4422 ) ;
  assign n4424 = ( ~x553 & x554 ) | ( ~x553 & x555 ) | ( x554 & x555 ) ;
  assign n4425 = ( x553 & ~n4421 ) | ( x553 & n4424 ) | ( ~n4421 & n4424 ) ;
  assign n4426 = n4423 & n4425 ;
  assign n4427 = ( n4420 & n4421 ) | ( n4420 & n4426 ) | ( n4421 & n4426 ) ;
  assign n4428 = ( x547 & x548 ) | ( x547 & x549 ) | ( x548 & x549 ) ;
  assign n4429 = ( x550 & x551 ) | ( x550 & x552 ) | ( x551 & x552 ) ;
  assign n4430 = ( ~x550 & x551 ) | ( ~x550 & x552 ) | ( x551 & x552 ) ;
  assign n4431 = ( x550 & ~n4429 ) | ( x550 & n4430 ) | ( ~n4429 & n4430 ) ;
  assign n4432 = ( ~x547 & x548 ) | ( ~x547 & x549 ) | ( x548 & x549 ) ;
  assign n4433 = ( x547 & ~n4428 ) | ( x547 & n4432 ) | ( ~n4428 & n4432 ) ;
  assign n4434 = n4431 & n4433 ;
  assign n4435 = ( n4428 & n4429 ) | ( n4428 & n4434 ) | ( n4429 & n4434 ) ;
  assign n4436 = ( ~n4420 & n4421 ) | ( ~n4420 & n4426 ) | ( n4421 & n4426 ) ;
  assign n4437 = ( n4420 & ~n4427 ) | ( n4420 & n4436 ) | ( ~n4427 & n4436 ) ;
  assign n4438 = ( ~n4428 & n4429 ) | ( ~n4428 & n4434 ) | ( n4429 & n4434 ) ;
  assign n4439 = ( n4428 & ~n4435 ) | ( n4428 & n4438 ) | ( ~n4435 & n4438 ) ;
  assign n4440 = n4423 | n4425 ;
  assign n4441 = ~n4426 & n4440 ;
  assign n4442 = n4431 | n4433 ;
  assign n4443 = ~n4434 & n4442 ;
  assign n4444 = n4441 & n4443 ;
  assign n4445 = ( n4437 & n4439 ) | ( n4437 & n4444 ) | ( n4439 & n4444 ) ;
  assign n4446 = ( n4427 & n4435 ) | ( n4427 & n4445 ) | ( n4435 & n4445 ) ;
  assign n4447 = ( x544 & x545 ) | ( x544 & x546 ) | ( x545 & x546 ) ;
  assign n4448 = ( x541 & x542 ) | ( x541 & x543 ) | ( x542 & x543 ) ;
  assign n4449 = ( ~x544 & x545 ) | ( ~x544 & x546 ) | ( x545 & x546 ) ;
  assign n4450 = ( x544 & ~n4447 ) | ( x544 & n4449 ) | ( ~n4447 & n4449 ) ;
  assign n4451 = ( ~x541 & x542 ) | ( ~x541 & x543 ) | ( x542 & x543 ) ;
  assign n4452 = ( x541 & ~n4448 ) | ( x541 & n4451 ) | ( ~n4448 & n4451 ) ;
  assign n4453 = n4450 & n4452 ;
  assign n4454 = ( n4447 & n4448 ) | ( n4447 & n4453 ) | ( n4448 & n4453 ) ;
  assign n4455 = ( x535 & x536 ) | ( x535 & x537 ) | ( x536 & x537 ) ;
  assign n4456 = ( x538 & x539 ) | ( x538 & x540 ) | ( x539 & x540 ) ;
  assign n4457 = ( ~x538 & x539 ) | ( ~x538 & x540 ) | ( x539 & x540 ) ;
  assign n4458 = ( x538 & ~n4456 ) | ( x538 & n4457 ) | ( ~n4456 & n4457 ) ;
  assign n4459 = ( ~x535 & x536 ) | ( ~x535 & x537 ) | ( x536 & x537 ) ;
  assign n4460 = ( x535 & ~n4455 ) | ( x535 & n4459 ) | ( ~n4455 & n4459 ) ;
  assign n4461 = n4458 & n4460 ;
  assign n4462 = ( n4455 & n4456 ) | ( n4455 & n4461 ) | ( n4456 & n4461 ) ;
  assign n4463 = ( ~n4447 & n4448 ) | ( ~n4447 & n4453 ) | ( n4448 & n4453 ) ;
  assign n4464 = ( n4447 & ~n4454 ) | ( n4447 & n4463 ) | ( ~n4454 & n4463 ) ;
  assign n4465 = ( ~n4455 & n4456 ) | ( ~n4455 & n4461 ) | ( n4456 & n4461 ) ;
  assign n4466 = ( n4455 & ~n4462 ) | ( n4455 & n4465 ) | ( ~n4462 & n4465 ) ;
  assign n4467 = n4458 | n4460 ;
  assign n4468 = ~n4461 & n4467 ;
  assign n4469 = ( n4450 & n4452 ) | ( n4450 & n4468 ) | ( n4452 & n4468 ) ;
  assign n4470 = ~n4453 & n4469 ;
  assign n4471 = ( n4464 & n4466 ) | ( n4464 & n4470 ) | ( n4466 & n4470 ) ;
  assign n4472 = ( n4454 & n4462 ) | ( n4454 & n4471 ) | ( n4462 & n4471 ) ;
  assign n4473 = ( ~n4454 & n4462 ) | ( ~n4454 & n4471 ) | ( n4462 & n4471 ) ;
  assign n4474 = ( n4454 & ~n4472 ) | ( n4454 & n4473 ) | ( ~n4472 & n4473 ) ;
  assign n4475 = ( ~n4427 & n4435 ) | ( ~n4427 & n4445 ) | ( n4435 & n4445 ) ;
  assign n4476 = ( n4427 & ~n4446 ) | ( n4427 & n4475 ) | ( ~n4446 & n4475 ) ;
  assign n4477 = ( ~n4437 & n4439 ) | ( ~n4437 & n4444 ) | ( n4439 & n4444 ) ;
  assign n4478 = ( n4437 & ~n4445 ) | ( n4437 & n4477 ) | ( ~n4445 & n4477 ) ;
  assign n4479 = ( ~n4464 & n4466 ) | ( ~n4464 & n4470 ) | ( n4466 & n4470 ) ;
  assign n4480 = ( n4464 & ~n4471 ) | ( n4464 & n4479 ) | ( ~n4471 & n4479 ) ;
  assign n4481 = ( ~n4450 & n4452 ) | ( ~n4450 & n4468 ) | ( n4452 & n4468 ) ;
  assign n4482 = ( n4450 & ~n4469 ) | ( n4450 & n4481 ) | ( ~n4469 & n4481 ) ;
  assign n4483 = ( n4441 & n4443 ) | ( n4441 & n4482 ) | ( n4443 & n4482 ) ;
  assign n4484 = ~n4444 & n4483 ;
  assign n4485 = ( n4478 & n4480 ) | ( n4478 & n4484 ) | ( n4480 & n4484 ) ;
  assign n4486 = ( n4474 & n4476 ) | ( n4474 & n4485 ) | ( n4476 & n4485 ) ;
  assign n4487 = ( n4446 & n4472 ) | ( n4446 & n4486 ) | ( n4472 & n4486 ) ;
  assign n4488 = ( x532 & x533 ) | ( x532 & x534 ) | ( x533 & x534 ) ;
  assign n4489 = ( x529 & x530 ) | ( x529 & x531 ) | ( x530 & x531 ) ;
  assign n4490 = ( ~x532 & x533 ) | ( ~x532 & x534 ) | ( x533 & x534 ) ;
  assign n4491 = ( x532 & ~n4488 ) | ( x532 & n4490 ) | ( ~n4488 & n4490 ) ;
  assign n4492 = ( ~x529 & x530 ) | ( ~x529 & x531 ) | ( x530 & x531 ) ;
  assign n4493 = ( x529 & ~n4489 ) | ( x529 & n4492 ) | ( ~n4489 & n4492 ) ;
  assign n4494 = n4491 & n4493 ;
  assign n4495 = ( n4488 & n4489 ) | ( n4488 & n4494 ) | ( n4489 & n4494 ) ;
  assign n4496 = ( x523 & x524 ) | ( x523 & x525 ) | ( x524 & x525 ) ;
  assign n4497 = ( x526 & x527 ) | ( x526 & x528 ) | ( x527 & x528 ) ;
  assign n4498 = ( ~x526 & x527 ) | ( ~x526 & x528 ) | ( x527 & x528 ) ;
  assign n4499 = ( x526 & ~n4497 ) | ( x526 & n4498 ) | ( ~n4497 & n4498 ) ;
  assign n4500 = ( ~x523 & x524 ) | ( ~x523 & x525 ) | ( x524 & x525 ) ;
  assign n4501 = ( x523 & ~n4496 ) | ( x523 & n4500 ) | ( ~n4496 & n4500 ) ;
  assign n4502 = n4499 & n4501 ;
  assign n4503 = ( n4496 & n4497 ) | ( n4496 & n4502 ) | ( n4497 & n4502 ) ;
  assign n4504 = ( ~n4488 & n4489 ) | ( ~n4488 & n4494 ) | ( n4489 & n4494 ) ;
  assign n4505 = ( n4488 & ~n4495 ) | ( n4488 & n4504 ) | ( ~n4495 & n4504 ) ;
  assign n4506 = ( ~n4496 & n4497 ) | ( ~n4496 & n4502 ) | ( n4497 & n4502 ) ;
  assign n4507 = ( n4496 & ~n4503 ) | ( n4496 & n4506 ) | ( ~n4503 & n4506 ) ;
  assign n4508 = n4491 | n4493 ;
  assign n4509 = ~n4494 & n4508 ;
  assign n4510 = n4499 | n4501 ;
  assign n4511 = ~n4502 & n4510 ;
  assign n4512 = n4509 & n4511 ;
  assign n4513 = ( n4505 & n4507 ) | ( n4505 & n4512 ) | ( n4507 & n4512 ) ;
  assign n4514 = ( n4495 & n4503 ) | ( n4495 & n4513 ) | ( n4503 & n4513 ) ;
  assign n4515 = ( x520 & x521 ) | ( x520 & x522 ) | ( x521 & x522 ) ;
  assign n4516 = ( x517 & x518 ) | ( x517 & x519 ) | ( x518 & x519 ) ;
  assign n4517 = ( ~x520 & x521 ) | ( ~x520 & x522 ) | ( x521 & x522 ) ;
  assign n4518 = ( x520 & ~n4515 ) | ( x520 & n4517 ) | ( ~n4515 & n4517 ) ;
  assign n4519 = ( ~x517 & x518 ) | ( ~x517 & x519 ) | ( x518 & x519 ) ;
  assign n4520 = ( x517 & ~n4516 ) | ( x517 & n4519 ) | ( ~n4516 & n4519 ) ;
  assign n4521 = n4518 & n4520 ;
  assign n4522 = ( n4515 & n4516 ) | ( n4515 & n4521 ) | ( n4516 & n4521 ) ;
  assign n4523 = ( x511 & x512 ) | ( x511 & x513 ) | ( x512 & x513 ) ;
  assign n4524 = ( x514 & x515 ) | ( x514 & x516 ) | ( x515 & x516 ) ;
  assign n4525 = ( ~x514 & x515 ) | ( ~x514 & x516 ) | ( x515 & x516 ) ;
  assign n4526 = ( x514 & ~n4524 ) | ( x514 & n4525 ) | ( ~n4524 & n4525 ) ;
  assign n4527 = ( ~x511 & x512 ) | ( ~x511 & x513 ) | ( x512 & x513 ) ;
  assign n4528 = ( x511 & ~n4523 ) | ( x511 & n4527 ) | ( ~n4523 & n4527 ) ;
  assign n4529 = n4526 & n4528 ;
  assign n4530 = ( n4523 & n4524 ) | ( n4523 & n4529 ) | ( n4524 & n4529 ) ;
  assign n4531 = ( ~n4515 & n4516 ) | ( ~n4515 & n4521 ) | ( n4516 & n4521 ) ;
  assign n4532 = ( n4515 & ~n4522 ) | ( n4515 & n4531 ) | ( ~n4522 & n4531 ) ;
  assign n4533 = ( ~n4523 & n4524 ) | ( ~n4523 & n4529 ) | ( n4524 & n4529 ) ;
  assign n4534 = ( n4523 & ~n4530 ) | ( n4523 & n4533 ) | ( ~n4530 & n4533 ) ;
  assign n4535 = n4526 | n4528 ;
  assign n4536 = ~n4529 & n4535 ;
  assign n4537 = ( n4518 & n4520 ) | ( n4518 & n4536 ) | ( n4520 & n4536 ) ;
  assign n4538 = ~n4521 & n4537 ;
  assign n4539 = ( n4532 & n4534 ) | ( n4532 & n4538 ) | ( n4534 & n4538 ) ;
  assign n4540 = ( n4522 & n4530 ) | ( n4522 & n4539 ) | ( n4530 & n4539 ) ;
  assign n4541 = ( ~n4522 & n4530 ) | ( ~n4522 & n4539 ) | ( n4530 & n4539 ) ;
  assign n4542 = ( n4522 & ~n4540 ) | ( n4522 & n4541 ) | ( ~n4540 & n4541 ) ;
  assign n4543 = ( ~n4495 & n4503 ) | ( ~n4495 & n4513 ) | ( n4503 & n4513 ) ;
  assign n4544 = ( n4495 & ~n4514 ) | ( n4495 & n4543 ) | ( ~n4514 & n4543 ) ;
  assign n4545 = ( ~n4505 & n4507 ) | ( ~n4505 & n4512 ) | ( n4507 & n4512 ) ;
  assign n4546 = ( n4505 & ~n4513 ) | ( n4505 & n4545 ) | ( ~n4513 & n4545 ) ;
  assign n4547 = ( ~n4532 & n4534 ) | ( ~n4532 & n4538 ) | ( n4534 & n4538 ) ;
  assign n4548 = ( n4532 & ~n4539 ) | ( n4532 & n4547 ) | ( ~n4539 & n4547 ) ;
  assign n4549 = ( ~n4518 & n4520 ) | ( ~n4518 & n4536 ) | ( n4520 & n4536 ) ;
  assign n4550 = ( n4518 & ~n4537 ) | ( n4518 & n4549 ) | ( ~n4537 & n4549 ) ;
  assign n4551 = ( n4509 & n4511 ) | ( n4509 & n4550 ) | ( n4511 & n4550 ) ;
  assign n4552 = ~n4512 & n4551 ;
  assign n4553 = ( n4546 & n4548 ) | ( n4546 & n4552 ) | ( n4548 & n4552 ) ;
  assign n4554 = ( n4542 & n4544 ) | ( n4542 & n4553 ) | ( n4544 & n4553 ) ;
  assign n4555 = ( n4514 & n4540 ) | ( n4514 & n4554 ) | ( n4540 & n4554 ) ;
  assign n4556 = ( ~n4446 & n4472 ) | ( ~n4446 & n4486 ) | ( n4472 & n4486 ) ;
  assign n4557 = ( n4446 & ~n4487 ) | ( n4446 & n4556 ) | ( ~n4487 & n4556 ) ;
  assign n4558 = ( ~n4514 & n4540 ) | ( ~n4514 & n4554 ) | ( n4540 & n4554 ) ;
  assign n4559 = ( n4514 & ~n4555 ) | ( n4514 & n4558 ) | ( ~n4555 & n4558 ) ;
  assign n4560 = ( ~n4542 & n4544 ) | ( ~n4542 & n4553 ) | ( n4544 & n4553 ) ;
  assign n4561 = ( n4542 & ~n4554 ) | ( n4542 & n4560 ) | ( ~n4554 & n4560 ) ;
  assign n4562 = ( ~n4474 & n4476 ) | ( ~n4474 & n4485 ) | ( n4476 & n4485 ) ;
  assign n4563 = ( n4474 & ~n4486 ) | ( n4474 & n4562 ) | ( ~n4486 & n4562 ) ;
  assign n4564 = ( n4478 & n4480 ) | ( n4478 & ~n4484 ) | ( n4480 & ~n4484 ) ;
  assign n4565 = ( n4484 & ~n4485 ) | ( n4484 & n4564 ) | ( ~n4485 & n4564 ) ;
  assign n4566 = ( n4546 & n4548 ) | ( n4546 & ~n4552 ) | ( n4548 & ~n4552 ) ;
  assign n4567 = ( n4552 & ~n4553 ) | ( n4552 & n4566 ) | ( ~n4553 & n4566 ) ;
  assign n4568 = ( ~n4441 & n4443 ) | ( ~n4441 & n4482 ) | ( n4443 & n4482 ) ;
  assign n4569 = ( n4441 & ~n4483 ) | ( n4441 & n4568 ) | ( ~n4483 & n4568 ) ;
  assign n4570 = ( ~n4509 & n4511 ) | ( ~n4509 & n4550 ) | ( n4511 & n4550 ) ;
  assign n4571 = ( n4509 & ~n4551 ) | ( n4509 & n4570 ) | ( ~n4551 & n4570 ) ;
  assign n4572 = n4569 & n4571 ;
  assign n4573 = ( n4565 & n4567 ) | ( n4565 & n4572 ) | ( n4567 & n4572 ) ;
  assign n4574 = ( n4561 & n4563 ) | ( n4561 & n4573 ) | ( n4563 & n4573 ) ;
  assign n4575 = ( n4557 & n4559 ) | ( n4557 & n4574 ) | ( n4559 & n4574 ) ;
  assign n4576 = ( n4487 & n4555 ) | ( n4487 & n4575 ) | ( n4555 & n4575 ) ;
  assign n4577 = ( x508 & x509 ) | ( x508 & x510 ) | ( x509 & x510 ) ;
  assign n4578 = ( x505 & x506 ) | ( x505 & x507 ) | ( x506 & x507 ) ;
  assign n4579 = ( ~x508 & x509 ) | ( ~x508 & x510 ) | ( x509 & x510 ) ;
  assign n4580 = ( x508 & ~n4577 ) | ( x508 & n4579 ) | ( ~n4577 & n4579 ) ;
  assign n4581 = ( ~x505 & x506 ) | ( ~x505 & x507 ) | ( x506 & x507 ) ;
  assign n4582 = ( x505 & ~n4578 ) | ( x505 & n4581 ) | ( ~n4578 & n4581 ) ;
  assign n4583 = n4580 & n4582 ;
  assign n4584 = ( n4577 & n4578 ) | ( n4577 & n4583 ) | ( n4578 & n4583 ) ;
  assign n4585 = ( x499 & x500 ) | ( x499 & x501 ) | ( x500 & x501 ) ;
  assign n4586 = ( x502 & x503 ) | ( x502 & x504 ) | ( x503 & x504 ) ;
  assign n4587 = ( ~x502 & x503 ) | ( ~x502 & x504 ) | ( x503 & x504 ) ;
  assign n4588 = ( x502 & ~n4586 ) | ( x502 & n4587 ) | ( ~n4586 & n4587 ) ;
  assign n4589 = ( ~x499 & x500 ) | ( ~x499 & x501 ) | ( x500 & x501 ) ;
  assign n4590 = ( x499 & ~n4585 ) | ( x499 & n4589 ) | ( ~n4585 & n4589 ) ;
  assign n4591 = n4588 & n4590 ;
  assign n4592 = ( n4585 & n4586 ) | ( n4585 & n4591 ) | ( n4586 & n4591 ) ;
  assign n4593 = ( ~n4577 & n4578 ) | ( ~n4577 & n4583 ) | ( n4578 & n4583 ) ;
  assign n4594 = ( n4577 & ~n4584 ) | ( n4577 & n4593 ) | ( ~n4584 & n4593 ) ;
  assign n4595 = ( ~n4585 & n4586 ) | ( ~n4585 & n4591 ) | ( n4586 & n4591 ) ;
  assign n4596 = ( n4585 & ~n4592 ) | ( n4585 & n4595 ) | ( ~n4592 & n4595 ) ;
  assign n4597 = n4580 | n4582 ;
  assign n4598 = ~n4583 & n4597 ;
  assign n4599 = n4588 | n4590 ;
  assign n4600 = ~n4591 & n4599 ;
  assign n4601 = n4598 & n4600 ;
  assign n4602 = ( n4594 & n4596 ) | ( n4594 & n4601 ) | ( n4596 & n4601 ) ;
  assign n4603 = ( n4584 & n4592 ) | ( n4584 & n4602 ) | ( n4592 & n4602 ) ;
  assign n4604 = ( x496 & x497 ) | ( x496 & x498 ) | ( x497 & x498 ) ;
  assign n4605 = ( x493 & x494 ) | ( x493 & x495 ) | ( x494 & x495 ) ;
  assign n4606 = ( ~x496 & x497 ) | ( ~x496 & x498 ) | ( x497 & x498 ) ;
  assign n4607 = ( x496 & ~n4604 ) | ( x496 & n4606 ) | ( ~n4604 & n4606 ) ;
  assign n4608 = ( ~x493 & x494 ) | ( ~x493 & x495 ) | ( x494 & x495 ) ;
  assign n4609 = ( x493 & ~n4605 ) | ( x493 & n4608 ) | ( ~n4605 & n4608 ) ;
  assign n4610 = n4607 & n4609 ;
  assign n4611 = ( n4604 & n4605 ) | ( n4604 & n4610 ) | ( n4605 & n4610 ) ;
  assign n4612 = ( x487 & x488 ) | ( x487 & x489 ) | ( x488 & x489 ) ;
  assign n4613 = ( x490 & x491 ) | ( x490 & x492 ) | ( x491 & x492 ) ;
  assign n4614 = ( ~x490 & x491 ) | ( ~x490 & x492 ) | ( x491 & x492 ) ;
  assign n4615 = ( x490 & ~n4613 ) | ( x490 & n4614 ) | ( ~n4613 & n4614 ) ;
  assign n4616 = ( ~x487 & x488 ) | ( ~x487 & x489 ) | ( x488 & x489 ) ;
  assign n4617 = ( x487 & ~n4612 ) | ( x487 & n4616 ) | ( ~n4612 & n4616 ) ;
  assign n4618 = n4615 & n4617 ;
  assign n4619 = ( n4612 & n4613 ) | ( n4612 & n4618 ) | ( n4613 & n4618 ) ;
  assign n4620 = ( ~n4604 & n4605 ) | ( ~n4604 & n4610 ) | ( n4605 & n4610 ) ;
  assign n4621 = ( n4604 & ~n4611 ) | ( n4604 & n4620 ) | ( ~n4611 & n4620 ) ;
  assign n4622 = ( ~n4612 & n4613 ) | ( ~n4612 & n4618 ) | ( n4613 & n4618 ) ;
  assign n4623 = ( n4612 & ~n4619 ) | ( n4612 & n4622 ) | ( ~n4619 & n4622 ) ;
  assign n4624 = n4615 | n4617 ;
  assign n4625 = ~n4618 & n4624 ;
  assign n4626 = ( n4607 & n4609 ) | ( n4607 & n4625 ) | ( n4609 & n4625 ) ;
  assign n4627 = ~n4610 & n4626 ;
  assign n4628 = ( n4621 & n4623 ) | ( n4621 & n4627 ) | ( n4623 & n4627 ) ;
  assign n4629 = ( n4611 & n4619 ) | ( n4611 & n4628 ) | ( n4619 & n4628 ) ;
  assign n4630 = ( ~n4611 & n4619 ) | ( ~n4611 & n4628 ) | ( n4619 & n4628 ) ;
  assign n4631 = ( n4611 & ~n4629 ) | ( n4611 & n4630 ) | ( ~n4629 & n4630 ) ;
  assign n4632 = ( ~n4584 & n4592 ) | ( ~n4584 & n4602 ) | ( n4592 & n4602 ) ;
  assign n4633 = ( n4584 & ~n4603 ) | ( n4584 & n4632 ) | ( ~n4603 & n4632 ) ;
  assign n4634 = ( ~n4594 & n4596 ) | ( ~n4594 & n4601 ) | ( n4596 & n4601 ) ;
  assign n4635 = ( n4594 & ~n4602 ) | ( n4594 & n4634 ) | ( ~n4602 & n4634 ) ;
  assign n4636 = ( ~n4621 & n4623 ) | ( ~n4621 & n4627 ) | ( n4623 & n4627 ) ;
  assign n4637 = ( n4621 & ~n4628 ) | ( n4621 & n4636 ) | ( ~n4628 & n4636 ) ;
  assign n4638 = ( ~n4607 & n4609 ) | ( ~n4607 & n4625 ) | ( n4609 & n4625 ) ;
  assign n4639 = ( n4607 & ~n4626 ) | ( n4607 & n4638 ) | ( ~n4626 & n4638 ) ;
  assign n4640 = ( n4598 & n4600 ) | ( n4598 & n4639 ) | ( n4600 & n4639 ) ;
  assign n4641 = ~n4601 & n4640 ;
  assign n4642 = ( n4635 & n4637 ) | ( n4635 & n4641 ) | ( n4637 & n4641 ) ;
  assign n4643 = ( n4631 & n4633 ) | ( n4631 & n4642 ) | ( n4633 & n4642 ) ;
  assign n4644 = ( n4603 & n4629 ) | ( n4603 & n4643 ) | ( n4629 & n4643 ) ;
  assign n4645 = ( x484 & x485 ) | ( x484 & x486 ) | ( x485 & x486 ) ;
  assign n4646 = ( x481 & x482 ) | ( x481 & x483 ) | ( x482 & x483 ) ;
  assign n4647 = ( ~x484 & x485 ) | ( ~x484 & x486 ) | ( x485 & x486 ) ;
  assign n4648 = ( x484 & ~n4645 ) | ( x484 & n4647 ) | ( ~n4645 & n4647 ) ;
  assign n4649 = ( ~x481 & x482 ) | ( ~x481 & x483 ) | ( x482 & x483 ) ;
  assign n4650 = ( x481 & ~n4646 ) | ( x481 & n4649 ) | ( ~n4646 & n4649 ) ;
  assign n4651 = n4648 & n4650 ;
  assign n4652 = ( n4645 & n4646 ) | ( n4645 & n4651 ) | ( n4646 & n4651 ) ;
  assign n4653 = ( x475 & x476 ) | ( x475 & x477 ) | ( x476 & x477 ) ;
  assign n4654 = ( x478 & x479 ) | ( x478 & x480 ) | ( x479 & x480 ) ;
  assign n4655 = ( ~x478 & x479 ) | ( ~x478 & x480 ) | ( x479 & x480 ) ;
  assign n4656 = ( x478 & ~n4654 ) | ( x478 & n4655 ) | ( ~n4654 & n4655 ) ;
  assign n4657 = ( ~x475 & x476 ) | ( ~x475 & x477 ) | ( x476 & x477 ) ;
  assign n4658 = ( x475 & ~n4653 ) | ( x475 & n4657 ) | ( ~n4653 & n4657 ) ;
  assign n4659 = n4656 & n4658 ;
  assign n4660 = ( n4653 & n4654 ) | ( n4653 & n4659 ) | ( n4654 & n4659 ) ;
  assign n4661 = ( ~n4645 & n4646 ) | ( ~n4645 & n4651 ) | ( n4646 & n4651 ) ;
  assign n4662 = ( n4645 & ~n4652 ) | ( n4645 & n4661 ) | ( ~n4652 & n4661 ) ;
  assign n4663 = ( ~n4653 & n4654 ) | ( ~n4653 & n4659 ) | ( n4654 & n4659 ) ;
  assign n4664 = ( n4653 & ~n4660 ) | ( n4653 & n4663 ) | ( ~n4660 & n4663 ) ;
  assign n4665 = n4656 | n4658 ;
  assign n4666 = ~n4659 & n4665 ;
  assign n4667 = n4648 | n4650 ;
  assign n4668 = ~n4651 & n4667 ;
  assign n4669 = n4666 & n4668 ;
  assign n4670 = ( n4662 & n4664 ) | ( n4662 & n4669 ) | ( n4664 & n4669 ) ;
  assign n4671 = ( n4652 & n4660 ) | ( n4652 & n4670 ) | ( n4660 & n4670 ) ;
  assign n4672 = ( x472 & x473 ) | ( x472 & x474 ) | ( x473 & x474 ) ;
  assign n4673 = ( x469 & x470 ) | ( x469 & x471 ) | ( x470 & x471 ) ;
  assign n4674 = ( ~x472 & x473 ) | ( ~x472 & x474 ) | ( x473 & x474 ) ;
  assign n4675 = ( x472 & ~n4672 ) | ( x472 & n4674 ) | ( ~n4672 & n4674 ) ;
  assign n4676 = ( ~x469 & x470 ) | ( ~x469 & x471 ) | ( x470 & x471 ) ;
  assign n4677 = ( x469 & ~n4673 ) | ( x469 & n4676 ) | ( ~n4673 & n4676 ) ;
  assign n4678 = n4675 & n4677 ;
  assign n4679 = ( n4672 & n4673 ) | ( n4672 & n4678 ) | ( n4673 & n4678 ) ;
  assign n4680 = ( x466 & x467 ) | ( x466 & x468 ) | ( x467 & x468 ) ;
  assign n4681 = ( x463 & x464 ) | ( x463 & x465 ) | ( x464 & x465 ) ;
  assign n4682 = ( ~x463 & x464 ) | ( ~x463 & x465 ) | ( x464 & x465 ) ;
  assign n4683 = ( x463 & ~n4681 ) | ( x463 & n4682 ) | ( ~n4681 & n4682 ) ;
  assign n4684 = ( ~x466 & x467 ) | ( ~x466 & x468 ) | ( x467 & x468 ) ;
  assign n4685 = ( x466 & ~n4680 ) | ( x466 & n4684 ) | ( ~n4680 & n4684 ) ;
  assign n4686 = n4683 & n4685 ;
  assign n4687 = ( n4680 & n4681 ) | ( n4680 & n4686 ) | ( n4681 & n4686 ) ;
  assign n4688 = ( ~n4672 & n4673 ) | ( ~n4672 & n4678 ) | ( n4673 & n4678 ) ;
  assign n4689 = ( n4672 & ~n4679 ) | ( n4672 & n4688 ) | ( ~n4679 & n4688 ) ;
  assign n4690 = ( ~n4680 & n4681 ) | ( ~n4680 & n4686 ) | ( n4681 & n4686 ) ;
  assign n4691 = ( n4680 & ~n4687 ) | ( n4680 & n4690 ) | ( ~n4687 & n4690 ) ;
  assign n4692 = n4675 | n4677 ;
  assign n4693 = ~n4678 & n4692 ;
  assign n4694 = ( n4683 & n4685 ) | ( n4683 & n4693 ) | ( n4685 & n4693 ) ;
  assign n4695 = ~n4686 & n4694 ;
  assign n4696 = ( n4689 & n4691 ) | ( n4689 & n4695 ) | ( n4691 & n4695 ) ;
  assign n4697 = ( n4679 & n4687 ) | ( n4679 & n4696 ) | ( n4687 & n4696 ) ;
  assign n4698 = ( ~n4679 & n4687 ) | ( ~n4679 & n4696 ) | ( n4687 & n4696 ) ;
  assign n4699 = ( n4679 & ~n4697 ) | ( n4679 & n4698 ) | ( ~n4697 & n4698 ) ;
  assign n4700 = ( ~n4652 & n4660 ) | ( ~n4652 & n4670 ) | ( n4660 & n4670 ) ;
  assign n4701 = ( n4652 & ~n4671 ) | ( n4652 & n4700 ) | ( ~n4671 & n4700 ) ;
  assign n4702 = ( ~n4662 & n4664 ) | ( ~n4662 & n4669 ) | ( n4664 & n4669 ) ;
  assign n4703 = ( n4662 & ~n4670 ) | ( n4662 & n4702 ) | ( ~n4670 & n4702 ) ;
  assign n4704 = ( ~n4689 & n4691 ) | ( ~n4689 & n4695 ) | ( n4691 & n4695 ) ;
  assign n4705 = ( n4689 & ~n4696 ) | ( n4689 & n4704 ) | ( ~n4696 & n4704 ) ;
  assign n4706 = ( ~n4683 & n4685 ) | ( ~n4683 & n4693 ) | ( n4685 & n4693 ) ;
  assign n4707 = ( n4683 & ~n4694 ) | ( n4683 & n4706 ) | ( ~n4694 & n4706 ) ;
  assign n4708 = ( n4666 & n4668 ) | ( n4666 & n4707 ) | ( n4668 & n4707 ) ;
  assign n4709 = ~n4669 & n4708 ;
  assign n4710 = ( n4703 & n4705 ) | ( n4703 & n4709 ) | ( n4705 & n4709 ) ;
  assign n4711 = ( n4699 & n4701 ) | ( n4699 & n4710 ) | ( n4701 & n4710 ) ;
  assign n4712 = ( n4671 & n4697 ) | ( n4671 & n4711 ) | ( n4697 & n4711 ) ;
  assign n4713 = ( ~n4603 & n4629 ) | ( ~n4603 & n4643 ) | ( n4629 & n4643 ) ;
  assign n4714 = ( n4603 & ~n4644 ) | ( n4603 & n4713 ) | ( ~n4644 & n4713 ) ;
  assign n4715 = ( ~n4671 & n4697 ) | ( ~n4671 & n4711 ) | ( n4697 & n4711 ) ;
  assign n4716 = ( n4671 & ~n4712 ) | ( n4671 & n4715 ) | ( ~n4712 & n4715 ) ;
  assign n4717 = ( ~n4699 & n4701 ) | ( ~n4699 & n4710 ) | ( n4701 & n4710 ) ;
  assign n4718 = ( n4699 & ~n4711 ) | ( n4699 & n4717 ) | ( ~n4711 & n4717 ) ;
  assign n4719 = ( ~n4631 & n4633 ) | ( ~n4631 & n4642 ) | ( n4633 & n4642 ) ;
  assign n4720 = ( n4631 & ~n4643 ) | ( n4631 & n4719 ) | ( ~n4643 & n4719 ) ;
  assign n4721 = ( n4635 & n4637 ) | ( n4635 & ~n4641 ) | ( n4637 & ~n4641 ) ;
  assign n4722 = ( n4641 & ~n4642 ) | ( n4641 & n4721 ) | ( ~n4642 & n4721 ) ;
  assign n4723 = ( n4703 & n4705 ) | ( n4703 & ~n4709 ) | ( n4705 & ~n4709 ) ;
  assign n4724 = ( n4709 & ~n4710 ) | ( n4709 & n4723 ) | ( ~n4710 & n4723 ) ;
  assign n4725 = ( ~n4666 & n4668 ) | ( ~n4666 & n4707 ) | ( n4668 & n4707 ) ;
  assign n4726 = ( n4666 & ~n4708 ) | ( n4666 & n4725 ) | ( ~n4708 & n4725 ) ;
  assign n4727 = ( ~n4598 & n4600 ) | ( ~n4598 & n4639 ) | ( n4600 & n4639 ) ;
  assign n4728 = ( n4598 & ~n4640 ) | ( n4598 & n4727 ) | ( ~n4640 & n4727 ) ;
  assign n4729 = n4726 & n4728 ;
  assign n4730 = ( n4722 & n4724 ) | ( n4722 & n4729 ) | ( n4724 & n4729 ) ;
  assign n4731 = ( n4718 & n4720 ) | ( n4718 & n4730 ) | ( n4720 & n4730 ) ;
  assign n4732 = ( n4714 & n4716 ) | ( n4714 & n4731 ) | ( n4716 & n4731 ) ;
  assign n4733 = ( n4644 & n4712 ) | ( n4644 & n4732 ) | ( n4712 & n4732 ) ;
  assign n4734 = ( ~n4644 & n4712 ) | ( ~n4644 & n4732 ) | ( n4712 & n4732 ) ;
  assign n4735 = ( n4644 & ~n4733 ) | ( n4644 & n4734 ) | ( ~n4733 & n4734 ) ;
  assign n4736 = ( ~n4487 & n4555 ) | ( ~n4487 & n4575 ) | ( n4555 & n4575 ) ;
  assign n4737 = ( n4487 & ~n4576 ) | ( n4487 & n4736 ) | ( ~n4576 & n4736 ) ;
  assign n4738 = ( ~n4557 & n4559 ) | ( ~n4557 & n4574 ) | ( n4559 & n4574 ) ;
  assign n4739 = ( n4557 & ~n4575 ) | ( n4557 & n4738 ) | ( ~n4575 & n4738 ) ;
  assign n4740 = ( ~n4714 & n4716 ) | ( ~n4714 & n4731 ) | ( n4716 & n4731 ) ;
  assign n4741 = ( n4714 & ~n4732 ) | ( n4714 & n4740 ) | ( ~n4732 & n4740 ) ;
  assign n4742 = ( ~n4718 & n4720 ) | ( ~n4718 & n4730 ) | ( n4720 & n4730 ) ;
  assign n4743 = ( n4718 & ~n4731 ) | ( n4718 & n4742 ) | ( ~n4731 & n4742 ) ;
  assign n4744 = ( ~n4561 & n4563 ) | ( ~n4561 & n4573 ) | ( n4563 & n4573 ) ;
  assign n4745 = ( n4561 & ~n4574 ) | ( n4561 & n4744 ) | ( ~n4574 & n4744 ) ;
  assign n4746 = ( ~n4565 & n4567 ) | ( ~n4565 & n4572 ) | ( n4567 & n4572 ) ;
  assign n4747 = ( n4565 & ~n4573 ) | ( n4565 & n4746 ) | ( ~n4573 & n4746 ) ;
  assign n4748 = ( ~n4722 & n4724 ) | ( ~n4722 & n4729 ) | ( n4724 & n4729 ) ;
  assign n4749 = ( n4722 & ~n4730 ) | ( n4722 & n4748 ) | ( ~n4730 & n4748 ) ;
  assign n4750 = n4726 | n4728 ;
  assign n4751 = ~n4729 & n4750 ;
  assign n4752 = ( n4569 & n4571 ) | ( n4569 & n4751 ) | ( n4571 & n4751 ) ;
  assign n4753 = ~n4572 & n4752 ;
  assign n4754 = ( n4747 & n4749 ) | ( n4747 & n4753 ) | ( n4749 & n4753 ) ;
  assign n4755 = ( n4743 & n4745 ) | ( n4743 & n4754 ) | ( n4745 & n4754 ) ;
  assign n4756 = ( n4739 & n4741 ) | ( n4739 & n4755 ) | ( n4741 & n4755 ) ;
  assign n4757 = ( n4735 & n4737 ) | ( n4735 & n4756 ) | ( n4737 & n4756 ) ;
  assign n4758 = ( n4576 & n4733 ) | ( n4576 & n4757 ) | ( n4733 & n4757 ) ;
  assign n4759 = ( ~n4237 & n4394 ) | ( ~n4237 & n4418 ) | ( n4394 & n4418 ) ;
  assign n4760 = ( n4237 & ~n4419 ) | ( n4237 & n4759 ) | ( ~n4419 & n4759 ) ;
  assign n4761 = ( ~n4576 & n4733 ) | ( ~n4576 & n4757 ) | ( n4733 & n4757 ) ;
  assign n4762 = ( n4576 & ~n4758 ) | ( n4576 & n4761 ) | ( ~n4758 & n4761 ) ;
  assign n4763 = ( ~n4735 & n4737 ) | ( ~n4735 & n4756 ) | ( n4737 & n4756 ) ;
  assign n4764 = ( n4735 & ~n4757 ) | ( n4735 & n4763 ) | ( ~n4757 & n4763 ) ;
  assign n4765 = ( ~n4396 & n4398 ) | ( ~n4396 & n4417 ) | ( n4398 & n4417 ) ;
  assign n4766 = ( n4396 & ~n4418 ) | ( n4396 & n4765 ) | ( ~n4418 & n4765 ) ;
  assign n4767 = ( ~n4400 & n4402 ) | ( ~n4400 & n4416 ) | ( n4402 & n4416 ) ;
  assign n4768 = ( n4400 & ~n4417 ) | ( n4400 & n4767 ) | ( ~n4417 & n4767 ) ;
  assign n4769 = ( ~n4739 & n4741 ) | ( ~n4739 & n4755 ) | ( n4741 & n4755 ) ;
  assign n4770 = ( n4739 & ~n4756 ) | ( n4739 & n4769 ) | ( ~n4756 & n4769 ) ;
  assign n4771 = ( ~n4743 & n4745 ) | ( ~n4743 & n4754 ) | ( n4745 & n4754 ) ;
  assign n4772 = ( n4743 & ~n4755 ) | ( n4743 & n4771 ) | ( ~n4755 & n4771 ) ;
  assign n4773 = ( ~n4404 & n4406 ) | ( ~n4404 & n4415 ) | ( n4406 & n4415 ) ;
  assign n4774 = ( n4404 & ~n4416 ) | ( n4404 & n4773 ) | ( ~n4416 & n4773 ) ;
  assign n4775 = ( n4408 & n4410 ) | ( n4408 & ~n4414 ) | ( n4410 & ~n4414 ) ;
  assign n4776 = ( n4414 & ~n4415 ) | ( n4414 & n4775 ) | ( ~n4415 & n4775 ) ;
  assign n4777 = ( n4747 & n4749 ) | ( n4747 & ~n4753 ) | ( n4749 & ~n4753 ) ;
  assign n4778 = ( n4753 & ~n4754 ) | ( n4753 & n4777 ) | ( ~n4754 & n4777 ) ;
  assign n4779 = ( ~n4569 & n4571 ) | ( ~n4569 & n4751 ) | ( n4571 & n4751 ) ;
  assign n4780 = ( n4569 & ~n4752 ) | ( n4569 & n4779 ) | ( ~n4752 & n4779 ) ;
  assign n4781 = ( ~n4230 & n4232 ) | ( ~n4230 & n4412 ) | ( n4232 & n4412 ) ;
  assign n4782 = ( n4230 & ~n4413 ) | ( n4230 & n4781 ) | ( ~n4413 & n4781 ) ;
  assign n4783 = n4780 & n4782 ;
  assign n4784 = ( n4776 & n4778 ) | ( n4776 & n4783 ) | ( n4778 & n4783 ) ;
  assign n4785 = ( n4772 & n4774 ) | ( n4772 & n4784 ) | ( n4774 & n4784 ) ;
  assign n4786 = ( n4768 & n4770 ) | ( n4768 & n4785 ) | ( n4770 & n4785 ) ;
  assign n4787 = ( n4764 & n4766 ) | ( n4764 & n4786 ) | ( n4766 & n4786 ) ;
  assign n4788 = ( n4760 & n4762 ) | ( n4760 & n4787 ) | ( n4762 & n4787 ) ;
  assign n4789 = ( n4419 & n4758 ) | ( n4419 & n4788 ) | ( n4758 & n4788 ) ;
  assign n4790 = ( ~n4419 & n4758 ) | ( ~n4419 & n4788 ) | ( n4758 & n4788 ) ;
  assign n4791 = ( n4419 & ~n4789 ) | ( n4419 & n4790 ) | ( ~n4789 & n4790 ) ;
  assign n4792 = ( ~n3710 & n4049 ) | ( ~n3710 & n4079 ) | ( n4049 & n4079 ) ;
  assign n4793 = ( n3710 & ~n4080 ) | ( n3710 & n4792 ) | ( ~n4080 & n4792 ) ;
  assign n4794 = ( ~n4051 & n4053 ) | ( ~n4051 & n4078 ) | ( n4053 & n4078 ) ;
  assign n4795 = ( n4051 & ~n4079 ) | ( n4051 & n4794 ) | ( ~n4079 & n4794 ) ;
  assign n4796 = ( ~n4760 & n4762 ) | ( ~n4760 & n4787 ) | ( n4762 & n4787 ) ;
  assign n4797 = ( n4760 & ~n4788 ) | ( n4760 & n4796 ) | ( ~n4788 & n4796 ) ;
  assign n4798 = ( ~n4764 & n4766 ) | ( ~n4764 & n4786 ) | ( n4766 & n4786 ) ;
  assign n4799 = ( n4764 & ~n4787 ) | ( n4764 & n4798 ) | ( ~n4787 & n4798 ) ;
  assign n4800 = ( ~n4055 & n4057 ) | ( ~n4055 & n4077 ) | ( n4057 & n4077 ) ;
  assign n4801 = ( n4055 & ~n4078 ) | ( n4055 & n4800 ) | ( ~n4078 & n4800 ) ;
  assign n4802 = ( ~n4059 & n4061 ) | ( ~n4059 & n4076 ) | ( n4061 & n4076 ) ;
  assign n4803 = ( n4059 & ~n4077 ) | ( n4059 & n4802 ) | ( ~n4077 & n4802 ) ;
  assign n4804 = ( ~n4768 & n4770 ) | ( ~n4768 & n4785 ) | ( n4770 & n4785 ) ;
  assign n4805 = ( n4768 & ~n4786 ) | ( n4768 & n4804 ) | ( ~n4786 & n4804 ) ;
  assign n4806 = ( ~n4772 & n4774 ) | ( ~n4772 & n4784 ) | ( n4774 & n4784 ) ;
  assign n4807 = ( n4772 & ~n4785 ) | ( n4772 & n4806 ) | ( ~n4785 & n4806 ) ;
  assign n4808 = ( ~n4063 & n4065 ) | ( ~n4063 & n4075 ) | ( n4065 & n4075 ) ;
  assign n4809 = ( n4063 & ~n4076 ) | ( n4063 & n4808 ) | ( ~n4076 & n4808 ) ;
  assign n4810 = ( ~n4067 & n4069 ) | ( ~n4067 & n4074 ) | ( n4069 & n4074 ) ;
  assign n4811 = ( n4067 & ~n4075 ) | ( n4067 & n4810 ) | ( ~n4075 & n4810 ) ;
  assign n4812 = ( ~n4776 & n4778 ) | ( ~n4776 & n4783 ) | ( n4778 & n4783 ) ;
  assign n4813 = ( n4776 & ~n4784 ) | ( n4776 & n4812 ) | ( ~n4784 & n4812 ) ;
  assign n4814 = n4780 | n4782 ;
  assign n4815 = ~n4783 & n4814 ;
  assign n4816 = ( n4071 & n4073 ) | ( n4071 & n4815 ) | ( n4073 & n4815 ) ;
  assign n4817 = ~n4074 & n4816 ;
  assign n4818 = ( n4811 & n4813 ) | ( n4811 & n4817 ) | ( n4813 & n4817 ) ;
  assign n4819 = ( n4807 & n4809 ) | ( n4807 & n4818 ) | ( n4809 & n4818 ) ;
  assign n4820 = ( n4803 & n4805 ) | ( n4803 & n4819 ) | ( n4805 & n4819 ) ;
  assign n4821 = ( n4799 & n4801 ) | ( n4799 & n4820 ) | ( n4801 & n4820 ) ;
  assign n4822 = ( n4795 & n4797 ) | ( n4795 & n4821 ) | ( n4797 & n4821 ) ;
  assign n4823 = ( n4791 & n4793 ) | ( n4791 & n4822 ) | ( n4793 & n4822 ) ;
  assign n4824 = ( n4080 & n4789 ) | ( n4080 & n4823 ) | ( n4789 & n4823 ) ;
  assign n4825 = ( ~n4080 & n4789 ) | ( ~n4080 & n4823 ) | ( n4789 & n4823 ) ;
  assign n4826 = ( n4080 & ~n4824 ) | ( n4080 & n4825 ) | ( ~n4824 & n4825 ) ;
  assign n4827 = ( ~n2457 & n3332 ) | ( ~n2457 & n3368 ) | ( n3332 & n3368 ) ;
  assign n4828 = ( n2457 & ~n3369 ) | ( n2457 & n4827 ) | ( ~n3369 & n4827 ) ;
  assign n4829 = n4826 & n4828 ;
  assign n4830 = ( ~n3334 & n3338 ) | ( ~n3334 & n3367 ) | ( n3338 & n3367 ) ;
  assign n4831 = ( n3334 & ~n3368 ) | ( n3334 & n4830 ) | ( ~n3368 & n4830 ) ;
  assign n4832 = ( ~n4791 & n4793 ) | ( ~n4791 & n4822 ) | ( n4793 & n4822 ) ;
  assign n4833 = ( n4791 & ~n4823 ) | ( n4791 & n4832 ) | ( ~n4823 & n4832 ) ;
  assign n4834 = ( ~n4071 & n4073 ) | ( ~n4071 & n4815 ) | ( n4073 & n4815 ) ;
  assign n4835 = ( n4071 & ~n4816 ) | ( n4071 & n4834 ) | ( ~n4816 & n4834 ) ;
  assign n4836 = ( ~n2445 & n2447 ) | ( ~n2445 & n3360 ) | ( n2447 & n3360 ) ;
  assign n4837 = ( n2445 & ~n3361 ) | ( n2445 & n4836 ) | ( ~n3361 & n4836 ) ;
  assign n4838 = n4835 & n4837 ;
  assign n4839 = ( ~n3356 & n3358 ) | ( ~n3356 & n3362 ) | ( n3358 & n3362 ) ;
  assign n4840 = ( n3356 & ~n3363 ) | ( n3356 & n4839 ) | ( ~n3363 & n4839 ) ;
  assign n4841 = ( n4811 & n4813 ) | ( n4811 & ~n4817 ) | ( n4813 & ~n4817 ) ;
  assign n4842 = ( n4817 & ~n4818 ) | ( n4817 & n4841 ) | ( ~n4818 & n4841 ) ;
  assign n4843 = ( n4838 & n4840 ) | ( n4838 & n4842 ) | ( n4840 & n4842 ) ;
  assign n4844 = ( ~n3352 & n3354 ) | ( ~n3352 & n3363 ) | ( n3354 & n3363 ) ;
  assign n4845 = ( n3352 & ~n3364 ) | ( n3352 & n4844 ) | ( ~n3364 & n4844 ) ;
  assign n4846 = ( ~n4807 & n4809 ) | ( ~n4807 & n4818 ) | ( n4809 & n4818 ) ;
  assign n4847 = ( n4807 & ~n4819 ) | ( n4807 & n4846 ) | ( ~n4819 & n4846 ) ;
  assign n4848 = ( n4843 & n4845 ) | ( n4843 & n4847 ) | ( n4845 & n4847 ) ;
  assign n4849 = ( ~n3348 & n3350 ) | ( ~n3348 & n3364 ) | ( n3350 & n3364 ) ;
  assign n4850 = ( n3348 & ~n3365 ) | ( n3348 & n4849 ) | ( ~n3365 & n4849 ) ;
  assign n4851 = ( ~n4803 & n4805 ) | ( ~n4803 & n4819 ) | ( n4805 & n4819 ) ;
  assign n4852 = ( n4803 & ~n4820 ) | ( n4803 & n4851 ) | ( ~n4820 & n4851 ) ;
  assign n4853 = ( n4848 & n4850 ) | ( n4848 & n4852 ) | ( n4850 & n4852 ) ;
  assign n4854 = ( ~n3344 & n3346 ) | ( ~n3344 & n3365 ) | ( n3346 & n3365 ) ;
  assign n4855 = ( n3344 & ~n3366 ) | ( n3344 & n4854 ) | ( ~n3366 & n4854 ) ;
  assign n4856 = ( ~n4799 & n4801 ) | ( ~n4799 & n4820 ) | ( n4801 & n4820 ) ;
  assign n4857 = ( n4799 & ~n4821 ) | ( n4799 & n4856 ) | ( ~n4821 & n4856 ) ;
  assign n4858 = ( n4853 & n4855 ) | ( n4853 & n4857 ) | ( n4855 & n4857 ) ;
  assign n4859 = ( ~n3340 & n3342 ) | ( ~n3340 & n3366 ) | ( n3342 & n3366 ) ;
  assign n4860 = ( n3340 & ~n3367 ) | ( n3340 & n4859 ) | ( ~n3367 & n4859 ) ;
  assign n4861 = ( ~n4795 & n4797 ) | ( ~n4795 & n4821 ) | ( n4797 & n4821 ) ;
  assign n4862 = ( n4795 & ~n4822 ) | ( n4795 & n4861 ) | ( ~n4822 & n4861 ) ;
  assign n4863 = ( n4858 & n4860 ) | ( n4858 & n4862 ) | ( n4860 & n4862 ) ;
  assign n4864 = ( n4831 & n4833 ) | ( n4831 & n4863 ) | ( n4833 & n4863 ) ;
  assign n4865 = ( ~n4858 & n4860 ) | ( ~n4858 & n4862 ) | ( n4860 & n4862 ) ;
  assign n4866 = ( n4858 & ~n4863 ) | ( n4858 & n4865 ) | ( ~n4863 & n4865 ) ;
  assign n4867 = ( ~n4848 & n4850 ) | ( ~n4848 & n4852 ) | ( n4850 & n4852 ) ;
  assign n4868 = ( n4848 & ~n4853 ) | ( n4848 & n4867 ) | ( ~n4853 & n4867 ) ;
  assign n4869 = ( ~n4843 & n4845 ) | ( ~n4843 & n4847 ) | ( n4845 & n4847 ) ;
  assign n4870 = ( n4843 & ~n4848 ) | ( n4843 & n4869 ) | ( ~n4848 & n4869 ) ;
  assign n4871 = n4835 | n4837 ;
  assign n4872 = ( x1000 & ~n4838 ) | ( x1000 & n4871 ) | ( ~n4838 & n4871 ) ;
  assign n4873 = ( ~n4838 & n4840 ) | ( ~n4838 & n4842 ) | ( n4840 & n4842 ) ;
  assign n4874 = ( n4838 & ~n4843 ) | ( n4838 & n4873 ) | ( ~n4843 & n4873 ) ;
  assign n4875 = n4872 | n4874 ;
  assign n4876 = n4870 & n4875 ;
  assign n4877 = n4868 | n4876 ;
  assign n4878 = ( ~n4853 & n4855 ) | ( ~n4853 & n4857 ) | ( n4855 & n4857 ) ;
  assign n4879 = ( n4853 & ~n4858 ) | ( n4853 & n4878 ) | ( ~n4858 & n4878 ) ;
  assign n4880 = n4877 & n4879 ;
  assign n4881 = n4866 & n4880 ;
  assign n4882 = ( n4831 & n4833 ) | ( n4831 & ~n4863 ) | ( n4833 & ~n4863 ) ;
  assign n4883 = ( n4863 & ~n4864 ) | ( n4863 & n4882 ) | ( ~n4864 & n4882 ) ;
  assign n4884 = n4881 & n4883 ;
  assign n4885 = n4826 | n4828 ;
  assign n4886 = ( n4864 & n4884 ) | ( n4864 & n4885 ) | ( n4884 & n4885 ) ;
  assign n4887 = n2455 | n3370 ;
  assign n4888 = ( n3369 & ~n3371 ) | ( n3369 & n4887 ) | ( ~n3371 & n4887 ) ;
  assign n4889 = ( n4824 & n4886 ) | ( n4824 & n4888 ) | ( n4886 & n4888 ) ;
  assign n4890 = n4829 | n4889 ;
  assign n4891 = ( n3369 & n4824 ) | ( n3369 & ~n4887 ) | ( n4824 & ~n4887 ) ;
  assign n4892 = n4887 | n4891 ;
  assign n4893 = n4864 & n4884 ;
  assign n4894 = n4892 | n4893 ;
  assign n4895 = ( n3371 & n4890 ) | ( n3371 & n4894 ) | ( n4890 & n4894 ) ;
  assign y0 = n4895 ;
endmodule
