module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 ;
  assign n257 = x126 & ~x254 ;
  assign n258 = x127 | n257 ;
  assign n259 = ~x255 & n258 ;
  assign n260 = x0 | n259 ;
  assign n428 = ~x123 & x250 ;
  assign n429 = x251 | n428 ;
  assign n430 = ~x124 & n429 ;
  assign n431 = x252 | n430 ;
  assign n432 = ~x125 & n431 ;
  assign n261 = x124 | x125 ;
  assign n262 = x123 | n261 ;
  assign n263 = x118 & ~x246 ;
  assign n264 = x119 | n263 ;
  assign n265 = ~x247 & n264 ;
  assign n266 = x120 | n265 ;
  assign n267 = ~x248 & n266 ;
  assign n268 = x121 | n267 ;
  assign n269 = ~x249 & n268 ;
  assign n270 = x122 | n269 ;
  assign n271 = n262 | n270 ;
  assign n272 = x248 | x249 ;
  assign n273 = x247 | n272 ;
  assign n274 = x246 | n273 ;
  assign n275 = x245 | n274 ;
  assign n433 = ~n271 & n275 ;
  assign n434 = n432 | n433 ;
  assign n435 = x253 | n434 ;
  assign n517 = x253 | x254 ;
  assign n518 = x255 | n517 ;
  assign n519 = ( ~x253 & n435 ) | ( ~x253 & n518 ) | ( n435 & n518 ) ;
  assign n276 = x241 | x242 ;
  assign n507 = x112 & ~x240 ;
  assign n508 = x113 | n507 ;
  assign n509 = ~n276 & n508 ;
  assign n510 = ( x114 & ~x242 ) | ( x114 & n509 ) | ( ~x242 & n509 ) ;
  assign n511 = x115 | n510 ;
  assign n277 = x240 | n276 ;
  assign n278 = x239 | n277 ;
  assign n279 = x101 | x102 ;
  assign n280 = x100 | n279 ;
  assign n281 = x99 | n280 ;
  assign n282 = x106 | n281 ;
  assign n283 = x105 | n282 ;
  assign n284 = x104 | n283 ;
  assign n285 = x103 | n284 ;
  assign n286 = x224 | x225 ;
  assign n331 = x95 & ~x223 ;
  assign n332 = x96 | n331 ;
  assign n333 = ~n286 & n332 ;
  assign n334 = ( x97 & ~x225 ) | ( x97 & n333 ) | ( ~x225 & n333 ) ;
  assign n335 = x98 | n334 ;
  assign n287 = x223 | n286 ;
  assign n288 = x222 | n287 ;
  assign n289 = x216 | x217 ;
  assign n319 = x86 & ~x214 ;
  assign n320 = x87 | n319 ;
  assign n321 = ~x215 & n320 ;
  assign n322 = x88 | n321 ;
  assign n323 = ~n289 & n322 ;
  assign n324 = ( x89 & ~x217 ) | ( x89 & n323 ) | ( ~x217 & n323 ) ;
  assign n325 = x90 | n324 ;
  assign n290 = x215 | n289 ;
  assign n291 = x214 | n290 ;
  assign n292 = x213 | n291 ;
  assign n293 = ~x78 & x205 ;
  assign n294 = x206 | n293 ;
  assign n295 = ~x79 & n294 ;
  assign n296 = x207 | n295 ;
  assign n297 = ~x80 & n296 ;
  assign n298 = x209 | n297 ;
  assign n299 = x208 | n298 ;
  assign n300 = ~x74 & x201 ;
  assign n301 = x202 | n300 ;
  assign n302 = ~x75 & n301 ;
  assign n303 = x203 | n302 ;
  assign n304 = ~x76 & n303 ;
  assign n305 = x204 | n304 ;
  assign n306 = x200 | n305 ;
  assign n307 = x199 | n306 ;
  assign n308 = x91 & ~x219 ;
  assign n309 = x92 | n308 ;
  assign n310 = ~x220 & n309 ;
  assign n311 = x93 | n310 ;
  assign n312 = ~x221 & n311 ;
  assign n313 = x220 | x221 ;
  assign n314 = x219 | n313 ;
  assign n315 = x218 | n314 ;
  assign n316 = x84 & ~x212 ;
  assign n317 = x85 | n316 ;
  assign n318 = ~n292 & n317 ;
  assign n326 = n318 | n325 ;
  assign n327 = ~n315 & n326 ;
  assign n328 = n312 | n327 ;
  assign n329 = x94 | n328 ;
  assign n330 = ~n288 & n329 ;
  assign n336 = n330 | n335 ;
  assign n337 = ~x226 & n336 ;
  assign n338 = n285 | n337 ;
  assign n339 = x36 | x37 ;
  assign n340 = x35 | n339 ;
  assign n341 = x34 | n340 ;
  assign n342 = x33 | n341 ;
  assign n343 = x32 | n342 ;
  assign n344 = x40 | x41 ;
  assign n345 = x39 | n344 ;
  assign n346 = x38 | n345 ;
  assign n347 = n343 | n346 ;
  assign n348 = x44 | n347 ;
  assign n349 = x43 | n348 ;
  assign n350 = x42 | n349 ;
  assign n351 = ~x26 & x153 ;
  assign n352 = x154 | n351 ;
  assign n353 = ~x27 & n352 ;
  assign n354 = x155 | n353 ;
  assign n355 = ~x28 & n354 ;
  assign n356 = x156 | n355 ;
  assign n357 = ~x29 & n356 ;
  assign n358 = x157 | n357 ;
  assign n359 = ~x30 & n358 ;
  assign n360 = x158 | n359 ;
  assign n361 = ~x31 & n360 ;
  assign n362 = x159 | n361 ;
  assign n363 = ~n350 & n362 ;
  assign n364 = x196 | x197 ;
  assign n365 = x198 | n364 ;
  assign n366 = x64 & ~x192 ;
  assign n367 = x65 | n366 ;
  assign n368 = ~x193 & n367 ;
  assign n369 = x66 | n368 ;
  assign n370 = x194 | x195 ;
  assign n371 = n369 & ~n370 ;
  assign n372 = ( x67 & ~x195 ) | ( x67 & n371 ) | ( ~x195 & n371 ) ;
  assign n373 = x68 | n372 ;
  assign n374 = ~x62 & x189 ;
  assign n375 = x190 | n374 ;
  assign n376 = ~x63 & n375 ;
  assign n377 = x193 | n370 ;
  assign n378 = x192 | n377 ;
  assign n379 = x191 | n378 ;
  assign n380 = n376 | n379 ;
  assign n381 = n365 | n380 ;
  assign n382 = ( n365 & ~n373 ) | ( n365 & n381 ) | ( ~n373 & n381 ) ;
  assign n383 = x176 | x177 ;
  assign n384 = x175 | n383 ;
  assign n385 = x174 | n384 ;
  assign n386 = x178 | x179 ;
  assign n387 = x173 | n386 ;
  assign n388 = x172 | n387 ;
  assign n389 = n385 | n388 ;
  assign n390 = x187 | x188 ;
  assign n391 = x183 | n390 ;
  assign n392 = x182 | n391 ;
  assign n393 = x181 | n392 ;
  assign n394 = x180 | n393 ;
  assign n395 = x186 | n394 ;
  assign n396 = x185 | n395 ;
  assign n397 = x184 | n396 ;
  assign n398 = n389 | n397 ;
  assign n399 = n382 | n398 ;
  assign n400 = x170 | x171 ;
  assign n401 = x169 | n400 ;
  assign n402 = x168 | n401 ;
  assign n403 = x167 | n402 ;
  assign n404 = ~x33 & x160 ;
  assign n405 = x161 | n404 ;
  assign n406 = ~x34 & n405 ;
  assign n407 = x165 | x166 ;
  assign n408 = x164 | n407 ;
  assign n409 = x163 | n408 ;
  assign n410 = x162 | n409 ;
  assign n411 = n406 | n410 ;
  assign n412 = ( ~x163 & n339 ) | ( ~x163 & n340 ) | ( n339 & n340 ) ;
  assign n413 = ( x37 & ~x164 ) | ( x37 & n412 ) | ( ~x164 & n412 ) ;
  assign n414 = ~n407 & n413 ;
  assign n415 = ( x38 & ~x166 ) | ( x38 & n414 ) | ( ~x166 & n414 ) ;
  assign n416 = x39 | n415 ;
  assign n417 = n411 & ~n416 ;
  assign n418 = n403 | n417 ;
  assign n419 = ( x41 & ~x168 ) | ( x41 & n344 ) | ( ~x168 & n344 ) ;
  assign n420 = ~x169 & n419 ;
  assign n421 = x42 | n420 ;
  assign n422 = ~n400 & n421 ;
  assign n423 = ( x43 & ~x171 ) | ( x43 & n422 ) | ( ~x171 & n422 ) ;
  assign n424 = x44 | n423 ;
  assign n425 = n418 & ~n424 ;
  assign n426 = n399 | n425 ;
  assign n427 = n363 | n426 ;
  assign n436 = ( x254 & ~n257 ) | ( x254 & n435 ) | ( ~n257 & n435 ) ;
  assign n437 = ~x127 & n436 ;
  assign n438 = x151 | x152 ;
  assign n439 = x150 | n438 ;
  assign n440 = x149 | n439 ;
  assign n441 = x148 | n440 ;
  assign n442 = x147 | n441 ;
  assign n443 = x141 | x142 ;
  assign n444 = x140 | n443 ;
  assign n445 = x145 | x146 ;
  assign n446 = x144 | n445 ;
  assign n447 = x143 | n446 ;
  assign n448 = x138 | x139 ;
  assign n449 = x137 | n448 ;
  assign n450 = x136 | n449 ;
  assign n451 = x135 | n450 ;
  assign n452 = x134 | n451 ;
  assign n453 = x132 | x133 ;
  assign n454 = x131 | n453 ;
  assign n455 = x130 | n454 ;
  assign n456 = x129 | n455 ;
  assign n457 = n452 | n456 ;
  assign n458 = n447 | n457 ;
  assign n459 = n444 | n458 ;
  assign n460 = n442 | n459 ;
  assign n461 = x237 | x238 ;
  assign n462 = x236 | n461 ;
  assign n463 = x235 | n462 ;
  assign n464 = x234 | n463 ;
  assign n465 = x128 | n464 ;
  assign n466 = n278 | n465 ;
  assign n467 = x255 | n466 ;
  assign n468 = x244 | n467 ;
  assign n469 = x243 | n468 ;
  assign n470 = x227 | x228 ;
  assign n471 = ( ~x100 & x228 ) | ( ~x100 & n470 ) | ( x228 & n470 ) ;
  assign n472 = ~x101 & n471 ;
  assign n473 = x229 | n472 ;
  assign n474 = ~x102 & n473 ;
  assign n475 = x230 | n474 ;
  assign n476 = ~x103 & n475 ;
  assign n477 = x231 | x232 ;
  assign n478 = n476 | n477 ;
  assign n479 = ( ~x104 & x232 ) | ( ~x104 & n478 ) | ( x232 & n478 ) ;
  assign n480 = ~x105 & n479 ;
  assign n481 = x233 | n480 ;
  assign n482 = ~x106 & n481 ;
  assign n483 = n469 | n482 ;
  assign n484 = n460 | n483 ;
  assign n485 = n437 | n484 ;
  assign n486 = n427 | n485 ;
  assign n487 = n338 & ~n486 ;
  assign n488 = x31 | n350 ;
  assign n489 = x30 | n488 ;
  assign n490 = x29 | n489 ;
  assign n491 = x28 | n490 ;
  assign n492 = x27 | n491 ;
  assign n493 = x121 | x122 ;
  assign n494 = x120 | n493 ;
  assign n495 = x119 | n494 ;
  assign n496 = x118 | n495 ;
  assign n497 = x117 | n496 ;
  assign n498 = n262 | n497 ;
  assign n499 = x107 & ~x235 ;
  assign n500 = x108 | n499 ;
  assign n501 = ~x236 & n500 ;
  assign n502 = x109 | n501 ;
  assign n503 = ~n461 & n502 ;
  assign n504 = ( x110 & ~x238 ) | ( x110 & n503 ) | ( ~x238 & n503 ) ;
  assign n505 = x111 | n504 ;
  assign n506 = ~n278 & n505 ;
  assign n512 = n506 | n511 ;
  assign n513 = ~x243 & n512 ;
  assign n514 = x116 | n513 ;
  assign n515 = ~x244 & n514 ;
  assign n516 = n498 | n515 ;
  assign n520 = n516 & ~n519 ;
  assign n521 = n260 | n520 ;
  assign n522 = ~x128 & n521 ;
  assign n523 = x1 | n522 ;
  assign n524 = ~n460 & n523 ;
  assign n525 = x20 & ~x148 ;
  assign n526 = x21 | n525 ;
  assign n527 = ~x149 & n526 ;
  assign n528 = x22 | n527 ;
  assign n529 = ~x150 & n528 ;
  assign n530 = x23 | n529 ;
  assign n531 = ~x151 & n530 ;
  assign n532 = x24 | n531 ;
  assign n533 = x13 & ~x141 ;
  assign n534 = x14 | n533 ;
  assign n535 = x2 & ~x130 ;
  assign n536 = x3 | n535 ;
  assign n537 = ~x131 & n536 ;
  assign n538 = x4 | n537 ;
  assign n539 = ~n453 & n538 ;
  assign n540 = ( x5 & ~x133 ) | ( x5 & n539 ) | ( ~x133 & n539 ) ;
  assign n541 = x6 | n540 ;
  assign n542 = ~n452 & n541 ;
  assign n543 = x7 & ~x135 ;
  assign n544 = x8 | n543 ;
  assign n545 = ~x136 & n544 ;
  assign n546 = x9 | n545 ;
  assign n547 = ~x137 & n546 ;
  assign n548 = x10 | n547 ;
  assign n549 = ~n448 & n548 ;
  assign n550 = ( x11 & ~x139 ) | ( x11 & n549 ) | ( ~x139 & n549 ) ;
  assign n551 = x12 | n550 ;
  assign n552 = n542 | n551 ;
  assign n553 = ~n444 & n552 ;
  assign n554 = ( ~x142 & n534 ) | ( ~x142 & n553 ) | ( n534 & n553 ) ;
  assign n555 = x15 | n554 ;
  assign n556 = ~n447 & n555 ;
  assign n557 = x16 & ~x144 ;
  assign n558 = x17 | n557 ;
  assign n559 = ~n445 & n558 ;
  assign n560 = ( x18 & ~x146 ) | ( x18 & n559 ) | ( ~x146 & n559 ) ;
  assign n561 = x19 | n560 ;
  assign n562 = n556 | n561 ;
  assign n563 = ~n442 & n562 ;
  assign n564 = ( ~x152 & n532 ) | ( ~x152 & n563 ) | ( n532 & n563 ) ;
  assign n565 = n524 | n564 ;
  assign n566 = x26 | n565 ;
  assign n567 = x25 | n566 ;
  assign n568 = n492 | n567 ;
  assign n569 = ~n427 & n568 ;
  assign n570 = x60 & ~x188 ;
  assign n571 = x64 | n570 ;
  assign n572 = x63 | n571 ;
  assign n573 = x62 | n572 ;
  assign n574 = x61 | n573 ;
  assign n575 = x68 | n574 ;
  assign n576 = x67 | n575 ;
  assign n577 = x66 | n576 ;
  assign n578 = x65 | n577 ;
  assign n579 = x53 & ~x181 ;
  assign n580 = x54 | n579 ;
  assign n581 = ~x182 & n580 ;
  assign n582 = x55 | n581 ;
  assign n583 = ~x183 & n582 ;
  assign n584 = x56 | n583 ;
  assign n585 = ~x184 & n584 ;
  assign n586 = x57 | n585 ;
  assign n587 = ~x185 & n586 ;
  assign n588 = x58 | n587 ;
  assign n589 = ~x186 & n588 ;
  assign n590 = x59 | n589 ;
  assign n591 = x45 & ~x173 ;
  assign n592 = x46 | n591 ;
  assign n593 = ~x174 & n592 ;
  assign n594 = x47 | n593 ;
  assign n595 = ~x175 & n594 ;
  assign n596 = x48 | n595 ;
  assign n597 = ~n383 & n596 ;
  assign n598 = ( x49 & ~x177 ) | ( x49 & n597 ) | ( ~x177 & n597 ) ;
  assign n599 = x50 | n598 ;
  assign n600 = ~n386 & n599 ;
  assign n601 = ( x51 & ~x179 ) | ( x51 & n600 ) | ( ~x179 & n600 ) ;
  assign n602 = x52 | n601 ;
  assign n603 = ~n397 & n602 ;
  assign n604 = ( ~n390 & n590 ) | ( ~n390 & n603 ) | ( n590 & n603 ) ;
  assign n605 = n578 | n604 ;
  assign n606 = ( ~n382 & n569 ) | ( ~n382 & n605 ) | ( n569 & n605 ) ;
  assign n607 = n487 | n606 ;
  assign n608 = ~n307 & n607 ;
  assign n609 = x79 | x80 ;
  assign n610 = x78 | n609 ;
  assign n611 = x77 | n610 ;
  assign n612 = x75 | x76 ;
  assign n613 = x74 | n612 ;
  assign n614 = x73 | n613 ;
  assign n615 = x69 & ~x197 ;
  assign n616 = x70 | n615 ;
  assign n617 = ~x198 & n616 ;
  assign n618 = x71 | n617 ;
  assign n619 = ~x199 & n618 ;
  assign n620 = x72 | n619 ;
  assign n621 = ~n306 & n620 ;
  assign n622 = ( ~n305 & n614 ) | ( ~n305 & n621 ) | ( n614 & n621 ) ;
  assign n623 = n611 | n622 ;
  assign n624 = n608 | n623 ;
  assign n625 = ~n299 & n624 ;
  assign n626 = ( x81 & ~x209 ) | ( x81 & n625 ) | ( ~x209 & n625 ) ;
  assign n627 = x82 | n626 ;
  assign n628 = ~x210 & n627 ;
  assign n629 = x83 | n628 ;
  assign n630 = ~x211 & n629 ;
  assign n631 = x84 | n630 ;
  assign n632 = ~x212 & n631 ;
  assign n633 = x85 | n632 ;
  assign n634 = ~n292 & n633 ;
  assign n635 = n325 | n634 ;
  assign n636 = ~x218 & n635 ;
  assign n637 = x91 | n636 ;
  assign n638 = ~x219 & n637 ;
  assign n639 = x92 | n638 ;
  assign n640 = ~x220 & n639 ;
  assign n641 = x93 | n640 ;
  assign n642 = ~x221 & n641 ;
  assign n643 = x94 | n642 ;
  assign n644 = ~n288 & n643 ;
  assign n645 = n335 | n644 ;
  assign n646 = ~x226 & n645 ;
  assign n647 = n285 | n646 ;
  assign n648 = x234 | n482 ;
  assign n649 = n647 & ~n648 ;
  assign n650 = x107 | n649 ;
  assign n651 = ~x235 & n650 ;
  assign n652 = x108 | n651 ;
  assign n653 = ~x236 & n652 ;
  assign n654 = x109 | n653 ;
  assign n655 = ~x237 & n654 ;
  assign n656 = x110 | n655 ;
  assign n657 = ~x238 & n656 ;
  assign n658 = x111 | n657 ;
  assign n659 = ~n278 & n658 ;
  assign n660 = n511 | n659 ;
  assign n661 = ~x243 & n660 ;
  assign n662 = x116 | n661 ;
  assign n663 = ~x244 & n662 ;
  assign n664 = x117 | n663 ;
  assign n665 = ~n275 & n664 ;
  assign n666 = n271 | n665 ;
  assign n667 = ~n519 & n666 ;
  assign n668 = n260 | n667 ;
  assign n669 = x128 & n668 ;
  assign n670 = ~x128 & n668 ;
  assign n671 = x1 | n670 ;
  assign n672 = x129 & n671 ;
  assign n673 = ~x129 & n671 ;
  assign n674 = x2 | n673 ;
  assign n675 = x130 & n674 ;
  assign n676 = ~x130 & n674 ;
  assign n677 = x3 | n676 ;
  assign n678 = x131 & n677 ;
  assign n679 = ~x131 & n677 ;
  assign n680 = x4 | n679 ;
  assign n681 = x132 & n680 ;
  assign n682 = ~x132 & n680 ;
  assign n683 = x5 | n682 ;
  assign n684 = x133 & n683 ;
  assign n685 = ~n456 & n671 ;
  assign n686 = n541 | n685 ;
  assign n687 = x134 & n686 ;
  assign n688 = ~x134 & n686 ;
  assign n689 = x7 | n688 ;
  assign n690 = x135 & n689 ;
  assign n691 = ~x135 & n689 ;
  assign n692 = x8 | n691 ;
  assign n693 = x136 & n692 ;
  assign n694 = ~x136 & n692 ;
  assign n695 = x9 | n694 ;
  assign n696 = x137 & n695 ;
  assign n697 = ~x137 & n695 ;
  assign n698 = x10 | n697 ;
  assign n699 = x138 & n698 ;
  assign n700 = ~x138 & n698 ;
  assign n701 = x11 | n700 ;
  assign n702 = x139 & n701 ;
  assign n703 = ~x139 & n701 ;
  assign n704 = x12 | n703 ;
  assign n705 = x140 & n704 ;
  assign n706 = ~x140 & n704 ;
  assign n707 = x13 | n706 ;
  assign n708 = x141 & n707 ;
  assign n709 = ~x141 & n707 ;
  assign n710 = x14 | n709 ;
  assign n711 = x142 & n710 ;
  assign n712 = ~x142 & n710 ;
  assign n713 = x15 | n712 ;
  assign n714 = x143 & n713 ;
  assign n715 = ~x143 & n713 ;
  assign n716 = x16 | n715 ;
  assign n717 = x144 & n716 ;
  assign n718 = ~x144 & n716 ;
  assign n719 = x17 | n718 ;
  assign n720 = x145 & n719 ;
  assign n721 = ~x145 & n719 ;
  assign n722 = x18 | n721 ;
  assign n723 = x146 & n722 ;
  assign n724 = ~n447 & n713 ;
  assign n725 = n561 | n724 ;
  assign n726 = x147 & n725 ;
  assign n727 = ~x147 & n725 ;
  assign n728 = x20 | n727 ;
  assign n729 = x148 & n728 ;
  assign n730 = ~x148 & n728 ;
  assign n731 = x21 | n730 ;
  assign n732 = x149 & n731 ;
  assign n733 = ~x149 & n731 ;
  assign n734 = x22 | n733 ;
  assign n735 = x150 & n734 ;
  assign n736 = ~x150 & n734 ;
  assign n737 = x23 | n736 ;
  assign n738 = x151 & n737 ;
  assign n739 = ~x151 & n737 ;
  assign n740 = x24 | n739 ;
  assign n741 = x152 & n740 ;
  assign n742 = ~x152 & n740 ;
  assign n743 = x25 | n742 ;
  assign n744 = x153 & n743 ;
  assign n745 = ( x26 & ~n351 ) | ( x26 & n743 ) | ( ~n351 & n743 ) ;
  assign n746 = x154 & n745 ;
  assign n747 = n352 | n485 ;
  assign n748 = n647 & ~n747 ;
  assign n749 = ( ~n352 & n567 ) | ( ~n352 & n748 ) | ( n567 & n748 ) ;
  assign n750 = x27 | n749 ;
  assign n751 = x155 & n750 ;
  assign n752 = ~x155 & n750 ;
  assign n753 = x28 | n752 ;
  assign n754 = x156 & n753 ;
  assign n755 = ~x156 & n753 ;
  assign n756 = x29 | n755 ;
  assign n757 = x157 & n756 ;
  assign n758 = ~x157 & n756 ;
  assign n759 = x30 | n758 ;
  assign n760 = x158 & n759 ;
  assign n761 = ~x158 & n759 ;
  assign n762 = x31 | n761 ;
  assign n763 = x159 & n762 ;
  assign n764 = ~x159 & n762 ;
  assign n765 = x32 | n764 ;
  assign n766 = x160 & n765 ;
  assign n767 = ( x33 & ~n404 ) | ( x33 & n765 ) | ( ~n404 & n765 ) ;
  assign n768 = x161 & n767 ;
  assign n769 = ( x34 & ~n406 ) | ( x34 & n767 ) | ( ~n406 & n767 ) ;
  assign n770 = x162 & n769 ;
  assign n771 = ~x162 & n769 ;
  assign n772 = x35 | n771 ;
  assign n773 = x163 & n772 ;
  assign n774 = ~x163 & n772 ;
  assign n775 = x36 | n774 ;
  assign n776 = x164 & n775 ;
  assign n777 = ~x164 & n775 ;
  assign n778 = x37 | n777 ;
  assign n779 = x165 & n778 ;
  assign n780 = ~x165 & n778 ;
  assign n781 = x38 | n780 ;
  assign n782 = x166 & n781 ;
  assign n783 = ( n416 & ~n417 ) | ( n416 & n769 ) | ( ~n417 & n769 ) ;
  assign n784 = x167 & n783 ;
  assign n785 = ~x167 & n783 ;
  assign n786 = x40 | n785 ;
  assign n787 = x168 & n786 ;
  assign n788 = ~x168 & n786 ;
  assign n789 = x41 | n788 ;
  assign n790 = x169 & n789 ;
  assign n791 = ~x169 & n789 ;
  assign n792 = x42 | n791 ;
  assign n793 = x170 & n792 ;
  assign n794 = ~x170 & n792 ;
  assign n795 = x43 | n794 ;
  assign n796 = x171 & n795 ;
  assign n797 = ( n424 & ~n425 ) | ( n424 & n783 ) | ( ~n425 & n783 ) ;
  assign n798 = x172 & n797 ;
  assign n799 = ~x172 & n797 ;
  assign n800 = x45 | n799 ;
  assign n801 = x173 & n800 ;
  assign n802 = ~x173 & n800 ;
  assign n803 = x46 | n802 ;
  assign n804 = x174 & n803 ;
  assign n805 = ~x174 & n803 ;
  assign n806 = x47 | n805 ;
  assign n807 = x175 & n806 ;
  assign n808 = ~x175 & n806 ;
  assign n809 = x48 | n808 ;
  assign n810 = x176 & n809 ;
  assign n811 = ~x176 & n809 ;
  assign n812 = x49 | n811 ;
  assign n813 = x177 & n812 ;
  assign n814 = ~x177 & n812 ;
  assign n815 = x50 | n814 ;
  assign n816 = x178 & n815 ;
  assign n817 = ~x178 & n815 ;
  assign n818 = x51 | n817 ;
  assign n819 = x179 & n818 ;
  assign n820 = ~n389 & n797 ;
  assign n821 = n602 | n820 ;
  assign n822 = x180 & n821 ;
  assign n823 = ~x180 & n821 ;
  assign n824 = x53 | n823 ;
  assign n825 = x181 & n824 ;
  assign n826 = ~x181 & n824 ;
  assign n827 = x54 | n826 ;
  assign n828 = x182 & n827 ;
  assign n829 = ~x182 & n827 ;
  assign n830 = x55 | n829 ;
  assign n831 = x183 & n830 ;
  assign n832 = ~x183 & n830 ;
  assign n833 = x56 | n832 ;
  assign n834 = x184 & n833 ;
  assign n835 = ~x184 & n833 ;
  assign n836 = x57 | n835 ;
  assign n837 = x185 & n836 ;
  assign n838 = ~x185 & n836 ;
  assign n839 = x58 | n838 ;
  assign n840 = x186 & n839 ;
  assign n841 = ~x186 & n839 ;
  assign n842 = x59 | n841 ;
  assign n843 = x187 & n842 ;
  assign n844 = ~x187 & n842 ;
  assign n845 = x60 | n844 ;
  assign n846 = x188 & n845 ;
  assign n847 = ~x188 & n845 ;
  assign n848 = x61 | n847 ;
  assign n849 = x189 & n848 ;
  assign n850 = ( x62 & ~n374 ) | ( x62 & n848 ) | ( ~n374 & n848 ) ;
  assign n851 = x190 & n850 ;
  assign n852 = ( x63 & ~n376 ) | ( x63 & n850 ) | ( ~n376 & n850 ) ;
  assign n853 = x191 & n852 ;
  assign n854 = ~x191 & n852 ;
  assign n855 = x64 | n854 ;
  assign n856 = x192 & n855 ;
  assign n857 = ~x192 & n855 ;
  assign n858 = x65 | n857 ;
  assign n859 = x193 & n858 ;
  assign n860 = ~x193 & n858 ;
  assign n861 = x66 | n860 ;
  assign n862 = x194 & n861 ;
  assign n863 = ~x194 & n861 ;
  assign n864 = x67 | n863 ;
  assign n865 = x195 & n864 ;
  assign n866 = ~n379 & n852 ;
  assign n867 = n373 | n866 ;
  assign n868 = x196 & n867 ;
  assign n869 = ~x196 & n867 ;
  assign n870 = x69 | n869 ;
  assign n871 = x197 & n870 ;
  assign n872 = ~x197 & n870 ;
  assign n873 = x70 | n872 ;
  assign n874 = x198 & n873 ;
  assign n875 = ~n486 & n646 ;
  assign n876 = n607 | n618 ;
  assign n877 = n875 | n876 ;
  assign n878 = x199 & n877 ;
  assign n879 = ~x199 & n877 ;
  assign n880 = x72 | n879 ;
  assign n881 = x200 & n880 ;
  assign n882 = ~x200 & n880 ;
  assign n883 = x73 | n882 ;
  assign n884 = x201 & n883 ;
  assign n885 = ( x74 & ~n300 ) | ( x74 & n883 ) | ( ~n300 & n883 ) ;
  assign n886 = x202 & n885 ;
  assign n887 = ( x75 & ~n302 ) | ( x75 & n885 ) | ( ~n302 & n885 ) ;
  assign n888 = x203 & n887 ;
  assign n889 = n614 | n882 ;
  assign n890 = ~n304 & n889 ;
  assign n891 = x204 & n890 ;
  assign n892 = ~x204 & n890 ;
  assign n893 = x77 | n892 ;
  assign n894 = x205 & n893 ;
  assign n895 = ( x78 & ~n293 ) | ( x78 & n893 ) | ( ~n293 & n893 ) ;
  assign n896 = x206 & n895 ;
  assign n897 = ( x79 & ~n295 ) | ( x79 & n895 ) | ( ~n295 & n895 ) ;
  assign n898 = x207 & n897 ;
  assign n899 = n623 | n892 ;
  assign n900 = ~n297 & n899 ;
  assign n901 = x208 & n900 ;
  assign n902 = ~x208 & n900 ;
  assign n903 = x81 | n902 ;
  assign n904 = x209 & n903 ;
  assign n905 = ~n299 & n893 ;
  assign n906 = n627 | n905 ;
  assign n907 = x210 & n906 ;
  assign n908 = x211 & n629 ;
  assign n909 = x212 & n631 ;
  assign n910 = x213 & n633 ;
  assign n911 = ~x213 & n633 ;
  assign n912 = x86 | n911 ;
  assign n913 = x214 & n912 ;
  assign n914 = ~x214 & n912 ;
  assign n915 = x87 | n914 ;
  assign n916 = x215 & n915 ;
  assign n917 = ~x215 & n915 ;
  assign n918 = x88 | n917 ;
  assign n919 = x216 & n918 ;
  assign n920 = ~x216 & n918 ;
  assign n921 = x89 | n920 ;
  assign n922 = x217 & n921 ;
  assign n923 = x218 & n635 ;
  assign n924 = x219 & n637 ;
  assign n925 = x220 & n639 ;
  assign n926 = x221 & n641 ;
  assign n927 = x222 & n643 ;
  assign n928 = ~x222 & n643 ;
  assign n929 = x95 | n928 ;
  assign n930 = x223 & n929 ;
  assign n931 = ~x223 & n929 ;
  assign n932 = x96 | n931 ;
  assign n933 = x224 & n932 ;
  assign n934 = ~x224 & n932 ;
  assign n935 = x97 | n934 ;
  assign n936 = x225 & n935 ;
  assign n937 = x226 & n645 ;
  assign n938 = x99 | n646 ;
  assign n939 = x227 & n938 ;
  assign n940 = ~x227 & n938 ;
  assign n941 = x100 | n940 ;
  assign n942 = x228 & n941 ;
  assign n943 = ( x101 & ~n472 ) | ( x101 & n941 ) | ( ~n472 & n941 ) ;
  assign n944 = x229 & n943 ;
  assign n945 = ( x102 & ~n474 ) | ( x102 & n943 ) | ( ~n474 & n943 ) ;
  assign n946 = x230 & n945 ;
  assign n947 = x102 | n943 ;
  assign n948 = ~n475 & n947 ;
  assign n949 = x103 | n948 ;
  assign n950 = x231 & n949 ;
  assign n951 = ~x231 & n949 ;
  assign n952 = x104 | n951 ;
  assign n953 = x232 & n952 ;
  assign n954 = ~x232 & n952 ;
  assign n955 = x105 | n954 ;
  assign n956 = x233 & n955 ;
  assign n957 = ~n482 & n647 ;
  assign n958 = x234 & n957 ;
  assign n959 = x235 & n650 ;
  assign n960 = x236 & n652 ;
  assign n961 = x237 & n654 ;
  assign n962 = x238 & n656 ;
  assign n963 = x239 & n658 ;
  assign n964 = ~x239 & n658 ;
  assign n965 = x112 | n964 ;
  assign n966 = x240 & n965 ;
  assign n967 = ~x240 & n965 ;
  assign n968 = x113 | n967 ;
  assign n969 = x241 & n968 ;
  assign n970 = ~x241 & n968 ;
  assign n971 = x114 | n970 ;
  assign n972 = x242 & n971 ;
  assign n973 = x243 & n660 ;
  assign n974 = x244 & n662 ;
  assign n975 = x245 & n664 ;
  assign n976 = ~x245 & n664 ;
  assign n977 = x118 | n976 ;
  assign n978 = x246 & n977 ;
  assign n979 = ~x246 & n977 ;
  assign n980 = x119 | n979 ;
  assign n981 = x247 & n980 ;
  assign n982 = ~x247 & n980 ;
  assign n983 = x120 | n982 ;
  assign n984 = x248 & n983 ;
  assign n985 = ~x248 & n983 ;
  assign n986 = x121 | n985 ;
  assign n987 = x249 & n986 ;
  assign n988 = n270 | n665 ;
  assign n989 = x250 & n988 ;
  assign n990 = ( x123 & ~n428 ) | ( x123 & n988 ) | ( ~n428 & n988 ) ;
  assign n991 = x251 & n990 ;
  assign n992 = ( x124 & ~n430 ) | ( x124 & n990 ) | ( ~n430 & n990 ) ;
  assign n993 = x252 & n992 ;
  assign n994 = ~n432 & n666 ;
  assign n995 = x253 & n994 ;
  assign n996 = ~x253 & n994 ;
  assign n997 = x126 | n996 ;
  assign n998 = x254 & n997 ;
  assign n999 = x127 | n498 ;
  assign n1000 = x126 | n999 ;
  assign n1001 = n988 | n1000 ;
  assign n1002 = ~n437 & n1001 ;
  assign n1003 = x255 & n1002 ;
  assign n1004 = x190 | x201 ;
  assign n1005 = x189 | n1004 ;
  assign n1006 = x161 | n1005 ;
  assign n1007 = x205 | n1006 ;
  assign n1008 = x204 | n1007 ;
  assign n1009 = x203 | n1008 ;
  assign n1010 = x202 | n1009 ;
  assign n1011 = x226 | n470 ;
  assign n1012 = x212 | n1011 ;
  assign n1013 = n1010 | n1012 ;
  assign n1014 = x211 | n1013 ;
  assign n1015 = x210 | n1014 ;
  assign n1016 = x207 | n1015 ;
  assign n1017 = x206 | n1016 ;
  assign n1018 = x209 | n517 ;
  assign n1019 = x208 | n1018 ;
  assign n1020 = x200 | n1019 ;
  assign n1021 = x199 | n1020 ;
  assign n1022 = x159 | x160 ;
  assign n1023 = x158 | n1022 ;
  assign n1024 = x157 | n1023 ;
  assign n1025 = n1021 | n1024 ;
  assign n1026 = x156 | n1025 ;
  assign n1027 = x155 | n1026 ;
  assign n1028 = x154 | n1027 ;
  assign n1029 = x153 | n1028 ;
  assign n1030 = x230 | n477 ;
  assign n1031 = x229 | n1030 ;
  assign n1032 = x252 | n1031 ;
  assign n1033 = x251 | n1032 ;
  assign n1034 = x250 | n1033 ;
  assign n1035 = x233 | n1034 ;
  assign n1036 = n288 | n1035 ;
  assign n1037 = n365 | n1036 ;
  assign n1038 = n315 | n1037 ;
  assign n1039 = n292 | n1038 ;
  assign n1040 = n379 | n398 ;
  assign n1041 = n403 | n1040 ;
  assign n1042 = n410 | n1041 ;
  assign n1043 = n275 | n1042 ;
  assign n1044 = n1039 | n1043 ;
  assign n1045 = n1029 | n1044 ;
  assign n1046 = n1017 | n1045 ;
  assign n1047 = n469 | n1046 ;
  assign n1048 = n460 | n1047 ;
  assign y0 = n669 ;
  assign y1 = n672 ;
  assign y2 = n675 ;
  assign y3 = n678 ;
  assign y4 = n681 ;
  assign y5 = n684 ;
  assign y6 = n687 ;
  assign y7 = n690 ;
  assign y8 = n693 ;
  assign y9 = n696 ;
  assign y10 = n699 ;
  assign y11 = n702 ;
  assign y12 = n705 ;
  assign y13 = n708 ;
  assign y14 = n711 ;
  assign y15 = n714 ;
  assign y16 = n717 ;
  assign y17 = n720 ;
  assign y18 = n723 ;
  assign y19 = n726 ;
  assign y20 = n729 ;
  assign y21 = n732 ;
  assign y22 = n735 ;
  assign y23 = n738 ;
  assign y24 = n741 ;
  assign y25 = n744 ;
  assign y26 = n746 ;
  assign y27 = n751 ;
  assign y28 = n754 ;
  assign y29 = n757 ;
  assign y30 = n760 ;
  assign y31 = n763 ;
  assign y32 = n766 ;
  assign y33 = n768 ;
  assign y34 = n770 ;
  assign y35 = n773 ;
  assign y36 = n776 ;
  assign y37 = n779 ;
  assign y38 = n782 ;
  assign y39 = n784 ;
  assign y40 = n787 ;
  assign y41 = n790 ;
  assign y42 = n793 ;
  assign y43 = n796 ;
  assign y44 = n798 ;
  assign y45 = n801 ;
  assign y46 = n804 ;
  assign y47 = n807 ;
  assign y48 = n810 ;
  assign y49 = n813 ;
  assign y50 = n816 ;
  assign y51 = n819 ;
  assign y52 = n822 ;
  assign y53 = n825 ;
  assign y54 = n828 ;
  assign y55 = n831 ;
  assign y56 = n834 ;
  assign y57 = n837 ;
  assign y58 = n840 ;
  assign y59 = n843 ;
  assign y60 = n846 ;
  assign y61 = n849 ;
  assign y62 = n851 ;
  assign y63 = n853 ;
  assign y64 = n856 ;
  assign y65 = n859 ;
  assign y66 = n862 ;
  assign y67 = n865 ;
  assign y68 = n868 ;
  assign y69 = n871 ;
  assign y70 = n874 ;
  assign y71 = n878 ;
  assign y72 = n881 ;
  assign y73 = n884 ;
  assign y74 = n886 ;
  assign y75 = n888 ;
  assign y76 = n891 ;
  assign y77 = n894 ;
  assign y78 = n896 ;
  assign y79 = n898 ;
  assign y80 = n901 ;
  assign y81 = n904 ;
  assign y82 = n907 ;
  assign y83 = n908 ;
  assign y84 = n909 ;
  assign y85 = n910 ;
  assign y86 = n913 ;
  assign y87 = n916 ;
  assign y88 = n919 ;
  assign y89 = n922 ;
  assign y90 = n923 ;
  assign y91 = n924 ;
  assign y92 = n925 ;
  assign y93 = n926 ;
  assign y94 = n927 ;
  assign y95 = n930 ;
  assign y96 = n933 ;
  assign y97 = n936 ;
  assign y98 = n937 ;
  assign y99 = n939 ;
  assign y100 = n942 ;
  assign y101 = n944 ;
  assign y102 = n946 ;
  assign y103 = n950 ;
  assign y104 = n953 ;
  assign y105 = n956 ;
  assign y106 = n958 ;
  assign y107 = n959 ;
  assign y108 = n960 ;
  assign y109 = n961 ;
  assign y110 = n962 ;
  assign y111 = n963 ;
  assign y112 = n966 ;
  assign y113 = n969 ;
  assign y114 = n972 ;
  assign y115 = n973 ;
  assign y116 = n974 ;
  assign y117 = n975 ;
  assign y118 = n978 ;
  assign y119 = n981 ;
  assign y120 = n984 ;
  assign y121 = n987 ;
  assign y122 = n989 ;
  assign y123 = n991 ;
  assign y124 = n993 ;
  assign y125 = n995 ;
  assign y126 = n998 ;
  assign y127 = n1003 ;
  assign y128 = n1048 ;
endmodule
