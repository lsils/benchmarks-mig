module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 ;
  assign n136 = x106 & ~x128 ;
  assign n137 = x105 & ~x128 ;
  assign n138 = ( x105 & n136 ) | ( x105 & ~n137 ) | ( n136 & ~n137 ) ;
  assign n139 = x129 & ~n138 ;
  assign n140 = x107 & x128 ;
  assign n141 = x108 & ~x128 ;
  assign n142 = ( x129 & ~n140 ) | ( x129 & n141 ) | ( ~n140 & n141 ) ;
  assign n143 = ( ~n139 & n140 ) | ( ~n139 & n142 ) | ( n140 & n142 ) ;
  assign n144 = x98 & ~x128 ;
  assign n145 = x97 & ~x128 ;
  assign n146 = ( x97 & n144 ) | ( x97 & ~n145 ) | ( n144 & ~n145 ) ;
  assign n147 = x129 & ~n146 ;
  assign n148 = x99 & x128 ;
  assign n149 = x100 & ~x128 ;
  assign n150 = ( x129 & ~n148 ) | ( x129 & n149 ) | ( ~n148 & n149 ) ;
  assign n151 = ( ~n147 & n148 ) | ( ~n147 & n150 ) | ( n148 & n150 ) ;
  assign n152 = x131 & ~n151 ;
  assign n153 = x131 & ~n143 ;
  assign n154 = ( n143 & ~n152 ) | ( n143 & n153 ) | ( ~n152 & n153 ) ;
  assign n155 = x130 & ~n154 ;
  assign n156 = x110 & ~x128 ;
  assign n157 = x109 & ~x128 ;
  assign n158 = ( x109 & n156 ) | ( x109 & ~n157 ) | ( n156 & ~n157 ) ;
  assign n159 = x129 & ~n158 ;
  assign n160 = x111 & x128 ;
  assign n161 = x112 & ~x128 ;
  assign n162 = ( x129 & ~n160 ) | ( x129 & n161 ) | ( ~n160 & n161 ) ;
  assign n163 = ( ~n159 & n160 ) | ( ~n159 & n162 ) | ( n160 & n162 ) ;
  assign n164 = x102 & ~x128 ;
  assign n165 = x101 & ~x128 ;
  assign n166 = ( x101 & n164 ) | ( x101 & ~n165 ) | ( n164 & ~n165 ) ;
  assign n167 = x129 & ~n166 ;
  assign n168 = x103 & x128 ;
  assign n169 = x104 & ~x128 ;
  assign n170 = ( x129 & ~n168 ) | ( x129 & n169 ) | ( ~n168 & n169 ) ;
  assign n171 = ( ~n167 & n168 ) | ( ~n167 & n170 ) | ( n168 & n170 ) ;
  assign n172 = x131 & ~n171 ;
  assign n173 = x131 & ~n163 ;
  assign n174 = ( n163 & ~n172 ) | ( n163 & n173 ) | ( ~n172 & n173 ) ;
  assign n175 = ~x130 & n174 ;
  assign n176 = ( x130 & ~n155 ) | ( x130 & n175 ) | ( ~n155 & n175 ) ;
  assign n177 = x74 & ~x128 ;
  assign n178 = x73 & ~x128 ;
  assign n179 = ( x73 & n177 ) | ( x73 & ~n178 ) | ( n177 & ~n178 ) ;
  assign n180 = x129 & ~n179 ;
  assign n181 = x75 & x128 ;
  assign n182 = x76 & ~x128 ;
  assign n183 = ( x129 & ~n181 ) | ( x129 & n182 ) | ( ~n181 & n182 ) ;
  assign n184 = ( ~n180 & n181 ) | ( ~n180 & n183 ) | ( n181 & n183 ) ;
  assign n185 = x66 & ~x128 ;
  assign n186 = x65 & ~x128 ;
  assign n187 = ( x65 & n185 ) | ( x65 & ~n186 ) | ( n185 & ~n186 ) ;
  assign n188 = x129 & ~n187 ;
  assign n189 = x67 & x128 ;
  assign n190 = x68 & ~x128 ;
  assign n191 = ( x129 & ~n189 ) | ( x129 & n190 ) | ( ~n189 & n190 ) ;
  assign n192 = ( ~n188 & n189 ) | ( ~n188 & n191 ) | ( n189 & n191 ) ;
  assign n193 = x131 & ~n192 ;
  assign n194 = x131 & ~n184 ;
  assign n195 = ( n184 & ~n193 ) | ( n184 & n194 ) | ( ~n193 & n194 ) ;
  assign n196 = x130 & ~n195 ;
  assign n197 = x78 & ~x128 ;
  assign n198 = x77 & ~x128 ;
  assign n199 = ( x77 & n197 ) | ( x77 & ~n198 ) | ( n197 & ~n198 ) ;
  assign n200 = x129 & ~n199 ;
  assign n201 = x79 & x128 ;
  assign n202 = x80 & ~x128 ;
  assign n203 = ( x129 & ~n201 ) | ( x129 & n202 ) | ( ~n201 & n202 ) ;
  assign n204 = ( ~n200 & n201 ) | ( ~n200 & n203 ) | ( n201 & n203 ) ;
  assign n205 = x70 & ~x128 ;
  assign n206 = x69 & ~x128 ;
  assign n207 = ( x69 & n205 ) | ( x69 & ~n206 ) | ( n205 & ~n206 ) ;
  assign n208 = x129 & ~n207 ;
  assign n209 = x71 & x128 ;
  assign n210 = x72 & ~x128 ;
  assign n211 = ( x129 & ~n209 ) | ( x129 & n210 ) | ( ~n209 & n210 ) ;
  assign n212 = ( ~n208 & n209 ) | ( ~n208 & n211 ) | ( n209 & n211 ) ;
  assign n213 = x131 & ~n212 ;
  assign n214 = x131 & ~n204 ;
  assign n215 = ( n204 & ~n213 ) | ( n204 & n214 ) | ( ~n213 & n214 ) ;
  assign n216 = ~x130 & n215 ;
  assign n217 = ( x130 & ~n196 ) | ( x130 & n216 ) | ( ~n196 & n216 ) ;
  assign n218 = x133 & ~n217 ;
  assign n219 = x133 & ~n176 ;
  assign n220 = ( n176 & ~n218 ) | ( n176 & n219 ) | ( ~n218 & n219 ) ;
  assign n221 = x132 & ~n220 ;
  assign n222 = x122 & ~x128 ;
  assign n223 = x121 & ~x128 ;
  assign n224 = ( x121 & n222 ) | ( x121 & ~n223 ) | ( n222 & ~n223 ) ;
  assign n225 = x129 & ~n224 ;
  assign n226 = x123 & x128 ;
  assign n227 = x124 & ~x128 ;
  assign n228 = ( x129 & ~n226 ) | ( x129 & n227 ) | ( ~n226 & n227 ) ;
  assign n229 = ( ~n225 & n226 ) | ( ~n225 & n228 ) | ( n226 & n228 ) ;
  assign n230 = x114 & ~x128 ;
  assign n231 = x113 & ~x128 ;
  assign n232 = ( x113 & n230 ) | ( x113 & ~n231 ) | ( n230 & ~n231 ) ;
  assign n233 = x129 & ~n232 ;
  assign n234 = x115 & x128 ;
  assign n235 = x116 & ~x128 ;
  assign n236 = ( x129 & ~n234 ) | ( x129 & n235 ) | ( ~n234 & n235 ) ;
  assign n237 = ( ~n233 & n234 ) | ( ~n233 & n236 ) | ( n234 & n236 ) ;
  assign n238 = x131 & ~n237 ;
  assign n239 = x131 & ~n229 ;
  assign n240 = ( n229 & ~n238 ) | ( n229 & n239 ) | ( ~n238 & n239 ) ;
  assign n241 = x130 & ~n240 ;
  assign n242 = x126 & ~x128 ;
  assign n243 = x125 & ~x128 ;
  assign n244 = ( x125 & n242 ) | ( x125 & ~n243 ) | ( n242 & ~n243 ) ;
  assign n245 = x129 & ~n244 ;
  assign n246 = x0 & ~x128 ;
  assign n247 = x127 & x128 ;
  assign n248 = ( x129 & ~n246 ) | ( x129 & n247 ) | ( ~n246 & n247 ) ;
  assign n249 = ( ~n245 & n246 ) | ( ~n245 & n248 ) | ( n246 & n248 ) ;
  assign n250 = x118 & ~x128 ;
  assign n251 = x117 & ~x128 ;
  assign n252 = ( x117 & n250 ) | ( x117 & ~n251 ) | ( n250 & ~n251 ) ;
  assign n253 = x129 & ~n252 ;
  assign n254 = x119 & x128 ;
  assign n255 = x120 & ~x128 ;
  assign n256 = ( x129 & ~n254 ) | ( x129 & n255 ) | ( ~n254 & n255 ) ;
  assign n257 = ( ~n253 & n254 ) | ( ~n253 & n256 ) | ( n254 & n256 ) ;
  assign n258 = x131 & ~n257 ;
  assign n259 = x131 & ~n249 ;
  assign n260 = ( n249 & ~n258 ) | ( n249 & n259 ) | ( ~n258 & n259 ) ;
  assign n261 = ~x130 & n260 ;
  assign n262 = ( x130 & ~n241 ) | ( x130 & n261 ) | ( ~n241 & n261 ) ;
  assign n263 = x90 & ~x128 ;
  assign n264 = x89 & ~x128 ;
  assign n265 = ( x89 & n263 ) | ( x89 & ~n264 ) | ( n263 & ~n264 ) ;
  assign n266 = x129 & ~n265 ;
  assign n267 = x91 & x128 ;
  assign n268 = x92 & ~x128 ;
  assign n269 = ( x129 & ~n267 ) | ( x129 & n268 ) | ( ~n267 & n268 ) ;
  assign n270 = ( ~n266 & n267 ) | ( ~n266 & n269 ) | ( n267 & n269 ) ;
  assign n271 = x82 & ~x128 ;
  assign n272 = x81 & ~x128 ;
  assign n273 = ( x81 & n271 ) | ( x81 & ~n272 ) | ( n271 & ~n272 ) ;
  assign n274 = x129 & ~n273 ;
  assign n275 = x83 & x128 ;
  assign n276 = x84 & ~x128 ;
  assign n277 = ( x129 & ~n275 ) | ( x129 & n276 ) | ( ~n275 & n276 ) ;
  assign n278 = ( ~n274 & n275 ) | ( ~n274 & n277 ) | ( n275 & n277 ) ;
  assign n279 = x131 & ~n278 ;
  assign n280 = x131 & ~n270 ;
  assign n281 = ( n270 & ~n279 ) | ( n270 & n280 ) | ( ~n279 & n280 ) ;
  assign n282 = x130 & ~n281 ;
  assign n283 = x94 & ~x128 ;
  assign n284 = x93 & ~x128 ;
  assign n285 = ( x93 & n283 ) | ( x93 & ~n284 ) | ( n283 & ~n284 ) ;
  assign n286 = x129 & ~n285 ;
  assign n287 = x95 & x128 ;
  assign n288 = x96 & ~x128 ;
  assign n289 = ( x129 & ~n287 ) | ( x129 & n288 ) | ( ~n287 & n288 ) ;
  assign n290 = ( ~n286 & n287 ) | ( ~n286 & n289 ) | ( n287 & n289 ) ;
  assign n291 = x86 & ~x128 ;
  assign n292 = x85 & ~x128 ;
  assign n293 = ( x85 & n291 ) | ( x85 & ~n292 ) | ( n291 & ~n292 ) ;
  assign n294 = x129 & ~n293 ;
  assign n295 = x87 & x128 ;
  assign n296 = x88 & ~x128 ;
  assign n297 = ( x129 & ~n295 ) | ( x129 & n296 ) | ( ~n295 & n296 ) ;
  assign n298 = ( ~n294 & n295 ) | ( ~n294 & n297 ) | ( n295 & n297 ) ;
  assign n299 = x131 & ~n298 ;
  assign n300 = x131 & ~n290 ;
  assign n301 = ( n290 & ~n299 ) | ( n290 & n300 ) | ( ~n299 & n300 ) ;
  assign n302 = ~x130 & n301 ;
  assign n303 = ( x130 & ~n282 ) | ( x130 & n302 ) | ( ~n282 & n302 ) ;
  assign n304 = x133 & ~n303 ;
  assign n305 = x133 & ~n262 ;
  assign n306 = ( n262 & ~n304 ) | ( n262 & n305 ) | ( ~n304 & n305 ) ;
  assign n307 = ~x132 & n306 ;
  assign n308 = ( x132 & ~n221 ) | ( x132 & n307 ) | ( ~n221 & n307 ) ;
  assign n309 = x42 & ~x128 ;
  assign n310 = x41 & ~x128 ;
  assign n311 = ( x41 & n309 ) | ( x41 & ~n310 ) | ( n309 & ~n310 ) ;
  assign n312 = x129 & ~n311 ;
  assign n313 = x43 & x128 ;
  assign n314 = x44 & ~x128 ;
  assign n315 = ( x129 & ~n313 ) | ( x129 & n314 ) | ( ~n313 & n314 ) ;
  assign n316 = ( ~n312 & n313 ) | ( ~n312 & n315 ) | ( n313 & n315 ) ;
  assign n317 = x34 & ~x128 ;
  assign n318 = x33 & ~x128 ;
  assign n319 = ( x33 & n317 ) | ( x33 & ~n318 ) | ( n317 & ~n318 ) ;
  assign n320 = x129 & ~n319 ;
  assign n321 = x35 & x128 ;
  assign n322 = x36 & ~x128 ;
  assign n323 = ( x129 & ~n321 ) | ( x129 & n322 ) | ( ~n321 & n322 ) ;
  assign n324 = ( ~n320 & n321 ) | ( ~n320 & n323 ) | ( n321 & n323 ) ;
  assign n325 = x131 & ~n324 ;
  assign n326 = x131 & ~n316 ;
  assign n327 = ( n316 & ~n325 ) | ( n316 & n326 ) | ( ~n325 & n326 ) ;
  assign n328 = x130 & ~n327 ;
  assign n329 = x46 & ~x128 ;
  assign n330 = x45 & ~x128 ;
  assign n331 = ( x45 & n329 ) | ( x45 & ~n330 ) | ( n329 & ~n330 ) ;
  assign n332 = x129 & ~n331 ;
  assign n333 = x47 & x128 ;
  assign n334 = x48 & ~x128 ;
  assign n335 = ( x129 & ~n333 ) | ( x129 & n334 ) | ( ~n333 & n334 ) ;
  assign n336 = ( ~n332 & n333 ) | ( ~n332 & n335 ) | ( n333 & n335 ) ;
  assign n337 = x38 & ~x128 ;
  assign n338 = x37 & ~x128 ;
  assign n339 = ( x37 & n337 ) | ( x37 & ~n338 ) | ( n337 & ~n338 ) ;
  assign n340 = x129 & ~n339 ;
  assign n341 = x39 & x128 ;
  assign n342 = x40 & ~x128 ;
  assign n343 = ( x129 & ~n341 ) | ( x129 & n342 ) | ( ~n341 & n342 ) ;
  assign n344 = ( ~n340 & n341 ) | ( ~n340 & n343 ) | ( n341 & n343 ) ;
  assign n345 = x131 & ~n344 ;
  assign n346 = x131 & ~n336 ;
  assign n347 = ( n336 & ~n345 ) | ( n336 & n346 ) | ( ~n345 & n346 ) ;
  assign n348 = ~x130 & n347 ;
  assign n349 = ( x130 & ~n328 ) | ( x130 & n348 ) | ( ~n328 & n348 ) ;
  assign n350 = x10 & ~x128 ;
  assign n351 = x9 & ~x128 ;
  assign n352 = ( x9 & n350 ) | ( x9 & ~n351 ) | ( n350 & ~n351 ) ;
  assign n353 = x129 & ~n352 ;
  assign n354 = x11 & x128 ;
  assign n355 = x12 & ~x128 ;
  assign n356 = ( x129 & ~n354 ) | ( x129 & n355 ) | ( ~n354 & n355 ) ;
  assign n357 = ( ~n353 & n354 ) | ( ~n353 & n356 ) | ( n354 & n356 ) ;
  assign n358 = x2 & ~x128 ;
  assign n359 = x1 & ~x128 ;
  assign n360 = ( x1 & n358 ) | ( x1 & ~n359 ) | ( n358 & ~n359 ) ;
  assign n361 = x129 & ~n360 ;
  assign n362 = x3 & x128 ;
  assign n363 = x4 & ~x128 ;
  assign n364 = ( x129 & ~n362 ) | ( x129 & n363 ) | ( ~n362 & n363 ) ;
  assign n365 = ( ~n361 & n362 ) | ( ~n361 & n364 ) | ( n362 & n364 ) ;
  assign n366 = x131 & ~n365 ;
  assign n367 = x131 & ~n357 ;
  assign n368 = ( n357 & ~n366 ) | ( n357 & n367 ) | ( ~n366 & n367 ) ;
  assign n369 = x130 & ~n368 ;
  assign n370 = x14 & ~x128 ;
  assign n371 = x13 & ~x128 ;
  assign n372 = ( x13 & n370 ) | ( x13 & ~n371 ) | ( n370 & ~n371 ) ;
  assign n373 = x129 & ~n372 ;
  assign n374 = x15 & x128 ;
  assign n375 = x16 & ~x128 ;
  assign n376 = ( x129 & ~n374 ) | ( x129 & n375 ) | ( ~n374 & n375 ) ;
  assign n377 = ( ~n373 & n374 ) | ( ~n373 & n376 ) | ( n374 & n376 ) ;
  assign n378 = x6 & ~x128 ;
  assign n379 = x5 & ~x128 ;
  assign n380 = ( x5 & n378 ) | ( x5 & ~n379 ) | ( n378 & ~n379 ) ;
  assign n381 = x129 & ~n380 ;
  assign n382 = x7 & x128 ;
  assign n383 = x8 & ~x128 ;
  assign n384 = ( x129 & ~n382 ) | ( x129 & n383 ) | ( ~n382 & n383 ) ;
  assign n385 = ( ~n381 & n382 ) | ( ~n381 & n384 ) | ( n382 & n384 ) ;
  assign n386 = x131 & ~n385 ;
  assign n387 = x131 & ~n377 ;
  assign n388 = ( n377 & ~n386 ) | ( n377 & n387 ) | ( ~n386 & n387 ) ;
  assign n389 = ~x130 & n388 ;
  assign n390 = ( x130 & ~n369 ) | ( x130 & n389 ) | ( ~n369 & n389 ) ;
  assign n391 = x133 & ~n390 ;
  assign n392 = x133 & ~n349 ;
  assign n393 = ( n349 & ~n391 ) | ( n349 & n392 ) | ( ~n391 & n392 ) ;
  assign n394 = x132 & ~n393 ;
  assign n395 = x58 & ~x128 ;
  assign n396 = x57 & ~x128 ;
  assign n397 = ( x57 & n395 ) | ( x57 & ~n396 ) | ( n395 & ~n396 ) ;
  assign n398 = x129 & ~n397 ;
  assign n399 = x59 & x128 ;
  assign n400 = x60 & ~x128 ;
  assign n401 = ( x129 & ~n399 ) | ( x129 & n400 ) | ( ~n399 & n400 ) ;
  assign n402 = ( ~n398 & n399 ) | ( ~n398 & n401 ) | ( n399 & n401 ) ;
  assign n403 = x50 & ~x128 ;
  assign n404 = x49 & ~x128 ;
  assign n405 = ( x49 & n403 ) | ( x49 & ~n404 ) | ( n403 & ~n404 ) ;
  assign n406 = x129 & ~n405 ;
  assign n407 = x51 & x128 ;
  assign n408 = x52 & ~x128 ;
  assign n409 = ( x129 & ~n407 ) | ( x129 & n408 ) | ( ~n407 & n408 ) ;
  assign n410 = ( ~n406 & n407 ) | ( ~n406 & n409 ) | ( n407 & n409 ) ;
  assign n411 = x131 & ~n410 ;
  assign n412 = x131 & ~n402 ;
  assign n413 = ( n402 & ~n411 ) | ( n402 & n412 ) | ( ~n411 & n412 ) ;
  assign n414 = x130 & ~n413 ;
  assign n415 = x62 & ~x128 ;
  assign n416 = x61 & ~x128 ;
  assign n417 = ( x61 & n415 ) | ( x61 & ~n416 ) | ( n415 & ~n416 ) ;
  assign n418 = x129 & ~n417 ;
  assign n419 = x63 & x128 ;
  assign n420 = x64 & ~x128 ;
  assign n421 = ( x129 & ~n419 ) | ( x129 & n420 ) | ( ~n419 & n420 ) ;
  assign n422 = ( ~n418 & n419 ) | ( ~n418 & n421 ) | ( n419 & n421 ) ;
  assign n423 = x54 & ~x128 ;
  assign n424 = x53 & ~x128 ;
  assign n425 = ( x53 & n423 ) | ( x53 & ~n424 ) | ( n423 & ~n424 ) ;
  assign n426 = x129 & ~n425 ;
  assign n427 = x55 & x128 ;
  assign n428 = x56 & ~x128 ;
  assign n429 = ( x129 & ~n427 ) | ( x129 & n428 ) | ( ~n427 & n428 ) ;
  assign n430 = ( ~n426 & n427 ) | ( ~n426 & n429 ) | ( n427 & n429 ) ;
  assign n431 = x131 & ~n430 ;
  assign n432 = x131 & ~n422 ;
  assign n433 = ( n422 & ~n431 ) | ( n422 & n432 ) | ( ~n431 & n432 ) ;
  assign n434 = ~x130 & n433 ;
  assign n435 = ( x130 & ~n414 ) | ( x130 & n434 ) | ( ~n414 & n434 ) ;
  assign n436 = x26 & ~x128 ;
  assign n437 = x25 & ~x128 ;
  assign n438 = ( x25 & n436 ) | ( x25 & ~n437 ) | ( n436 & ~n437 ) ;
  assign n439 = x129 & ~n438 ;
  assign n440 = x27 & x128 ;
  assign n441 = x28 & ~x128 ;
  assign n442 = ( x129 & ~n440 ) | ( x129 & n441 ) | ( ~n440 & n441 ) ;
  assign n443 = ( ~n439 & n440 ) | ( ~n439 & n442 ) | ( n440 & n442 ) ;
  assign n444 = x18 & ~x128 ;
  assign n445 = x17 & ~x128 ;
  assign n446 = ( x17 & n444 ) | ( x17 & ~n445 ) | ( n444 & ~n445 ) ;
  assign n447 = x129 & ~n446 ;
  assign n448 = x19 & x128 ;
  assign n449 = x20 & ~x128 ;
  assign n450 = ( x129 & ~n448 ) | ( x129 & n449 ) | ( ~n448 & n449 ) ;
  assign n451 = ( ~n447 & n448 ) | ( ~n447 & n450 ) | ( n448 & n450 ) ;
  assign n452 = x131 & ~n451 ;
  assign n453 = x131 & ~n443 ;
  assign n454 = ( n443 & ~n452 ) | ( n443 & n453 ) | ( ~n452 & n453 ) ;
  assign n455 = x130 & ~n454 ;
  assign n456 = x30 & ~x128 ;
  assign n457 = x29 & ~x128 ;
  assign n458 = ( x29 & n456 ) | ( x29 & ~n457 ) | ( n456 & ~n457 ) ;
  assign n459 = x129 & ~n458 ;
  assign n460 = x31 & x128 ;
  assign n461 = x32 & ~x128 ;
  assign n462 = ( x129 & ~n460 ) | ( x129 & n461 ) | ( ~n460 & n461 ) ;
  assign n463 = ( ~n459 & n460 ) | ( ~n459 & n462 ) | ( n460 & n462 ) ;
  assign n464 = x22 & ~x128 ;
  assign n465 = x21 & ~x128 ;
  assign n466 = ( x21 & n464 ) | ( x21 & ~n465 ) | ( n464 & ~n465 ) ;
  assign n467 = x129 & ~n466 ;
  assign n468 = x23 & x128 ;
  assign n469 = x24 & ~x128 ;
  assign n470 = ( x129 & ~n468 ) | ( x129 & n469 ) | ( ~n468 & n469 ) ;
  assign n471 = ( ~n467 & n468 ) | ( ~n467 & n470 ) | ( n468 & n470 ) ;
  assign n472 = x131 & ~n471 ;
  assign n473 = x131 & ~n463 ;
  assign n474 = ( n463 & ~n472 ) | ( n463 & n473 ) | ( ~n472 & n473 ) ;
  assign n475 = ~x130 & n474 ;
  assign n476 = ( x130 & ~n455 ) | ( x130 & n475 ) | ( ~n455 & n475 ) ;
  assign n477 = x133 & ~n476 ;
  assign n478 = x133 & ~n435 ;
  assign n479 = ( n435 & ~n477 ) | ( n435 & n478 ) | ( ~n477 & n478 ) ;
  assign n480 = ~x132 & n479 ;
  assign n481 = ( x132 & ~n394 ) | ( x132 & n480 ) | ( ~n394 & n480 ) ;
  assign n482 = x134 & ~n481 ;
  assign n483 = x134 & ~n308 ;
  assign n484 = ( n308 & ~n482 ) | ( n308 & n483 ) | ( ~n482 & n483 ) ;
  assign n485 = x99 & ~x128 ;
  assign n486 = ( x98 & ~n144 ) | ( x98 & n485 ) | ( ~n144 & n485 ) ;
  assign n487 = x129 & ~n486 ;
  assign n488 = ( x100 & ~n149 ) | ( x100 & n165 ) | ( ~n149 & n165 ) ;
  assign n489 = x129 & ~n488 ;
  assign n490 = ( ~n487 & n488 ) | ( ~n487 & n489 ) | ( n488 & n489 ) ;
  assign n491 = x131 & ~n490 ;
  assign n492 = x107 & ~x128 ;
  assign n493 = ( x106 & ~n136 ) | ( x106 & n492 ) | ( ~n136 & n492 ) ;
  assign n494 = x129 & ~n493 ;
  assign n495 = ( x108 & ~n141 ) | ( x108 & n157 ) | ( ~n141 & n157 ) ;
  assign n496 = x129 & ~n495 ;
  assign n497 = ( ~n494 & n495 ) | ( ~n494 & n496 ) | ( n495 & n496 ) ;
  assign n498 = x131 & ~n497 ;
  assign n499 = ( ~n491 & n497 ) | ( ~n491 & n498 ) | ( n497 & n498 ) ;
  assign n500 = x130 & ~n499 ;
  assign n501 = x103 & ~x128 ;
  assign n502 = ( x102 & ~n164 ) | ( x102 & n501 ) | ( ~n164 & n501 ) ;
  assign n503 = x129 & ~n502 ;
  assign n504 = ( x104 & n137 ) | ( x104 & ~n169 ) | ( n137 & ~n169 ) ;
  assign n505 = x129 & ~n504 ;
  assign n506 = ( ~n503 & n504 ) | ( ~n503 & n505 ) | ( n504 & n505 ) ;
  assign n507 = x131 & ~n506 ;
  assign n508 = x111 & ~x128 ;
  assign n509 = ( x110 & ~n156 ) | ( x110 & n508 ) | ( ~n156 & n508 ) ;
  assign n510 = x129 & ~n509 ;
  assign n511 = ( x112 & ~n161 ) | ( x112 & n231 ) | ( ~n161 & n231 ) ;
  assign n512 = x129 & ~n511 ;
  assign n513 = ( ~n510 & n511 ) | ( ~n510 & n512 ) | ( n511 & n512 ) ;
  assign n514 = x131 & ~n513 ;
  assign n515 = ( ~n507 & n513 ) | ( ~n507 & n514 ) | ( n513 & n514 ) ;
  assign n516 = ~x130 & n515 ;
  assign n517 = ( x130 & ~n500 ) | ( x130 & n516 ) | ( ~n500 & n516 ) ;
  assign n518 = x67 & ~x128 ;
  assign n519 = ( x66 & ~n185 ) | ( x66 & n518 ) | ( ~n185 & n518 ) ;
  assign n520 = x129 & ~n519 ;
  assign n521 = ( x68 & ~n190 ) | ( x68 & n206 ) | ( ~n190 & n206 ) ;
  assign n522 = x129 & ~n521 ;
  assign n523 = ( ~n520 & n521 ) | ( ~n520 & n522 ) | ( n521 & n522 ) ;
  assign n524 = x131 & ~n523 ;
  assign n525 = x75 & ~x128 ;
  assign n526 = ( x74 & ~n177 ) | ( x74 & n525 ) | ( ~n177 & n525 ) ;
  assign n527 = x129 & ~n526 ;
  assign n528 = ( x76 & ~n182 ) | ( x76 & n198 ) | ( ~n182 & n198 ) ;
  assign n529 = x129 & ~n528 ;
  assign n530 = ( ~n527 & n528 ) | ( ~n527 & n529 ) | ( n528 & n529 ) ;
  assign n531 = x131 & ~n530 ;
  assign n532 = ( ~n524 & n530 ) | ( ~n524 & n531 ) | ( n530 & n531 ) ;
  assign n533 = x130 & ~n532 ;
  assign n534 = x71 & ~x128 ;
  assign n535 = ( x70 & ~n205 ) | ( x70 & n534 ) | ( ~n205 & n534 ) ;
  assign n536 = x129 & ~n535 ;
  assign n537 = ( x72 & n178 ) | ( x72 & ~n210 ) | ( n178 & ~n210 ) ;
  assign n538 = x129 & ~n537 ;
  assign n539 = ( ~n536 & n537 ) | ( ~n536 & n538 ) | ( n537 & n538 ) ;
  assign n540 = x131 & ~n539 ;
  assign n541 = x79 & ~x128 ;
  assign n542 = ( x78 & ~n197 ) | ( x78 & n541 ) | ( ~n197 & n541 ) ;
  assign n543 = x129 & ~n542 ;
  assign n544 = ( x80 & ~n202 ) | ( x80 & n272 ) | ( ~n202 & n272 ) ;
  assign n545 = x129 & ~n544 ;
  assign n546 = ( ~n543 & n544 ) | ( ~n543 & n545 ) | ( n544 & n545 ) ;
  assign n547 = x131 & ~n546 ;
  assign n548 = ( ~n540 & n546 ) | ( ~n540 & n547 ) | ( n546 & n547 ) ;
  assign n549 = ~x130 & n548 ;
  assign n550 = ( x130 & ~n533 ) | ( x130 & n549 ) | ( ~n533 & n549 ) ;
  assign n551 = x133 & ~n550 ;
  assign n552 = x133 & ~n517 ;
  assign n553 = ( n517 & ~n551 ) | ( n517 & n552 ) | ( ~n551 & n552 ) ;
  assign n554 = x132 & ~n553 ;
  assign n555 = x115 & ~x128 ;
  assign n556 = ( x114 & ~n230 ) | ( x114 & n555 ) | ( ~n230 & n555 ) ;
  assign n557 = x129 & ~n556 ;
  assign n558 = ( x116 & ~n235 ) | ( x116 & n251 ) | ( ~n235 & n251 ) ;
  assign n559 = x129 & ~n558 ;
  assign n560 = ( ~n557 & n558 ) | ( ~n557 & n559 ) | ( n558 & n559 ) ;
  assign n561 = x131 & ~n560 ;
  assign n562 = x123 & ~x128 ;
  assign n563 = ( x122 & ~n222 ) | ( x122 & n562 ) | ( ~n222 & n562 ) ;
  assign n564 = x129 & ~n563 ;
  assign n565 = ( x124 & ~n227 ) | ( x124 & n243 ) | ( ~n227 & n243 ) ;
  assign n566 = x129 & ~n565 ;
  assign n567 = ( ~n564 & n565 ) | ( ~n564 & n566 ) | ( n565 & n566 ) ;
  assign n568 = x131 & ~n567 ;
  assign n569 = ( ~n561 & n567 ) | ( ~n561 & n568 ) | ( n567 & n568 ) ;
  assign n570 = x130 & ~n569 ;
  assign n571 = x119 & ~x128 ;
  assign n572 = ( x118 & ~n250 ) | ( x118 & n571 ) | ( ~n250 & n571 ) ;
  assign n573 = x129 & ~n572 ;
  assign n574 = ( x120 & n223 ) | ( x120 & ~n255 ) | ( n223 & ~n255 ) ;
  assign n575 = x129 & ~n574 ;
  assign n576 = ( ~n573 & n574 ) | ( ~n573 & n575 ) | ( n574 & n575 ) ;
  assign n577 = x131 & ~n576 ;
  assign n578 = x127 & ~x128 ;
  assign n579 = ( x126 & ~n242 ) | ( x126 & n578 ) | ( ~n242 & n578 ) ;
  assign n580 = x129 & ~n579 ;
  assign n581 = ( x0 & ~n246 ) | ( x0 & n359 ) | ( ~n246 & n359 ) ;
  assign n582 = x129 & ~n581 ;
  assign n583 = ( ~n580 & n581 ) | ( ~n580 & n582 ) | ( n581 & n582 ) ;
  assign n584 = x131 & ~n583 ;
  assign n585 = ( ~n577 & n583 ) | ( ~n577 & n584 ) | ( n583 & n584 ) ;
  assign n586 = ~x130 & n585 ;
  assign n587 = ( x130 & ~n570 ) | ( x130 & n586 ) | ( ~n570 & n586 ) ;
  assign n588 = x83 & ~x128 ;
  assign n589 = ( x82 & ~n271 ) | ( x82 & n588 ) | ( ~n271 & n588 ) ;
  assign n590 = x129 & ~n589 ;
  assign n591 = ( x84 & ~n276 ) | ( x84 & n292 ) | ( ~n276 & n292 ) ;
  assign n592 = x129 & ~n591 ;
  assign n593 = ( ~n590 & n591 ) | ( ~n590 & n592 ) | ( n591 & n592 ) ;
  assign n594 = x131 & ~n593 ;
  assign n595 = x91 & ~x128 ;
  assign n596 = ( x90 & ~n263 ) | ( x90 & n595 ) | ( ~n263 & n595 ) ;
  assign n597 = x129 & ~n596 ;
  assign n598 = ( x92 & ~n268 ) | ( x92 & n284 ) | ( ~n268 & n284 ) ;
  assign n599 = x129 & ~n598 ;
  assign n600 = ( ~n597 & n598 ) | ( ~n597 & n599 ) | ( n598 & n599 ) ;
  assign n601 = x131 & ~n600 ;
  assign n602 = ( ~n594 & n600 ) | ( ~n594 & n601 ) | ( n600 & n601 ) ;
  assign n603 = x130 & ~n602 ;
  assign n604 = x87 & ~x128 ;
  assign n605 = ( x86 & ~n291 ) | ( x86 & n604 ) | ( ~n291 & n604 ) ;
  assign n606 = x129 & ~n605 ;
  assign n607 = ( x88 & n264 ) | ( x88 & ~n296 ) | ( n264 & ~n296 ) ;
  assign n608 = x129 & ~n607 ;
  assign n609 = ( ~n606 & n607 ) | ( ~n606 & n608 ) | ( n607 & n608 ) ;
  assign n610 = x131 & ~n609 ;
  assign n611 = x95 & ~x128 ;
  assign n612 = ( x94 & ~n283 ) | ( x94 & n611 ) | ( ~n283 & n611 ) ;
  assign n613 = x129 & ~n612 ;
  assign n614 = ( x96 & n145 ) | ( x96 & ~n288 ) | ( n145 & ~n288 ) ;
  assign n615 = x129 & ~n614 ;
  assign n616 = ( ~n613 & n614 ) | ( ~n613 & n615 ) | ( n614 & n615 ) ;
  assign n617 = x131 & ~n616 ;
  assign n618 = ( ~n610 & n616 ) | ( ~n610 & n617 ) | ( n616 & n617 ) ;
  assign n619 = ~x130 & n618 ;
  assign n620 = ( x130 & ~n603 ) | ( x130 & n619 ) | ( ~n603 & n619 ) ;
  assign n621 = x133 & ~n620 ;
  assign n622 = x133 & ~n587 ;
  assign n623 = ( n587 & ~n621 ) | ( n587 & n622 ) | ( ~n621 & n622 ) ;
  assign n624 = ~x132 & n623 ;
  assign n625 = ( x132 & ~n554 ) | ( x132 & n624 ) | ( ~n554 & n624 ) ;
  assign n626 = x35 & ~x128 ;
  assign n627 = ( x34 & ~n317 ) | ( x34 & n626 ) | ( ~n317 & n626 ) ;
  assign n628 = x129 & ~n627 ;
  assign n629 = ( x36 & ~n322 ) | ( x36 & n338 ) | ( ~n322 & n338 ) ;
  assign n630 = x129 & ~n629 ;
  assign n631 = ( ~n628 & n629 ) | ( ~n628 & n630 ) | ( n629 & n630 ) ;
  assign n632 = x131 & ~n631 ;
  assign n633 = x43 & ~x128 ;
  assign n634 = ( x42 & ~n309 ) | ( x42 & n633 ) | ( ~n309 & n633 ) ;
  assign n635 = x129 & ~n634 ;
  assign n636 = ( x44 & ~n314 ) | ( x44 & n330 ) | ( ~n314 & n330 ) ;
  assign n637 = x129 & ~n636 ;
  assign n638 = ( ~n635 & n636 ) | ( ~n635 & n637 ) | ( n636 & n637 ) ;
  assign n639 = x131 & ~n638 ;
  assign n640 = ( ~n632 & n638 ) | ( ~n632 & n639 ) | ( n638 & n639 ) ;
  assign n641 = x130 & ~n640 ;
  assign n642 = x39 & ~x128 ;
  assign n643 = ( x38 & ~n337 ) | ( x38 & n642 ) | ( ~n337 & n642 ) ;
  assign n644 = x129 & ~n643 ;
  assign n645 = ( x40 & n310 ) | ( x40 & ~n342 ) | ( n310 & ~n342 ) ;
  assign n646 = x129 & ~n645 ;
  assign n647 = ( ~n644 & n645 ) | ( ~n644 & n646 ) | ( n645 & n646 ) ;
  assign n648 = x131 & ~n647 ;
  assign n649 = x47 & ~x128 ;
  assign n650 = ( x46 & ~n329 ) | ( x46 & n649 ) | ( ~n329 & n649 ) ;
  assign n651 = x129 & ~n650 ;
  assign n652 = ( x48 & ~n334 ) | ( x48 & n404 ) | ( ~n334 & n404 ) ;
  assign n653 = x129 & ~n652 ;
  assign n654 = ( ~n651 & n652 ) | ( ~n651 & n653 ) | ( n652 & n653 ) ;
  assign n655 = x131 & ~n654 ;
  assign n656 = ( ~n648 & n654 ) | ( ~n648 & n655 ) | ( n654 & n655 ) ;
  assign n657 = ~x130 & n656 ;
  assign n658 = ( x130 & ~n641 ) | ( x130 & n657 ) | ( ~n641 & n657 ) ;
  assign n659 = x3 & ~x128 ;
  assign n660 = ( x2 & ~n358 ) | ( x2 & n659 ) | ( ~n358 & n659 ) ;
  assign n661 = x129 & ~n660 ;
  assign n662 = ( x4 & ~n363 ) | ( x4 & n379 ) | ( ~n363 & n379 ) ;
  assign n663 = x129 & ~n662 ;
  assign n664 = ( ~n661 & n662 ) | ( ~n661 & n663 ) | ( n662 & n663 ) ;
  assign n665 = x131 & ~n664 ;
  assign n666 = x11 & ~x128 ;
  assign n667 = ( x10 & ~n350 ) | ( x10 & n666 ) | ( ~n350 & n666 ) ;
  assign n668 = x129 & ~n667 ;
  assign n669 = ( x12 & ~n355 ) | ( x12 & n371 ) | ( ~n355 & n371 ) ;
  assign n670 = x129 & ~n669 ;
  assign n671 = ( ~n668 & n669 ) | ( ~n668 & n670 ) | ( n669 & n670 ) ;
  assign n672 = x131 & ~n671 ;
  assign n673 = ( ~n665 & n671 ) | ( ~n665 & n672 ) | ( n671 & n672 ) ;
  assign n674 = x130 & ~n673 ;
  assign n675 = x7 & ~x128 ;
  assign n676 = ( x6 & ~n378 ) | ( x6 & n675 ) | ( ~n378 & n675 ) ;
  assign n677 = x129 & ~n676 ;
  assign n678 = ( x8 & n351 ) | ( x8 & ~n383 ) | ( n351 & ~n383 ) ;
  assign n679 = x129 & ~n678 ;
  assign n680 = ( ~n677 & n678 ) | ( ~n677 & n679 ) | ( n678 & n679 ) ;
  assign n681 = x131 & ~n680 ;
  assign n682 = x15 & ~x128 ;
  assign n683 = ( x14 & ~n370 ) | ( x14 & n682 ) | ( ~n370 & n682 ) ;
  assign n684 = x129 & ~n683 ;
  assign n685 = ( x16 & ~n375 ) | ( x16 & n445 ) | ( ~n375 & n445 ) ;
  assign n686 = x129 & ~n685 ;
  assign n687 = ( ~n684 & n685 ) | ( ~n684 & n686 ) | ( n685 & n686 ) ;
  assign n688 = x131 & ~n687 ;
  assign n689 = ( ~n681 & n687 ) | ( ~n681 & n688 ) | ( n687 & n688 ) ;
  assign n690 = ~x130 & n689 ;
  assign n691 = ( x130 & ~n674 ) | ( x130 & n690 ) | ( ~n674 & n690 ) ;
  assign n692 = x133 & ~n691 ;
  assign n693 = x133 & ~n658 ;
  assign n694 = ( n658 & ~n692 ) | ( n658 & n693 ) | ( ~n692 & n693 ) ;
  assign n695 = x132 & ~n694 ;
  assign n696 = x51 & ~x128 ;
  assign n697 = ( x50 & ~n403 ) | ( x50 & n696 ) | ( ~n403 & n696 ) ;
  assign n698 = x129 & ~n697 ;
  assign n699 = ( x52 & ~n408 ) | ( x52 & n424 ) | ( ~n408 & n424 ) ;
  assign n700 = x129 & ~n699 ;
  assign n701 = ( ~n698 & n699 ) | ( ~n698 & n700 ) | ( n699 & n700 ) ;
  assign n702 = x131 & ~n701 ;
  assign n703 = x59 & ~x128 ;
  assign n704 = ( x58 & ~n395 ) | ( x58 & n703 ) | ( ~n395 & n703 ) ;
  assign n705 = x129 & ~n704 ;
  assign n706 = ( x60 & ~n400 ) | ( x60 & n416 ) | ( ~n400 & n416 ) ;
  assign n707 = x129 & ~n706 ;
  assign n708 = ( ~n705 & n706 ) | ( ~n705 & n707 ) | ( n706 & n707 ) ;
  assign n709 = x131 & ~n708 ;
  assign n710 = ( ~n702 & n708 ) | ( ~n702 & n709 ) | ( n708 & n709 ) ;
  assign n711 = x130 & ~n710 ;
  assign n712 = x55 & ~x128 ;
  assign n713 = ( x54 & ~n423 ) | ( x54 & n712 ) | ( ~n423 & n712 ) ;
  assign n714 = x129 & ~n713 ;
  assign n715 = ( x56 & n396 ) | ( x56 & ~n428 ) | ( n396 & ~n428 ) ;
  assign n716 = x129 & ~n715 ;
  assign n717 = ( ~n714 & n715 ) | ( ~n714 & n716 ) | ( n715 & n716 ) ;
  assign n718 = x131 & ~n717 ;
  assign n719 = x63 & ~x128 ;
  assign n720 = ( x62 & ~n415 ) | ( x62 & n719 ) | ( ~n415 & n719 ) ;
  assign n721 = x129 & ~n720 ;
  assign n722 = ( x64 & n186 ) | ( x64 & ~n420 ) | ( n186 & ~n420 ) ;
  assign n723 = x129 & ~n722 ;
  assign n724 = ( ~n721 & n722 ) | ( ~n721 & n723 ) | ( n722 & n723 ) ;
  assign n725 = x131 & ~n724 ;
  assign n726 = ( ~n718 & n724 ) | ( ~n718 & n725 ) | ( n724 & n725 ) ;
  assign n727 = ~x130 & n726 ;
  assign n728 = ( x130 & ~n711 ) | ( x130 & n727 ) | ( ~n711 & n727 ) ;
  assign n729 = x19 & ~x128 ;
  assign n730 = ( x18 & ~n444 ) | ( x18 & n729 ) | ( ~n444 & n729 ) ;
  assign n731 = x129 & ~n730 ;
  assign n732 = ( x20 & ~n449 ) | ( x20 & n465 ) | ( ~n449 & n465 ) ;
  assign n733 = x129 & ~n732 ;
  assign n734 = ( ~n731 & n732 ) | ( ~n731 & n733 ) | ( n732 & n733 ) ;
  assign n735 = x131 & ~n734 ;
  assign n736 = x27 & ~x128 ;
  assign n737 = ( x26 & ~n436 ) | ( x26 & n736 ) | ( ~n436 & n736 ) ;
  assign n738 = x129 & ~n737 ;
  assign n739 = ( x28 & ~n441 ) | ( x28 & n457 ) | ( ~n441 & n457 ) ;
  assign n740 = x129 & ~n739 ;
  assign n741 = ( ~n738 & n739 ) | ( ~n738 & n740 ) | ( n739 & n740 ) ;
  assign n742 = x131 & ~n741 ;
  assign n743 = ( ~n735 & n741 ) | ( ~n735 & n742 ) | ( n741 & n742 ) ;
  assign n744 = x130 & ~n743 ;
  assign n745 = x23 & ~x128 ;
  assign n746 = ( x22 & ~n464 ) | ( x22 & n745 ) | ( ~n464 & n745 ) ;
  assign n747 = x129 & ~n746 ;
  assign n748 = ( x24 & n437 ) | ( x24 & ~n469 ) | ( n437 & ~n469 ) ;
  assign n749 = x129 & ~n748 ;
  assign n750 = ( ~n747 & n748 ) | ( ~n747 & n749 ) | ( n748 & n749 ) ;
  assign n751 = x131 & ~n750 ;
  assign n752 = x31 & ~x128 ;
  assign n753 = ( x30 & ~n456 ) | ( x30 & n752 ) | ( ~n456 & n752 ) ;
  assign n754 = x129 & ~n753 ;
  assign n755 = ( x32 & n318 ) | ( x32 & ~n461 ) | ( n318 & ~n461 ) ;
  assign n756 = x129 & ~n755 ;
  assign n757 = ( ~n754 & n755 ) | ( ~n754 & n756 ) | ( n755 & n756 ) ;
  assign n758 = x131 & ~n757 ;
  assign n759 = ( ~n751 & n757 ) | ( ~n751 & n758 ) | ( n757 & n758 ) ;
  assign n760 = ~x130 & n759 ;
  assign n761 = ( x130 & ~n744 ) | ( x130 & n760 ) | ( ~n744 & n760 ) ;
  assign n762 = x133 & ~n761 ;
  assign n763 = x133 & ~n728 ;
  assign n764 = ( n728 & ~n762 ) | ( n728 & n763 ) | ( ~n762 & n763 ) ;
  assign n765 = ~x132 & n764 ;
  assign n766 = ( x132 & ~n695 ) | ( x132 & n765 ) | ( ~n695 & n765 ) ;
  assign n767 = x134 & ~n766 ;
  assign n768 = x134 & ~n625 ;
  assign n769 = ( n625 & ~n767 ) | ( n625 & n768 ) | ( ~n767 & n768 ) ;
  assign n770 = x129 | n158 ;
  assign n771 = ( n141 & ~n142 ) | ( n141 & n770 ) | ( ~n142 & n770 ) ;
  assign n772 = x129 | n166 ;
  assign n773 = ( n149 & ~n150 ) | ( n149 & n772 ) | ( ~n150 & n772 ) ;
  assign n774 = x131 & ~n773 ;
  assign n775 = x131 & ~n771 ;
  assign n776 = ( n771 & ~n774 ) | ( n771 & n775 ) | ( ~n774 & n775 ) ;
  assign n777 = x130 & ~n776 ;
  assign n778 = x129 | n232 ;
  assign n779 = ( n161 & ~n162 ) | ( n161 & n778 ) | ( ~n162 & n778 ) ;
  assign n780 = x129 | n138 ;
  assign n781 = ( n169 & ~n170 ) | ( n169 & n780 ) | ( ~n170 & n780 ) ;
  assign n782 = x131 & ~n781 ;
  assign n783 = x131 & ~n779 ;
  assign n784 = ( n779 & ~n782 ) | ( n779 & n783 ) | ( ~n782 & n783 ) ;
  assign n785 = ~x130 & n784 ;
  assign n786 = ( x130 & ~n777 ) | ( x130 & n785 ) | ( ~n777 & n785 ) ;
  assign n787 = ~x133 & n786 ;
  assign n788 = x129 | n199 ;
  assign n789 = ( n182 & ~n183 ) | ( n182 & n788 ) | ( ~n183 & n788 ) ;
  assign n790 = x129 | n207 ;
  assign n791 = ( n190 & ~n191 ) | ( n190 & n790 ) | ( ~n191 & n790 ) ;
  assign n792 = x131 & ~n791 ;
  assign n793 = x131 & ~n789 ;
  assign n794 = ( n789 & ~n792 ) | ( n789 & n793 ) | ( ~n792 & n793 ) ;
  assign n795 = x130 & ~n794 ;
  assign n796 = x129 | n273 ;
  assign n797 = ( n202 & ~n203 ) | ( n202 & n796 ) | ( ~n203 & n796 ) ;
  assign n798 = x129 | n179 ;
  assign n799 = ( n210 & ~n211 ) | ( n210 & n798 ) | ( ~n211 & n798 ) ;
  assign n800 = x131 & ~n799 ;
  assign n801 = x131 & ~n797 ;
  assign n802 = ( n797 & ~n800 ) | ( n797 & n801 ) | ( ~n800 & n801 ) ;
  assign n803 = ~x130 & n802 ;
  assign n804 = ( x130 & ~n795 ) | ( x130 & n803 ) | ( ~n795 & n803 ) ;
  assign n805 = x133 & n804 ;
  assign n806 = ( x132 & n787 ) | ( x132 & n805 ) | ( n787 & n805 ) ;
  assign n807 = x129 | n244 ;
  assign n808 = ( n227 & ~n228 ) | ( n227 & n807 ) | ( ~n228 & n807 ) ;
  assign n809 = x129 | n252 ;
  assign n810 = ( n235 & ~n236 ) | ( n235 & n809 ) | ( ~n236 & n809 ) ;
  assign n811 = x131 & ~n810 ;
  assign n812 = x131 & ~n808 ;
  assign n813 = ( n808 & ~n811 ) | ( n808 & n812 ) | ( ~n811 & n812 ) ;
  assign n814 = x130 & ~n813 ;
  assign n815 = x129 | n360 ;
  assign n816 = ( n247 & ~n248 ) | ( n247 & n815 ) | ( ~n248 & n815 ) ;
  assign n817 = x129 | n224 ;
  assign n818 = ( n255 & ~n256 ) | ( n255 & n817 ) | ( ~n256 & n817 ) ;
  assign n819 = x131 & ~n818 ;
  assign n820 = x131 & ~n816 ;
  assign n821 = ( n816 & ~n819 ) | ( n816 & n820 ) | ( ~n819 & n820 ) ;
  assign n822 = ~x130 & n821 ;
  assign n823 = ( x130 & ~n814 ) | ( x130 & n822 ) | ( ~n814 & n822 ) ;
  assign n824 = ~x133 & n823 ;
  assign n825 = x129 | n285 ;
  assign n826 = ( n268 & ~n269 ) | ( n268 & n825 ) | ( ~n269 & n825 ) ;
  assign n827 = x129 | n293 ;
  assign n828 = ( n276 & ~n277 ) | ( n276 & n827 ) | ( ~n277 & n827 ) ;
  assign n829 = x131 & ~n828 ;
  assign n830 = x131 & ~n826 ;
  assign n831 = ( n826 & ~n829 ) | ( n826 & n830 ) | ( ~n829 & n830 ) ;
  assign n832 = x130 & ~n831 ;
  assign n833 = x129 | n146 ;
  assign n834 = ( n288 & ~n289 ) | ( n288 & n833 ) | ( ~n289 & n833 ) ;
  assign n835 = x129 | n265 ;
  assign n836 = ( n296 & ~n297 ) | ( n296 & n835 ) | ( ~n297 & n835 ) ;
  assign n837 = x131 & ~n836 ;
  assign n838 = x131 & ~n834 ;
  assign n839 = ( n834 & ~n837 ) | ( n834 & n838 ) | ( ~n837 & n838 ) ;
  assign n840 = ~x130 & n839 ;
  assign n841 = ( x130 & ~n832 ) | ( x130 & n840 ) | ( ~n832 & n840 ) ;
  assign n842 = x133 & n841 ;
  assign n843 = ( ~x132 & n824 ) | ( ~x132 & n842 ) | ( n824 & n842 ) ;
  assign n844 = n806 | n843 ;
  assign n845 = x129 | n331 ;
  assign n846 = ( n314 & ~n315 ) | ( n314 & n845 ) | ( ~n315 & n845 ) ;
  assign n847 = x129 | n339 ;
  assign n848 = ( n322 & ~n323 ) | ( n322 & n847 ) | ( ~n323 & n847 ) ;
  assign n849 = x131 & ~n848 ;
  assign n850 = x131 & ~n846 ;
  assign n851 = ( n846 & ~n849 ) | ( n846 & n850 ) | ( ~n849 & n850 ) ;
  assign n852 = x130 & ~n851 ;
  assign n853 = x129 | n405 ;
  assign n854 = ( n334 & ~n335 ) | ( n334 & n853 ) | ( ~n335 & n853 ) ;
  assign n855 = x129 | n311 ;
  assign n856 = ( n342 & ~n343 ) | ( n342 & n855 ) | ( ~n343 & n855 ) ;
  assign n857 = x131 & ~n856 ;
  assign n858 = x131 & ~n854 ;
  assign n859 = ( n854 & ~n857 ) | ( n854 & n858 ) | ( ~n857 & n858 ) ;
  assign n860 = ~x130 & n859 ;
  assign n861 = ( x130 & ~n852 ) | ( x130 & n860 ) | ( ~n852 & n860 ) ;
  assign n862 = x132 & ~n861 ;
  assign n863 = x129 | n417 ;
  assign n864 = ( n400 & ~n401 ) | ( n400 & n863 ) | ( ~n401 & n863 ) ;
  assign n865 = x129 | n425 ;
  assign n866 = ( n408 & ~n409 ) | ( n408 & n865 ) | ( ~n409 & n865 ) ;
  assign n867 = x131 & ~n866 ;
  assign n868 = x131 & ~n864 ;
  assign n869 = ( n864 & ~n867 ) | ( n864 & n868 ) | ( ~n867 & n868 ) ;
  assign n870 = x130 & ~n869 ;
  assign n871 = x129 | n187 ;
  assign n872 = ( n420 & ~n421 ) | ( n420 & n871 ) | ( ~n421 & n871 ) ;
  assign n873 = x129 | n397 ;
  assign n874 = ( n428 & ~n429 ) | ( n428 & n873 ) | ( ~n429 & n873 ) ;
  assign n875 = x131 & ~n874 ;
  assign n876 = x131 & ~n872 ;
  assign n877 = ( n872 & ~n875 ) | ( n872 & n876 ) | ( ~n875 & n876 ) ;
  assign n878 = ~x130 & n877 ;
  assign n879 = ( x130 & ~n870 ) | ( x130 & n878 ) | ( ~n870 & n878 ) ;
  assign n880 = x132 | n879 ;
  assign n881 = ( x133 & ~n862 ) | ( x133 & n880 ) | ( ~n862 & n880 ) ;
  assign n882 = x129 | n372 ;
  assign n883 = ( n355 & ~n356 ) | ( n355 & n882 ) | ( ~n356 & n882 ) ;
  assign n884 = x129 | n380 ;
  assign n885 = ( n363 & ~n364 ) | ( n363 & n884 ) | ( ~n364 & n884 ) ;
  assign n886 = x131 & ~n885 ;
  assign n887 = x131 & ~n883 ;
  assign n888 = ( n883 & ~n886 ) | ( n883 & n887 ) | ( ~n886 & n887 ) ;
  assign n889 = x130 & ~n888 ;
  assign n890 = x129 | n446 ;
  assign n891 = ( n375 & ~n376 ) | ( n375 & n890 ) | ( ~n376 & n890 ) ;
  assign n892 = x129 | n352 ;
  assign n893 = ( n383 & ~n384 ) | ( n383 & n892 ) | ( ~n384 & n892 ) ;
  assign n894 = x131 & ~n893 ;
  assign n895 = x131 & ~n891 ;
  assign n896 = ( n891 & ~n894 ) | ( n891 & n895 ) | ( ~n894 & n895 ) ;
  assign n897 = ~x130 & n896 ;
  assign n898 = ( x130 & ~n889 ) | ( x130 & n897 ) | ( ~n889 & n897 ) ;
  assign n899 = x132 & ~n898 ;
  assign n900 = x129 | n458 ;
  assign n901 = ( n441 & ~n442 ) | ( n441 & n900 ) | ( ~n442 & n900 ) ;
  assign n902 = x129 | n466 ;
  assign n903 = ( n449 & ~n450 ) | ( n449 & n902 ) | ( ~n450 & n902 ) ;
  assign n904 = x131 & ~n903 ;
  assign n905 = x131 & ~n901 ;
  assign n906 = ( n901 & ~n904 ) | ( n901 & n905 ) | ( ~n904 & n905 ) ;
  assign n907 = x130 & ~n906 ;
  assign n908 = x129 | n319 ;
  assign n909 = ( n461 & ~n462 ) | ( n461 & n908 ) | ( ~n462 & n908 ) ;
  assign n910 = x129 | n438 ;
  assign n911 = ( n469 & ~n470 ) | ( n469 & n910 ) | ( ~n470 & n910 ) ;
  assign n912 = x131 & ~n911 ;
  assign n913 = x131 & ~n909 ;
  assign n914 = ( n909 & ~n912 ) | ( n909 & n913 ) | ( ~n912 & n913 ) ;
  assign n915 = ~x130 & n914 ;
  assign n916 = ( x130 & ~n907 ) | ( x130 & n915 ) | ( ~n907 & n915 ) ;
  assign n917 = x132 | n916 ;
  assign n918 = ( x133 & n899 ) | ( x133 & ~n917 ) | ( n899 & ~n917 ) ;
  assign n919 = n881 & ~n918 ;
  assign n920 = x134 & ~n919 ;
  assign n921 = x134 & ~n844 ;
  assign n922 = ( n844 & ~n920 ) | ( n844 & n921 ) | ( ~n920 & n921 ) ;
  assign n923 = ( ~n496 & n509 ) | ( ~n496 & n510 ) | ( n509 & n510 ) ;
  assign n924 = ( ~n489 & n502 ) | ( ~n489 & n503 ) | ( n502 & n503 ) ;
  assign n925 = x131 & ~n924 ;
  assign n926 = x131 & ~n923 ;
  assign n927 = ( n923 & ~n925 ) | ( n923 & n926 ) | ( ~n925 & n926 ) ;
  assign n928 = x130 & ~n927 ;
  assign n929 = ( ~n512 & n556 ) | ( ~n512 & n557 ) | ( n556 & n557 ) ;
  assign n930 = ( n493 & n494 ) | ( n493 & ~n505 ) | ( n494 & ~n505 ) ;
  assign n931 = x131 & ~n930 ;
  assign n932 = x131 & ~n929 ;
  assign n933 = ( n929 & ~n931 ) | ( n929 & n932 ) | ( ~n931 & n932 ) ;
  assign n934 = ~x130 & n933 ;
  assign n935 = ( x130 & ~n928 ) | ( x130 & n934 ) | ( ~n928 & n934 ) ;
  assign n936 = ( ~n529 & n542 ) | ( ~n529 & n543 ) | ( n542 & n543 ) ;
  assign n937 = ( ~n522 & n535 ) | ( ~n522 & n536 ) | ( n535 & n536 ) ;
  assign n938 = x131 & ~n937 ;
  assign n939 = x131 & ~n936 ;
  assign n940 = ( n936 & ~n938 ) | ( n936 & n939 ) | ( ~n938 & n939 ) ;
  assign n941 = x130 & ~n940 ;
  assign n942 = ( ~n545 & n589 ) | ( ~n545 & n590 ) | ( n589 & n590 ) ;
  assign n943 = ( n526 & n527 ) | ( n526 & ~n538 ) | ( n527 & ~n538 ) ;
  assign n944 = x131 & ~n943 ;
  assign n945 = x131 & ~n942 ;
  assign n946 = ( n942 & ~n944 ) | ( n942 & n945 ) | ( ~n944 & n945 ) ;
  assign n947 = ~x130 & n946 ;
  assign n948 = ( x130 & ~n941 ) | ( x130 & n947 ) | ( ~n941 & n947 ) ;
  assign n949 = x133 & ~n948 ;
  assign n950 = x133 & ~n935 ;
  assign n951 = ( n935 & ~n949 ) | ( n935 & n950 ) | ( ~n949 & n950 ) ;
  assign n952 = x132 & ~n951 ;
  assign n953 = ( ~n566 & n579 ) | ( ~n566 & n580 ) | ( n579 & n580 ) ;
  assign n954 = ( ~n559 & n572 ) | ( ~n559 & n573 ) | ( n572 & n573 ) ;
  assign n955 = x131 & ~n954 ;
  assign n956 = x131 & ~n953 ;
  assign n957 = ( n953 & ~n955 ) | ( n953 & n956 ) | ( ~n955 & n956 ) ;
  assign n958 = x130 & ~n957 ;
  assign n959 = ( ~n582 & n660 ) | ( ~n582 & n661 ) | ( n660 & n661 ) ;
  assign n960 = ( n563 & n564 ) | ( n563 & ~n575 ) | ( n564 & ~n575 ) ;
  assign n961 = x131 & ~n960 ;
  assign n962 = x131 & ~n959 ;
  assign n963 = ( n959 & ~n961 ) | ( n959 & n962 ) | ( ~n961 & n962 ) ;
  assign n964 = ~x130 & n963 ;
  assign n965 = ( x130 & ~n958 ) | ( x130 & n964 ) | ( ~n958 & n964 ) ;
  assign n966 = ( ~n599 & n612 ) | ( ~n599 & n613 ) | ( n612 & n613 ) ;
  assign n967 = ( ~n592 & n605 ) | ( ~n592 & n606 ) | ( n605 & n606 ) ;
  assign n968 = x131 & ~n967 ;
  assign n969 = x131 & ~n966 ;
  assign n970 = ( n966 & ~n968 ) | ( n966 & n969 ) | ( ~n968 & n969 ) ;
  assign n971 = x130 & ~n970 ;
  assign n972 = ( n486 & n487 ) | ( n486 & ~n615 ) | ( n487 & ~n615 ) ;
  assign n973 = ( n596 & n597 ) | ( n596 & ~n608 ) | ( n597 & ~n608 ) ;
  assign n974 = x131 & ~n973 ;
  assign n975 = x131 & ~n972 ;
  assign n976 = ( n972 & ~n974 ) | ( n972 & n975 ) | ( ~n974 & n975 ) ;
  assign n977 = ~x130 & n976 ;
  assign n978 = ( x130 & ~n971 ) | ( x130 & n977 ) | ( ~n971 & n977 ) ;
  assign n979 = x133 & ~n978 ;
  assign n980 = x133 & ~n965 ;
  assign n981 = ( n965 & ~n979 ) | ( n965 & n980 ) | ( ~n979 & n980 ) ;
  assign n982 = ~x132 & n981 ;
  assign n983 = ( x132 & ~n952 ) | ( x132 & n982 ) | ( ~n952 & n982 ) ;
  assign n984 = ( ~n637 & n650 ) | ( ~n637 & n651 ) | ( n650 & n651 ) ;
  assign n985 = ( ~n630 & n643 ) | ( ~n630 & n644 ) | ( n643 & n644 ) ;
  assign n986 = x131 & ~n985 ;
  assign n987 = x131 & ~n984 ;
  assign n988 = ( n984 & ~n986 ) | ( n984 & n987 ) | ( ~n986 & n987 ) ;
  assign n989 = x130 & ~n988 ;
  assign n990 = ( ~n653 & n697 ) | ( ~n653 & n698 ) | ( n697 & n698 ) ;
  assign n991 = ( n634 & n635 ) | ( n634 & ~n646 ) | ( n635 & ~n646 ) ;
  assign n992 = x131 & ~n991 ;
  assign n993 = x131 & ~n990 ;
  assign n994 = ( n990 & ~n992 ) | ( n990 & n993 ) | ( ~n992 & n993 ) ;
  assign n995 = ~x130 & n994 ;
  assign n996 = ( x130 & ~n989 ) | ( x130 & n995 ) | ( ~n989 & n995 ) ;
  assign n997 = ( ~n670 & n683 ) | ( ~n670 & n684 ) | ( n683 & n684 ) ;
  assign n998 = ( ~n663 & n676 ) | ( ~n663 & n677 ) | ( n676 & n677 ) ;
  assign n999 = x131 & ~n998 ;
  assign n1000 = x131 & ~n997 ;
  assign n1001 = ( n997 & ~n999 ) | ( n997 & n1000 ) | ( ~n999 & n1000 ) ;
  assign n1002 = x130 & ~n1001 ;
  assign n1003 = ( ~n686 & n730 ) | ( ~n686 & n731 ) | ( n730 & n731 ) ;
  assign n1004 = ( n667 & n668 ) | ( n667 & ~n679 ) | ( n668 & ~n679 ) ;
  assign n1005 = x131 & ~n1004 ;
  assign n1006 = x131 & ~n1003 ;
  assign n1007 = ( n1003 & ~n1005 ) | ( n1003 & n1006 ) | ( ~n1005 & n1006 ) ;
  assign n1008 = ~x130 & n1007 ;
  assign n1009 = ( x130 & ~n1002 ) | ( x130 & n1008 ) | ( ~n1002 & n1008 ) ;
  assign n1010 = x133 & ~n1009 ;
  assign n1011 = x133 & ~n996 ;
  assign n1012 = ( n996 & ~n1010 ) | ( n996 & n1011 ) | ( ~n1010 & n1011 ) ;
  assign n1013 = x132 & ~n1012 ;
  assign n1014 = ( ~n707 & n720 ) | ( ~n707 & n721 ) | ( n720 & n721 ) ;
  assign n1015 = ( ~n700 & n713 ) | ( ~n700 & n714 ) | ( n713 & n714 ) ;
  assign n1016 = x131 & ~n1015 ;
  assign n1017 = x131 & ~n1014 ;
  assign n1018 = ( n1014 & ~n1016 ) | ( n1014 & n1017 ) | ( ~n1016 & n1017 ) ;
  assign n1019 = x130 & ~n1018 ;
  assign n1020 = ( n519 & n520 ) | ( n519 & ~n723 ) | ( n520 & ~n723 ) ;
  assign n1021 = ( n704 & n705 ) | ( n704 & ~n716 ) | ( n705 & ~n716 ) ;
  assign n1022 = x131 & ~n1021 ;
  assign n1023 = x131 & ~n1020 ;
  assign n1024 = ( n1020 & ~n1022 ) | ( n1020 & n1023 ) | ( ~n1022 & n1023 ) ;
  assign n1025 = ~x130 & n1024 ;
  assign n1026 = ( x130 & ~n1019 ) | ( x130 & n1025 ) | ( ~n1019 & n1025 ) ;
  assign n1027 = ( ~n740 & n753 ) | ( ~n740 & n754 ) | ( n753 & n754 ) ;
  assign n1028 = ( ~n733 & n746 ) | ( ~n733 & n747 ) | ( n746 & n747 ) ;
  assign n1029 = x131 & ~n1028 ;
  assign n1030 = x131 & ~n1027 ;
  assign n1031 = ( n1027 & ~n1029 ) | ( n1027 & n1030 ) | ( ~n1029 & n1030 ) ;
  assign n1032 = x130 & ~n1031 ;
  assign n1033 = ( n627 & n628 ) | ( n627 & ~n756 ) | ( n628 & ~n756 ) ;
  assign n1034 = ( n737 & n738 ) | ( n737 & ~n749 ) | ( n738 & ~n749 ) ;
  assign n1035 = x131 & ~n1034 ;
  assign n1036 = x131 & ~n1033 ;
  assign n1037 = ( n1033 & ~n1035 ) | ( n1033 & n1036 ) | ( ~n1035 & n1036 ) ;
  assign n1038 = ~x130 & n1037 ;
  assign n1039 = ( x130 & ~n1032 ) | ( x130 & n1038 ) | ( ~n1032 & n1038 ) ;
  assign n1040 = x133 & ~n1039 ;
  assign n1041 = x133 & ~n1026 ;
  assign n1042 = ( n1026 & ~n1040 ) | ( n1026 & n1041 ) | ( ~n1040 & n1041 ) ;
  assign n1043 = ~x132 & n1042 ;
  assign n1044 = ( x132 & ~n1013 ) | ( x132 & n1043 ) | ( ~n1013 & n1043 ) ;
  assign n1045 = x134 & ~n1044 ;
  assign n1046 = x134 & ~n983 ;
  assign n1047 = ( n983 & ~n1045 ) | ( n983 & n1046 ) | ( ~n1045 & n1046 ) ;
  assign n1048 = ( ~n153 & n237 ) | ( ~n153 & n238 ) | ( n237 & n238 ) ;
  assign n1049 = ~x130 & n1048 ;
  assign n1050 = ( n174 & ~n175 ) | ( n174 & n1049 ) | ( ~n175 & n1049 ) ;
  assign n1051 = ( ~n194 & n278 ) | ( ~n194 & n279 ) | ( n278 & n279 ) ;
  assign n1052 = ~x130 & n1051 ;
  assign n1053 = ( n215 & ~n216 ) | ( n215 & n1052 ) | ( ~n216 & n1052 ) ;
  assign n1054 = x133 & ~n1053 ;
  assign n1055 = x133 & ~n1050 ;
  assign n1056 = ( n1050 & ~n1054 ) | ( n1050 & n1055 ) | ( ~n1054 & n1055 ) ;
  assign n1057 = x132 & ~n1056 ;
  assign n1058 = ( ~n239 & n365 ) | ( ~n239 & n366 ) | ( n365 & n366 ) ;
  assign n1059 = ~x130 & n1058 ;
  assign n1060 = ( n260 & ~n261 ) | ( n260 & n1059 ) | ( ~n261 & n1059 ) ;
  assign n1061 = ( n151 & n152 ) | ( n151 & ~n280 ) | ( n152 & ~n280 ) ;
  assign n1062 = ~x130 & n1061 ;
  assign n1063 = ( n301 & ~n302 ) | ( n301 & n1062 ) | ( ~n302 & n1062 ) ;
  assign n1064 = x133 & ~n1063 ;
  assign n1065 = x133 & ~n1060 ;
  assign n1066 = ( n1060 & ~n1064 ) | ( n1060 & n1065 ) | ( ~n1064 & n1065 ) ;
  assign n1067 = ~x132 & n1066 ;
  assign n1068 = ( x132 & ~n1057 ) | ( x132 & n1067 ) | ( ~n1057 & n1067 ) ;
  assign n1069 = ( ~n326 & n410 ) | ( ~n326 & n411 ) | ( n410 & n411 ) ;
  assign n1070 = ~x130 & n1069 ;
  assign n1071 = ( n347 & ~n348 ) | ( n347 & n1070 ) | ( ~n348 & n1070 ) ;
  assign n1072 = ( ~n367 & n451 ) | ( ~n367 & n452 ) | ( n451 & n452 ) ;
  assign n1073 = ~x130 & n1072 ;
  assign n1074 = ( n388 & ~n389 ) | ( n388 & n1073 ) | ( ~n389 & n1073 ) ;
  assign n1075 = x133 & ~n1074 ;
  assign n1076 = x133 & ~n1071 ;
  assign n1077 = ( n1071 & ~n1075 ) | ( n1071 & n1076 ) | ( ~n1075 & n1076 ) ;
  assign n1078 = x132 & ~n1077 ;
  assign n1079 = ( n192 & n193 ) | ( n192 & ~n412 ) | ( n193 & ~n412 ) ;
  assign n1080 = ~x130 & n1079 ;
  assign n1081 = ( n433 & ~n434 ) | ( n433 & n1080 ) | ( ~n434 & n1080 ) ;
  assign n1082 = ( n324 & n325 ) | ( n324 & ~n453 ) | ( n325 & ~n453 ) ;
  assign n1083 = ~x130 & n1082 ;
  assign n1084 = ( n474 & ~n475 ) | ( n474 & n1083 ) | ( ~n475 & n1083 ) ;
  assign n1085 = x133 & ~n1084 ;
  assign n1086 = x133 & ~n1081 ;
  assign n1087 = ( n1081 & ~n1085 ) | ( n1081 & n1086 ) | ( ~n1085 & n1086 ) ;
  assign n1088 = ~x132 & n1087 ;
  assign n1089 = ( x132 & ~n1078 ) | ( x132 & n1088 ) | ( ~n1078 & n1088 ) ;
  assign n1090 = x134 & ~n1089 ;
  assign n1091 = x134 & ~n1068 ;
  assign n1092 = ( n1068 & ~n1090 ) | ( n1068 & n1091 ) | ( ~n1090 & n1091 ) ;
  assign n1093 = ( ~n498 & n560 ) | ( ~n498 & n561 ) | ( n560 & n561 ) ;
  assign n1094 = ~x130 & n1093 ;
  assign n1095 = ( n515 & ~n516 ) | ( n515 & n1094 ) | ( ~n516 & n1094 ) ;
  assign n1096 = ( ~n531 & n593 ) | ( ~n531 & n594 ) | ( n593 & n594 ) ;
  assign n1097 = ~x130 & n1096 ;
  assign n1098 = ( n548 & ~n549 ) | ( n548 & n1097 ) | ( ~n549 & n1097 ) ;
  assign n1099 = x133 & ~n1098 ;
  assign n1100 = x133 & ~n1095 ;
  assign n1101 = ( n1095 & ~n1099 ) | ( n1095 & n1100 ) | ( ~n1099 & n1100 ) ;
  assign n1102 = x132 & ~n1101 ;
  assign n1103 = ( ~n568 & n664 ) | ( ~n568 & n665 ) | ( n664 & n665 ) ;
  assign n1104 = ~x130 & n1103 ;
  assign n1105 = ( n585 & ~n586 ) | ( n585 & n1104 ) | ( ~n586 & n1104 ) ;
  assign n1106 = ( n490 & n491 ) | ( n490 & ~n601 ) | ( n491 & ~n601 ) ;
  assign n1107 = ~x130 & n1106 ;
  assign n1108 = ( n618 & ~n619 ) | ( n618 & n1107 ) | ( ~n619 & n1107 ) ;
  assign n1109 = x133 & ~n1108 ;
  assign n1110 = x133 & ~n1105 ;
  assign n1111 = ( n1105 & ~n1109 ) | ( n1105 & n1110 ) | ( ~n1109 & n1110 ) ;
  assign n1112 = ~x132 & n1111 ;
  assign n1113 = ( x132 & ~n1102 ) | ( x132 & n1112 ) | ( ~n1102 & n1112 ) ;
  assign n1114 = ( ~n639 & n701 ) | ( ~n639 & n702 ) | ( n701 & n702 ) ;
  assign n1115 = ~x130 & n1114 ;
  assign n1116 = ( n656 & ~n657 ) | ( n656 & n1115 ) | ( ~n657 & n1115 ) ;
  assign n1117 = ( ~n672 & n734 ) | ( ~n672 & n735 ) | ( n734 & n735 ) ;
  assign n1118 = ~x130 & n1117 ;
  assign n1119 = ( n689 & ~n690 ) | ( n689 & n1118 ) | ( ~n690 & n1118 ) ;
  assign n1120 = x133 & ~n1119 ;
  assign n1121 = x133 & ~n1116 ;
  assign n1122 = ( n1116 & ~n1120 ) | ( n1116 & n1121 ) | ( ~n1120 & n1121 ) ;
  assign n1123 = x132 & ~n1122 ;
  assign n1124 = ( n523 & n524 ) | ( n523 & ~n709 ) | ( n524 & ~n709 ) ;
  assign n1125 = ~x130 & n1124 ;
  assign n1126 = ( n726 & ~n727 ) | ( n726 & n1125 ) | ( ~n727 & n1125 ) ;
  assign n1127 = ( n631 & n632 ) | ( n631 & ~n742 ) | ( n632 & ~n742 ) ;
  assign n1128 = ~x130 & n1127 ;
  assign n1129 = ( n759 & ~n760 ) | ( n759 & n1128 ) | ( ~n760 & n1128 ) ;
  assign n1130 = x133 & ~n1129 ;
  assign n1131 = x133 & ~n1126 ;
  assign n1132 = ( n1126 & ~n1130 ) | ( n1126 & n1131 ) | ( ~n1130 & n1131 ) ;
  assign n1133 = ~x132 & n1132 ;
  assign n1134 = ( x132 & ~n1123 ) | ( x132 & n1133 ) | ( ~n1123 & n1133 ) ;
  assign n1135 = x134 & ~n1134 ;
  assign n1136 = x134 & ~n1113 ;
  assign n1137 = ( n1113 & ~n1135 ) | ( n1113 & n1136 ) | ( ~n1135 & n1136 ) ;
  assign n1138 = ( ~n775 & n810 ) | ( ~n775 & n811 ) | ( n810 & n811 ) ;
  assign n1139 = ~x130 & n1138 ;
  assign n1140 = ( n784 & ~n785 ) | ( n784 & n1139 ) | ( ~n785 & n1139 ) ;
  assign n1141 = ( ~n793 & n828 ) | ( ~n793 & n829 ) | ( n828 & n829 ) ;
  assign n1142 = ~x130 & n1141 ;
  assign n1143 = ( n802 & ~n803 ) | ( n802 & n1142 ) | ( ~n803 & n1142 ) ;
  assign n1144 = x133 & ~n1143 ;
  assign n1145 = x133 & ~n1140 ;
  assign n1146 = ( n1140 & ~n1144 ) | ( n1140 & n1145 ) | ( ~n1144 & n1145 ) ;
  assign n1147 = x132 & ~n1146 ;
  assign n1148 = ( ~n812 & n885 ) | ( ~n812 & n886 ) | ( n885 & n886 ) ;
  assign n1149 = ~x130 & n1148 ;
  assign n1150 = ( n821 & ~n822 ) | ( n821 & n1149 ) | ( ~n822 & n1149 ) ;
  assign n1151 = ( n773 & n774 ) | ( n773 & ~n830 ) | ( n774 & ~n830 ) ;
  assign n1152 = ~x130 & n1151 ;
  assign n1153 = ( n839 & ~n840 ) | ( n839 & n1152 ) | ( ~n840 & n1152 ) ;
  assign n1154 = x133 & ~n1153 ;
  assign n1155 = x133 & ~n1150 ;
  assign n1156 = ( n1150 & ~n1154 ) | ( n1150 & n1155 ) | ( ~n1154 & n1155 ) ;
  assign n1157 = ~x132 & n1156 ;
  assign n1158 = ( x132 & ~n1147 ) | ( x132 & n1157 ) | ( ~n1147 & n1157 ) ;
  assign n1159 = ( ~n850 & n866 ) | ( ~n850 & n867 ) | ( n866 & n867 ) ;
  assign n1160 = ~x130 & n1159 ;
  assign n1161 = ( n859 & ~n860 ) | ( n859 & n1160 ) | ( ~n860 & n1160 ) ;
  assign n1162 = ( ~n887 & n903 ) | ( ~n887 & n904 ) | ( n903 & n904 ) ;
  assign n1163 = ~x130 & n1162 ;
  assign n1164 = ( n896 & ~n897 ) | ( n896 & n1163 ) | ( ~n897 & n1163 ) ;
  assign n1165 = x133 & ~n1164 ;
  assign n1166 = x133 & ~n1161 ;
  assign n1167 = ( n1161 & ~n1165 ) | ( n1161 & n1166 ) | ( ~n1165 & n1166 ) ;
  assign n1168 = x132 & ~n1167 ;
  assign n1169 = ( n791 & n792 ) | ( n791 & ~n868 ) | ( n792 & ~n868 ) ;
  assign n1170 = ~x130 & n1169 ;
  assign n1171 = ( n877 & ~n878 ) | ( n877 & n1170 ) | ( ~n878 & n1170 ) ;
  assign n1172 = ( n848 & n849 ) | ( n848 & ~n905 ) | ( n849 & ~n905 ) ;
  assign n1173 = ~x130 & n1172 ;
  assign n1174 = ( n914 & ~n915 ) | ( n914 & n1173 ) | ( ~n915 & n1173 ) ;
  assign n1175 = x133 & ~n1174 ;
  assign n1176 = x133 & ~n1171 ;
  assign n1177 = ( n1171 & ~n1175 ) | ( n1171 & n1176 ) | ( ~n1175 & n1176 ) ;
  assign n1178 = ~x132 & n1177 ;
  assign n1179 = ( x132 & ~n1168 ) | ( x132 & n1178 ) | ( ~n1168 & n1178 ) ;
  assign n1180 = x134 & ~n1179 ;
  assign n1181 = x134 & ~n1158 ;
  assign n1182 = ( n1158 & ~n1180 ) | ( n1158 & n1181 ) | ( ~n1180 & n1181 ) ;
  assign n1183 = ( ~n956 & n998 ) | ( ~n956 & n999 ) | ( n998 & n999 ) ;
  assign n1184 = ~x130 & n1183 ;
  assign n1185 = ( n963 & ~n964 ) | ( n963 & n1184 ) | ( ~n964 & n1184 ) ;
  assign n1186 = ( n924 & n925 ) | ( n924 & ~n969 ) | ( n925 & ~n969 ) ;
  assign n1187 = ~x130 & n1186 ;
  assign n1188 = ( n976 & ~n977 ) | ( n976 & n1187 ) | ( ~n977 & n1187 ) ;
  assign n1189 = x133 & ~n1188 ;
  assign n1190 = x133 & ~n1185 ;
  assign n1191 = ( n1185 & ~n1189 ) | ( n1185 & n1190 ) | ( ~n1189 & n1190 ) ;
  assign n1192 = ~x132 & n1191 ;
  assign n1193 = ( ~n926 & n954 ) | ( ~n926 & n955 ) | ( n954 & n955 ) ;
  assign n1194 = ~x130 & n1193 ;
  assign n1195 = ( n933 & ~n934 ) | ( n933 & n1194 ) | ( ~n934 & n1194 ) ;
  assign n1196 = ( ~n939 & n967 ) | ( ~n939 & n968 ) | ( n967 & n968 ) ;
  assign n1197 = ~x130 & n1196 ;
  assign n1198 = ( n946 & ~n947 ) | ( n946 & n1197 ) | ( ~n947 & n1197 ) ;
  assign n1199 = x133 & ~n1198 ;
  assign n1200 = x133 & ~n1195 ;
  assign n1201 = ( n1195 & ~n1199 ) | ( n1195 & n1200 ) | ( ~n1199 & n1200 ) ;
  assign n1202 = x132 & n1201 ;
  assign n1203 = n1192 | n1202 ;
  assign n1204 = ( ~n987 & n1015 ) | ( ~n987 & n1016 ) | ( n1015 & n1016 ) ;
  assign n1205 = ~x130 & n1204 ;
  assign n1206 = ( n994 & ~n995 ) | ( n994 & n1205 ) | ( ~n995 & n1205 ) ;
  assign n1207 = ~x133 & n1206 ;
  assign n1208 = ( ~n1000 & n1028 ) | ( ~n1000 & n1029 ) | ( n1028 & n1029 ) ;
  assign n1209 = ~x130 & n1208 ;
  assign n1210 = ( n1007 & ~n1008 ) | ( n1007 & n1209 ) | ( ~n1008 & n1209 ) ;
  assign n1211 = x133 & ~n1210 ;
  assign n1212 = ( x133 & n1207 ) | ( x133 & ~n1211 ) | ( n1207 & ~n1211 ) ;
  assign n1213 = x132 & ~n1212 ;
  assign n1214 = ( n937 & n938 ) | ( n937 & ~n1017 ) | ( n938 & ~n1017 ) ;
  assign n1215 = ~x130 & n1214 ;
  assign n1216 = ( n1024 & ~n1025 ) | ( n1024 & n1215 ) | ( ~n1025 & n1215 ) ;
  assign n1217 = ~x133 & n1216 ;
  assign n1218 = ( n985 & n986 ) | ( n985 & ~n1030 ) | ( n986 & ~n1030 ) ;
  assign n1219 = ~x130 & n1218 ;
  assign n1220 = ( n1037 & ~n1038 ) | ( n1037 & n1219 ) | ( ~n1038 & n1219 ) ;
  assign n1221 = x133 & ~n1220 ;
  assign n1222 = ( x133 & n1217 ) | ( x133 & ~n1221 ) | ( n1217 & ~n1221 ) ;
  assign n1223 = ~x132 & n1222 ;
  assign n1224 = ( x132 & ~n1213 ) | ( x132 & n1223 ) | ( ~n1213 & n1223 ) ;
  assign n1225 = x134 & ~n1224 ;
  assign n1226 = x134 & ~n1203 ;
  assign n1227 = ( n1203 & ~n1225 ) | ( n1203 & n1226 ) | ( ~n1225 & n1226 ) ;
  assign n1228 = ( ~n173 & n257 ) | ( ~n173 & n258 ) | ( n257 & n258 ) ;
  assign n1229 = ~x130 & n1228 ;
  assign n1230 = ( n1048 & ~n1049 ) | ( n1048 & n1229 ) | ( ~n1049 & n1229 ) ;
  assign n1231 = ( ~n214 & n298 ) | ( ~n214 & n299 ) | ( n298 & n299 ) ;
  assign n1232 = ~x130 & n1231 ;
  assign n1233 = ( n1051 & ~n1052 ) | ( n1051 & n1232 ) | ( ~n1052 & n1232 ) ;
  assign n1234 = x133 & ~n1233 ;
  assign n1235 = x133 & ~n1230 ;
  assign n1236 = ( n1230 & ~n1234 ) | ( n1230 & n1235 ) | ( ~n1234 & n1235 ) ;
  assign n1237 = x132 & ~n1236 ;
  assign n1238 = ( ~n259 & n385 ) | ( ~n259 & n386 ) | ( n385 & n386 ) ;
  assign n1239 = ~x130 & n1238 ;
  assign n1240 = ( n1058 & ~n1059 ) | ( n1058 & n1239 ) | ( ~n1059 & n1239 ) ;
  assign n1241 = ( n171 & n172 ) | ( n171 & ~n300 ) | ( n172 & ~n300 ) ;
  assign n1242 = ~x130 & n1241 ;
  assign n1243 = ( n1061 & ~n1062 ) | ( n1061 & n1242 ) | ( ~n1062 & n1242 ) ;
  assign n1244 = x133 & ~n1243 ;
  assign n1245 = x133 & ~n1240 ;
  assign n1246 = ( n1240 & ~n1244 ) | ( n1240 & n1245 ) | ( ~n1244 & n1245 ) ;
  assign n1247 = ~x132 & n1246 ;
  assign n1248 = ( x132 & ~n1237 ) | ( x132 & n1247 ) | ( ~n1237 & n1247 ) ;
  assign n1249 = ( ~n346 & n430 ) | ( ~n346 & n431 ) | ( n430 & n431 ) ;
  assign n1250 = ~x130 & n1249 ;
  assign n1251 = ( n1069 & ~n1070 ) | ( n1069 & n1250 ) | ( ~n1070 & n1250 ) ;
  assign n1252 = ( ~n387 & n471 ) | ( ~n387 & n472 ) | ( n471 & n472 ) ;
  assign n1253 = ~x130 & n1252 ;
  assign n1254 = ( n1072 & ~n1073 ) | ( n1072 & n1253 ) | ( ~n1073 & n1253 ) ;
  assign n1255 = x133 & ~n1254 ;
  assign n1256 = x133 & ~n1251 ;
  assign n1257 = ( n1251 & ~n1255 ) | ( n1251 & n1256 ) | ( ~n1255 & n1256 ) ;
  assign n1258 = x132 & ~n1257 ;
  assign n1259 = ( n212 & n213 ) | ( n212 & ~n432 ) | ( n213 & ~n432 ) ;
  assign n1260 = ~x130 & n1259 ;
  assign n1261 = ( n1079 & ~n1080 ) | ( n1079 & n1260 ) | ( ~n1080 & n1260 ) ;
  assign n1262 = ( n344 & n345 ) | ( n344 & ~n473 ) | ( n345 & ~n473 ) ;
  assign n1263 = ~x130 & n1262 ;
  assign n1264 = ( n1082 & ~n1083 ) | ( n1082 & n1263 ) | ( ~n1083 & n1263 ) ;
  assign n1265 = x133 & ~n1264 ;
  assign n1266 = x133 & ~n1261 ;
  assign n1267 = ( n1261 & ~n1265 ) | ( n1261 & n1266 ) | ( ~n1265 & n1266 ) ;
  assign n1268 = ~x132 & n1267 ;
  assign n1269 = ( x132 & ~n1258 ) | ( x132 & n1268 ) | ( ~n1258 & n1268 ) ;
  assign n1270 = x134 & ~n1269 ;
  assign n1271 = x134 & ~n1248 ;
  assign n1272 = ( n1248 & ~n1270 ) | ( n1248 & n1271 ) | ( ~n1270 & n1271 ) ;
  assign n1273 = ( ~n514 & n576 ) | ( ~n514 & n577 ) | ( n576 & n577 ) ;
  assign n1274 = ~x130 & n1273 ;
  assign n1275 = ( n1093 & ~n1094 ) | ( n1093 & n1274 ) | ( ~n1094 & n1274 ) ;
  assign n1276 = ( ~n547 & n609 ) | ( ~n547 & n610 ) | ( n609 & n610 ) ;
  assign n1277 = ~x130 & n1276 ;
  assign n1278 = ( n1096 & ~n1097 ) | ( n1096 & n1277 ) | ( ~n1097 & n1277 ) ;
  assign n1279 = x133 & ~n1278 ;
  assign n1280 = x133 & ~n1275 ;
  assign n1281 = ( n1275 & ~n1279 ) | ( n1275 & n1280 ) | ( ~n1279 & n1280 ) ;
  assign n1282 = x132 & ~n1281 ;
  assign n1283 = ( ~n584 & n680 ) | ( ~n584 & n681 ) | ( n680 & n681 ) ;
  assign n1284 = ~x130 & n1283 ;
  assign n1285 = ( n1103 & ~n1104 ) | ( n1103 & n1284 ) | ( ~n1104 & n1284 ) ;
  assign n1286 = ( n506 & n507 ) | ( n506 & ~n617 ) | ( n507 & ~n617 ) ;
  assign n1287 = ~x130 & n1286 ;
  assign n1288 = ( n1106 & ~n1107 ) | ( n1106 & n1287 ) | ( ~n1107 & n1287 ) ;
  assign n1289 = x133 & ~n1288 ;
  assign n1290 = x133 & ~n1285 ;
  assign n1291 = ( n1285 & ~n1289 ) | ( n1285 & n1290 ) | ( ~n1289 & n1290 ) ;
  assign n1292 = ~x132 & n1291 ;
  assign n1293 = ( x132 & ~n1282 ) | ( x132 & n1292 ) | ( ~n1282 & n1292 ) ;
  assign n1294 = ( ~n655 & n717 ) | ( ~n655 & n718 ) | ( n717 & n718 ) ;
  assign n1295 = ~x130 & n1294 ;
  assign n1296 = ( n1114 & ~n1115 ) | ( n1114 & n1295 ) | ( ~n1115 & n1295 ) ;
  assign n1297 = ( ~n688 & n750 ) | ( ~n688 & n751 ) | ( n750 & n751 ) ;
  assign n1298 = ~x130 & n1297 ;
  assign n1299 = ( n1117 & ~n1118 ) | ( n1117 & n1298 ) | ( ~n1118 & n1298 ) ;
  assign n1300 = x133 & ~n1299 ;
  assign n1301 = x133 & ~n1296 ;
  assign n1302 = ( n1296 & ~n1300 ) | ( n1296 & n1301 ) | ( ~n1300 & n1301 ) ;
  assign n1303 = x132 & ~n1302 ;
  assign n1304 = ( n539 & n540 ) | ( n539 & ~n725 ) | ( n540 & ~n725 ) ;
  assign n1305 = ~x130 & n1304 ;
  assign n1306 = ( n1124 & ~n1125 ) | ( n1124 & n1305 ) | ( ~n1125 & n1305 ) ;
  assign n1307 = ( n647 & n648 ) | ( n647 & ~n758 ) | ( n648 & ~n758 ) ;
  assign n1308 = ~x130 & n1307 ;
  assign n1309 = ( n1127 & ~n1128 ) | ( n1127 & n1308 ) | ( ~n1128 & n1308 ) ;
  assign n1310 = x133 & ~n1309 ;
  assign n1311 = x133 & ~n1306 ;
  assign n1312 = ( n1306 & ~n1310 ) | ( n1306 & n1311 ) | ( ~n1310 & n1311 ) ;
  assign n1313 = ~x132 & n1312 ;
  assign n1314 = ( x132 & ~n1303 ) | ( x132 & n1313 ) | ( ~n1303 & n1313 ) ;
  assign n1315 = x134 & ~n1314 ;
  assign n1316 = x134 & ~n1293 ;
  assign n1317 = ( n1293 & ~n1315 ) | ( n1293 & n1316 ) | ( ~n1315 & n1316 ) ;
  assign n1318 = ( ~n783 & n818 ) | ( ~n783 & n819 ) | ( n818 & n819 ) ;
  assign n1319 = ~x130 & n1318 ;
  assign n1320 = ( n1138 & ~n1139 ) | ( n1138 & n1319 ) | ( ~n1139 & n1319 ) ;
  assign n1321 = ( ~n801 & n836 ) | ( ~n801 & n837 ) | ( n836 & n837 ) ;
  assign n1322 = ~x130 & n1321 ;
  assign n1323 = ( n1141 & ~n1142 ) | ( n1141 & n1322 ) | ( ~n1142 & n1322 ) ;
  assign n1324 = x133 & ~n1323 ;
  assign n1325 = x133 & ~n1320 ;
  assign n1326 = ( n1320 & ~n1324 ) | ( n1320 & n1325 ) | ( ~n1324 & n1325 ) ;
  assign n1327 = x132 & ~n1326 ;
  assign n1328 = ( ~n820 & n893 ) | ( ~n820 & n894 ) | ( n893 & n894 ) ;
  assign n1329 = ~x130 & n1328 ;
  assign n1330 = ( n1148 & ~n1149 ) | ( n1148 & n1329 ) | ( ~n1149 & n1329 ) ;
  assign n1331 = ( n781 & n782 ) | ( n781 & ~n838 ) | ( n782 & ~n838 ) ;
  assign n1332 = ~x130 & n1331 ;
  assign n1333 = ( n1151 & ~n1152 ) | ( n1151 & n1332 ) | ( ~n1152 & n1332 ) ;
  assign n1334 = x133 & ~n1333 ;
  assign n1335 = x133 & ~n1330 ;
  assign n1336 = ( n1330 & ~n1334 ) | ( n1330 & n1335 ) | ( ~n1334 & n1335 ) ;
  assign n1337 = ~x132 & n1336 ;
  assign n1338 = ( x132 & ~n1327 ) | ( x132 & n1337 ) | ( ~n1327 & n1337 ) ;
  assign n1339 = ( ~n858 & n874 ) | ( ~n858 & n875 ) | ( n874 & n875 ) ;
  assign n1340 = ~x130 & n1339 ;
  assign n1341 = ( n1159 & ~n1160 ) | ( n1159 & n1340 ) | ( ~n1160 & n1340 ) ;
  assign n1342 = ( ~n895 & n911 ) | ( ~n895 & n912 ) | ( n911 & n912 ) ;
  assign n1343 = ~x130 & n1342 ;
  assign n1344 = ( n1162 & ~n1163 ) | ( n1162 & n1343 ) | ( ~n1163 & n1343 ) ;
  assign n1345 = x133 & ~n1344 ;
  assign n1346 = x133 & ~n1341 ;
  assign n1347 = ( n1341 & ~n1345 ) | ( n1341 & n1346 ) | ( ~n1345 & n1346 ) ;
  assign n1348 = x132 & ~n1347 ;
  assign n1349 = ( n799 & n800 ) | ( n799 & ~n876 ) | ( n800 & ~n876 ) ;
  assign n1350 = ~x130 & n1349 ;
  assign n1351 = ( n1169 & ~n1170 ) | ( n1169 & n1350 ) | ( ~n1170 & n1350 ) ;
  assign n1352 = ( n856 & n857 ) | ( n856 & ~n913 ) | ( n857 & ~n913 ) ;
  assign n1353 = ~x130 & n1352 ;
  assign n1354 = ( n1172 & ~n1173 ) | ( n1172 & n1353 ) | ( ~n1173 & n1353 ) ;
  assign n1355 = x133 & ~n1354 ;
  assign n1356 = x133 & ~n1351 ;
  assign n1357 = ( n1351 & ~n1355 ) | ( n1351 & n1356 ) | ( ~n1355 & n1356 ) ;
  assign n1358 = ~x132 & n1357 ;
  assign n1359 = ( x132 & ~n1348 ) | ( x132 & n1358 ) | ( ~n1348 & n1358 ) ;
  assign n1360 = x134 & ~n1359 ;
  assign n1361 = x134 & ~n1338 ;
  assign n1362 = ( n1338 & ~n1360 ) | ( n1338 & n1361 ) | ( ~n1360 & n1361 ) ;
  assign n1363 = ( ~n932 & n960 ) | ( ~n932 & n961 ) | ( n960 & n961 ) ;
  assign n1364 = ~x130 & n1363 ;
  assign n1365 = ( n1193 & ~n1194 ) | ( n1193 & n1364 ) | ( ~n1194 & n1364 ) ;
  assign n1366 = ( ~n945 & n973 ) | ( ~n945 & n974 ) | ( n973 & n974 ) ;
  assign n1367 = ~x130 & n1366 ;
  assign n1368 = ( n1196 & ~n1197 ) | ( n1196 & n1367 ) | ( ~n1197 & n1367 ) ;
  assign n1369 = x133 & ~n1368 ;
  assign n1370 = x133 & ~n1365 ;
  assign n1371 = ( n1365 & ~n1369 ) | ( n1365 & n1370 ) | ( ~n1369 & n1370 ) ;
  assign n1372 = x132 & ~n1371 ;
  assign n1373 = ( ~n962 & n1004 ) | ( ~n962 & n1005 ) | ( n1004 & n1005 ) ;
  assign n1374 = ~x130 & n1373 ;
  assign n1375 = ( n1183 & ~n1184 ) | ( n1183 & n1374 ) | ( ~n1184 & n1374 ) ;
  assign n1376 = ( n930 & n931 ) | ( n930 & ~n975 ) | ( n931 & ~n975 ) ;
  assign n1377 = ~x130 & n1376 ;
  assign n1378 = ( n1186 & ~n1187 ) | ( n1186 & n1377 ) | ( ~n1187 & n1377 ) ;
  assign n1379 = x133 & ~n1378 ;
  assign n1380 = x133 & ~n1375 ;
  assign n1381 = ( n1375 & ~n1379 ) | ( n1375 & n1380 ) | ( ~n1379 & n1380 ) ;
  assign n1382 = ~x132 & n1381 ;
  assign n1383 = ( x132 & ~n1372 ) | ( x132 & n1382 ) | ( ~n1372 & n1382 ) ;
  assign n1384 = ( ~n993 & n1021 ) | ( ~n993 & n1022 ) | ( n1021 & n1022 ) ;
  assign n1385 = ~x130 & n1384 ;
  assign n1386 = ( n1204 & ~n1205 ) | ( n1204 & n1385 ) | ( ~n1205 & n1385 ) ;
  assign n1387 = ( ~n1006 & n1034 ) | ( ~n1006 & n1035 ) | ( n1034 & n1035 ) ;
  assign n1388 = ~x130 & n1387 ;
  assign n1389 = ( n1208 & ~n1209 ) | ( n1208 & n1388 ) | ( ~n1209 & n1388 ) ;
  assign n1390 = x133 & ~n1389 ;
  assign n1391 = x133 & ~n1386 ;
  assign n1392 = ( n1386 & ~n1390 ) | ( n1386 & n1391 ) | ( ~n1390 & n1391 ) ;
  assign n1393 = x132 & ~n1392 ;
  assign n1394 = ( n943 & n944 ) | ( n943 & ~n1023 ) | ( n944 & ~n1023 ) ;
  assign n1395 = ~x130 & n1394 ;
  assign n1396 = ( n1214 & ~n1215 ) | ( n1214 & n1395 ) | ( ~n1215 & n1395 ) ;
  assign n1397 = ( n991 & n992 ) | ( n991 & ~n1036 ) | ( n992 & ~n1036 ) ;
  assign n1398 = ~x130 & n1397 ;
  assign n1399 = ( n1218 & ~n1219 ) | ( n1218 & n1398 ) | ( ~n1219 & n1398 ) ;
  assign n1400 = x133 & ~n1399 ;
  assign n1401 = x133 & ~n1396 ;
  assign n1402 = ( n1396 & ~n1400 ) | ( n1396 & n1401 ) | ( ~n1400 & n1401 ) ;
  assign n1403 = ~x132 & n1402 ;
  assign n1404 = ( x132 & ~n1393 ) | ( x132 & n1403 ) | ( ~n1393 & n1403 ) ;
  assign n1405 = x134 & ~n1404 ;
  assign n1406 = x134 & ~n1383 ;
  assign n1407 = ( n1383 & ~n1405 ) | ( n1383 & n1406 ) | ( ~n1405 & n1406 ) ;
  assign n1408 = x130 & ~n1228 ;
  assign n1409 = ( n240 & n241 ) | ( n240 & ~n1408 ) | ( n241 & ~n1408 ) ;
  assign n1410 = x130 & ~n1231 ;
  assign n1411 = ( n281 & n282 ) | ( n281 & ~n1410 ) | ( n282 & ~n1410 ) ;
  assign n1412 = x133 & ~n1411 ;
  assign n1413 = x133 & ~n1409 ;
  assign n1414 = ( n1409 & ~n1412 ) | ( n1409 & n1413 ) | ( ~n1412 & n1413 ) ;
  assign n1415 = x132 & ~n1414 ;
  assign n1416 = x130 & ~n1238 ;
  assign n1417 = ( n368 & n369 ) | ( n368 & ~n1416 ) | ( n369 & ~n1416 ) ;
  assign n1418 = x130 & ~n1241 ;
  assign n1419 = ( n154 & n155 ) | ( n154 & ~n1418 ) | ( n155 & ~n1418 ) ;
  assign n1420 = x133 & ~n1419 ;
  assign n1421 = x133 & ~n1417 ;
  assign n1422 = ( n1417 & ~n1420 ) | ( n1417 & n1421 ) | ( ~n1420 & n1421 ) ;
  assign n1423 = ~x132 & n1422 ;
  assign n1424 = ( x132 & ~n1415 ) | ( x132 & n1423 ) | ( ~n1415 & n1423 ) ;
  assign n1425 = x130 & ~n1249 ;
  assign n1426 = ( n413 & n414 ) | ( n413 & ~n1425 ) | ( n414 & ~n1425 ) ;
  assign n1427 = x130 & ~n1252 ;
  assign n1428 = ( n454 & n455 ) | ( n454 & ~n1427 ) | ( n455 & ~n1427 ) ;
  assign n1429 = x133 & ~n1428 ;
  assign n1430 = x133 & ~n1426 ;
  assign n1431 = ( n1426 & ~n1429 ) | ( n1426 & n1430 ) | ( ~n1429 & n1430 ) ;
  assign n1432 = x132 & ~n1431 ;
  assign n1433 = x130 & ~n1259 ;
  assign n1434 = ( n195 & n196 ) | ( n195 & ~n1433 ) | ( n196 & ~n1433 ) ;
  assign n1435 = x130 & ~n1262 ;
  assign n1436 = ( n327 & n328 ) | ( n327 & ~n1435 ) | ( n328 & ~n1435 ) ;
  assign n1437 = x133 & ~n1436 ;
  assign n1438 = x133 & ~n1434 ;
  assign n1439 = ( n1434 & ~n1437 ) | ( n1434 & n1438 ) | ( ~n1437 & n1438 ) ;
  assign n1440 = ~x132 & n1439 ;
  assign n1441 = ( x132 & ~n1432 ) | ( x132 & n1440 ) | ( ~n1432 & n1440 ) ;
  assign n1442 = x134 & ~n1441 ;
  assign n1443 = x134 & ~n1424 ;
  assign n1444 = ( n1424 & ~n1442 ) | ( n1424 & n1443 ) | ( ~n1442 & n1443 ) ;
  assign n1445 = x130 & ~n1273 ;
  assign n1446 = ( n569 & n570 ) | ( n569 & ~n1445 ) | ( n570 & ~n1445 ) ;
  assign n1447 = x130 & ~n1276 ;
  assign n1448 = ( n602 & n603 ) | ( n602 & ~n1447 ) | ( n603 & ~n1447 ) ;
  assign n1449 = x133 & ~n1448 ;
  assign n1450 = x133 & ~n1446 ;
  assign n1451 = ( n1446 & ~n1449 ) | ( n1446 & n1450 ) | ( ~n1449 & n1450 ) ;
  assign n1452 = x132 & ~n1451 ;
  assign n1453 = x130 & ~n1283 ;
  assign n1454 = ( n673 & n674 ) | ( n673 & ~n1453 ) | ( n674 & ~n1453 ) ;
  assign n1455 = x130 & ~n1286 ;
  assign n1456 = ( n499 & n500 ) | ( n499 & ~n1455 ) | ( n500 & ~n1455 ) ;
  assign n1457 = x133 & ~n1456 ;
  assign n1458 = x133 & ~n1454 ;
  assign n1459 = ( n1454 & ~n1457 ) | ( n1454 & n1458 ) | ( ~n1457 & n1458 ) ;
  assign n1460 = ~x132 & n1459 ;
  assign n1461 = ( x132 & ~n1452 ) | ( x132 & n1460 ) | ( ~n1452 & n1460 ) ;
  assign n1462 = x130 & ~n1294 ;
  assign n1463 = ( n710 & n711 ) | ( n710 & ~n1462 ) | ( n711 & ~n1462 ) ;
  assign n1464 = x130 & ~n1297 ;
  assign n1465 = ( n743 & n744 ) | ( n743 & ~n1464 ) | ( n744 & ~n1464 ) ;
  assign n1466 = x133 & ~n1465 ;
  assign n1467 = x133 & ~n1463 ;
  assign n1468 = ( n1463 & ~n1466 ) | ( n1463 & n1467 ) | ( ~n1466 & n1467 ) ;
  assign n1469 = x132 & ~n1468 ;
  assign n1470 = x130 & ~n1304 ;
  assign n1471 = ( n532 & n533 ) | ( n532 & ~n1470 ) | ( n533 & ~n1470 ) ;
  assign n1472 = x130 & ~n1307 ;
  assign n1473 = ( n640 & n641 ) | ( n640 & ~n1472 ) | ( n641 & ~n1472 ) ;
  assign n1474 = x133 & ~n1473 ;
  assign n1475 = x133 & ~n1471 ;
  assign n1476 = ( n1471 & ~n1474 ) | ( n1471 & n1475 ) | ( ~n1474 & n1475 ) ;
  assign n1477 = ~x132 & n1476 ;
  assign n1478 = ( x132 & ~n1469 ) | ( x132 & n1477 ) | ( ~n1469 & n1477 ) ;
  assign n1479 = x134 & ~n1478 ;
  assign n1480 = x134 & ~n1461 ;
  assign n1481 = ( n1461 & ~n1479 ) | ( n1461 & n1480 ) | ( ~n1479 & n1480 ) ;
  assign n1482 = x130 & ~n1318 ;
  assign n1483 = ( n813 & n814 ) | ( n813 & ~n1482 ) | ( n814 & ~n1482 ) ;
  assign n1484 = x130 & ~n1321 ;
  assign n1485 = ( n831 & n832 ) | ( n831 & ~n1484 ) | ( n832 & ~n1484 ) ;
  assign n1486 = x133 & ~n1485 ;
  assign n1487 = x133 & ~n1483 ;
  assign n1488 = ( n1483 & ~n1486 ) | ( n1483 & n1487 ) | ( ~n1486 & n1487 ) ;
  assign n1489 = x132 & ~n1488 ;
  assign n1490 = x130 & ~n1328 ;
  assign n1491 = ( n888 & n889 ) | ( n888 & ~n1490 ) | ( n889 & ~n1490 ) ;
  assign n1492 = x130 & ~n1331 ;
  assign n1493 = ( n776 & n777 ) | ( n776 & ~n1492 ) | ( n777 & ~n1492 ) ;
  assign n1494 = x133 & ~n1493 ;
  assign n1495 = x133 & ~n1491 ;
  assign n1496 = ( n1491 & ~n1494 ) | ( n1491 & n1495 ) | ( ~n1494 & n1495 ) ;
  assign n1497 = ~x132 & n1496 ;
  assign n1498 = ( x132 & ~n1489 ) | ( x132 & n1497 ) | ( ~n1489 & n1497 ) ;
  assign n1499 = x130 & ~n1339 ;
  assign n1500 = ( n869 & n870 ) | ( n869 & ~n1499 ) | ( n870 & ~n1499 ) ;
  assign n1501 = x130 & ~n1342 ;
  assign n1502 = ( n906 & n907 ) | ( n906 & ~n1501 ) | ( n907 & ~n1501 ) ;
  assign n1503 = x133 & ~n1502 ;
  assign n1504 = x133 & ~n1500 ;
  assign n1505 = ( n1500 & ~n1503 ) | ( n1500 & n1504 ) | ( ~n1503 & n1504 ) ;
  assign n1506 = x132 & ~n1505 ;
  assign n1507 = x130 & ~n1349 ;
  assign n1508 = ( n794 & n795 ) | ( n794 & ~n1507 ) | ( n795 & ~n1507 ) ;
  assign n1509 = x130 & ~n1352 ;
  assign n1510 = ( n851 & n852 ) | ( n851 & ~n1509 ) | ( n852 & ~n1509 ) ;
  assign n1511 = x133 & ~n1510 ;
  assign n1512 = x133 & ~n1508 ;
  assign n1513 = ( n1508 & ~n1511 ) | ( n1508 & n1512 ) | ( ~n1511 & n1512 ) ;
  assign n1514 = ~x132 & n1513 ;
  assign n1515 = ( x132 & ~n1506 ) | ( x132 & n1514 ) | ( ~n1506 & n1514 ) ;
  assign n1516 = x134 & ~n1515 ;
  assign n1517 = x134 & ~n1498 ;
  assign n1518 = ( n1498 & ~n1516 ) | ( n1498 & n1517 ) | ( ~n1516 & n1517 ) ;
  assign n1519 = x130 & ~n1363 ;
  assign n1520 = ( n957 & n958 ) | ( n957 & ~n1519 ) | ( n958 & ~n1519 ) ;
  assign n1521 = x130 & ~n1366 ;
  assign n1522 = ( n970 & n971 ) | ( n970 & ~n1521 ) | ( n971 & ~n1521 ) ;
  assign n1523 = x133 & ~n1522 ;
  assign n1524 = x133 & ~n1520 ;
  assign n1525 = ( n1520 & ~n1523 ) | ( n1520 & n1524 ) | ( ~n1523 & n1524 ) ;
  assign n1526 = x132 & ~n1525 ;
  assign n1527 = x130 & ~n1373 ;
  assign n1528 = ( n1001 & n1002 ) | ( n1001 & ~n1527 ) | ( n1002 & ~n1527 ) ;
  assign n1529 = x130 & ~n1376 ;
  assign n1530 = ( n927 & n928 ) | ( n927 & ~n1529 ) | ( n928 & ~n1529 ) ;
  assign n1531 = x133 & ~n1530 ;
  assign n1532 = x133 & ~n1528 ;
  assign n1533 = ( n1528 & ~n1531 ) | ( n1528 & n1532 ) | ( ~n1531 & n1532 ) ;
  assign n1534 = ~x132 & n1533 ;
  assign n1535 = ( x132 & ~n1526 ) | ( x132 & n1534 ) | ( ~n1526 & n1534 ) ;
  assign n1536 = x130 & ~n1384 ;
  assign n1537 = ( n1018 & n1019 ) | ( n1018 & ~n1536 ) | ( n1019 & ~n1536 ) ;
  assign n1538 = x130 & ~n1387 ;
  assign n1539 = ( n1031 & n1032 ) | ( n1031 & ~n1538 ) | ( n1032 & ~n1538 ) ;
  assign n1540 = x133 & ~n1539 ;
  assign n1541 = x133 & ~n1537 ;
  assign n1542 = ( n1537 & ~n1540 ) | ( n1537 & n1541 ) | ( ~n1540 & n1541 ) ;
  assign n1543 = x132 & ~n1542 ;
  assign n1544 = x130 & ~n1394 ;
  assign n1545 = ( n940 & n941 ) | ( n940 & ~n1544 ) | ( n941 & ~n1544 ) ;
  assign n1546 = x130 & ~n1397 ;
  assign n1547 = ( n988 & n989 ) | ( n988 & ~n1546 ) | ( n989 & ~n1546 ) ;
  assign n1548 = x133 & ~n1547 ;
  assign n1549 = x133 & ~n1545 ;
  assign n1550 = ( n1545 & ~n1548 ) | ( n1545 & n1549 ) | ( ~n1548 & n1549 ) ;
  assign n1551 = ~x132 & n1550 ;
  assign n1552 = ( x132 & ~n1543 ) | ( x132 & n1551 ) | ( ~n1543 & n1551 ) ;
  assign n1553 = x134 & ~n1552 ;
  assign n1554 = x134 & ~n1535 ;
  assign n1555 = ( n1535 & ~n1553 ) | ( n1535 & n1554 ) | ( ~n1553 & n1554 ) ;
  assign n1556 = ( ~n219 & n390 ) | ( ~n219 & n391 ) | ( n390 & n391 ) ;
  assign n1557 = ~x132 & n1556 ;
  assign n1558 = ( n306 & ~n307 ) | ( n306 & n1557 ) | ( ~n307 & n1557 ) ;
  assign n1559 = ( n217 & n218 ) | ( n217 & ~n392 ) | ( n218 & ~n392 ) ;
  assign n1560 = ~x132 & n1559 ;
  assign n1561 = ( n479 & ~n480 ) | ( n479 & n1560 ) | ( ~n480 & n1560 ) ;
  assign n1562 = x134 & ~n1561 ;
  assign n1563 = x134 & ~n1558 ;
  assign n1564 = ( n1558 & ~n1562 ) | ( n1558 & n1563 ) | ( ~n1562 & n1563 ) ;
  assign n1565 = ( ~n552 & n691 ) | ( ~n552 & n692 ) | ( n691 & n692 ) ;
  assign n1566 = ~x132 & n1565 ;
  assign n1567 = ( n623 & ~n624 ) | ( n623 & n1566 ) | ( ~n624 & n1566 ) ;
  assign n1568 = ( n550 & n551 ) | ( n550 & ~n693 ) | ( n551 & ~n693 ) ;
  assign n1569 = ~x132 & n1568 ;
  assign n1570 = ( n764 & ~n765 ) | ( n764 & n1569 ) | ( ~n765 & n1569 ) ;
  assign n1571 = x134 & ~n1570 ;
  assign n1572 = x134 & ~n1567 ;
  assign n1573 = ( n1567 & ~n1571 ) | ( n1567 & n1572 ) | ( ~n1571 & n1572 ) ;
  assign n1574 = ~x133 & n879 ;
  assign n1575 = x133 & n861 ;
  assign n1576 = ( n804 & ~n805 ) | ( n804 & n1575 ) | ( ~n805 & n1575 ) ;
  assign n1577 = x132 | n1576 ;
  assign n1578 = x133 & n916 ;
  assign n1579 = ( x132 & n1574 ) | ( x132 & ~n1578 ) | ( n1574 & ~n1578 ) ;
  assign n1580 = ( n1574 & n1577 ) | ( n1574 & ~n1579 ) | ( n1577 & ~n1579 ) ;
  assign n1581 = x134 & ~n1580 ;
  assign n1582 = n824 | n842 ;
  assign n1583 = ~x133 & n898 ;
  assign n1584 = ( n786 & ~n787 ) | ( n786 & n1583 ) | ( ~n787 & n1583 ) ;
  assign n1585 = ~x132 & n1584 ;
  assign n1586 = ( ~n843 & n1582 ) | ( ~n843 & n1585 ) | ( n1582 & n1585 ) ;
  assign n1587 = x134 & ~n1586 ;
  assign n1588 = ( ~n1581 & n1586 ) | ( ~n1581 & n1587 ) | ( n1586 & n1587 ) ;
  assign n1589 = ( ~n950 & n1009 ) | ( ~n950 & n1010 ) | ( n1009 & n1010 ) ;
  assign n1590 = ~x132 & n1589 ;
  assign n1591 = ( n981 & ~n982 ) | ( n981 & n1590 ) | ( ~n982 & n1590 ) ;
  assign n1592 = ( n948 & n949 ) | ( n948 & ~n1011 ) | ( n949 & ~n1011 ) ;
  assign n1593 = ~x132 & n1592 ;
  assign n1594 = ( n1042 & ~n1043 ) | ( n1042 & n1593 ) | ( ~n1043 & n1593 ) ;
  assign n1595 = x134 & ~n1594 ;
  assign n1596 = x134 & ~n1591 ;
  assign n1597 = ( n1591 & ~n1595 ) | ( n1591 & n1596 ) | ( ~n1595 & n1596 ) ;
  assign n1598 = ( ~n1055 & n1074 ) | ( ~n1055 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1599 = ~x132 & n1598 ;
  assign n1600 = ( n1066 & ~n1067 ) | ( n1066 & n1599 ) | ( ~n1067 & n1599 ) ;
  assign n1601 = ( n1053 & n1054 ) | ( n1053 & ~n1076 ) | ( n1054 & ~n1076 ) ;
  assign n1602 = ~x132 & n1601 ;
  assign n1603 = ( n1087 & ~n1088 ) | ( n1087 & n1602 ) | ( ~n1088 & n1602 ) ;
  assign n1604 = x134 & ~n1603 ;
  assign n1605 = x134 & ~n1600 ;
  assign n1606 = ( n1600 & ~n1604 ) | ( n1600 & n1605 ) | ( ~n1604 & n1605 ) ;
  assign n1607 = ( ~n1100 & n1119 ) | ( ~n1100 & n1120 ) | ( n1119 & n1120 ) ;
  assign n1608 = ~x132 & n1607 ;
  assign n1609 = ( n1111 & ~n1112 ) | ( n1111 & n1608 ) | ( ~n1112 & n1608 ) ;
  assign n1610 = ( n1098 & n1099 ) | ( n1098 & ~n1121 ) | ( n1099 & ~n1121 ) ;
  assign n1611 = ~x132 & n1610 ;
  assign n1612 = ( n1132 & ~n1133 ) | ( n1132 & n1611 ) | ( ~n1133 & n1611 ) ;
  assign n1613 = x134 & ~n1612 ;
  assign n1614 = x134 & ~n1609 ;
  assign n1615 = ( n1609 & ~n1613 ) | ( n1609 & n1614 ) | ( ~n1613 & n1614 ) ;
  assign n1616 = ( ~n1145 & n1164 ) | ( ~n1145 & n1165 ) | ( n1164 & n1165 ) ;
  assign n1617 = ~x132 & n1616 ;
  assign n1618 = ( n1156 & ~n1157 ) | ( n1156 & n1617 ) | ( ~n1157 & n1617 ) ;
  assign n1619 = ( n1143 & n1144 ) | ( n1143 & ~n1166 ) | ( n1144 & ~n1166 ) ;
  assign n1620 = ~x132 & n1619 ;
  assign n1621 = ( n1177 & ~n1178 ) | ( n1177 & n1620 ) | ( ~n1178 & n1620 ) ;
  assign n1622 = x134 & ~n1621 ;
  assign n1623 = x134 & ~n1618 ;
  assign n1624 = ( n1618 & ~n1622 ) | ( n1618 & n1623 ) | ( ~n1622 & n1623 ) ;
  assign n1625 = ~x133 & n1198 ;
  assign n1626 = x133 & n1206 ;
  assign n1627 = ( ~x132 & n1625 ) | ( ~x132 & n1626 ) | ( n1625 & n1626 ) ;
  assign n1628 = ( n1222 & ~n1223 ) | ( n1222 & n1627 ) | ( ~n1223 & n1627 ) ;
  assign n1629 = x134 & ~n1628 ;
  assign n1630 = ( ~n1200 & n1210 ) | ( ~n1200 & n1211 ) | ( n1210 & n1211 ) ;
  assign n1631 = ~x132 & n1630 ;
  assign n1632 = ( n1191 & ~n1192 ) | ( n1191 & n1631 ) | ( ~n1192 & n1631 ) ;
  assign n1633 = x134 & ~n1632 ;
  assign n1634 = ( ~n1629 & n1632 ) | ( ~n1629 & n1633 ) | ( n1632 & n1633 ) ;
  assign n1635 = ( ~n1235 & n1254 ) | ( ~n1235 & n1255 ) | ( n1254 & n1255 ) ;
  assign n1636 = ~x132 & n1635 ;
  assign n1637 = ( n1246 & ~n1247 ) | ( n1246 & n1636 ) | ( ~n1247 & n1636 ) ;
  assign n1638 = ( n1233 & n1234 ) | ( n1233 & ~n1256 ) | ( n1234 & ~n1256 ) ;
  assign n1639 = ~x132 & n1638 ;
  assign n1640 = ( n1267 & ~n1268 ) | ( n1267 & n1639 ) | ( ~n1268 & n1639 ) ;
  assign n1641 = x134 & ~n1640 ;
  assign n1642 = x134 & ~n1637 ;
  assign n1643 = ( n1637 & ~n1641 ) | ( n1637 & n1642 ) | ( ~n1641 & n1642 ) ;
  assign n1644 = ( ~n1280 & n1299 ) | ( ~n1280 & n1300 ) | ( n1299 & n1300 ) ;
  assign n1645 = ~x132 & n1644 ;
  assign n1646 = ( n1291 & ~n1292 ) | ( n1291 & n1645 ) | ( ~n1292 & n1645 ) ;
  assign n1647 = ( n1278 & n1279 ) | ( n1278 & ~n1301 ) | ( n1279 & ~n1301 ) ;
  assign n1648 = ~x132 & n1647 ;
  assign n1649 = ( n1312 & ~n1313 ) | ( n1312 & n1648 ) | ( ~n1313 & n1648 ) ;
  assign n1650 = x134 & ~n1649 ;
  assign n1651 = x134 & ~n1646 ;
  assign n1652 = ( n1646 & ~n1650 ) | ( n1646 & n1651 ) | ( ~n1650 & n1651 ) ;
  assign n1653 = ( ~n1325 & n1344 ) | ( ~n1325 & n1345 ) | ( n1344 & n1345 ) ;
  assign n1654 = ~x132 & n1653 ;
  assign n1655 = ( n1336 & ~n1337 ) | ( n1336 & n1654 ) | ( ~n1337 & n1654 ) ;
  assign n1656 = ( n1323 & n1324 ) | ( n1323 & ~n1346 ) | ( n1324 & ~n1346 ) ;
  assign n1657 = ~x132 & n1656 ;
  assign n1658 = ( n1357 & ~n1358 ) | ( n1357 & n1657 ) | ( ~n1358 & n1657 ) ;
  assign n1659 = x134 & ~n1658 ;
  assign n1660 = x134 & ~n1655 ;
  assign n1661 = ( n1655 & ~n1659 ) | ( n1655 & n1660 ) | ( ~n1659 & n1660 ) ;
  assign n1662 = ( ~n1370 & n1389 ) | ( ~n1370 & n1390 ) | ( n1389 & n1390 ) ;
  assign n1663 = ~x132 & n1662 ;
  assign n1664 = ( n1381 & ~n1382 ) | ( n1381 & n1663 ) | ( ~n1382 & n1663 ) ;
  assign n1665 = ( n1368 & n1369 ) | ( n1368 & ~n1391 ) | ( n1369 & ~n1391 ) ;
  assign n1666 = ~x132 & n1665 ;
  assign n1667 = ( n1402 & ~n1403 ) | ( n1402 & n1666 ) | ( ~n1403 & n1666 ) ;
  assign n1668 = x134 & ~n1667 ;
  assign n1669 = x134 & ~n1664 ;
  assign n1670 = ( n1664 & ~n1668 ) | ( n1664 & n1669 ) | ( ~n1668 & n1669 ) ;
  assign n1671 = ( ~n1413 & n1428 ) | ( ~n1413 & n1429 ) | ( n1428 & n1429 ) ;
  assign n1672 = ~x132 & n1671 ;
  assign n1673 = ( n1422 & ~n1423 ) | ( n1422 & n1672 ) | ( ~n1423 & n1672 ) ;
  assign n1674 = ( n1411 & n1412 ) | ( n1411 & ~n1430 ) | ( n1412 & ~n1430 ) ;
  assign n1675 = ~x132 & n1674 ;
  assign n1676 = ( n1439 & ~n1440 ) | ( n1439 & n1675 ) | ( ~n1440 & n1675 ) ;
  assign n1677 = x134 & ~n1676 ;
  assign n1678 = x134 & ~n1673 ;
  assign n1679 = ( n1673 & ~n1677 ) | ( n1673 & n1678 ) | ( ~n1677 & n1678 ) ;
  assign n1680 = ( ~n1450 & n1465 ) | ( ~n1450 & n1466 ) | ( n1465 & n1466 ) ;
  assign n1681 = ~x132 & n1680 ;
  assign n1682 = ( n1459 & ~n1460 ) | ( n1459 & n1681 ) | ( ~n1460 & n1681 ) ;
  assign n1683 = ( n1448 & n1449 ) | ( n1448 & ~n1467 ) | ( n1449 & ~n1467 ) ;
  assign n1684 = ~x132 & n1683 ;
  assign n1685 = ( n1476 & ~n1477 ) | ( n1476 & n1684 ) | ( ~n1477 & n1684 ) ;
  assign n1686 = x134 & ~n1685 ;
  assign n1687 = x134 & ~n1682 ;
  assign n1688 = ( n1682 & ~n1686 ) | ( n1682 & n1687 ) | ( ~n1686 & n1687 ) ;
  assign n1689 = ( ~n1487 & n1502 ) | ( ~n1487 & n1503 ) | ( n1502 & n1503 ) ;
  assign n1690 = ~x132 & n1689 ;
  assign n1691 = ( n1496 & ~n1497 ) | ( n1496 & n1690 ) | ( ~n1497 & n1690 ) ;
  assign n1692 = ( n1485 & n1486 ) | ( n1485 & ~n1504 ) | ( n1486 & ~n1504 ) ;
  assign n1693 = ~x132 & n1692 ;
  assign n1694 = ( n1513 & ~n1514 ) | ( n1513 & n1693 ) | ( ~n1514 & n1693 ) ;
  assign n1695 = x134 & ~n1694 ;
  assign n1696 = x134 & ~n1691 ;
  assign n1697 = ( n1691 & ~n1695 ) | ( n1691 & n1696 ) | ( ~n1695 & n1696 ) ;
  assign n1698 = ( ~n1524 & n1539 ) | ( ~n1524 & n1540 ) | ( n1539 & n1540 ) ;
  assign n1699 = ~x132 & n1698 ;
  assign n1700 = ( n1533 & ~n1534 ) | ( n1533 & n1699 ) | ( ~n1534 & n1699 ) ;
  assign n1701 = ( n1522 & n1523 ) | ( n1522 & ~n1541 ) | ( n1523 & ~n1541 ) ;
  assign n1702 = ~x132 & n1701 ;
  assign n1703 = ( n1550 & ~n1551 ) | ( n1550 & n1702 ) | ( ~n1551 & n1702 ) ;
  assign n1704 = x134 & ~n1703 ;
  assign n1705 = x134 & ~n1700 ;
  assign n1706 = ( n1700 & ~n1704 ) | ( n1700 & n1705 ) | ( ~n1704 & n1705 ) ;
  assign n1707 = ( ~n305 & n476 ) | ( ~n305 & n477 ) | ( n476 & n477 ) ;
  assign n1708 = ~x132 & n1707 ;
  assign n1709 = ( n1556 & ~n1557 ) | ( n1556 & n1708 ) | ( ~n1557 & n1708 ) ;
  assign n1710 = ( n303 & n304 ) | ( n303 & ~n478 ) | ( n304 & ~n478 ) ;
  assign n1711 = ~x132 & n1710 ;
  assign n1712 = ( n1559 & ~n1560 ) | ( n1559 & n1711 ) | ( ~n1560 & n1711 ) ;
  assign n1713 = x134 & ~n1712 ;
  assign n1714 = x134 & ~n1709 ;
  assign n1715 = ( n1709 & ~n1713 ) | ( n1709 & n1714 ) | ( ~n1713 & n1714 ) ;
  assign n1716 = ( ~n622 & n761 ) | ( ~n622 & n762 ) | ( n761 & n762 ) ;
  assign n1717 = ~x132 & n1716 ;
  assign n1718 = ( n1565 & ~n1566 ) | ( n1565 & n1717 ) | ( ~n1566 & n1717 ) ;
  assign n1719 = ( n620 & n621 ) | ( n620 & ~n763 ) | ( n621 & ~n763 ) ;
  assign n1720 = ~x132 & n1719 ;
  assign n1721 = ( n1568 & ~n1569 ) | ( n1568 & n1720 ) | ( ~n1569 & n1720 ) ;
  assign n1722 = x134 & ~n1721 ;
  assign n1723 = x134 & ~n1718 ;
  assign n1724 = ( n1718 & ~n1722 ) | ( n1718 & n1723 ) | ( ~n1722 & n1723 ) ;
  assign n1725 = ~x133 & n916 ;
  assign n1726 = ( n823 & ~n824 ) | ( n823 & n1725 ) | ( ~n824 & n1725 ) ;
  assign n1727 = ~x132 & n1726 ;
  assign n1728 = ( n1584 & ~n1585 ) | ( n1584 & n1727 ) | ( ~n1585 & n1727 ) ;
  assign n1729 = ~x133 & n841 ;
  assign n1730 = ( n879 & ~n1574 ) | ( n879 & n1729 ) | ( ~n1574 & n1729 ) ;
  assign n1731 = x132 | n1730 ;
  assign n1732 = ( n1576 & ~n1577 ) | ( n1576 & n1731 ) | ( ~n1577 & n1731 ) ;
  assign n1733 = x134 & ~n1732 ;
  assign n1734 = x134 & ~n1728 ;
  assign n1735 = ( n1728 & ~n1733 ) | ( n1728 & n1734 ) | ( ~n1733 & n1734 ) ;
  assign n1736 = ( ~n980 & n1039 ) | ( ~n980 & n1040 ) | ( n1039 & n1040 ) ;
  assign n1737 = ~x132 & n1736 ;
  assign n1738 = ( n1589 & ~n1590 ) | ( n1589 & n1737 ) | ( ~n1590 & n1737 ) ;
  assign n1739 = ( n978 & n979 ) | ( n978 & ~n1041 ) | ( n979 & ~n1041 ) ;
  assign n1740 = ~x132 & n1739 ;
  assign n1741 = ( n1592 & ~n1593 ) | ( n1592 & n1740 ) | ( ~n1593 & n1740 ) ;
  assign n1742 = x134 & ~n1741 ;
  assign n1743 = x134 & ~n1738 ;
  assign n1744 = ( n1738 & ~n1742 ) | ( n1738 & n1743 ) | ( ~n1742 & n1743 ) ;
  assign n1745 = ( ~n1065 & n1084 ) | ( ~n1065 & n1085 ) | ( n1084 & n1085 ) ;
  assign n1746 = ~x132 & n1745 ;
  assign n1747 = ( n1598 & ~n1599 ) | ( n1598 & n1746 ) | ( ~n1599 & n1746 ) ;
  assign n1748 = ( n1063 & n1064 ) | ( n1063 & ~n1086 ) | ( n1064 & ~n1086 ) ;
  assign n1749 = ~x132 & n1748 ;
  assign n1750 = ( n1601 & ~n1602 ) | ( n1601 & n1749 ) | ( ~n1602 & n1749 ) ;
  assign n1751 = x134 & ~n1750 ;
  assign n1752 = x134 & ~n1747 ;
  assign n1753 = ( n1747 & ~n1751 ) | ( n1747 & n1752 ) | ( ~n1751 & n1752 ) ;
  assign n1754 = ( ~n1110 & n1129 ) | ( ~n1110 & n1130 ) | ( n1129 & n1130 ) ;
  assign n1755 = ~x132 & n1754 ;
  assign n1756 = ( n1607 & ~n1608 ) | ( n1607 & n1755 ) | ( ~n1608 & n1755 ) ;
  assign n1757 = ( n1108 & n1109 ) | ( n1108 & ~n1131 ) | ( n1109 & ~n1131 ) ;
  assign n1758 = ~x132 & n1757 ;
  assign n1759 = ( n1610 & ~n1611 ) | ( n1610 & n1758 ) | ( ~n1611 & n1758 ) ;
  assign n1760 = x134 & ~n1759 ;
  assign n1761 = x134 & ~n1756 ;
  assign n1762 = ( n1756 & ~n1760 ) | ( n1756 & n1761 ) | ( ~n1760 & n1761 ) ;
  assign n1763 = ( ~n1155 & n1174 ) | ( ~n1155 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1764 = ~x132 & n1763 ;
  assign n1765 = ( n1616 & ~n1617 ) | ( n1616 & n1764 ) | ( ~n1617 & n1764 ) ;
  assign n1766 = ( n1153 & n1154 ) | ( n1153 & ~n1176 ) | ( n1154 & ~n1176 ) ;
  assign n1767 = ~x132 & n1766 ;
  assign n1768 = ( n1619 & ~n1620 ) | ( n1619 & n1767 ) | ( ~n1620 & n1767 ) ;
  assign n1769 = x134 & ~n1768 ;
  assign n1770 = x134 & ~n1765 ;
  assign n1771 = ( n1765 & ~n1769 ) | ( n1765 & n1770 ) | ( ~n1769 & n1770 ) ;
  assign n1772 = ( ~n1190 & n1220 ) | ( ~n1190 & n1221 ) | ( n1220 & n1221 ) ;
  assign n1773 = ~x132 & n1772 ;
  assign n1774 = ( n1630 & ~n1631 ) | ( n1630 & n1773 ) | ( ~n1631 & n1773 ) ;
  assign n1775 = x132 & x133 ;
  assign n1776 = n1206 & n1775 ;
  assign n1777 = x132 & ~x133 ;
  assign n1778 = n1198 & n1777 ;
  assign n1779 = x132 | x133 ;
  assign n1780 = n1188 & ~n1779 ;
  assign n1781 = ~x132 & x133 ;
  assign n1782 = n1216 & n1781 ;
  assign n1783 = ( ~n1776 & n1780 ) | ( ~n1776 & n1782 ) | ( n1780 & n1782 ) ;
  assign n1784 = ( ~n1776 & n1778 ) | ( ~n1776 & n1783 ) | ( n1778 & n1783 ) ;
  assign n1785 = n1776 | n1784 ;
  assign n1786 = x134 & ~n1785 ;
  assign n1787 = x134 & ~n1774 ;
  assign n1788 = ( n1774 & ~n1786 ) | ( n1774 & n1787 ) | ( ~n1786 & n1787 ) ;
  assign n1789 = ( ~n1245 & n1264 ) | ( ~n1245 & n1265 ) | ( n1264 & n1265 ) ;
  assign n1790 = ~x132 & n1789 ;
  assign n1791 = ( n1635 & ~n1636 ) | ( n1635 & n1790 ) | ( ~n1636 & n1790 ) ;
  assign n1792 = ( n1243 & n1244 ) | ( n1243 & ~n1266 ) | ( n1244 & ~n1266 ) ;
  assign n1793 = ~x132 & n1792 ;
  assign n1794 = ( n1638 & ~n1639 ) | ( n1638 & n1793 ) | ( ~n1639 & n1793 ) ;
  assign n1795 = x134 & ~n1794 ;
  assign n1796 = x134 & ~n1791 ;
  assign n1797 = ( n1791 & ~n1795 ) | ( n1791 & n1796 ) | ( ~n1795 & n1796 ) ;
  assign n1798 = ( ~n1290 & n1309 ) | ( ~n1290 & n1310 ) | ( n1309 & n1310 ) ;
  assign n1799 = ~x132 & n1798 ;
  assign n1800 = ( n1644 & ~n1645 ) | ( n1644 & n1799 ) | ( ~n1645 & n1799 ) ;
  assign n1801 = ( n1288 & n1289 ) | ( n1288 & ~n1311 ) | ( n1289 & ~n1311 ) ;
  assign n1802 = ~x132 & n1801 ;
  assign n1803 = ( n1647 & ~n1648 ) | ( n1647 & n1802 ) | ( ~n1648 & n1802 ) ;
  assign n1804 = x134 & ~n1803 ;
  assign n1805 = x134 & ~n1800 ;
  assign n1806 = ( n1800 & ~n1804 ) | ( n1800 & n1805 ) | ( ~n1804 & n1805 ) ;
  assign n1807 = ( ~n1335 & n1354 ) | ( ~n1335 & n1355 ) | ( n1354 & n1355 ) ;
  assign n1808 = ~x132 & n1807 ;
  assign n1809 = ( n1653 & ~n1654 ) | ( n1653 & n1808 ) | ( ~n1654 & n1808 ) ;
  assign n1810 = ( n1333 & n1334 ) | ( n1333 & ~n1356 ) | ( n1334 & ~n1356 ) ;
  assign n1811 = ~x132 & n1810 ;
  assign n1812 = ( n1656 & ~n1657 ) | ( n1656 & n1811 ) | ( ~n1657 & n1811 ) ;
  assign n1813 = x134 & ~n1812 ;
  assign n1814 = x134 & ~n1809 ;
  assign n1815 = ( n1809 & ~n1813 ) | ( n1809 & n1814 ) | ( ~n1813 & n1814 ) ;
  assign n1816 = ( ~n1380 & n1399 ) | ( ~n1380 & n1400 ) | ( n1399 & n1400 ) ;
  assign n1817 = ~x132 & n1816 ;
  assign n1818 = ( n1662 & ~n1663 ) | ( n1662 & n1817 ) | ( ~n1663 & n1817 ) ;
  assign n1819 = ( n1378 & n1379 ) | ( n1378 & ~n1401 ) | ( n1379 & ~n1401 ) ;
  assign n1820 = ~x132 & n1819 ;
  assign n1821 = ( n1665 & ~n1666 ) | ( n1665 & n1820 ) | ( ~n1666 & n1820 ) ;
  assign n1822 = x134 & ~n1821 ;
  assign n1823 = x134 & ~n1818 ;
  assign n1824 = ( n1818 & ~n1822 ) | ( n1818 & n1823 ) | ( ~n1822 & n1823 ) ;
  assign n1825 = ( ~n1421 & n1436 ) | ( ~n1421 & n1437 ) | ( n1436 & n1437 ) ;
  assign n1826 = ~x132 & n1825 ;
  assign n1827 = ( n1671 & ~n1672 ) | ( n1671 & n1826 ) | ( ~n1672 & n1826 ) ;
  assign n1828 = ( n1419 & n1420 ) | ( n1419 & ~n1438 ) | ( n1420 & ~n1438 ) ;
  assign n1829 = ~x132 & n1828 ;
  assign n1830 = ( n1674 & ~n1675 ) | ( n1674 & n1829 ) | ( ~n1675 & n1829 ) ;
  assign n1831 = x134 & ~n1830 ;
  assign n1832 = x134 & ~n1827 ;
  assign n1833 = ( n1827 & ~n1831 ) | ( n1827 & n1832 ) | ( ~n1831 & n1832 ) ;
  assign n1834 = ( ~n1458 & n1473 ) | ( ~n1458 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1835 = ~x132 & n1834 ;
  assign n1836 = ( n1680 & ~n1681 ) | ( n1680 & n1835 ) | ( ~n1681 & n1835 ) ;
  assign n1837 = ( n1456 & n1457 ) | ( n1456 & ~n1475 ) | ( n1457 & ~n1475 ) ;
  assign n1838 = ~x132 & n1837 ;
  assign n1839 = ( n1683 & ~n1684 ) | ( n1683 & n1838 ) | ( ~n1684 & n1838 ) ;
  assign n1840 = x134 & ~n1839 ;
  assign n1841 = x134 & ~n1836 ;
  assign n1842 = ( n1836 & ~n1840 ) | ( n1836 & n1841 ) | ( ~n1840 & n1841 ) ;
  assign n1843 = ( ~n1495 & n1510 ) | ( ~n1495 & n1511 ) | ( n1510 & n1511 ) ;
  assign n1844 = ~x132 & n1843 ;
  assign n1845 = ( n1689 & ~n1690 ) | ( n1689 & n1844 ) | ( ~n1690 & n1844 ) ;
  assign n1846 = ( n1493 & n1494 ) | ( n1493 & ~n1512 ) | ( n1494 & ~n1512 ) ;
  assign n1847 = ~x132 & n1846 ;
  assign n1848 = ( n1692 & ~n1693 ) | ( n1692 & n1847 ) | ( ~n1693 & n1847 ) ;
  assign n1849 = x134 & ~n1848 ;
  assign n1850 = x134 & ~n1845 ;
  assign n1851 = ( n1845 & ~n1849 ) | ( n1845 & n1850 ) | ( ~n1849 & n1850 ) ;
  assign n1852 = ( ~n1532 & n1547 ) | ( ~n1532 & n1548 ) | ( n1547 & n1548 ) ;
  assign n1853 = ~x132 & n1852 ;
  assign n1854 = ( n1698 & ~n1699 ) | ( n1698 & n1853 ) | ( ~n1699 & n1853 ) ;
  assign n1855 = ( n1530 & n1531 ) | ( n1530 & ~n1549 ) | ( n1531 & ~n1549 ) ;
  assign n1856 = ~x132 & n1855 ;
  assign n1857 = ( n1701 & ~n1702 ) | ( n1701 & n1856 ) | ( ~n1702 & n1856 ) ;
  assign n1858 = x134 & ~n1857 ;
  assign n1859 = x134 & ~n1854 ;
  assign n1860 = ( n1854 & ~n1858 ) | ( n1854 & n1859 ) | ( ~n1858 & n1859 ) ;
  assign n1861 = x132 & ~n1707 ;
  assign n1862 = ( n393 & n394 ) | ( n393 & ~n1861 ) | ( n394 & ~n1861 ) ;
  assign n1863 = x132 & ~n1710 ;
  assign n1864 = ( n220 & n221 ) | ( n220 & ~n1863 ) | ( n221 & ~n1863 ) ;
  assign n1865 = x134 & ~n1864 ;
  assign n1866 = x134 & ~n1862 ;
  assign n1867 = ( n1862 & ~n1865 ) | ( n1862 & n1866 ) | ( ~n1865 & n1866 ) ;
  assign n1868 = x132 & ~n1716 ;
  assign n1869 = ( n694 & n695 ) | ( n694 & ~n1868 ) | ( n695 & ~n1868 ) ;
  assign n1870 = x132 & ~n1719 ;
  assign n1871 = ( n553 & n554 ) | ( n553 & ~n1870 ) | ( n554 & ~n1870 ) ;
  assign n1872 = x134 & ~n1871 ;
  assign n1873 = x134 & ~n1869 ;
  assign n1874 = ( n1869 & ~n1872 ) | ( n1869 & n1873 ) | ( ~n1872 & n1873 ) ;
  assign n1875 = n861 & ~n1779 ;
  assign n1876 = n898 & n1781 ;
  assign n1877 = ( n1726 & ~n1727 ) | ( n1726 & n1876 ) | ( ~n1727 & n1876 ) ;
  assign n1878 = n1875 | n1877 ;
  assign n1879 = ( x132 & n787 ) | ( x132 & ~n805 ) | ( n787 & ~n805 ) ;
  assign n1880 = x132 & ~n1730 ;
  assign n1881 = ( n805 & n1879 ) | ( n805 & ~n1880 ) | ( n1879 & ~n1880 ) ;
  assign n1882 = x134 & ~n1881 ;
  assign n1883 = x134 & ~n1878 ;
  assign n1884 = ( n1878 & ~n1882 ) | ( n1878 & n1883 ) | ( ~n1882 & n1883 ) ;
  assign n1885 = x132 & ~n1736 ;
  assign n1886 = ( n1012 & n1013 ) | ( n1012 & ~n1885 ) | ( n1013 & ~n1885 ) ;
  assign n1887 = x132 & ~n1739 ;
  assign n1888 = ( n951 & n952 ) | ( n951 & ~n1887 ) | ( n952 & ~n1887 ) ;
  assign n1889 = x134 & ~n1888 ;
  assign n1890 = x134 & ~n1886 ;
  assign n1891 = ( n1886 & ~n1889 ) | ( n1886 & n1890 ) | ( ~n1889 & n1890 ) ;
  assign n1892 = x132 & ~n1745 ;
  assign n1893 = ( n1077 & n1078 ) | ( n1077 & ~n1892 ) | ( n1078 & ~n1892 ) ;
  assign n1894 = x132 & ~n1748 ;
  assign n1895 = ( n1056 & n1057 ) | ( n1056 & ~n1894 ) | ( n1057 & ~n1894 ) ;
  assign n1896 = x134 & ~n1895 ;
  assign n1897 = x134 & ~n1893 ;
  assign n1898 = ( n1893 & ~n1896 ) | ( n1893 & n1897 ) | ( ~n1896 & n1897 ) ;
  assign n1899 = x132 & ~n1754 ;
  assign n1900 = ( n1122 & n1123 ) | ( n1122 & ~n1899 ) | ( n1123 & ~n1899 ) ;
  assign n1901 = x132 & ~n1757 ;
  assign n1902 = ( n1101 & n1102 ) | ( n1101 & ~n1901 ) | ( n1102 & ~n1901 ) ;
  assign n1903 = x134 & ~n1902 ;
  assign n1904 = x134 & ~n1900 ;
  assign n1905 = ( n1900 & ~n1903 ) | ( n1900 & n1904 ) | ( ~n1903 & n1904 ) ;
  assign n1906 = x132 & ~n1763 ;
  assign n1907 = ( n1167 & n1168 ) | ( n1167 & ~n1906 ) | ( n1168 & ~n1906 ) ;
  assign n1908 = x132 & ~n1766 ;
  assign n1909 = ( n1146 & n1147 ) | ( n1146 & ~n1908 ) | ( n1147 & ~n1908 ) ;
  assign n1910 = x134 & ~n1909 ;
  assign n1911 = x134 & ~n1907 ;
  assign n1912 = ( n1907 & ~n1910 ) | ( n1907 & n1911 ) | ( ~n1910 & n1911 ) ;
  assign n1913 = n1216 & n1775 ;
  assign n1914 = n1188 & n1777 ;
  assign n1915 = ( n1201 & ~n1202 ) | ( n1201 & n1914 ) | ( ~n1202 & n1914 ) ;
  assign n1916 = n1913 | n1915 ;
  assign n1917 = x132 & ~n1772 ;
  assign n1918 = ( n1212 & n1213 ) | ( n1212 & ~n1917 ) | ( n1213 & ~n1917 ) ;
  assign n1919 = x134 | n1918 ;
  assign n1920 = x134 | n1916 ;
  assign n1921 = ( n1916 & n1919 ) | ( n1916 & ~n1920 ) | ( n1919 & ~n1920 ) ;
  assign n1922 = x132 & ~n1789 ;
  assign n1923 = ( n1257 & n1258 ) | ( n1257 & ~n1922 ) | ( n1258 & ~n1922 ) ;
  assign n1924 = x132 & ~n1792 ;
  assign n1925 = ( n1236 & n1237 ) | ( n1236 & ~n1924 ) | ( n1237 & ~n1924 ) ;
  assign n1926 = x134 & ~n1925 ;
  assign n1927 = x134 & ~n1923 ;
  assign n1928 = ( n1923 & ~n1926 ) | ( n1923 & n1927 ) | ( ~n1926 & n1927 ) ;
  assign n1929 = x132 & ~n1798 ;
  assign n1930 = ( n1302 & n1303 ) | ( n1302 & ~n1929 ) | ( n1303 & ~n1929 ) ;
  assign n1931 = x132 & ~n1801 ;
  assign n1932 = ( n1281 & n1282 ) | ( n1281 & ~n1931 ) | ( n1282 & ~n1931 ) ;
  assign n1933 = x134 & ~n1932 ;
  assign n1934 = x134 & ~n1930 ;
  assign n1935 = ( n1930 & ~n1933 ) | ( n1930 & n1934 ) | ( ~n1933 & n1934 ) ;
  assign n1936 = x132 & ~n1807 ;
  assign n1937 = ( n1347 & n1348 ) | ( n1347 & ~n1936 ) | ( n1348 & ~n1936 ) ;
  assign n1938 = x132 & ~n1810 ;
  assign n1939 = ( n1326 & n1327 ) | ( n1326 & ~n1938 ) | ( n1327 & ~n1938 ) ;
  assign n1940 = x134 & ~n1939 ;
  assign n1941 = x134 & ~n1937 ;
  assign n1942 = ( n1937 & ~n1940 ) | ( n1937 & n1941 ) | ( ~n1940 & n1941 ) ;
  assign n1943 = x132 & ~n1816 ;
  assign n1944 = ( n1392 & n1393 ) | ( n1392 & ~n1943 ) | ( n1393 & ~n1943 ) ;
  assign n1945 = x132 & ~n1819 ;
  assign n1946 = ( n1371 & n1372 ) | ( n1371 & ~n1945 ) | ( n1372 & ~n1945 ) ;
  assign n1947 = x134 & ~n1946 ;
  assign n1948 = x134 & ~n1944 ;
  assign n1949 = ( n1944 & ~n1947 ) | ( n1944 & n1948 ) | ( ~n1947 & n1948 ) ;
  assign n1950 = x132 & ~n1825 ;
  assign n1951 = ( n1431 & n1432 ) | ( n1431 & ~n1950 ) | ( n1432 & ~n1950 ) ;
  assign n1952 = x132 & ~n1828 ;
  assign n1953 = ( n1414 & n1415 ) | ( n1414 & ~n1952 ) | ( n1415 & ~n1952 ) ;
  assign n1954 = x134 & ~n1953 ;
  assign n1955 = x134 & ~n1951 ;
  assign n1956 = ( n1951 & ~n1954 ) | ( n1951 & n1955 ) | ( ~n1954 & n1955 ) ;
  assign n1957 = x132 & ~n1834 ;
  assign n1958 = ( n1468 & n1469 ) | ( n1468 & ~n1957 ) | ( n1469 & ~n1957 ) ;
  assign n1959 = x132 & ~n1837 ;
  assign n1960 = ( n1451 & n1452 ) | ( n1451 & ~n1959 ) | ( n1452 & ~n1959 ) ;
  assign n1961 = x134 & ~n1960 ;
  assign n1962 = x134 & ~n1958 ;
  assign n1963 = ( n1958 & ~n1961 ) | ( n1958 & n1962 ) | ( ~n1961 & n1962 ) ;
  assign n1964 = x132 & ~n1843 ;
  assign n1965 = ( n1505 & n1506 ) | ( n1505 & ~n1964 ) | ( n1506 & ~n1964 ) ;
  assign n1966 = x132 & ~n1846 ;
  assign n1967 = ( n1488 & n1489 ) | ( n1488 & ~n1966 ) | ( n1489 & ~n1966 ) ;
  assign n1968 = x134 & ~n1967 ;
  assign n1969 = x134 & ~n1965 ;
  assign n1970 = ( n1965 & ~n1968 ) | ( n1965 & n1969 ) | ( ~n1968 & n1969 ) ;
  assign n1971 = x132 & ~n1852 ;
  assign n1972 = ( n1542 & n1543 ) | ( n1542 & ~n1971 ) | ( n1543 & ~n1971 ) ;
  assign n1973 = x132 & ~n1855 ;
  assign n1974 = ( n1525 & n1526 ) | ( n1525 & ~n1973 ) | ( n1526 & ~n1973 ) ;
  assign n1975 = x134 & ~n1974 ;
  assign n1976 = x134 & ~n1972 ;
  assign n1977 = ( n1972 & ~n1975 ) | ( n1972 & n1976 ) | ( ~n1975 & n1976 ) ;
  assign n1978 = ( n481 & n482 ) | ( n481 & ~n483 ) | ( n482 & ~n483 ) ;
  assign n1979 = ( n766 & n767 ) | ( n766 & ~n768 ) | ( n767 & ~n768 ) ;
  assign n1980 = ( n919 & n920 ) | ( n919 & ~n921 ) | ( n920 & ~n921 ) ;
  assign n1981 = ( n1044 & n1045 ) | ( n1044 & ~n1046 ) | ( n1045 & ~n1046 ) ;
  assign n1982 = ( n1089 & n1090 ) | ( n1089 & ~n1091 ) | ( n1090 & ~n1091 ) ;
  assign n1983 = ( n1134 & n1135 ) | ( n1134 & ~n1136 ) | ( n1135 & ~n1136 ) ;
  assign n1984 = ( n1179 & n1180 ) | ( n1179 & ~n1181 ) | ( n1180 & ~n1181 ) ;
  assign n1985 = ( n1224 & n1225 ) | ( n1224 & ~n1226 ) | ( n1225 & ~n1226 ) ;
  assign n1986 = ( n1269 & n1270 ) | ( n1269 & ~n1271 ) | ( n1270 & ~n1271 ) ;
  assign n1987 = ( n1314 & n1315 ) | ( n1314 & ~n1316 ) | ( n1315 & ~n1316 ) ;
  assign n1988 = ( n1359 & n1360 ) | ( n1359 & ~n1361 ) | ( n1360 & ~n1361 ) ;
  assign n1989 = ( n1404 & n1405 ) | ( n1404 & ~n1406 ) | ( n1405 & ~n1406 ) ;
  assign n1990 = ( n1441 & n1442 ) | ( n1441 & ~n1443 ) | ( n1442 & ~n1443 ) ;
  assign n1991 = ( n1478 & n1479 ) | ( n1478 & ~n1480 ) | ( n1479 & ~n1480 ) ;
  assign n1992 = ( n1515 & n1516 ) | ( n1515 & ~n1517 ) | ( n1516 & ~n1517 ) ;
  assign n1993 = ( n1552 & n1553 ) | ( n1552 & ~n1554 ) | ( n1553 & ~n1554 ) ;
  assign n1994 = ( n1561 & n1562 ) | ( n1561 & ~n1563 ) | ( n1562 & ~n1563 ) ;
  assign n1995 = ( n1570 & n1571 ) | ( n1570 & ~n1572 ) | ( n1571 & ~n1572 ) ;
  assign n1996 = ( n1580 & n1581 ) | ( n1580 & ~n1587 ) | ( n1581 & ~n1587 ) ;
  assign n1997 = ( n1594 & n1595 ) | ( n1594 & ~n1596 ) | ( n1595 & ~n1596 ) ;
  assign n1998 = ( n1603 & n1604 ) | ( n1603 & ~n1605 ) | ( n1604 & ~n1605 ) ;
  assign n1999 = ( n1612 & n1613 ) | ( n1612 & ~n1614 ) | ( n1613 & ~n1614 ) ;
  assign n2000 = ( n1621 & n1622 ) | ( n1621 & ~n1623 ) | ( n1622 & ~n1623 ) ;
  assign n2001 = ( n1628 & n1629 ) | ( n1628 & ~n1633 ) | ( n1629 & ~n1633 ) ;
  assign n2002 = ( n1640 & n1641 ) | ( n1640 & ~n1642 ) | ( n1641 & ~n1642 ) ;
  assign n2003 = ( n1649 & n1650 ) | ( n1649 & ~n1651 ) | ( n1650 & ~n1651 ) ;
  assign n2004 = ( n1658 & n1659 ) | ( n1658 & ~n1660 ) | ( n1659 & ~n1660 ) ;
  assign n2005 = ( n1667 & n1668 ) | ( n1667 & ~n1669 ) | ( n1668 & ~n1669 ) ;
  assign n2006 = ( n1676 & n1677 ) | ( n1676 & ~n1678 ) | ( n1677 & ~n1678 ) ;
  assign n2007 = ( n1685 & n1686 ) | ( n1685 & ~n1687 ) | ( n1686 & ~n1687 ) ;
  assign n2008 = ( n1694 & n1695 ) | ( n1694 & ~n1696 ) | ( n1695 & ~n1696 ) ;
  assign n2009 = ( n1703 & n1704 ) | ( n1703 & ~n1705 ) | ( n1704 & ~n1705 ) ;
  assign n2010 = ( n1712 & n1713 ) | ( n1712 & ~n1714 ) | ( n1713 & ~n1714 ) ;
  assign n2011 = ( n1721 & n1722 ) | ( n1721 & ~n1723 ) | ( n1722 & ~n1723 ) ;
  assign n2012 = ( n1732 & n1733 ) | ( n1732 & ~n1734 ) | ( n1733 & ~n1734 ) ;
  assign n2013 = ( n1741 & n1742 ) | ( n1741 & ~n1743 ) | ( n1742 & ~n1743 ) ;
  assign n2014 = ( n1750 & n1751 ) | ( n1750 & ~n1752 ) | ( n1751 & ~n1752 ) ;
  assign n2015 = ( n1759 & n1760 ) | ( n1759 & ~n1761 ) | ( n1760 & ~n1761 ) ;
  assign n2016 = ( n1768 & n1769 ) | ( n1768 & ~n1770 ) | ( n1769 & ~n1770 ) ;
  assign n2017 = ( n1785 & n1786 ) | ( n1785 & ~n1787 ) | ( n1786 & ~n1787 ) ;
  assign n2018 = ( n1794 & n1795 ) | ( n1794 & ~n1796 ) | ( n1795 & ~n1796 ) ;
  assign n2019 = ( n1803 & n1804 ) | ( n1803 & ~n1805 ) | ( n1804 & ~n1805 ) ;
  assign n2020 = ( n1812 & n1813 ) | ( n1812 & ~n1814 ) | ( n1813 & ~n1814 ) ;
  assign n2021 = ( n1821 & n1822 ) | ( n1821 & ~n1823 ) | ( n1822 & ~n1823 ) ;
  assign n2022 = ( n1830 & n1831 ) | ( n1830 & ~n1832 ) | ( n1831 & ~n1832 ) ;
  assign n2023 = ( n1839 & n1840 ) | ( n1839 & ~n1841 ) | ( n1840 & ~n1841 ) ;
  assign n2024 = ( n1848 & n1849 ) | ( n1848 & ~n1850 ) | ( n1849 & ~n1850 ) ;
  assign n2025 = ( n1857 & n1858 ) | ( n1857 & ~n1859 ) | ( n1858 & ~n1859 ) ;
  assign n2026 = ( n1864 & n1865 ) | ( n1864 & ~n1866 ) | ( n1865 & ~n1866 ) ;
  assign n2027 = ( n1871 & n1872 ) | ( n1871 & ~n1873 ) | ( n1872 & ~n1873 ) ;
  assign n2028 = ( n1881 & n1882 ) | ( n1881 & ~n1883 ) | ( n1882 & ~n1883 ) ;
  assign n2029 = ( n1888 & n1889 ) | ( n1888 & ~n1890 ) | ( n1889 & ~n1890 ) ;
  assign n2030 = ( n1895 & n1896 ) | ( n1895 & ~n1897 ) | ( n1896 & ~n1897 ) ;
  assign n2031 = ( n1902 & n1903 ) | ( n1902 & ~n1904 ) | ( n1903 & ~n1904 ) ;
  assign n2032 = ( n1909 & n1910 ) | ( n1909 & ~n1911 ) | ( n1910 & ~n1911 ) ;
  assign n2033 = ( n1918 & ~n1919 ) | ( n1918 & n1920 ) | ( ~n1919 & n1920 ) ;
  assign n2034 = ( n1925 & n1926 ) | ( n1925 & ~n1927 ) | ( n1926 & ~n1927 ) ;
  assign n2035 = ( n1932 & n1933 ) | ( n1932 & ~n1934 ) | ( n1933 & ~n1934 ) ;
  assign n2036 = ( n1939 & n1940 ) | ( n1939 & ~n1941 ) | ( n1940 & ~n1941 ) ;
  assign n2037 = ( n1946 & n1947 ) | ( n1946 & ~n1948 ) | ( n1947 & ~n1948 ) ;
  assign n2038 = ( n1953 & n1954 ) | ( n1953 & ~n1955 ) | ( n1954 & ~n1955 ) ;
  assign n2039 = ( n1960 & n1961 ) | ( n1960 & ~n1962 ) | ( n1961 & ~n1962 ) ;
  assign n2040 = ( n1967 & n1968 ) | ( n1967 & ~n1969 ) | ( n1968 & ~n1969 ) ;
  assign n2041 = ( n1974 & n1975 ) | ( n1974 & ~n1976 ) | ( n1975 & ~n1976 ) ;
  assign y0 = n484 ;
  assign y1 = n769 ;
  assign y2 = n922 ;
  assign y3 = n1047 ;
  assign y4 = n1092 ;
  assign y5 = n1137 ;
  assign y6 = n1182 ;
  assign y7 = n1227 ;
  assign y8 = n1272 ;
  assign y9 = n1317 ;
  assign y10 = n1362 ;
  assign y11 = n1407 ;
  assign y12 = n1444 ;
  assign y13 = n1481 ;
  assign y14 = n1518 ;
  assign y15 = n1555 ;
  assign y16 = n1564 ;
  assign y17 = n1573 ;
  assign y18 = n1588 ;
  assign y19 = n1597 ;
  assign y20 = n1606 ;
  assign y21 = n1615 ;
  assign y22 = n1624 ;
  assign y23 = n1634 ;
  assign y24 = n1643 ;
  assign y25 = n1652 ;
  assign y26 = n1661 ;
  assign y27 = n1670 ;
  assign y28 = n1679 ;
  assign y29 = n1688 ;
  assign y30 = n1697 ;
  assign y31 = n1706 ;
  assign y32 = n1715 ;
  assign y33 = n1724 ;
  assign y34 = n1735 ;
  assign y35 = n1744 ;
  assign y36 = n1753 ;
  assign y37 = n1762 ;
  assign y38 = n1771 ;
  assign y39 = n1788 ;
  assign y40 = n1797 ;
  assign y41 = n1806 ;
  assign y42 = n1815 ;
  assign y43 = n1824 ;
  assign y44 = n1833 ;
  assign y45 = n1842 ;
  assign y46 = n1851 ;
  assign y47 = n1860 ;
  assign y48 = n1867 ;
  assign y49 = n1874 ;
  assign y50 = n1884 ;
  assign y51 = n1891 ;
  assign y52 = n1898 ;
  assign y53 = n1905 ;
  assign y54 = n1912 ;
  assign y55 = n1921 ;
  assign y56 = n1928 ;
  assign y57 = n1935 ;
  assign y58 = n1942 ;
  assign y59 = n1949 ;
  assign y60 = n1956 ;
  assign y61 = n1963 ;
  assign y62 = n1970 ;
  assign y63 = n1977 ;
  assign y64 = n1978 ;
  assign y65 = n1979 ;
  assign y66 = n1980 ;
  assign y67 = n1981 ;
  assign y68 = n1982 ;
  assign y69 = n1983 ;
  assign y70 = n1984 ;
  assign y71 = n1985 ;
  assign y72 = n1986 ;
  assign y73 = n1987 ;
  assign y74 = n1988 ;
  assign y75 = n1989 ;
  assign y76 = n1990 ;
  assign y77 = n1991 ;
  assign y78 = n1992 ;
  assign y79 = n1993 ;
  assign y80 = n1994 ;
  assign y81 = n1995 ;
  assign y82 = n1996 ;
  assign y83 = n1997 ;
  assign y84 = n1998 ;
  assign y85 = n1999 ;
  assign y86 = n2000 ;
  assign y87 = n2001 ;
  assign y88 = n2002 ;
  assign y89 = n2003 ;
  assign y90 = n2004 ;
  assign y91 = n2005 ;
  assign y92 = n2006 ;
  assign y93 = n2007 ;
  assign y94 = n2008 ;
  assign y95 = n2009 ;
  assign y96 = n2010 ;
  assign y97 = n2011 ;
  assign y98 = n2012 ;
  assign y99 = n2013 ;
  assign y100 = n2014 ;
  assign y101 = n2015 ;
  assign y102 = n2016 ;
  assign y103 = n2017 ;
  assign y104 = n2018 ;
  assign y105 = n2019 ;
  assign y106 = n2020 ;
  assign y107 = n2021 ;
  assign y108 = n2022 ;
  assign y109 = n2023 ;
  assign y110 = n2024 ;
  assign y111 = n2025 ;
  assign y112 = n2026 ;
  assign y113 = n2027 ;
  assign y114 = n2028 ;
  assign y115 = n2029 ;
  assign y116 = n2030 ;
  assign y117 = n2031 ;
  assign y118 = n2032 ;
  assign y119 = n2033 ;
  assign y120 = n2034 ;
  assign y121 = n2035 ;
  assign y122 = n2036 ;
  assign y123 = n2037 ;
  assign y124 = n2038 ;
  assign y125 = n2039 ;
  assign y126 = n2040 ;
  assign y127 = n2041 ;
endmodule
